magic
tech ihp-sg13g2
magscale 1 2
timestamp 1743692330
<< metal1 >>
rect 1152 9848 45216 9872
rect 1152 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 45216 9848
rect 1152 9784 45216 9808
rect 1851 9680 1893 9689
rect 1851 9640 1852 9680
rect 1892 9640 1893 9680
rect 1851 9631 1893 9640
rect 3003 9680 3045 9689
rect 3003 9640 3004 9680
rect 3044 9640 3045 9680
rect 3003 9631 3045 9640
rect 9627 9680 9669 9689
rect 9627 9640 9628 9680
rect 9668 9640 9669 9680
rect 9627 9631 9669 9640
rect 11163 9680 11205 9689
rect 11163 9640 11164 9680
rect 11204 9640 11205 9680
rect 11163 9631 11205 9640
rect 12699 9680 12741 9689
rect 12699 9640 12700 9680
rect 12740 9640 12741 9680
rect 12699 9631 12741 9640
rect 13851 9680 13893 9689
rect 13851 9640 13852 9680
rect 13892 9640 13893 9680
rect 13851 9631 13893 9640
rect 16155 9680 16197 9689
rect 16155 9640 16156 9680
rect 16196 9640 16197 9680
rect 16155 9631 16197 9640
rect 17307 9680 17349 9689
rect 17307 9640 17308 9680
rect 17348 9640 17349 9680
rect 17307 9631 17349 9640
rect 17691 9680 17733 9689
rect 17691 9640 17692 9680
rect 17732 9640 17733 9680
rect 17691 9631 17733 9640
rect 18459 9680 18501 9689
rect 18459 9640 18460 9680
rect 18500 9640 18501 9680
rect 18459 9631 18501 9640
rect 18843 9680 18885 9689
rect 18843 9640 18844 9680
rect 18884 9640 18885 9680
rect 18843 9631 18885 9640
rect 19611 9680 19653 9689
rect 19611 9640 19612 9680
rect 19652 9640 19653 9680
rect 19611 9631 19653 9640
rect 21531 9680 21573 9689
rect 21531 9640 21532 9680
rect 21572 9640 21573 9680
rect 21531 9631 21573 9640
rect 22683 9680 22725 9689
rect 22683 9640 22684 9680
rect 22724 9640 22725 9680
rect 22683 9631 22725 9640
rect 26619 9680 26661 9689
rect 26619 9640 26620 9680
rect 26660 9640 26661 9680
rect 26619 9631 26661 9640
rect 30075 9680 30117 9689
rect 30075 9640 30076 9680
rect 30116 9640 30117 9680
rect 30075 9631 30117 9640
rect 31227 9680 31269 9689
rect 31227 9640 31228 9680
rect 31268 9640 31269 9680
rect 31227 9631 31269 9640
rect 31995 9680 32037 9689
rect 31995 9640 31996 9680
rect 32036 9640 32037 9680
rect 31995 9631 32037 9640
rect 32763 9680 32805 9689
rect 32763 9640 32764 9680
rect 32804 9640 32805 9680
rect 32763 9631 32805 9640
rect 33531 9680 33573 9689
rect 33531 9640 33532 9680
rect 33572 9640 33573 9680
rect 33531 9631 33573 9640
rect 35451 9680 35493 9689
rect 35451 9640 35452 9680
rect 35492 9640 35493 9680
rect 35451 9631 35493 9640
rect 36219 9680 36261 9689
rect 36219 9640 36220 9680
rect 36260 9640 36261 9680
rect 36219 9631 36261 9640
rect 42843 9680 42885 9689
rect 42843 9640 42844 9680
rect 42884 9640 42885 9680
rect 42843 9631 42885 9640
rect 43227 9680 43269 9689
rect 43227 9640 43228 9680
rect 43268 9640 43269 9680
rect 43227 9631 43269 9640
rect 43611 9680 43653 9689
rect 43611 9640 43612 9680
rect 43652 9640 43653 9680
rect 43611 9631 43653 9640
rect 43995 9680 44037 9689
rect 43995 9640 43996 9680
rect 44036 9640 44037 9680
rect 43995 9631 44037 9640
rect 10011 9596 10053 9605
rect 10011 9556 10012 9596
rect 10052 9556 10053 9596
rect 10011 9547 10053 9556
rect 13083 9596 13125 9605
rect 13083 9556 13084 9596
rect 13124 9556 13125 9596
rect 13083 9547 13125 9556
rect 18075 9596 18117 9605
rect 18075 9556 18076 9596
rect 18116 9556 18117 9596
rect 18075 9547 18117 9556
rect 19227 9596 19269 9605
rect 19227 9556 19228 9596
rect 19268 9556 19269 9596
rect 19227 9547 19269 9556
rect 28923 9596 28965 9605
rect 28923 9556 28924 9596
rect 28964 9556 28965 9596
rect 28923 9547 28965 9556
rect 31611 9596 31653 9605
rect 31611 9556 31612 9596
rect 31652 9556 31653 9596
rect 31611 9547 31653 9556
rect 32379 9596 32421 9605
rect 32379 9556 32380 9596
rect 32420 9556 32421 9596
rect 32379 9547 32421 9556
rect 35835 9596 35877 9605
rect 35835 9556 35836 9596
rect 35876 9556 35877 9596
rect 35835 9547 35877 9556
rect 1227 9512 1269 9521
rect 1227 9472 1228 9512
rect 1268 9472 1269 9512
rect 1227 9463 1269 9472
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2379 9512 2421 9521
rect 2379 9472 2380 9512
rect 2420 9472 2421 9512
rect 2379 9463 2421 9472
rect 2763 9512 2805 9521
rect 2763 9472 2764 9512
rect 2804 9472 2805 9512
rect 2763 9463 2805 9472
rect 3147 9512 3189 9521
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 9387 9512 9429 9521
rect 9387 9472 9388 9512
rect 9428 9472 9429 9512
rect 9387 9463 9429 9472
rect 9771 9512 9813 9521
rect 9771 9472 9772 9512
rect 9812 9472 9813 9512
rect 9771 9463 9813 9472
rect 10155 9512 10197 9521
rect 10155 9472 10156 9512
rect 10196 9472 10197 9512
rect 10155 9463 10197 9472
rect 10395 9512 10437 9521
rect 10395 9472 10396 9512
rect 10436 9472 10437 9512
rect 10395 9463 10437 9472
rect 10539 9512 10581 9521
rect 10539 9472 10540 9512
rect 10580 9472 10581 9512
rect 10539 9463 10581 9472
rect 10923 9512 10965 9521
rect 10923 9472 10924 9512
rect 10964 9472 10965 9512
rect 10923 9463 10965 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11691 9512 11733 9521
rect 11691 9472 11692 9512
rect 11732 9472 11733 9512
rect 11691 9463 11733 9472
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 12459 9512 12501 9521
rect 12459 9472 12460 9512
rect 12500 9472 12501 9512
rect 12459 9463 12501 9472
rect 12843 9512 12885 9521
rect 12843 9472 12844 9512
rect 12884 9472 12885 9512
rect 12843 9463 12885 9472
rect 13227 9512 13269 9521
rect 13227 9472 13228 9512
rect 13268 9472 13269 9512
rect 13227 9463 13269 9472
rect 13467 9512 13509 9521
rect 13467 9472 13468 9512
rect 13508 9472 13509 9512
rect 13467 9463 13509 9472
rect 13611 9512 13653 9521
rect 13611 9472 13612 9512
rect 13652 9472 13653 9512
rect 13611 9463 13653 9472
rect 13995 9512 14037 9521
rect 13995 9472 13996 9512
rect 14036 9472 14037 9512
rect 13995 9463 14037 9472
rect 14379 9512 14421 9521
rect 14379 9472 14380 9512
rect 14420 9472 14421 9512
rect 14379 9463 14421 9472
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 14763 9463 14805 9472
rect 15003 9512 15045 9521
rect 15003 9472 15004 9512
rect 15044 9472 15045 9512
rect 15003 9463 15045 9472
rect 15147 9512 15189 9521
rect 15147 9472 15148 9512
rect 15188 9472 15189 9512
rect 15147 9463 15189 9472
rect 15531 9512 15573 9521
rect 15531 9472 15532 9512
rect 15572 9472 15573 9512
rect 15531 9463 15573 9472
rect 15915 9512 15957 9521
rect 15915 9472 15916 9512
rect 15956 9472 15957 9512
rect 15915 9463 15957 9472
rect 16299 9512 16341 9521
rect 16299 9472 16300 9512
rect 16340 9472 16341 9512
rect 16299 9463 16341 9472
rect 16683 9512 16725 9521
rect 16683 9472 16684 9512
rect 16724 9472 16725 9512
rect 16683 9463 16725 9472
rect 16923 9512 16965 9521
rect 16923 9472 16924 9512
rect 16964 9472 16965 9512
rect 16923 9463 16965 9472
rect 17067 9512 17109 9521
rect 17067 9472 17068 9512
rect 17108 9472 17109 9512
rect 17067 9463 17109 9472
rect 17451 9512 17493 9521
rect 17451 9472 17452 9512
rect 17492 9472 17493 9512
rect 17451 9463 17493 9472
rect 17835 9512 17877 9521
rect 17835 9472 17836 9512
rect 17876 9472 17877 9512
rect 17835 9463 17877 9472
rect 18219 9512 18261 9521
rect 18219 9472 18220 9512
rect 18260 9472 18261 9512
rect 18219 9463 18261 9472
rect 18603 9512 18645 9521
rect 18603 9472 18604 9512
rect 18644 9472 18645 9512
rect 18603 9463 18645 9472
rect 18987 9512 19029 9521
rect 18987 9472 18988 9512
rect 19028 9472 19029 9512
rect 18987 9463 19029 9472
rect 19371 9512 19413 9521
rect 19371 9472 19372 9512
rect 19412 9472 19413 9512
rect 19371 9463 19413 9472
rect 19755 9512 19797 9521
rect 19755 9472 19756 9512
rect 19796 9472 19797 9512
rect 19755 9463 19797 9472
rect 20523 9512 20565 9521
rect 20523 9472 20524 9512
rect 20564 9472 20565 9512
rect 20523 9463 20565 9472
rect 20763 9512 20805 9521
rect 20763 9472 20764 9512
rect 20804 9472 20805 9512
rect 20763 9463 20805 9472
rect 21099 9512 21141 9521
rect 21099 9472 21100 9512
rect 21140 9472 21141 9512
rect 21099 9463 21141 9472
rect 21291 9512 21333 9521
rect 21291 9472 21292 9512
rect 21332 9472 21333 9512
rect 21291 9463 21333 9472
rect 21867 9512 21909 9521
rect 21867 9472 21868 9512
rect 21908 9472 21909 9512
rect 21867 9463 21909 9472
rect 22251 9512 22293 9521
rect 22251 9472 22252 9512
rect 22292 9472 22293 9512
rect 22251 9463 22293 9472
rect 22443 9512 22485 9521
rect 22443 9472 22444 9512
rect 22484 9472 22485 9512
rect 22443 9463 22485 9472
rect 23019 9512 23061 9521
rect 23019 9472 23020 9512
rect 23060 9472 23061 9512
rect 23019 9463 23061 9472
rect 23403 9512 23445 9521
rect 23403 9472 23404 9512
rect 23444 9472 23445 9512
rect 23403 9463 23445 9472
rect 23787 9512 23829 9521
rect 23787 9472 23788 9512
rect 23828 9472 23829 9512
rect 23787 9463 23829 9472
rect 23979 9512 24021 9521
rect 23979 9472 23980 9512
rect 24020 9472 24021 9512
rect 23979 9463 24021 9472
rect 24363 9512 24405 9521
rect 24363 9472 24364 9512
rect 24404 9472 24405 9512
rect 24363 9463 24405 9472
rect 24939 9512 24981 9521
rect 24939 9472 24940 9512
rect 24980 9472 24981 9512
rect 24939 9463 24981 9472
rect 25323 9512 25365 9521
rect 25323 9472 25324 9512
rect 25364 9472 25365 9512
rect 25323 9463 25365 9472
rect 25515 9512 25557 9521
rect 25515 9472 25516 9512
rect 25556 9472 25557 9512
rect 25515 9463 25557 9472
rect 25851 9512 25893 9521
rect 25851 9472 25852 9512
rect 25892 9472 25893 9512
rect 25851 9463 25893 9472
rect 26091 9512 26133 9521
rect 26091 9472 26092 9512
rect 26132 9472 26133 9512
rect 26091 9463 26133 9472
rect 26475 9512 26517 9521
rect 26475 9472 26476 9512
rect 26516 9472 26517 9512
rect 26475 9463 26517 9472
rect 26859 9512 26901 9521
rect 26859 9472 26860 9512
rect 26900 9472 26901 9512
rect 26859 9463 26901 9472
rect 27243 9512 27285 9521
rect 27243 9472 27244 9512
rect 27284 9472 27285 9512
rect 27243 9463 27285 9472
rect 28395 9512 28437 9521
rect 28395 9472 28396 9512
rect 28436 9472 28437 9512
rect 28395 9463 28437 9472
rect 28539 9512 28581 9521
rect 28539 9472 28540 9512
rect 28580 9472 28581 9512
rect 28539 9463 28581 9472
rect 28779 9512 28821 9521
rect 28779 9472 28780 9512
rect 28820 9472 28821 9512
rect 28779 9463 28821 9472
rect 29163 9512 29205 9521
rect 29163 9472 29164 9512
rect 29204 9472 29205 9512
rect 29163 9463 29205 9472
rect 29355 9512 29397 9521
rect 29355 9472 29356 9512
rect 29396 9472 29397 9512
rect 29355 9463 29397 9472
rect 29691 9512 29733 9521
rect 29691 9472 29692 9512
rect 29732 9472 29733 9512
rect 29691 9463 29733 9472
rect 29931 9512 29973 9521
rect 29931 9472 29932 9512
rect 29972 9472 29973 9512
rect 29931 9463 29973 9472
rect 30315 9512 30357 9521
rect 30315 9472 30316 9512
rect 30356 9472 30357 9512
rect 30315 9463 30357 9472
rect 30699 9512 30741 9521
rect 30699 9472 30700 9512
rect 30740 9472 30741 9512
rect 30699 9463 30741 9472
rect 31467 9512 31509 9521
rect 31467 9472 31468 9512
rect 31508 9472 31509 9512
rect 31467 9463 31509 9472
rect 31851 9512 31893 9521
rect 31851 9472 31852 9512
rect 31892 9472 31893 9512
rect 31851 9463 31893 9472
rect 32235 9512 32277 9521
rect 32235 9472 32236 9512
rect 32276 9472 32277 9512
rect 32235 9463 32277 9472
rect 32619 9512 32661 9521
rect 32619 9472 32620 9512
rect 32660 9472 32661 9512
rect 32619 9463 32661 9472
rect 33003 9512 33045 9521
rect 33003 9472 33004 9512
rect 33044 9472 33045 9512
rect 33003 9463 33045 9472
rect 33387 9512 33429 9521
rect 33387 9472 33388 9512
rect 33428 9472 33429 9512
rect 33387 9463 33429 9472
rect 33771 9512 33813 9521
rect 33771 9472 33772 9512
rect 33812 9472 33813 9512
rect 33771 9463 33813 9472
rect 34155 9512 34197 9521
rect 34155 9472 34156 9512
rect 34196 9472 34197 9512
rect 34155 9463 34197 9472
rect 34474 9512 34532 9513
rect 34474 9472 34483 9512
rect 34523 9472 34532 9512
rect 34474 9471 34532 9472
rect 34683 9512 34725 9521
rect 34683 9472 34684 9512
rect 34724 9472 34725 9512
rect 34683 9463 34725 9472
rect 34971 9512 35013 9521
rect 34971 9472 34972 9512
rect 35012 9472 35013 9512
rect 34971 9463 35013 9472
rect 35307 9512 35349 9521
rect 35307 9472 35308 9512
rect 35348 9472 35349 9512
rect 35307 9463 35349 9472
rect 35691 9512 35733 9521
rect 35691 9472 35692 9512
rect 35732 9472 35733 9512
rect 35691 9463 35733 9472
rect 36075 9512 36117 9521
rect 36075 9472 36076 9512
rect 36116 9472 36117 9512
rect 36075 9463 36117 9472
rect 36459 9512 36501 9521
rect 36459 9472 36460 9512
rect 36500 9472 36501 9512
rect 36459 9463 36501 9472
rect 41835 9512 41877 9521
rect 41835 9472 41836 9512
rect 41876 9472 41877 9512
rect 41835 9463 41877 9472
rect 42219 9512 42261 9521
rect 42219 9472 42220 9512
rect 42260 9472 42261 9512
rect 42219 9463 42261 9472
rect 42603 9512 42645 9521
rect 42603 9472 42604 9512
rect 42644 9472 42645 9512
rect 42603 9463 42645 9472
rect 42987 9512 43029 9521
rect 42987 9472 42988 9512
rect 43028 9472 43029 9512
rect 42987 9463 43029 9472
rect 43371 9512 43413 9521
rect 43371 9472 43372 9512
rect 43412 9472 43413 9512
rect 43371 9463 43413 9472
rect 43755 9512 43797 9521
rect 43755 9472 43756 9512
rect 43796 9472 43797 9512
rect 43755 9463 43797 9472
rect 44139 9512 44181 9521
rect 44139 9472 44140 9512
rect 44180 9472 44181 9512
rect 44139 9463 44181 9472
rect 44907 9512 44949 9521
rect 44907 9472 44908 9512
rect 44948 9472 44949 9512
rect 44907 9463 44949 9472
rect 44619 9428 44661 9437
rect 44619 9388 44620 9428
rect 44660 9388 44661 9428
rect 44619 9379 44661 9388
rect 2235 9344 2277 9353
rect 2235 9304 2236 9344
rect 2276 9304 2277 9344
rect 2235 9295 2277 9304
rect 3387 9344 3429 9353
rect 3387 9304 3388 9344
rect 3428 9304 3429 9344
rect 3387 9295 3429 9304
rect 11547 9344 11589 9353
rect 11547 9304 11548 9344
rect 11588 9304 11589 9344
rect 11547 9295 11589 9304
rect 11931 9344 11973 9353
rect 11931 9304 11932 9344
rect 11972 9304 11973 9344
rect 11931 9295 11973 9304
rect 14235 9344 14277 9353
rect 14235 9304 14236 9344
rect 14276 9304 14277 9344
rect 14235 9295 14277 9304
rect 14619 9344 14661 9353
rect 14619 9304 14620 9344
rect 14660 9304 14661 9344
rect 14619 9295 14661 9304
rect 16539 9344 16581 9353
rect 16539 9304 16540 9344
rect 16580 9304 16581 9344
rect 16539 9295 16581 9304
rect 19995 9344 20037 9353
rect 19995 9304 19996 9344
rect 20036 9304 20037 9344
rect 19995 9295 20037 9304
rect 20859 9344 20901 9353
rect 20859 9304 20860 9344
rect 20900 9304 20901 9344
rect 20859 9295 20901 9304
rect 22011 9344 22053 9353
rect 22011 9304 22012 9344
rect 22052 9304 22053 9344
rect 22011 9295 22053 9304
rect 23547 9344 23589 9353
rect 23547 9304 23548 9344
rect 23588 9304 23589 9344
rect 23547 9295 23589 9304
rect 24219 9344 24261 9353
rect 24219 9304 24220 9344
rect 24260 9304 24261 9344
rect 24219 9295 24261 9304
rect 24603 9344 24645 9353
rect 24603 9304 24604 9344
rect 24644 9304 24645 9344
rect 24603 9295 24645 9304
rect 25083 9344 25125 9353
rect 25083 9304 25084 9344
rect 25124 9304 25125 9344
rect 25083 9295 25125 9304
rect 25755 9344 25797 9353
rect 25755 9304 25756 9344
rect 25796 9304 25797 9344
rect 25755 9295 25797 9304
rect 29595 9344 29637 9353
rect 29595 9304 29596 9344
rect 29636 9304 29637 9344
rect 29595 9295 29637 9304
rect 33147 9344 33189 9353
rect 33147 9304 33148 9344
rect 33188 9304 33189 9344
rect 33147 9295 33189 9304
rect 35067 9344 35109 9353
rect 35067 9304 35068 9344
rect 35108 9304 35109 9344
rect 35067 9295 35109 9304
rect 42459 9344 42501 9353
rect 42459 9304 42460 9344
rect 42500 9304 42501 9344
rect 42459 9295 42501 9304
rect 44379 9344 44421 9353
rect 44379 9304 44380 9344
rect 44420 9304 44421 9344
rect 44379 9295 44421 9304
rect 1467 9260 1509 9269
rect 1467 9220 1468 9260
rect 1508 9220 1509 9260
rect 1467 9211 1509 9220
rect 2619 9260 2661 9269
rect 2619 9220 2620 9260
rect 2660 9220 2661 9260
rect 2619 9211 2661 9220
rect 10779 9260 10821 9269
rect 10779 9220 10780 9260
rect 10820 9220 10821 9260
rect 10779 9211 10821 9220
rect 12315 9260 12357 9269
rect 12315 9220 12316 9260
rect 12356 9220 12357 9260
rect 12315 9211 12357 9220
rect 15387 9260 15429 9269
rect 15387 9220 15388 9260
rect 15428 9220 15429 9260
rect 15387 9211 15429 9220
rect 15771 9260 15813 9269
rect 15771 9220 15772 9260
rect 15812 9220 15813 9260
rect 15771 9211 15813 9220
rect 20331 9260 20373 9269
rect 20331 9220 20332 9260
rect 20372 9220 20373 9260
rect 20331 9211 20373 9220
rect 21627 9260 21669 9269
rect 21627 9220 21628 9260
rect 21668 9220 21669 9260
rect 21627 9211 21669 9220
rect 22779 9260 22821 9269
rect 22779 9220 22780 9260
rect 22820 9220 22821 9260
rect 22779 9211 22821 9220
rect 23163 9260 23205 9269
rect 23163 9220 23164 9260
rect 23204 9220 23205 9260
rect 23163 9211 23205 9220
rect 24699 9260 24741 9269
rect 24699 9220 24700 9260
rect 24740 9220 24741 9260
rect 24699 9211 24741 9220
rect 26235 9260 26277 9269
rect 26235 9220 26236 9260
rect 26276 9220 26277 9260
rect 26235 9211 26277 9220
rect 27003 9260 27045 9269
rect 27003 9220 27004 9260
rect 27044 9220 27045 9260
rect 27003 9211 27045 9220
rect 28155 9260 28197 9269
rect 28155 9220 28156 9260
rect 28196 9220 28197 9260
rect 28155 9211 28197 9220
rect 30459 9260 30501 9269
rect 30459 9220 30460 9260
rect 30500 9220 30501 9260
rect 30459 9211 30501 9220
rect 33915 9260 33957 9269
rect 33915 9220 33916 9260
rect 33956 9220 33957 9260
rect 33915 9211 33957 9220
rect 34299 9260 34341 9269
rect 34299 9220 34300 9260
rect 34340 9220 34341 9260
rect 34299 9211 34341 9220
rect 40474 9260 40532 9261
rect 40474 9220 40483 9260
rect 40523 9220 40532 9260
rect 40474 9219 40532 9220
rect 40666 9260 40724 9261
rect 40666 9220 40675 9260
rect 40715 9220 40724 9260
rect 40666 9219 40724 9220
rect 40954 9260 41012 9261
rect 40954 9220 40963 9260
rect 41003 9220 41012 9260
rect 40954 9219 41012 9220
rect 41242 9260 41300 9261
rect 41242 9220 41251 9260
rect 41291 9220 41300 9260
rect 41242 9219 41300 9220
rect 41530 9260 41588 9261
rect 41530 9220 41539 9260
rect 41579 9220 41588 9260
rect 41530 9219 41588 9220
rect 42075 9260 42117 9269
rect 42075 9220 42076 9260
rect 42116 9220 42117 9260
rect 42075 9211 42117 9220
rect 45147 9260 45189 9269
rect 45147 9220 45148 9260
rect 45188 9220 45189 9260
rect 45147 9211 45189 9220
rect 1152 9092 45216 9116
rect 1152 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 45216 9092
rect 1152 9028 45216 9052
rect 1467 8924 1509 8933
rect 1467 8884 1468 8924
rect 1508 8884 1509 8924
rect 1467 8875 1509 8884
rect 3195 8924 3237 8933
rect 3195 8884 3196 8924
rect 3236 8884 3237 8924
rect 3195 8875 3237 8884
rect 10299 8924 10341 8933
rect 10299 8884 10300 8924
rect 10340 8884 10341 8924
rect 10299 8875 10341 8884
rect 11067 8924 11109 8933
rect 11067 8884 11068 8924
rect 11108 8884 11109 8924
rect 11067 8875 11109 8884
rect 12603 8924 12645 8933
rect 12603 8884 12604 8924
rect 12644 8884 12645 8924
rect 12603 8875 12645 8884
rect 14139 8924 14181 8933
rect 14139 8884 14140 8924
rect 14180 8884 14181 8924
rect 14139 8875 14181 8884
rect 15147 8924 15189 8933
rect 15147 8884 15148 8924
rect 15188 8884 15189 8924
rect 15147 8875 15189 8884
rect 15867 8924 15909 8933
rect 15867 8884 15868 8924
rect 15908 8884 15909 8924
rect 15867 8875 15909 8884
rect 16251 8924 16293 8933
rect 16251 8884 16252 8924
rect 16292 8884 16293 8924
rect 16251 8875 16293 8884
rect 18459 8924 18501 8933
rect 18459 8884 18460 8924
rect 18500 8884 18501 8924
rect 18459 8875 18501 8884
rect 18843 8924 18885 8933
rect 18843 8884 18844 8924
rect 18884 8884 18885 8924
rect 18843 8875 18885 8884
rect 19227 8924 19269 8933
rect 19227 8884 19228 8924
rect 19268 8884 19269 8924
rect 19227 8875 19269 8884
rect 19611 8924 19653 8933
rect 19611 8884 19612 8924
rect 19652 8884 19653 8924
rect 19611 8875 19653 8884
rect 19995 8924 20037 8933
rect 19995 8884 19996 8924
rect 20036 8884 20037 8924
rect 19995 8875 20037 8884
rect 20379 8924 20421 8933
rect 20379 8884 20380 8924
rect 20420 8884 20421 8924
rect 20379 8875 20421 8884
rect 20763 8924 20805 8933
rect 20763 8884 20764 8924
rect 20804 8884 20805 8924
rect 20763 8875 20805 8884
rect 21435 8924 21477 8933
rect 21435 8884 21436 8924
rect 21476 8884 21477 8924
rect 21435 8875 21477 8884
rect 29595 8924 29637 8933
rect 29595 8884 29596 8924
rect 29636 8884 29637 8924
rect 29595 8875 29637 8884
rect 32187 8924 32229 8933
rect 32187 8884 32188 8924
rect 32228 8884 32229 8924
rect 32187 8875 32229 8884
rect 32571 8924 32613 8933
rect 32571 8884 32572 8924
rect 32612 8884 32613 8924
rect 32571 8875 32613 8884
rect 32955 8924 32997 8933
rect 32955 8884 32956 8924
rect 32996 8884 32997 8924
rect 32955 8875 32997 8884
rect 33339 8924 33381 8933
rect 33339 8884 33340 8924
rect 33380 8884 33381 8924
rect 33339 8875 33381 8884
rect 33723 8924 33765 8933
rect 33723 8884 33724 8924
rect 33764 8884 33765 8924
rect 33723 8875 33765 8884
rect 34107 8924 34149 8933
rect 34107 8884 34108 8924
rect 34148 8884 34149 8924
rect 34107 8875 34149 8884
rect 35739 8924 35781 8933
rect 35739 8884 35740 8924
rect 35780 8884 35781 8924
rect 35739 8875 35781 8884
rect 43035 8924 43077 8933
rect 43035 8884 43036 8924
rect 43076 8884 43077 8924
rect 43035 8875 43077 8884
rect 43419 8924 43461 8933
rect 43419 8884 43420 8924
rect 43460 8884 43461 8924
rect 43419 8875 43461 8884
rect 1851 8840 1893 8849
rect 1851 8800 1852 8840
rect 1892 8800 1893 8840
rect 1851 8791 1893 8800
rect 3579 8840 3621 8849
rect 3579 8800 3580 8840
rect 3620 8800 3621 8840
rect 3579 8791 3621 8800
rect 11451 8840 11493 8849
rect 11451 8800 11452 8840
rect 11492 8800 11493 8840
rect 11451 8791 11493 8800
rect 12219 8840 12261 8849
rect 12219 8800 12220 8840
rect 12260 8800 12261 8840
rect 12219 8791 12261 8800
rect 12987 8840 13029 8849
rect 12987 8800 12988 8840
rect 13028 8800 13029 8840
rect 12987 8791 13029 8800
rect 17979 8840 18021 8849
rect 17979 8800 17980 8840
rect 18020 8800 18021 8840
rect 17979 8791 18021 8800
rect 23163 8840 23205 8849
rect 23163 8800 23164 8840
rect 23204 8800 23205 8840
rect 23163 8791 23205 8800
rect 25275 8840 25317 8849
rect 25275 8800 25276 8840
rect 25316 8800 25317 8840
rect 25275 8791 25317 8800
rect 25947 8840 25989 8849
rect 25947 8800 25948 8840
rect 25988 8800 25989 8840
rect 25947 8791 25989 8800
rect 34491 8840 34533 8849
rect 34491 8800 34492 8840
rect 34532 8800 34533 8840
rect 34491 8791 34533 8800
rect 35355 8840 35397 8849
rect 35355 8800 35356 8840
rect 35396 8800 35397 8840
rect 35355 8791 35397 8800
rect 38091 8840 38133 8849
rect 38091 8800 38092 8840
rect 38132 8800 38133 8840
rect 38091 8791 38133 8800
rect 38523 8840 38565 8849
rect 38523 8800 38524 8840
rect 38564 8800 38565 8840
rect 38523 8791 38565 8800
rect 44379 8840 44421 8849
rect 44379 8800 44380 8840
rect 44420 8800 44421 8840
rect 44379 8791 44421 8800
rect 15051 8756 15093 8765
rect 15051 8716 15052 8756
rect 15092 8716 15093 8756
rect 15051 8707 15093 8716
rect 15226 8756 15284 8757
rect 15226 8716 15235 8756
rect 15275 8716 15284 8756
rect 15226 8715 15284 8716
rect 17643 8756 17685 8765
rect 17643 8716 17644 8756
rect 17684 8716 17685 8756
rect 17643 8707 17685 8716
rect 17835 8756 17877 8765
rect 17835 8716 17836 8756
rect 17876 8716 17877 8756
rect 17835 8707 17877 8716
rect 41259 8756 41301 8765
rect 41259 8716 41260 8756
rect 41300 8716 41301 8756
rect 41259 8707 41301 8716
rect 41643 8756 41685 8765
rect 41643 8716 41644 8756
rect 41684 8716 41685 8756
rect 41643 8707 41685 8716
rect 41931 8756 41973 8765
rect 41931 8716 41932 8756
rect 41972 8716 41973 8756
rect 41931 8707 41973 8716
rect 42219 8756 42261 8765
rect 42219 8716 42220 8756
rect 42260 8716 42261 8756
rect 42219 8707 42261 8716
rect 42507 8756 42549 8765
rect 42507 8716 42508 8756
rect 42548 8716 42549 8756
rect 42507 8707 42549 8716
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 1611 8672 1653 8681
rect 1611 8632 1612 8672
rect 1652 8632 1653 8672
rect 1611 8623 1653 8632
rect 1995 8672 2037 8681
rect 1995 8632 1996 8672
rect 2036 8632 2037 8672
rect 1995 8623 2037 8632
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 2619 8672 2661 8681
rect 2619 8632 2620 8672
rect 2660 8632 2661 8672
rect 2619 8623 2661 8632
rect 2955 8672 2997 8681
rect 2955 8632 2956 8672
rect 2996 8632 2997 8672
rect 2955 8623 2997 8632
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 10059 8672 10101 8681
rect 10059 8632 10060 8672
rect 10100 8632 10101 8672
rect 10059 8623 10101 8632
rect 10443 8672 10485 8681
rect 10443 8632 10444 8672
rect 10484 8632 10485 8672
rect 10443 8623 10485 8632
rect 10827 8672 10869 8681
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 11211 8672 11253 8681
rect 11211 8632 11212 8672
rect 11252 8632 11253 8672
rect 11211 8623 11253 8632
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 11979 8672 12021 8681
rect 11979 8632 11980 8672
rect 12020 8632 12021 8672
rect 11979 8623 12021 8632
rect 12363 8672 12405 8681
rect 12363 8632 12364 8672
rect 12404 8632 12405 8672
rect 12363 8623 12405 8632
rect 12747 8672 12789 8681
rect 12747 8632 12748 8672
rect 12788 8632 12789 8672
rect 12747 8623 12789 8632
rect 13131 8672 13173 8681
rect 13131 8632 13132 8672
rect 13172 8632 13173 8672
rect 13131 8623 13173 8632
rect 13515 8672 13557 8681
rect 13515 8632 13516 8672
rect 13556 8632 13557 8672
rect 13515 8623 13557 8632
rect 13755 8672 13797 8681
rect 13755 8632 13756 8672
rect 13796 8632 13797 8672
rect 13755 8623 13797 8632
rect 13899 8672 13941 8681
rect 13899 8632 13900 8672
rect 13940 8632 13941 8672
rect 13899 8623 13941 8632
rect 14283 8672 14325 8681
rect 14283 8632 14284 8672
rect 14324 8632 14325 8672
rect 14283 8623 14325 8632
rect 14523 8672 14565 8681
rect 14523 8632 14524 8672
rect 14564 8632 14565 8672
rect 14523 8623 14565 8632
rect 14667 8672 14709 8681
rect 14667 8632 14668 8672
rect 14708 8632 14709 8672
rect 14667 8623 14709 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 16011 8672 16053 8681
rect 16011 8632 16012 8672
rect 16052 8632 16053 8672
rect 16011 8623 16053 8632
rect 16395 8672 16437 8681
rect 16395 8632 16396 8672
rect 16436 8632 16437 8672
rect 16395 8623 16437 8632
rect 16635 8672 16677 8681
rect 16635 8632 16636 8672
rect 16676 8632 16677 8672
rect 16635 8623 16677 8632
rect 17259 8672 17301 8681
rect 17259 8632 17260 8672
rect 17300 8632 17301 8672
rect 17259 8623 17301 8632
rect 18219 8672 18261 8681
rect 18219 8632 18220 8672
rect 18260 8632 18261 8672
rect 18219 8623 18261 8632
rect 18699 8672 18741 8681
rect 18699 8632 18700 8672
rect 18740 8632 18741 8672
rect 18699 8623 18741 8632
rect 19083 8672 19125 8681
rect 19083 8632 19084 8672
rect 19124 8632 19125 8672
rect 19083 8623 19125 8632
rect 19467 8672 19509 8681
rect 19467 8632 19468 8672
rect 19508 8632 19509 8672
rect 19467 8623 19509 8632
rect 19851 8672 19893 8681
rect 19851 8632 19852 8672
rect 19892 8632 19893 8672
rect 19851 8623 19893 8632
rect 20235 8672 20277 8681
rect 20235 8632 20236 8672
rect 20276 8632 20277 8672
rect 20235 8623 20277 8632
rect 20619 8672 20661 8681
rect 20619 8632 20620 8672
rect 20660 8632 20661 8672
rect 20619 8623 20661 8632
rect 21003 8672 21045 8681
rect 21003 8632 21004 8672
rect 21044 8632 21045 8672
rect 21003 8623 21045 8632
rect 21195 8672 21237 8681
rect 21195 8632 21196 8672
rect 21236 8632 21237 8672
rect 21195 8623 21237 8632
rect 21867 8672 21909 8681
rect 21867 8632 21868 8672
rect 21908 8632 21909 8672
rect 21867 8623 21909 8632
rect 22059 8672 22101 8681
rect 22059 8632 22060 8672
rect 22100 8632 22101 8672
rect 22059 8623 22101 8632
rect 22299 8672 22341 8681
rect 22299 8632 22300 8672
rect 22340 8632 22341 8672
rect 22299 8623 22341 8632
rect 22779 8672 22821 8681
rect 22779 8632 22780 8672
rect 22820 8632 22821 8672
rect 22779 8623 22821 8632
rect 23019 8672 23061 8681
rect 23019 8632 23020 8672
rect 23060 8632 23061 8672
rect 23019 8623 23061 8632
rect 23403 8672 23445 8681
rect 23403 8632 23404 8672
rect 23444 8632 23445 8672
rect 23403 8623 23445 8632
rect 23547 8672 23589 8681
rect 23547 8632 23548 8672
rect 23588 8632 23589 8672
rect 23547 8623 23589 8632
rect 23787 8672 23829 8681
rect 23787 8632 23788 8672
rect 23828 8632 23829 8672
rect 23787 8623 23829 8632
rect 25515 8672 25557 8681
rect 25515 8632 25516 8672
rect 25556 8632 25557 8672
rect 25515 8623 25557 8632
rect 25707 8672 25749 8681
rect 25707 8632 25708 8672
rect 25748 8632 25749 8672
rect 25707 8623 25749 8632
rect 26283 8672 26325 8681
rect 26283 8632 26284 8672
rect 26324 8632 26325 8672
rect 26283 8623 26325 8632
rect 26475 8672 26517 8681
rect 26475 8632 26476 8672
rect 26516 8632 26517 8672
rect 26475 8623 26517 8632
rect 26715 8672 26757 8681
rect 26715 8632 26716 8672
rect 26756 8632 26757 8672
rect 26715 8623 26757 8632
rect 29355 8672 29397 8681
rect 29355 8632 29356 8672
rect 29396 8632 29397 8672
rect 29355 8623 29397 8632
rect 29835 8672 29877 8681
rect 29835 8632 29836 8672
rect 29876 8632 29877 8672
rect 29835 8623 29877 8632
rect 32427 8672 32469 8681
rect 32427 8632 32428 8672
rect 32468 8632 32469 8672
rect 32427 8623 32469 8632
rect 32811 8672 32853 8681
rect 32811 8632 32812 8672
rect 32852 8632 32853 8672
rect 32811 8623 32853 8632
rect 33195 8672 33237 8681
rect 33195 8632 33196 8672
rect 33236 8632 33237 8672
rect 33195 8623 33237 8632
rect 33579 8672 33621 8681
rect 33579 8632 33580 8672
rect 33620 8632 33621 8672
rect 33579 8623 33621 8632
rect 33963 8672 34005 8681
rect 33963 8632 33964 8672
rect 34004 8632 34005 8672
rect 33963 8623 34005 8632
rect 34347 8672 34389 8681
rect 34347 8632 34348 8672
rect 34388 8632 34389 8672
rect 34347 8623 34389 8632
rect 34731 8672 34773 8681
rect 34731 8632 34732 8672
rect 34772 8632 34773 8672
rect 34731 8623 34773 8632
rect 35115 8672 35157 8681
rect 35115 8632 35116 8672
rect 35156 8632 35157 8672
rect 35115 8623 35157 8632
rect 35530 8672 35588 8673
rect 35530 8632 35539 8672
rect 35579 8632 35588 8672
rect 35530 8631 35588 8632
rect 38091 8672 38133 8681
rect 38091 8632 38092 8672
rect 38132 8632 38133 8672
rect 38091 8623 38133 8632
rect 38283 8672 38325 8681
rect 38283 8632 38284 8672
rect 38324 8632 38325 8672
rect 38283 8623 38325 8632
rect 38763 8672 38805 8681
rect 38763 8632 38764 8672
rect 38804 8632 38805 8672
rect 38763 8623 38805 8632
rect 39051 8672 39093 8681
rect 39051 8632 39052 8672
rect 39092 8632 39093 8672
rect 39051 8623 39093 8632
rect 39339 8672 39381 8681
rect 39339 8632 39340 8672
rect 39380 8632 39381 8672
rect 39339 8623 39381 8632
rect 39627 8672 39669 8681
rect 39627 8632 39628 8672
rect 39668 8632 39669 8672
rect 39627 8623 39669 8632
rect 39915 8672 39957 8681
rect 39915 8632 39916 8672
rect 39956 8632 39957 8672
rect 39915 8623 39957 8632
rect 40203 8672 40245 8681
rect 40203 8632 40204 8672
rect 40244 8632 40245 8672
rect 40203 8623 40245 8632
rect 40491 8672 40533 8681
rect 40491 8632 40492 8672
rect 40532 8632 40533 8672
rect 40491 8623 40533 8632
rect 40779 8672 40821 8681
rect 40779 8632 40780 8672
rect 40820 8632 40821 8672
rect 40779 8623 40821 8632
rect 40971 8672 41013 8681
rect 40971 8632 40972 8672
rect 41012 8632 41013 8672
rect 40971 8623 41013 8632
rect 42651 8672 42693 8681
rect 42651 8632 42652 8672
rect 42692 8632 42693 8672
rect 42651 8623 42693 8632
rect 42891 8672 42933 8681
rect 42891 8632 42892 8672
rect 42932 8632 42933 8672
rect 42891 8623 42933 8632
rect 43275 8672 43317 8681
rect 43275 8632 43276 8672
rect 43316 8632 43317 8672
rect 43275 8623 43317 8632
rect 43659 8672 43701 8681
rect 43659 8632 43660 8672
rect 43700 8632 43701 8672
rect 43659 8623 43701 8632
rect 43947 8672 43989 8681
rect 43947 8632 43948 8672
rect 43988 8632 43989 8672
rect 43947 8623 43989 8632
rect 44139 8672 44181 8681
rect 44139 8632 44140 8672
rect 44180 8632 44181 8672
rect 44139 8623 44181 8632
rect 44523 8672 44565 8681
rect 44523 8632 44524 8672
rect 44564 8632 44565 8672
rect 44523 8623 44565 8632
rect 44907 8672 44949 8681
rect 44907 8632 44908 8672
rect 44948 8632 44949 8672
rect 44907 8623 44949 8632
rect 2235 8588 2277 8597
rect 2235 8548 2236 8588
rect 2276 8548 2277 8588
rect 2235 8539 2277 8548
rect 10683 8588 10725 8597
rect 10683 8548 10684 8588
rect 10724 8548 10725 8588
rect 10683 8539 10725 8548
rect 13371 8588 13413 8597
rect 13371 8548 13372 8588
rect 13412 8548 13413 8588
rect 13371 8539 13413 8548
rect 14907 8588 14949 8597
rect 14907 8548 14908 8588
rect 14948 8548 14949 8588
rect 14907 8539 14949 8548
rect 17019 8588 17061 8597
rect 17019 8548 17020 8588
rect 17060 8548 17061 8588
rect 17019 8539 17061 8548
rect 21627 8588 21669 8597
rect 21627 8548 21628 8588
rect 21668 8548 21669 8588
rect 21627 8539 21669 8548
rect 44763 8588 44805 8597
rect 44763 8548 44764 8588
rect 44804 8548 44805 8588
rect 44763 8539 44805 8548
rect 11835 8504 11877 8513
rect 11835 8464 11836 8504
rect 11876 8464 11877 8504
rect 11835 8455 11877 8464
rect 17643 8504 17685 8513
rect 17643 8464 17644 8504
rect 17684 8464 17685 8504
rect 17643 8455 17685 8464
rect 26043 8504 26085 8513
rect 26043 8464 26044 8504
rect 26084 8464 26085 8504
rect 26043 8455 26085 8464
rect 29115 8504 29157 8513
rect 29115 8464 29116 8504
rect 29156 8464 29157 8504
rect 29115 8455 29157 8464
rect 45147 8504 45189 8513
rect 45147 8464 45148 8504
rect 45188 8464 45189 8504
rect 45147 8455 45189 8464
rect 1152 8336 45216 8360
rect 1152 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 45216 8336
rect 1152 8272 45216 8296
rect 11163 8168 11205 8177
rect 11163 8128 11164 8168
rect 11204 8128 11205 8168
rect 11163 8119 11205 8128
rect 14235 8168 14277 8177
rect 14235 8128 14236 8168
rect 14276 8128 14277 8168
rect 14235 8119 14277 8128
rect 18603 8168 18645 8177
rect 18603 8128 18604 8168
rect 18644 8128 18645 8168
rect 18603 8119 18645 8128
rect 28539 8168 28581 8177
rect 28539 8128 28540 8168
rect 28580 8128 28581 8168
rect 28539 8119 28581 8128
rect 28923 8168 28965 8177
rect 28923 8128 28924 8168
rect 28964 8128 28965 8168
rect 28923 8119 28965 8128
rect 31227 8168 31269 8177
rect 31227 8128 31228 8168
rect 31268 8128 31269 8168
rect 31227 8119 31269 8128
rect 31995 8168 32037 8177
rect 31995 8128 31996 8168
rect 32036 8128 32037 8168
rect 31995 8119 32037 8128
rect 34875 8168 34917 8177
rect 34875 8128 34876 8168
rect 34916 8128 34917 8168
rect 34875 8119 34917 8128
rect 35355 8168 35397 8177
rect 35355 8128 35356 8168
rect 35396 8128 35397 8168
rect 35355 8119 35397 8128
rect 43227 8168 43269 8177
rect 43227 8128 43228 8168
rect 43268 8128 43269 8168
rect 43227 8119 43269 8128
rect 15339 8084 15381 8093
rect 15339 8044 15340 8084
rect 15380 8044 15381 8084
rect 15339 8035 15381 8044
rect 19899 8084 19941 8093
rect 19899 8044 19900 8084
rect 19940 8044 19941 8084
rect 19899 8035 19941 8044
rect 29835 8084 29877 8093
rect 29835 8044 29836 8084
rect 29876 8044 29877 8084
rect 29835 8035 29877 8044
rect 31611 8084 31653 8093
rect 31611 8044 31612 8084
rect 31652 8044 31653 8084
rect 31611 8035 31653 8044
rect 34971 8084 35013 8093
rect 34971 8044 34972 8084
rect 35012 8044 35013 8084
rect 34971 8035 35013 8044
rect 43611 8084 43653 8093
rect 43611 8044 43612 8084
rect 43652 8044 43653 8084
rect 43611 8035 43653 8044
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 10923 8000 10965 8009
rect 10923 7960 10924 8000
rect 10964 7960 10965 8000
rect 10923 7951 10965 7960
rect 11307 8000 11349 8009
rect 11307 7960 11308 8000
rect 11348 7960 11349 8000
rect 11307 7951 11349 7960
rect 11787 8000 11829 8009
rect 11787 7960 11788 8000
rect 11828 7960 11829 8000
rect 11787 7951 11829 7960
rect 13899 8000 13941 8009
rect 13899 7960 13900 8000
rect 13940 7960 13941 8000
rect 13899 7951 13941 7960
rect 14475 8000 14517 8009
rect 14475 7960 14476 8000
rect 14516 7960 14517 8000
rect 14475 7951 14517 7960
rect 15706 8000 15764 8001
rect 15706 7960 15715 8000
rect 15755 7960 15764 8000
rect 15706 7959 15764 7960
rect 16186 8000 16244 8001
rect 16186 7960 16195 8000
rect 16235 7960 16244 8000
rect 16186 7959 16244 7960
rect 17163 8000 17205 8009
rect 17163 7960 17164 8000
rect 17204 7960 17205 8000
rect 17163 7951 17205 7960
rect 19659 8000 19701 8009
rect 19659 7960 19660 8000
rect 19700 7960 19701 8000
rect 19659 7951 19701 7960
rect 25995 8000 26037 8009
rect 25995 7960 25996 8000
rect 26036 7960 26037 8000
rect 25995 7951 26037 7960
rect 28779 8000 28821 8009
rect 28779 7960 28780 8000
rect 28820 7960 28821 8000
rect 28779 7951 28821 7960
rect 29163 8000 29205 8009
rect 29163 7960 29164 8000
rect 29204 7960 29205 8000
rect 29163 7951 29205 7960
rect 29434 8000 29492 8001
rect 29434 7960 29443 8000
rect 29483 7960 29492 8000
rect 29434 7959 29492 7960
rect 31467 8000 31509 8009
rect 31467 7960 31468 8000
rect 31508 7960 31509 8000
rect 31467 7951 31509 7960
rect 31851 8000 31893 8009
rect 31851 7960 31852 8000
rect 31892 7960 31893 8000
rect 31851 7951 31893 7960
rect 32235 8000 32277 8009
rect 32235 7960 32236 8000
rect 32276 7960 32277 8000
rect 32235 7951 32277 7960
rect 34635 8000 34677 8009
rect 34635 7960 34636 8000
rect 34676 7960 34677 8000
rect 34635 7951 34677 7960
rect 35211 8000 35253 8009
rect 35211 7960 35212 8000
rect 35252 7960 35253 8000
rect 35211 7951 35253 7960
rect 35595 8000 35637 8009
rect 35595 7960 35596 8000
rect 35636 7960 35637 8000
rect 35595 7951 35637 7960
rect 38379 8000 38421 8009
rect 38379 7960 38380 8000
rect 38420 7960 38421 8000
rect 38379 7951 38421 7960
rect 38955 8000 38997 8009
rect 38955 7960 38956 8000
rect 38996 7960 38997 8000
rect 38955 7951 38997 7960
rect 39819 8000 39861 8009
rect 39819 7960 39820 8000
rect 39860 7960 39861 8000
rect 39819 7951 39861 7960
rect 40155 8000 40197 8009
rect 40155 7960 40156 8000
rect 40196 7960 40197 8000
rect 40155 7951 40197 7960
rect 40395 8000 40437 8009
rect 40395 7960 40396 8000
rect 40436 7960 40437 8000
rect 40395 7951 40437 7960
rect 42315 8000 42357 8009
rect 42315 7960 42316 8000
rect 42356 7960 42357 8000
rect 42315 7951 42357 7960
rect 42699 8000 42741 8009
rect 42699 7960 42700 8000
rect 42740 7960 42741 8000
rect 42699 7951 42741 7960
rect 43083 8000 43125 8009
rect 43083 7960 43084 8000
rect 43124 7960 43125 8000
rect 43083 7951 43125 7960
rect 43467 8000 43509 8009
rect 43467 7960 43468 8000
rect 43508 7960 43509 8000
rect 43467 7951 43509 7960
rect 43851 8000 43893 8009
rect 43851 7960 43852 8000
rect 43892 7960 43893 8000
rect 43851 7951 43893 7960
rect 44235 8000 44277 8009
rect 44235 7960 44236 8000
rect 44276 7960 44277 8000
rect 44235 7951 44277 7960
rect 44619 8000 44661 8009
rect 44619 7960 44620 8000
rect 44660 7960 44661 8000
rect 44619 7951 44661 7960
rect 44907 8000 44949 8009
rect 44907 7960 44908 8000
rect 44948 7960 44949 8000
rect 44907 7951 44949 7960
rect 16674 7934 16720 7943
rect 12171 7916 12213 7925
rect 12171 7876 12172 7916
rect 12212 7876 12213 7916
rect 12171 7867 12213 7876
rect 13411 7916 13469 7917
rect 13411 7876 13420 7916
rect 13460 7876 13469 7916
rect 13411 7875 13469 7876
rect 14650 7916 14708 7917
rect 14650 7876 14659 7916
rect 14699 7876 14708 7916
rect 14650 7875 14708 7876
rect 14955 7916 14997 7925
rect 14955 7876 14956 7916
rect 14996 7876 14997 7916
rect 14955 7867 14997 7876
rect 15133 7916 15175 7925
rect 15133 7876 15134 7916
rect 15174 7876 15175 7916
rect 15133 7867 15175 7876
rect 15243 7916 15285 7925
rect 15243 7876 15244 7916
rect 15284 7876 15285 7916
rect 15243 7867 15285 7876
rect 15436 7916 15478 7925
rect 15436 7876 15437 7916
rect 15477 7876 15478 7916
rect 15436 7867 15478 7876
rect 15574 7916 15616 7925
rect 15574 7876 15575 7916
rect 15615 7876 15616 7916
rect 15574 7867 15616 7876
rect 15819 7916 15861 7925
rect 15819 7876 15820 7916
rect 15860 7876 15861 7916
rect 15819 7867 15861 7876
rect 16059 7916 16101 7925
rect 16059 7876 16060 7916
rect 16100 7876 16101 7916
rect 16059 7867 16101 7876
rect 16299 7916 16341 7925
rect 16299 7876 16300 7916
rect 16340 7876 16341 7916
rect 16674 7894 16675 7934
rect 16715 7894 16720 7934
rect 16674 7885 16720 7894
rect 16779 7916 16821 7925
rect 16299 7867 16341 7876
rect 16779 7876 16780 7916
rect 16820 7876 16821 7916
rect 16779 7867 16821 7876
rect 17259 7916 17301 7925
rect 17259 7876 17260 7916
rect 17300 7876 17301 7916
rect 17259 7867 17301 7876
rect 17731 7916 17789 7917
rect 17731 7876 17740 7916
rect 17780 7876 17789 7916
rect 17731 7875 17789 7876
rect 18219 7916 18277 7917
rect 18219 7876 18228 7916
rect 18268 7876 18277 7916
rect 18219 7875 18277 7876
rect 18603 7916 18645 7925
rect 18603 7876 18604 7916
rect 18644 7876 18645 7916
rect 18603 7867 18645 7876
rect 18795 7916 18837 7925
rect 18795 7876 18796 7916
rect 18836 7876 18837 7916
rect 18795 7867 18837 7876
rect 20227 7916 20285 7917
rect 20227 7876 20236 7916
rect 20276 7876 20285 7916
rect 20227 7875 20285 7876
rect 21483 7916 21525 7925
rect 21483 7876 21484 7916
rect 21524 7876 21525 7916
rect 21483 7867 21525 7876
rect 29307 7916 29349 7925
rect 29307 7876 29308 7916
rect 29348 7876 29349 7916
rect 29307 7867 29349 7876
rect 29547 7916 29589 7925
rect 29547 7876 29548 7916
rect 29588 7876 29589 7916
rect 29547 7867 29589 7876
rect 29835 7916 29877 7925
rect 29835 7876 29836 7916
rect 29876 7876 29877 7916
rect 29835 7867 29877 7876
rect 29950 7916 29992 7925
rect 29950 7876 29951 7916
rect 29991 7876 29992 7916
rect 29950 7867 29992 7876
rect 30123 7916 30165 7925
rect 30123 7876 30124 7916
rect 30164 7876 30165 7916
rect 30123 7867 30165 7876
rect 30315 7916 30357 7925
rect 30315 7876 30316 7916
rect 30356 7876 30357 7916
rect 30315 7867 30357 7876
rect 30507 7916 30549 7925
rect 30507 7876 30508 7916
rect 30548 7876 30549 7916
rect 30507 7867 30549 7876
rect 12027 7832 12069 7841
rect 12027 7792 12028 7832
rect 12068 7792 12069 7832
rect 12027 7783 12069 7792
rect 14139 7832 14181 7841
rect 14139 7792 14140 7832
rect 14180 7792 14181 7832
rect 14139 7783 14181 7792
rect 14859 7832 14901 7841
rect 14859 7792 14860 7832
rect 14900 7792 14901 7832
rect 14859 7783 14901 7792
rect 16378 7832 16436 7833
rect 16378 7792 16387 7832
rect 16427 7792 16436 7832
rect 16378 7791 16436 7792
rect 37227 7832 37269 7841
rect 37227 7792 37228 7832
rect 37268 7792 37269 7832
rect 37227 7783 37269 7792
rect 37515 7832 37557 7841
rect 37515 7792 37516 7832
rect 37556 7792 37557 7832
rect 37515 7783 37557 7792
rect 37803 7832 37845 7841
rect 37803 7792 37804 7832
rect 37844 7792 37845 7832
rect 37803 7783 37845 7792
rect 38091 7832 38133 7841
rect 38091 7792 38092 7832
rect 38132 7792 38133 7832
rect 38091 7783 38133 7792
rect 40059 7832 40101 7841
rect 40059 7792 40060 7832
rect 40100 7792 40101 7832
rect 40059 7783 40101 7792
rect 42843 7832 42885 7841
rect 42843 7792 42844 7832
rect 42884 7792 42885 7832
rect 42843 7783 42885 7792
rect 43995 7832 44037 7841
rect 43995 7792 43996 7832
rect 44036 7792 44037 7832
rect 43995 7783 44037 7792
rect 1467 7748 1509 7757
rect 1467 7708 1468 7748
rect 1508 7708 1509 7748
rect 1467 7699 1509 7708
rect 1851 7748 1893 7757
rect 1851 7708 1852 7748
rect 1892 7708 1893 7748
rect 1851 7699 1893 7708
rect 11547 7748 11589 7757
rect 11547 7708 11548 7748
rect 11588 7708 11589 7748
rect 11547 7699 11589 7708
rect 13611 7748 13653 7757
rect 13611 7708 13612 7748
rect 13652 7708 13653 7748
rect 13611 7699 13653 7708
rect 15898 7748 15956 7749
rect 15898 7708 15907 7748
rect 15947 7708 15956 7748
rect 15898 7707 15956 7708
rect 18411 7748 18453 7757
rect 18411 7708 18412 7748
rect 18452 7708 18453 7748
rect 18411 7699 18453 7708
rect 20043 7748 20085 7757
rect 20043 7708 20044 7748
rect 20084 7708 20085 7748
rect 20043 7699 20085 7708
rect 26235 7748 26277 7757
rect 26235 7708 26236 7748
rect 26276 7708 26277 7748
rect 26235 7699 26277 7708
rect 29626 7748 29684 7749
rect 29626 7708 29635 7748
rect 29675 7708 29684 7748
rect 29626 7707 29684 7708
rect 30411 7748 30453 7757
rect 30411 7708 30412 7748
rect 30452 7708 30453 7748
rect 30411 7699 30453 7708
rect 38619 7748 38661 7757
rect 38619 7708 38620 7748
rect 38660 7708 38661 7748
rect 38619 7699 38661 7708
rect 39195 7748 39237 7757
rect 39195 7708 39196 7748
rect 39236 7708 39237 7748
rect 39195 7699 39237 7708
rect 42075 7748 42117 7757
rect 42075 7708 42076 7748
rect 42116 7708 42117 7748
rect 42075 7699 42117 7708
rect 42459 7748 42501 7757
rect 42459 7708 42460 7748
rect 42500 7708 42501 7748
rect 42459 7699 42501 7708
rect 44379 7748 44421 7757
rect 44379 7708 44380 7748
rect 44420 7708 44421 7748
rect 44379 7699 44421 7708
rect 45147 7748 45189 7757
rect 45147 7708 45148 7748
rect 45188 7708 45189 7748
rect 45147 7699 45189 7708
rect 1152 7580 45216 7604
rect 1152 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 45216 7580
rect 1152 7516 45216 7540
rect 16954 7412 17012 7413
rect 16954 7372 16963 7412
rect 17003 7372 17012 7412
rect 16954 7371 17012 7372
rect 42778 7412 42836 7413
rect 42778 7372 42787 7412
rect 42827 7372 42836 7412
rect 42778 7371 42836 7372
rect 44218 7412 44276 7413
rect 44218 7372 44227 7412
rect 44267 7372 44276 7412
rect 44218 7371 44276 7372
rect 13035 7328 13077 7337
rect 13035 7288 13036 7328
rect 13076 7288 13077 7328
rect 13035 7279 13077 7288
rect 16107 7328 16149 7337
rect 16107 7288 16108 7328
rect 16148 7288 16149 7328
rect 16107 7279 16149 7288
rect 27339 7328 27381 7337
rect 27339 7288 27340 7328
rect 27380 7288 27381 7328
rect 27339 7279 27381 7288
rect 29067 7328 29109 7337
rect 29067 7288 29068 7328
rect 29108 7288 29109 7328
rect 29067 7279 29109 7288
rect 11595 7244 11637 7253
rect 15898 7244 15956 7245
rect 11595 7204 11596 7244
rect 11636 7204 11637 7244
rect 11595 7195 11637 7204
rect 12843 7235 12885 7244
rect 12843 7195 12844 7235
rect 12884 7195 12885 7235
rect 15898 7204 15907 7244
rect 15947 7204 15956 7244
rect 15898 7203 15956 7204
rect 16203 7244 16245 7253
rect 16203 7204 16204 7244
rect 16244 7204 16245 7244
rect 16203 7195 16245 7204
rect 16630 7244 16672 7253
rect 16630 7204 16631 7244
rect 16671 7204 16672 7244
rect 16630 7195 16672 7204
rect 16875 7244 16917 7253
rect 16875 7204 16876 7244
rect 16916 7204 16917 7244
rect 16875 7195 16917 7204
rect 25899 7244 25941 7253
rect 28491 7244 28533 7253
rect 25899 7204 25900 7244
rect 25940 7204 25941 7244
rect 25899 7195 25941 7204
rect 27147 7235 27189 7244
rect 27147 7195 27148 7235
rect 27188 7195 27189 7235
rect 28491 7204 28492 7244
rect 28532 7204 28533 7244
rect 28491 7195 28533 7204
rect 28666 7244 28724 7245
rect 28666 7204 28675 7244
rect 28715 7204 28724 7244
rect 28666 7203 28724 7204
rect 28854 7244 28896 7253
rect 28854 7204 28855 7244
rect 28895 7204 28896 7244
rect 28854 7195 28896 7204
rect 29163 7244 29205 7253
rect 29163 7204 29164 7244
rect 29204 7204 29205 7244
rect 29163 7195 29205 7204
rect 29354 7244 29396 7253
rect 29354 7204 29355 7244
rect 29395 7204 29396 7244
rect 29354 7195 29396 7204
rect 29643 7244 29685 7253
rect 29643 7204 29644 7244
rect 29684 7204 29685 7244
rect 29643 7195 29685 7204
rect 29930 7244 29972 7253
rect 29930 7204 29931 7244
rect 29971 7204 29972 7244
rect 29930 7195 29972 7204
rect 30160 7244 30218 7245
rect 30160 7204 30169 7244
rect 30209 7204 30218 7244
rect 30160 7203 30218 7204
rect 30490 7244 30548 7245
rect 31467 7244 31509 7253
rect 30490 7204 30499 7244
rect 30539 7204 30548 7244
rect 30490 7203 30548 7204
rect 30987 7235 31029 7244
rect 30987 7195 30988 7235
rect 31028 7195 31029 7235
rect 31467 7204 31468 7244
rect 31508 7204 31509 7244
rect 31467 7195 31509 7204
rect 31947 7244 31989 7253
rect 31947 7204 31948 7244
rect 31988 7204 31989 7244
rect 31947 7195 31989 7204
rect 32057 7244 32115 7245
rect 32057 7204 32066 7244
rect 32106 7204 32115 7244
rect 32057 7203 32115 7204
rect 12843 7186 12885 7195
rect 27147 7186 27189 7195
rect 30987 7186 31029 7195
rect 3435 7160 3477 7169
rect 3435 7120 3436 7160
rect 3476 7120 3477 7160
rect 3435 7111 3477 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 4059 7160 4101 7169
rect 4059 7120 4060 7160
rect 4100 7120 4101 7160
rect 4059 7111 4101 7120
rect 15051 7160 15093 7169
rect 15051 7120 15052 7160
rect 15092 7120 15093 7160
rect 15051 7111 15093 7120
rect 15483 7160 15525 7169
rect 15483 7120 15484 7160
rect 15524 7120 15525 7160
rect 15483 7111 15525 7120
rect 15723 7160 15765 7169
rect 15723 7120 15724 7160
rect 15764 7120 15765 7160
rect 15723 7111 15765 7120
rect 16762 7160 16820 7161
rect 16762 7120 16771 7160
rect 16811 7120 16820 7160
rect 16762 7119 16820 7120
rect 17499 7160 17541 7169
rect 17499 7120 17500 7160
rect 17540 7120 17541 7160
rect 17499 7111 17541 7120
rect 17739 7160 17781 7169
rect 17739 7120 17740 7160
rect 17780 7120 17781 7160
rect 17739 7111 17781 7120
rect 18123 7160 18165 7169
rect 18123 7120 18124 7160
rect 18164 7120 18165 7160
rect 18123 7111 18165 7120
rect 21867 7160 21909 7169
rect 21867 7120 21868 7160
rect 21908 7120 21909 7160
rect 21867 7111 21909 7120
rect 22155 7160 22197 7169
rect 22155 7120 22156 7160
rect 22196 7120 22197 7160
rect 22155 7111 22197 7120
rect 25515 7160 25557 7169
rect 25515 7120 25516 7160
rect 25556 7120 25557 7160
rect 25515 7111 25557 7120
rect 29835 7160 29877 7169
rect 31563 7160 31605 7169
rect 29835 7120 29836 7160
rect 29876 7120 29877 7160
rect 29835 7111 29877 7120
rect 30066 7151 30112 7160
rect 30066 7111 30067 7151
rect 30107 7111 30112 7151
rect 31563 7120 31564 7160
rect 31604 7120 31605 7160
rect 31563 7111 31605 7120
rect 35691 7160 35733 7169
rect 35691 7120 35692 7160
rect 35732 7120 35733 7160
rect 35691 7111 35733 7120
rect 38091 7160 38133 7169
rect 38091 7120 38092 7160
rect 38132 7120 38133 7160
rect 38091 7111 38133 7120
rect 38379 7160 38421 7169
rect 38379 7120 38380 7160
rect 38420 7120 38421 7160
rect 38379 7111 38421 7120
rect 38667 7160 38709 7169
rect 38667 7120 38668 7160
rect 38708 7120 38709 7160
rect 38667 7111 38709 7120
rect 39003 7160 39045 7169
rect 39003 7120 39004 7160
rect 39044 7120 39045 7160
rect 39003 7111 39045 7120
rect 39435 7160 39477 7169
rect 39435 7120 39436 7160
rect 39476 7120 39477 7160
rect 39435 7111 39477 7120
rect 39723 7160 39765 7169
rect 39723 7120 39724 7160
rect 39764 7120 39765 7160
rect 39723 7111 39765 7120
rect 40011 7160 40053 7169
rect 40011 7120 40012 7160
rect 40052 7120 40053 7160
rect 40011 7111 40053 7120
rect 40635 7160 40677 7169
rect 40635 7120 40636 7160
rect 40676 7120 40677 7160
rect 40635 7111 40677 7120
rect 40875 7160 40917 7169
rect 40875 7120 40876 7160
rect 40916 7120 40917 7160
rect 40875 7111 40917 7120
rect 42939 7160 42981 7169
rect 42939 7120 42940 7160
rect 42980 7120 42981 7160
rect 42939 7111 42981 7120
rect 43179 7160 43221 7169
rect 43179 7120 43180 7160
rect 43220 7120 43221 7160
rect 43179 7111 43221 7120
rect 43563 7160 43605 7169
rect 43563 7120 43564 7160
rect 43604 7120 43605 7160
rect 43563 7111 43605 7120
rect 43947 7160 43989 7169
rect 43947 7120 43948 7160
rect 43988 7120 43989 7160
rect 43947 7111 43989 7120
rect 44523 7160 44565 7169
rect 44523 7120 44524 7160
rect 44564 7120 44565 7160
rect 44523 7111 44565 7120
rect 44907 7160 44949 7169
rect 44907 7120 44908 7160
rect 44948 7120 44949 7160
rect 44907 7111 44949 7120
rect 30066 7102 30112 7111
rect 15291 7076 15333 7085
rect 15291 7036 15292 7076
rect 15332 7036 15333 7076
rect 15291 7027 15333 7036
rect 25755 7076 25797 7085
rect 25755 7036 25756 7076
rect 25796 7036 25797 7076
rect 25755 7027 25797 7036
rect 35451 7076 35493 7085
rect 35451 7036 35452 7076
rect 35492 7036 35493 7076
rect 35451 7027 35493 7036
rect 43323 7076 43365 7085
rect 43323 7036 43324 7076
rect 43364 7036 43365 7076
rect 43323 7027 43365 7036
rect 3675 6992 3717 7001
rect 3675 6952 3676 6992
rect 3716 6952 3717 6992
rect 3675 6943 3717 6952
rect 17883 6992 17925 7001
rect 17883 6952 17884 6992
rect 17924 6952 17925 6992
rect 17883 6943 17925 6952
rect 21627 6992 21669 7001
rect 21627 6952 21628 6992
rect 21668 6952 21669 6992
rect 21627 6943 21669 6952
rect 22395 6992 22437 7001
rect 22395 6952 22396 6992
rect 22436 6952 22437 6992
rect 22395 6943 22437 6952
rect 28666 6992 28724 6993
rect 28666 6952 28675 6992
rect 28715 6952 28724 6992
rect 28666 6951 28724 6952
rect 29355 6992 29397 7001
rect 29355 6952 29356 6992
rect 29396 6952 29397 6992
rect 29355 6943 29397 6952
rect 30267 6992 30309 7001
rect 30267 6952 30268 6992
rect 30308 6952 30309 6992
rect 30267 6943 30309 6952
rect 39291 6992 39333 7001
rect 39291 6952 39292 6992
rect 39332 6952 39333 6992
rect 39291 6943 39333 6952
rect 43707 6992 43749 7001
rect 43707 6952 43708 6992
rect 43748 6952 43749 6992
rect 43707 6943 43749 6952
rect 44763 6992 44805 7001
rect 44763 6952 44764 6992
rect 44804 6952 44805 6992
rect 44763 6943 44805 6952
rect 45147 6992 45189 7001
rect 45147 6952 45148 6992
rect 45188 6952 45189 6992
rect 45147 6943 45189 6952
rect 1152 6824 45216 6848
rect 1152 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 45216 6824
rect 1152 6760 45216 6784
rect 27627 6656 27669 6665
rect 27627 6616 27628 6656
rect 27668 6616 27669 6656
rect 27627 6607 27669 6616
rect 30010 6656 30068 6657
rect 30010 6616 30019 6656
rect 30059 6616 30068 6656
rect 30010 6615 30068 6616
rect 29403 6488 29445 6497
rect 29010 6479 29056 6488
rect 29010 6439 29011 6479
rect 29051 6439 29056 6479
rect 29403 6448 29404 6488
rect 29444 6448 29445 6488
rect 29403 6439 29445 6448
rect 29643 6488 29685 6497
rect 29643 6448 29644 6488
rect 29684 6448 29685 6488
rect 29643 6439 29685 6448
rect 31179 6488 31221 6497
rect 31179 6448 31180 6488
rect 31220 6448 31221 6488
rect 31179 6439 31221 6448
rect 34635 6488 34677 6497
rect 34635 6448 34636 6488
rect 34676 6448 34677 6488
rect 34635 6439 34677 6448
rect 34875 6488 34917 6497
rect 34875 6448 34876 6488
rect 34916 6448 34917 6488
rect 34875 6439 34917 6448
rect 35307 6488 35349 6497
rect 35307 6448 35308 6488
rect 35348 6448 35349 6488
rect 35307 6439 35349 6448
rect 35691 6488 35733 6497
rect 35691 6448 35692 6488
rect 35732 6448 35733 6488
rect 35691 6439 35733 6448
rect 37035 6488 37077 6497
rect 37035 6448 37036 6488
rect 37076 6448 37077 6488
rect 37035 6439 37077 6448
rect 41643 6488 41685 6497
rect 41643 6448 41644 6488
rect 41684 6448 41685 6488
rect 41643 6439 41685 6448
rect 44523 6488 44565 6497
rect 44523 6448 44524 6488
rect 44564 6448 44565 6488
rect 44523 6439 44565 6448
rect 44907 6488 44949 6497
rect 44907 6448 44908 6488
rect 44948 6448 44949 6488
rect 44907 6439 44949 6448
rect 29010 6430 29056 6439
rect 26187 6404 26229 6413
rect 26187 6364 26188 6404
rect 26228 6364 26229 6404
rect 26187 6355 26229 6364
rect 27427 6404 27485 6405
rect 27427 6364 27436 6404
rect 27476 6364 27485 6404
rect 27427 6363 27485 6364
rect 28875 6404 28917 6413
rect 28875 6364 28876 6404
rect 28916 6364 28917 6404
rect 28875 6355 28917 6364
rect 29104 6404 29162 6405
rect 29104 6364 29113 6404
rect 29153 6364 29162 6404
rect 29104 6363 29162 6364
rect 29842 6404 29884 6413
rect 29842 6364 29843 6404
rect 29883 6364 29884 6404
rect 29842 6355 29884 6364
rect 30010 6404 30068 6405
rect 30010 6364 30019 6404
rect 30059 6364 30068 6404
rect 30010 6363 30068 6364
rect 41883 6320 41925 6329
rect 41883 6280 41884 6320
rect 41924 6280 41925 6320
rect 41883 6271 41925 6280
rect 45147 6320 45189 6329
rect 45147 6280 45148 6320
rect 45188 6280 45189 6320
rect 45147 6271 45189 6280
rect 28779 6236 28821 6245
rect 28779 6196 28780 6236
rect 28820 6196 28821 6236
rect 28779 6187 28821 6196
rect 30939 6236 30981 6245
rect 30939 6196 30940 6236
rect 30980 6196 30981 6236
rect 30939 6187 30981 6196
rect 35547 6236 35589 6245
rect 35547 6196 35548 6236
rect 35588 6196 35589 6236
rect 35547 6187 35589 6196
rect 35931 6236 35973 6245
rect 35931 6196 35932 6236
rect 35972 6196 35973 6236
rect 35931 6187 35973 6196
rect 37275 6236 37317 6245
rect 37275 6196 37276 6236
rect 37316 6196 37317 6236
rect 37275 6187 37317 6196
rect 43546 6236 43604 6237
rect 43546 6196 43555 6236
rect 43595 6196 43604 6236
rect 43546 6195 43604 6196
rect 43834 6236 43892 6237
rect 43834 6196 43843 6236
rect 43883 6196 43892 6236
rect 43834 6195 43892 6196
rect 44122 6236 44180 6237
rect 44122 6196 44131 6236
rect 44171 6196 44180 6236
rect 44122 6195 44180 6196
rect 44763 6236 44805 6245
rect 44763 6196 44764 6236
rect 44804 6196 44805 6236
rect 44763 6187 44805 6196
rect 1152 6068 45216 6092
rect 1152 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 45216 6068
rect 1152 6004 45216 6028
rect 34635 5648 34677 5657
rect 34635 5608 34636 5648
rect 34676 5608 34677 5648
rect 34635 5599 34677 5608
rect 34875 5648 34917 5657
rect 34875 5608 34876 5648
rect 34916 5608 34917 5648
rect 34875 5599 34917 5608
rect 43131 5648 43173 5657
rect 43131 5608 43132 5648
rect 43172 5608 43173 5648
rect 43131 5599 43173 5608
rect 43371 5648 43413 5657
rect 43371 5608 43372 5648
rect 43412 5608 43413 5648
rect 43371 5599 43413 5608
rect 43563 5648 43605 5657
rect 43563 5608 43564 5648
rect 43604 5608 43605 5648
rect 43563 5599 43605 5608
rect 43851 5648 43893 5657
rect 43851 5608 43852 5648
rect 43892 5608 43893 5648
rect 43851 5599 43893 5608
rect 44139 5648 44181 5657
rect 44139 5608 44140 5648
rect 44180 5608 44181 5648
rect 44139 5599 44181 5608
rect 44523 5648 44565 5657
rect 44523 5608 44524 5648
rect 44564 5608 44565 5648
rect 44523 5599 44565 5608
rect 44907 5648 44949 5657
rect 44907 5608 44908 5648
rect 44948 5608 44949 5648
rect 44907 5599 44949 5608
rect 45147 5648 45189 5657
rect 45147 5608 45148 5648
rect 45188 5608 45189 5648
rect 45147 5599 45189 5608
rect 44763 5480 44805 5489
rect 44763 5440 44764 5480
rect 44804 5440 44805 5480
rect 44763 5431 44805 5440
rect 1152 5312 45216 5336
rect 1152 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 45216 5312
rect 1152 5248 45216 5272
rect 29067 5144 29109 5153
rect 29067 5104 29068 5144
rect 29108 5104 29109 5144
rect 29067 5095 29109 5104
rect 20811 4976 20853 4985
rect 20811 4936 20812 4976
rect 20852 4936 20853 4976
rect 20811 4927 20853 4936
rect 34731 4976 34773 4985
rect 34731 4936 34732 4976
rect 34772 4936 34773 4976
rect 34731 4927 34773 4936
rect 35019 4976 35061 4985
rect 35019 4936 35020 4976
rect 35060 4936 35061 4976
rect 35019 4927 35061 4936
rect 35307 4976 35349 4985
rect 35307 4936 35308 4976
rect 35348 4936 35349 4976
rect 35307 4927 35349 4936
rect 35499 4976 35541 4985
rect 35499 4936 35500 4976
rect 35540 4936 35541 4976
rect 35499 4927 35541 4936
rect 44523 4976 44565 4985
rect 44523 4936 44524 4976
rect 44564 4936 44565 4976
rect 44523 4927 44565 4936
rect 44907 4976 44949 4985
rect 44907 4936 44908 4976
rect 44948 4936 44949 4976
rect 44907 4927 44949 4936
rect 45147 4976 45189 4985
rect 45147 4936 45148 4976
rect 45188 4936 45189 4976
rect 45147 4927 45189 4936
rect 12843 4892 12885 4901
rect 12843 4852 12844 4892
rect 12884 4852 12885 4892
rect 12843 4843 12885 4852
rect 13018 4892 13076 4893
rect 13018 4852 13027 4892
rect 13067 4852 13076 4892
rect 13018 4851 13076 4852
rect 21195 4892 21237 4901
rect 21195 4852 21196 4892
rect 21236 4852 21237 4892
rect 21195 4843 21237 4852
rect 22435 4892 22493 4893
rect 22435 4852 22444 4892
rect 22484 4852 22493 4892
rect 22435 4851 22493 4852
rect 23307 4892 23349 4901
rect 23307 4852 23308 4892
rect 23348 4852 23349 4892
rect 23307 4843 23349 4852
rect 23482 4892 23540 4893
rect 23482 4852 23491 4892
rect 23531 4852 23540 4892
rect 23482 4851 23540 4852
rect 27627 4892 27669 4901
rect 27627 4852 27628 4892
rect 27668 4852 27669 4892
rect 27627 4843 27669 4852
rect 28867 4892 28925 4893
rect 28867 4852 28876 4892
rect 28916 4852 28925 4892
rect 28867 4851 28925 4852
rect 12939 4724 12981 4733
rect 12939 4684 12940 4724
rect 12980 4684 12981 4724
rect 12939 4675 12981 4684
rect 21051 4724 21093 4733
rect 21051 4684 21052 4724
rect 21092 4684 21093 4724
rect 21051 4675 21093 4684
rect 22635 4724 22677 4733
rect 22635 4684 22636 4724
rect 22676 4684 22677 4724
rect 22635 4675 22677 4684
rect 23403 4724 23445 4733
rect 23403 4684 23404 4724
rect 23444 4684 23445 4724
rect 23403 4675 23445 4684
rect 44763 4724 44805 4733
rect 44763 4684 44764 4724
rect 44804 4684 44805 4724
rect 44763 4675 44805 4684
rect 1152 4556 45216 4580
rect 1152 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 45216 4556
rect 1152 4492 45216 4516
rect 12123 4388 12165 4397
rect 12123 4348 12124 4388
rect 12164 4348 12165 4388
rect 12123 4339 12165 4348
rect 12843 4304 12885 4313
rect 12843 4264 12844 4304
rect 12884 4264 12885 4304
rect 12843 4255 12885 4264
rect 17595 4304 17637 4313
rect 17595 4264 17596 4304
rect 17636 4264 17637 4304
rect 17595 4255 17637 4264
rect 19275 4304 19317 4313
rect 19275 4264 19276 4304
rect 19316 4264 19317 4304
rect 19275 4255 19317 4264
rect 23482 4304 23540 4305
rect 23482 4264 23491 4304
rect 23531 4264 23540 4304
rect 23482 4263 23540 4264
rect 23691 4304 23733 4313
rect 23691 4264 23692 4304
rect 23732 4264 23733 4304
rect 23691 4255 23733 4264
rect 45147 4304 45189 4313
rect 45147 4264 45148 4304
rect 45188 4264 45189 4304
rect 45147 4255 45189 4264
rect 12634 4220 12692 4221
rect 12634 4180 12643 4220
rect 12683 4180 12692 4220
rect 12634 4179 12692 4180
rect 12939 4220 12981 4229
rect 12939 4180 12940 4220
rect 12980 4180 12981 4220
rect 12939 4171 12981 4180
rect 13129 4220 13171 4229
rect 13129 4180 13130 4220
rect 13170 4180 13171 4220
rect 13129 4171 13171 4180
rect 13246 4220 13288 4229
rect 13246 4180 13247 4220
rect 13287 4180 13288 4220
rect 13246 4171 13288 4180
rect 13419 4220 13461 4229
rect 13419 4180 13420 4220
rect 13460 4180 13461 4220
rect 13419 4171 13461 4180
rect 15094 4220 15136 4229
rect 15094 4180 15095 4220
rect 15135 4180 15136 4220
rect 15094 4171 15136 4180
rect 15339 4220 15381 4229
rect 15339 4180 15340 4220
rect 15380 4180 15381 4220
rect 15339 4171 15381 4180
rect 17835 4220 17877 4229
rect 22234 4220 22292 4221
rect 17835 4180 17836 4220
rect 17876 4180 17877 4220
rect 17835 4171 17877 4180
rect 19083 4211 19125 4220
rect 19083 4171 19084 4211
rect 19124 4171 19125 4211
rect 22234 4180 22243 4220
rect 22283 4180 22292 4220
rect 22234 4179 22292 4180
rect 22539 4220 22581 4229
rect 22539 4180 22540 4220
rect 22580 4180 22581 4220
rect 22539 4171 22581 4180
rect 22714 4220 22772 4221
rect 22714 4180 22723 4220
rect 22763 4180 22772 4220
rect 22714 4179 22772 4180
rect 22998 4220 23040 4229
rect 22998 4180 22999 4220
rect 23039 4180 23040 4220
rect 22998 4171 23040 4180
rect 23163 4220 23205 4229
rect 23163 4180 23164 4220
rect 23204 4180 23205 4220
rect 23163 4171 23205 4180
rect 23403 4220 23445 4229
rect 23403 4180 23404 4220
rect 23444 4180 23445 4220
rect 23403 4171 23445 4180
rect 23787 4220 23829 4229
rect 23787 4180 23788 4220
rect 23828 4180 23829 4220
rect 24171 4220 24213 4229
rect 23787 4171 23829 4180
rect 24027 4178 24069 4187
rect 19083 4162 19125 4171
rect 11883 4136 11925 4145
rect 11883 4096 11884 4136
rect 11924 4096 11925 4136
rect 11883 4087 11925 4096
rect 12267 4136 12309 4145
rect 12267 4096 12268 4136
rect 12308 4096 12309 4136
rect 12267 4087 12309 4096
rect 12507 4136 12549 4145
rect 12507 4096 12508 4136
rect 12548 4096 12549 4136
rect 12507 4087 12549 4096
rect 13611 4136 13653 4145
rect 13611 4096 13612 4136
rect 13652 4096 13653 4136
rect 13611 4087 13653 4096
rect 15226 4136 15284 4137
rect 15226 4096 15235 4136
rect 15275 4096 15284 4136
rect 15226 4095 15284 4096
rect 15435 4136 15477 4145
rect 15435 4096 15436 4136
rect 15476 4096 15477 4136
rect 15435 4087 15477 4096
rect 17355 4136 17397 4145
rect 17355 4096 17356 4136
rect 17396 4096 17397 4136
rect 17355 4087 17397 4096
rect 23290 4136 23348 4137
rect 23290 4096 23299 4136
rect 23339 4096 23348 4136
rect 23290 4095 23348 4096
rect 23906 4136 23948 4145
rect 23906 4096 23907 4136
rect 23947 4096 23948 4136
rect 24027 4138 24028 4178
rect 24068 4138 24069 4178
rect 24171 4180 24172 4220
rect 24212 4180 24213 4220
rect 24171 4171 24213 4180
rect 24346 4220 24404 4221
rect 24346 4180 24355 4220
rect 24395 4180 24404 4220
rect 24346 4179 24404 4180
rect 24562 4220 24620 4221
rect 24562 4180 24571 4220
rect 24611 4180 24620 4220
rect 24562 4179 24620 4180
rect 24747 4220 24789 4229
rect 24747 4180 24748 4220
rect 24788 4180 24789 4220
rect 24747 4171 24789 4180
rect 24027 4129 24069 4138
rect 27723 4136 27765 4145
rect 23906 4087 23948 4096
rect 27723 4096 27724 4136
rect 27764 4096 27765 4136
rect 27723 4087 27765 4096
rect 33291 4136 33333 4145
rect 33291 4096 33292 4136
rect 33332 4096 33333 4136
rect 33291 4087 33333 4096
rect 33531 4136 33573 4145
rect 33531 4096 33532 4136
rect 33572 4096 33573 4136
rect 33531 4087 33573 4096
rect 38571 4136 38613 4145
rect 38571 4096 38572 4136
rect 38612 4096 38613 4136
rect 38571 4087 38613 4096
rect 40491 4136 40533 4145
rect 40491 4096 40492 4136
rect 40532 4096 40533 4136
rect 40491 4087 40533 4096
rect 40875 4136 40917 4145
rect 40875 4096 40876 4136
rect 40916 4096 40917 4136
rect 40875 4087 40917 4096
rect 41259 4136 41301 4145
rect 41259 4096 41260 4136
rect 41300 4096 41301 4136
rect 41259 4087 41301 4096
rect 42123 4136 42165 4145
rect 42123 4096 42124 4136
rect 42164 4096 42165 4136
rect 42123 4087 42165 4096
rect 44523 4136 44565 4145
rect 44523 4096 44524 4136
rect 44564 4096 44565 4136
rect 44523 4087 44565 4096
rect 44907 4136 44949 4145
rect 44907 4096 44908 4136
rect 44948 4096 44949 4136
rect 44907 4087 44949 4096
rect 13323 4052 13365 4061
rect 13323 4012 13324 4052
rect 13364 4012 13365 4052
rect 13323 4003 13365 4012
rect 22539 4052 22581 4061
rect 22539 4012 22540 4052
rect 22580 4012 22581 4052
rect 22539 4003 22581 4012
rect 24346 4052 24404 4053
rect 24346 4012 24355 4052
rect 24395 4012 24404 4052
rect 24346 4011 24404 4012
rect 40251 4052 40293 4061
rect 40251 4012 40252 4052
rect 40292 4012 40293 4052
rect 40251 4003 40293 4012
rect 40635 4052 40677 4061
rect 40635 4012 40636 4052
rect 40676 4012 40677 4052
rect 40635 4003 40677 4012
rect 41019 4052 41061 4061
rect 41019 4012 41020 4052
rect 41060 4012 41061 4052
rect 41019 4003 41061 4012
rect 44763 4052 44805 4061
rect 44763 4012 44764 4052
rect 44804 4012 44805 4052
rect 44763 4003 44805 4012
rect 13851 3968 13893 3977
rect 13851 3928 13852 3968
rect 13892 3928 13893 3968
rect 13851 3919 13893 3928
rect 23019 3968 23061 3977
rect 23019 3928 23020 3968
rect 23060 3928 23061 3968
rect 23019 3919 23061 3928
rect 24555 3968 24597 3977
rect 24555 3928 24556 3968
rect 24596 3928 24597 3968
rect 24555 3919 24597 3928
rect 27963 3968 28005 3977
rect 27963 3928 27964 3968
rect 28004 3928 28005 3968
rect 27963 3919 28005 3928
rect 38331 3968 38373 3977
rect 38331 3928 38332 3968
rect 38372 3928 38373 3968
rect 38331 3919 38373 3928
rect 42363 3968 42405 3977
rect 42363 3928 42364 3968
rect 42404 3928 42405 3968
rect 42363 3919 42405 3928
rect 1152 3800 45216 3824
rect 1152 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 45216 3800
rect 1152 3736 45216 3760
rect 8955 3632 8997 3641
rect 8955 3592 8956 3632
rect 8996 3592 8997 3632
rect 8955 3583 8997 3592
rect 11547 3632 11589 3641
rect 11547 3592 11548 3632
rect 11588 3592 11589 3632
rect 11547 3583 11589 3592
rect 24075 3632 24117 3641
rect 24075 3592 24076 3632
rect 24116 3592 24117 3632
rect 24075 3583 24117 3592
rect 24891 3632 24933 3641
rect 24891 3592 24892 3632
rect 24932 3592 24933 3632
rect 24891 3583 24933 3592
rect 38715 3632 38757 3641
rect 38715 3592 38716 3632
rect 38756 3592 38757 3632
rect 38715 3583 38757 3592
rect 40539 3632 40581 3641
rect 40539 3592 40540 3632
rect 40580 3592 40581 3632
rect 40539 3583 40581 3592
rect 45147 3632 45189 3641
rect 45147 3592 45148 3632
rect 45188 3592 45189 3632
rect 45147 3583 45189 3592
rect 16203 3548 16245 3557
rect 16203 3508 16204 3548
rect 16244 3508 16245 3548
rect 16203 3499 16245 3508
rect 25851 3548 25893 3557
rect 25851 3508 25852 3548
rect 25892 3508 25893 3548
rect 25851 3499 25893 3508
rect 42363 3548 42405 3557
rect 42363 3508 42364 3548
rect 42404 3508 42405 3548
rect 42363 3499 42405 3508
rect 8715 3464 8757 3473
rect 8715 3424 8716 3464
rect 8756 3424 8757 3464
rect 8715 3415 8757 3424
rect 9387 3464 9429 3473
rect 9387 3424 9388 3464
rect 9428 3424 9429 3464
rect 9387 3415 9429 3424
rect 11787 3464 11829 3473
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 12555 3464 12597 3473
rect 12555 3424 12556 3464
rect 12596 3424 12597 3464
rect 12555 3415 12597 3424
rect 14746 3464 14804 3465
rect 14746 3424 14755 3464
rect 14795 3424 14804 3464
rect 14746 3423 14804 3424
rect 14955 3464 14997 3473
rect 14955 3424 14956 3464
rect 14996 3424 14997 3464
rect 14955 3415 14997 3424
rect 15819 3464 15861 3473
rect 15819 3424 15820 3464
rect 15860 3424 15861 3464
rect 15819 3415 15861 3424
rect 21243 3464 21285 3473
rect 21243 3424 21244 3464
rect 21284 3424 21285 3464
rect 21243 3415 21285 3424
rect 21483 3464 21525 3473
rect 21483 3424 21484 3464
rect 21524 3424 21525 3464
rect 21483 3415 21525 3424
rect 21867 3464 21909 3473
rect 21867 3424 21868 3464
rect 21908 3424 21909 3464
rect 21867 3415 21909 3424
rect 22635 3464 22677 3473
rect 22635 3424 22636 3464
rect 22676 3424 22677 3464
rect 22635 3415 22677 3424
rect 24747 3464 24789 3473
rect 24747 3424 24748 3464
rect 24788 3424 24789 3464
rect 24747 3415 24789 3424
rect 25131 3464 25173 3473
rect 25131 3424 25132 3464
rect 25172 3424 25173 3464
rect 25131 3415 25173 3424
rect 25611 3464 25653 3473
rect 25611 3424 25612 3464
rect 25652 3424 25653 3464
rect 25611 3415 25653 3424
rect 25978 3464 26036 3465
rect 25978 3424 25987 3464
rect 26027 3424 26036 3464
rect 25978 3423 26036 3424
rect 37851 3464 37893 3473
rect 37851 3424 37852 3464
rect 37892 3424 37893 3464
rect 37851 3415 37893 3424
rect 38091 3464 38133 3473
rect 38091 3424 38092 3464
rect 38132 3424 38133 3464
rect 38091 3415 38133 3424
rect 38475 3464 38517 3473
rect 38475 3424 38476 3464
rect 38516 3424 38517 3464
rect 38475 3415 38517 3424
rect 38955 3464 38997 3473
rect 38955 3424 38956 3464
rect 38996 3424 38997 3464
rect 38955 3415 38997 3424
rect 39435 3464 39477 3473
rect 39435 3424 39436 3464
rect 39476 3424 39477 3464
rect 39435 3415 39477 3424
rect 39723 3464 39765 3473
rect 39723 3424 39724 3464
rect 39764 3424 39765 3464
rect 39723 3415 39765 3424
rect 40011 3464 40053 3473
rect 40011 3424 40012 3464
rect 40052 3424 40053 3464
rect 40011 3415 40053 3424
rect 40299 3464 40341 3473
rect 40299 3424 40300 3464
rect 40340 3424 40341 3464
rect 40299 3415 40341 3424
rect 40875 3464 40917 3473
rect 40875 3424 40876 3464
rect 40916 3424 40917 3464
rect 40875 3415 40917 3424
rect 41355 3464 41397 3473
rect 41355 3424 41356 3464
rect 41396 3424 41397 3464
rect 41355 3415 41397 3424
rect 41739 3464 41781 3473
rect 41739 3424 41740 3464
rect 41780 3424 41781 3464
rect 41739 3415 41781 3424
rect 42123 3464 42165 3473
rect 42123 3424 42124 3464
rect 42164 3424 42165 3464
rect 42123 3415 42165 3424
rect 42507 3464 42549 3473
rect 42507 3424 42508 3464
rect 42548 3424 42549 3464
rect 42507 3415 42549 3424
rect 42891 3464 42933 3473
rect 42891 3424 42892 3464
rect 42932 3424 42933 3464
rect 42891 3415 42933 3424
rect 44523 3464 44565 3473
rect 44523 3424 44524 3464
rect 44564 3424 44565 3464
rect 44523 3415 44565 3424
rect 44907 3464 44949 3473
rect 44907 3424 44908 3464
rect 44948 3424 44949 3464
rect 44907 3415 44949 3424
rect 9771 3380 9813 3389
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 11011 3380 11069 3381
rect 11011 3340 11020 3380
rect 11060 3340 11069 3380
rect 11011 3339 11069 3340
rect 12058 3380 12116 3381
rect 12058 3340 12067 3380
rect 12107 3340 12116 3380
rect 12058 3339 12116 3340
rect 12171 3380 12213 3389
rect 12171 3340 12172 3380
rect 12212 3340 12213 3380
rect 12171 3331 12213 3340
rect 12651 3380 12693 3389
rect 12651 3340 12652 3380
rect 12692 3340 12693 3380
rect 12651 3331 12693 3340
rect 13123 3380 13181 3381
rect 13123 3340 13132 3380
rect 13172 3340 13181 3380
rect 13123 3339 13181 3340
rect 13611 3380 13669 3381
rect 13611 3340 13620 3380
rect 13660 3340 13669 3380
rect 13611 3339 13669 3340
rect 13978 3380 14036 3381
rect 13978 3340 13987 3380
rect 14027 3340 14036 3380
rect 13978 3339 14036 3340
rect 14283 3380 14325 3389
rect 14283 3340 14284 3380
rect 14324 3340 14325 3380
rect 14283 3331 14325 3340
rect 14614 3380 14656 3389
rect 14614 3340 14615 3380
rect 14655 3340 14656 3380
rect 14614 3331 14656 3340
rect 14859 3380 14901 3389
rect 14859 3340 14860 3380
rect 14900 3340 14901 3380
rect 14859 3331 14901 3340
rect 15243 3380 15285 3389
rect 15243 3340 15244 3380
rect 15284 3340 15285 3380
rect 15243 3331 15285 3340
rect 15418 3380 15476 3381
rect 15418 3340 15427 3380
rect 15467 3340 15476 3380
rect 15418 3339 15476 3340
rect 16387 3380 16445 3381
rect 16387 3340 16396 3380
rect 16436 3340 16445 3380
rect 16387 3339 16445 3340
rect 17603 3380 17645 3389
rect 17603 3340 17604 3380
rect 17644 3340 17645 3380
rect 17603 3331 17645 3340
rect 22125 3380 22167 3389
rect 22125 3340 22126 3380
rect 22166 3340 22167 3380
rect 22125 3331 22167 3340
rect 22251 3380 22293 3389
rect 22251 3340 22252 3380
rect 22292 3340 22293 3380
rect 22251 3331 22293 3340
rect 22731 3380 22773 3389
rect 22731 3340 22732 3380
rect 22772 3340 22773 3380
rect 22731 3331 22773 3340
rect 23203 3380 23261 3381
rect 23203 3340 23212 3380
rect 23252 3340 23261 3380
rect 23203 3339 23261 3340
rect 23691 3380 23749 3381
rect 23691 3340 23700 3380
rect 23740 3340 23749 3380
rect 23691 3339 23749 3340
rect 24075 3380 24117 3389
rect 24075 3340 24076 3380
rect 24116 3340 24117 3380
rect 24075 3331 24117 3340
rect 24190 3380 24232 3389
rect 24190 3340 24191 3380
rect 24231 3340 24232 3380
rect 24190 3331 24232 3340
rect 24363 3380 24405 3389
rect 24363 3340 24364 3380
rect 24404 3340 24405 3380
rect 24363 3331 24405 3340
rect 26179 3380 26237 3381
rect 26179 3340 26188 3380
rect 26228 3340 26237 3380
rect 26179 3339 26237 3340
rect 27435 3380 27477 3389
rect 27435 3340 27436 3380
rect 27476 3340 27477 3380
rect 27435 3331 27477 3340
rect 11211 3296 11253 3305
rect 11211 3256 11212 3296
rect 11252 3256 11253 3296
rect 11211 3247 11253 3256
rect 14187 3296 14229 3305
rect 14187 3256 14188 3296
rect 14228 3256 14229 3296
rect 14187 3247 14229 3256
rect 16059 3296 16101 3305
rect 16059 3256 16060 3296
rect 16100 3256 16101 3296
rect 16059 3247 16101 3256
rect 24507 3296 24549 3305
rect 24507 3256 24508 3296
rect 24548 3256 24549 3296
rect 24507 3247 24549 3256
rect 40635 3296 40677 3305
rect 40635 3256 40636 3296
rect 40676 3256 40677 3296
rect 40635 3247 40677 3256
rect 41979 3296 42021 3305
rect 41979 3256 41980 3296
rect 42020 3256 42021 3296
rect 41979 3247 42021 3256
rect 42747 3296 42789 3305
rect 42747 3256 42748 3296
rect 42788 3256 42789 3296
rect 42747 3247 42789 3256
rect 44763 3296 44805 3305
rect 44763 3256 44764 3296
rect 44804 3256 44805 3296
rect 44763 3247 44805 3256
rect 9627 3212 9669 3221
rect 9627 3172 9628 3212
rect 9668 3172 9669 3212
rect 9627 3163 9669 3172
rect 13803 3212 13845 3221
rect 13803 3172 13804 3212
rect 13844 3172 13845 3212
rect 13803 3163 13845 3172
rect 15339 3212 15381 3221
rect 15339 3172 15340 3212
rect 15380 3172 15381 3212
rect 15339 3163 15381 3172
rect 21627 3212 21669 3221
rect 21627 3172 21628 3212
rect 21668 3172 21669 3212
rect 21627 3163 21669 3172
rect 23883 3212 23925 3221
rect 23883 3172 23884 3212
rect 23924 3172 23925 3212
rect 23883 3163 23925 3172
rect 38235 3212 38277 3221
rect 38235 3172 38236 3212
rect 38276 3172 38277 3212
rect 38235 3163 38277 3172
rect 41595 3212 41637 3221
rect 41595 3172 41596 3212
rect 41636 3172 41637 3212
rect 41595 3163 41637 3172
rect 43131 3212 43173 3221
rect 43131 3172 43132 3212
rect 43172 3172 43173 3212
rect 43131 3163 43173 3172
rect 1152 3044 45216 3068
rect 1152 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 45216 3044
rect 1152 2980 45216 3004
rect 38907 2876 38949 2885
rect 38907 2836 38908 2876
rect 38948 2836 38949 2876
rect 38907 2827 38949 2836
rect 40090 2876 40148 2877
rect 40090 2836 40099 2876
rect 40139 2836 40148 2876
rect 40090 2835 40148 2836
rect 40299 2876 40341 2885
rect 40299 2836 40300 2876
rect 40340 2836 40341 2876
rect 40299 2827 40341 2836
rect 40587 2876 40629 2885
rect 40587 2836 40588 2876
rect 40628 2836 40629 2876
rect 40587 2827 40629 2836
rect 40875 2876 40917 2885
rect 40875 2836 40876 2876
rect 40916 2836 40917 2876
rect 40875 2827 40917 2836
rect 41163 2876 41205 2885
rect 41163 2836 41164 2876
rect 41204 2836 41205 2876
rect 41163 2827 41205 2836
rect 41451 2876 41493 2885
rect 41451 2836 41452 2876
rect 41492 2836 41493 2876
rect 41451 2827 41493 2836
rect 41722 2876 41780 2877
rect 41722 2836 41731 2876
rect 41771 2836 41780 2876
rect 41722 2835 41780 2836
rect 45147 2876 45189 2885
rect 45147 2836 45148 2876
rect 45188 2836 45189 2876
rect 45147 2827 45189 2836
rect 10539 2792 10581 2801
rect 10539 2752 10540 2792
rect 10580 2752 10581 2792
rect 10539 2743 10581 2752
rect 12027 2792 12069 2801
rect 12027 2752 12028 2792
rect 12068 2752 12069 2792
rect 12027 2743 12069 2752
rect 12891 2792 12933 2801
rect 12891 2752 12892 2792
rect 12932 2752 12933 2792
rect 12891 2743 12933 2752
rect 13786 2792 13844 2793
rect 13786 2752 13795 2792
rect 13835 2752 13844 2792
rect 13786 2751 13844 2752
rect 15051 2792 15093 2801
rect 15051 2752 15052 2792
rect 15092 2752 15093 2792
rect 15051 2743 15093 2752
rect 22683 2792 22725 2801
rect 22683 2752 22684 2792
rect 22724 2752 22725 2792
rect 22683 2743 22725 2752
rect 23386 2792 23444 2793
rect 23386 2752 23395 2792
rect 23435 2752 23444 2792
rect 23386 2751 23444 2752
rect 39291 2792 39333 2801
rect 39291 2752 39292 2792
rect 39332 2752 39333 2792
rect 39291 2743 39333 2752
rect 42747 2792 42789 2801
rect 42747 2752 42748 2792
rect 42788 2752 42789 2792
rect 42747 2743 42789 2752
rect 9099 2708 9141 2717
rect 13474 2708 13532 2709
rect 9099 2668 9100 2708
rect 9140 2668 9141 2708
rect 9099 2659 9141 2668
rect 10347 2699 10389 2708
rect 10347 2659 10348 2699
rect 10388 2659 10389 2699
rect 13474 2668 13483 2708
rect 13523 2668 13532 2708
rect 13474 2667 13532 2668
rect 13707 2708 13749 2717
rect 13707 2668 13708 2708
rect 13748 2668 13749 2708
rect 13707 2659 13749 2668
rect 14955 2708 14997 2717
rect 14955 2668 14956 2708
rect 14996 2668 14997 2708
rect 14955 2659 14997 2668
rect 15147 2708 15189 2717
rect 15147 2668 15148 2708
rect 15188 2668 15189 2708
rect 15147 2659 15189 2668
rect 23062 2708 23104 2717
rect 23062 2668 23063 2708
rect 23103 2668 23104 2708
rect 23062 2659 23104 2668
rect 23308 2708 23350 2717
rect 23308 2668 23309 2708
rect 23349 2668 23350 2708
rect 23308 2659 23350 2668
rect 10347 2650 10389 2659
rect 12267 2624 12309 2633
rect 12267 2584 12268 2624
rect 12308 2584 12309 2624
rect 12267 2575 12309 2584
rect 12651 2624 12693 2633
rect 12651 2584 12652 2624
rect 12692 2584 12693 2624
rect 12651 2575 12693 2584
rect 13594 2624 13652 2625
rect 13594 2584 13603 2624
rect 13643 2584 13652 2624
rect 13594 2583 13652 2584
rect 14187 2624 14229 2633
rect 14187 2584 14188 2624
rect 14228 2584 14229 2624
rect 14187 2575 14229 2584
rect 14475 2624 14517 2633
rect 14475 2584 14476 2624
rect 14516 2584 14517 2624
rect 14475 2575 14517 2584
rect 14715 2624 14757 2633
rect 14715 2584 14716 2624
rect 14756 2584 14757 2624
rect 14715 2575 14757 2584
rect 22539 2624 22581 2633
rect 22539 2584 22540 2624
rect 22580 2584 22581 2624
rect 22539 2575 22581 2584
rect 22923 2624 22965 2633
rect 22923 2584 22924 2624
rect 22964 2584 22965 2624
rect 22923 2575 22965 2584
rect 23194 2624 23252 2625
rect 23194 2584 23203 2624
rect 23243 2584 23252 2624
rect 23194 2583 23252 2584
rect 23787 2624 23829 2633
rect 23787 2584 23788 2624
rect 23828 2584 23829 2624
rect 23787 2575 23829 2584
rect 24171 2624 24213 2633
rect 24171 2584 24172 2624
rect 24212 2584 24213 2624
rect 24171 2575 24213 2584
rect 39147 2624 39189 2633
rect 39147 2584 39148 2624
rect 39188 2584 39189 2624
rect 39147 2575 39189 2584
rect 39531 2624 39573 2633
rect 39531 2584 39532 2624
rect 39572 2584 39573 2624
rect 39531 2575 39573 2584
rect 42123 2624 42165 2633
rect 42123 2584 42124 2624
rect 42164 2584 42165 2624
rect 42123 2575 42165 2584
rect 42507 2624 42549 2633
rect 42507 2584 42508 2624
rect 42548 2584 42549 2624
rect 42507 2575 42549 2584
rect 44139 2624 44181 2633
rect 44139 2584 44140 2624
rect 44180 2584 44181 2624
rect 44139 2575 44181 2584
rect 44523 2624 44565 2633
rect 44523 2584 44524 2624
rect 44564 2584 44565 2624
rect 44523 2575 44565 2584
rect 44907 2624 44949 2633
rect 44907 2584 44908 2624
rect 44948 2584 44949 2624
rect 44907 2575 44949 2584
rect 42363 2540 42405 2549
rect 42363 2500 42364 2540
rect 42404 2500 42405 2540
rect 42363 2491 42405 2500
rect 44763 2540 44805 2549
rect 44763 2500 44764 2540
rect 44804 2500 44805 2540
rect 44763 2491 44805 2500
rect 13947 2456 13989 2465
rect 13947 2416 13948 2456
rect 13988 2416 13989 2456
rect 13947 2407 13989 2416
rect 22299 2456 22341 2465
rect 22299 2416 22300 2456
rect 22340 2416 22341 2456
rect 22299 2407 22341 2416
rect 23547 2456 23589 2465
rect 23547 2416 23548 2456
rect 23588 2416 23589 2456
rect 23547 2407 23589 2416
rect 23931 2456 23973 2465
rect 23931 2416 23932 2456
rect 23972 2416 23973 2456
rect 23931 2407 23973 2416
rect 44379 2456 44421 2465
rect 44379 2416 44380 2456
rect 44420 2416 44421 2456
rect 44379 2407 44421 2416
rect 1152 2288 45216 2312
rect 1152 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 45216 2288
rect 1152 2224 45216 2248
rect 1755 2120 1797 2129
rect 1755 2080 1756 2120
rect 1796 2080 1797 2120
rect 1755 2071 1797 2080
rect 45147 2120 45189 2129
rect 45147 2080 45148 2120
rect 45188 2080 45189 2120
rect 45147 2071 45189 2080
rect 1515 1952 1557 1961
rect 1515 1912 1516 1952
rect 1556 1912 1557 1952
rect 1515 1903 1557 1912
rect 3435 1952 3477 1961
rect 3435 1912 3436 1952
rect 3476 1912 3477 1952
rect 3435 1903 3477 1912
rect 5163 1952 5205 1961
rect 5163 1912 5164 1952
rect 5204 1912 5205 1952
rect 5163 1903 5205 1912
rect 6891 1952 6933 1961
rect 6891 1912 6892 1952
rect 6932 1912 6933 1952
rect 6891 1903 6933 1912
rect 8619 1952 8661 1961
rect 8619 1912 8620 1952
rect 8660 1912 8661 1952
rect 8619 1903 8661 1912
rect 43371 1952 43413 1961
rect 43371 1912 43372 1952
rect 43412 1912 43413 1952
rect 43371 1903 43413 1912
rect 43755 1952 43797 1961
rect 43755 1912 43756 1952
rect 43796 1912 43797 1952
rect 43755 1903 43797 1912
rect 44139 1952 44181 1961
rect 44139 1912 44140 1952
rect 44180 1912 44181 1952
rect 44139 1903 44181 1912
rect 44523 1952 44565 1961
rect 44523 1912 44524 1952
rect 44564 1912 44565 1952
rect 44523 1903 44565 1912
rect 44907 1952 44949 1961
rect 44907 1912 44908 1952
rect 44948 1912 44949 1952
rect 44907 1903 44949 1912
rect 43995 1784 44037 1793
rect 43995 1744 43996 1784
rect 44036 1744 44037 1784
rect 43995 1735 44037 1744
rect 3195 1700 3237 1709
rect 3195 1660 3196 1700
rect 3236 1660 3237 1700
rect 3195 1651 3237 1660
rect 4923 1700 4965 1709
rect 4923 1660 4924 1700
rect 4964 1660 4965 1700
rect 4923 1651 4965 1660
rect 6651 1700 6693 1709
rect 6651 1660 6652 1700
rect 6692 1660 6693 1700
rect 6651 1651 6693 1660
rect 8379 1700 8421 1709
rect 8379 1660 8380 1700
rect 8420 1660 8421 1700
rect 8379 1651 8421 1660
rect 43611 1700 43653 1709
rect 43611 1660 43612 1700
rect 43652 1660 43653 1700
rect 43611 1651 43653 1660
rect 44379 1700 44421 1709
rect 44379 1660 44380 1700
rect 44420 1660 44421 1700
rect 44379 1651 44421 1660
rect 44763 1700 44805 1709
rect 44763 1660 44764 1700
rect 44804 1660 44805 1700
rect 44763 1651 44805 1660
rect 1152 1532 45216 1556
rect 1152 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 45216 1532
rect 1152 1468 45216 1492
<< via1 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 1852 9640 1892 9680
rect 3004 9640 3044 9680
rect 9628 9640 9668 9680
rect 11164 9640 11204 9680
rect 12700 9640 12740 9680
rect 13852 9640 13892 9680
rect 16156 9640 16196 9680
rect 17308 9640 17348 9680
rect 17692 9640 17732 9680
rect 18460 9640 18500 9680
rect 18844 9640 18884 9680
rect 19612 9640 19652 9680
rect 21532 9640 21572 9680
rect 22684 9640 22724 9680
rect 26620 9640 26660 9680
rect 30076 9640 30116 9680
rect 31228 9640 31268 9680
rect 31996 9640 32036 9680
rect 32764 9640 32804 9680
rect 33532 9640 33572 9680
rect 35452 9640 35492 9680
rect 36220 9640 36260 9680
rect 42844 9640 42884 9680
rect 43228 9640 43268 9680
rect 43612 9640 43652 9680
rect 43996 9640 44036 9680
rect 10012 9556 10052 9596
rect 13084 9556 13124 9596
rect 18076 9556 18116 9596
rect 19228 9556 19268 9596
rect 28924 9556 28964 9596
rect 31612 9556 31652 9596
rect 32380 9556 32420 9596
rect 35836 9556 35876 9596
rect 1228 9472 1268 9512
rect 1612 9472 1652 9512
rect 1996 9472 2036 9512
rect 2380 9472 2420 9512
rect 2764 9472 2804 9512
rect 3148 9472 3188 9512
rect 9388 9472 9428 9512
rect 9772 9472 9812 9512
rect 10156 9472 10196 9512
rect 10396 9472 10436 9512
rect 10540 9472 10580 9512
rect 10924 9472 10964 9512
rect 11308 9472 11348 9512
rect 11692 9472 11732 9512
rect 12076 9472 12116 9512
rect 12460 9472 12500 9512
rect 12844 9472 12884 9512
rect 13228 9472 13268 9512
rect 13468 9472 13508 9512
rect 13612 9472 13652 9512
rect 13996 9472 14036 9512
rect 14380 9472 14420 9512
rect 14764 9472 14804 9512
rect 15004 9472 15044 9512
rect 15148 9472 15188 9512
rect 15532 9472 15572 9512
rect 15916 9472 15956 9512
rect 16300 9472 16340 9512
rect 16684 9472 16724 9512
rect 16924 9472 16964 9512
rect 17068 9472 17108 9512
rect 17452 9472 17492 9512
rect 17836 9472 17876 9512
rect 18220 9472 18260 9512
rect 18604 9472 18644 9512
rect 18988 9472 19028 9512
rect 19372 9472 19412 9512
rect 19756 9472 19796 9512
rect 20524 9472 20564 9512
rect 20764 9472 20804 9512
rect 21100 9472 21140 9512
rect 21292 9472 21332 9512
rect 21868 9472 21908 9512
rect 22252 9472 22292 9512
rect 22444 9472 22484 9512
rect 23020 9472 23060 9512
rect 23404 9472 23444 9512
rect 23788 9472 23828 9512
rect 23980 9472 24020 9512
rect 24364 9472 24404 9512
rect 24940 9472 24980 9512
rect 25324 9472 25364 9512
rect 25516 9472 25556 9512
rect 25852 9472 25892 9512
rect 26092 9472 26132 9512
rect 26476 9472 26516 9512
rect 26860 9472 26900 9512
rect 27244 9472 27284 9512
rect 28396 9472 28436 9512
rect 28540 9472 28580 9512
rect 28780 9472 28820 9512
rect 29164 9472 29204 9512
rect 29356 9472 29396 9512
rect 29692 9472 29732 9512
rect 29932 9472 29972 9512
rect 30316 9472 30356 9512
rect 30700 9472 30740 9512
rect 31468 9472 31508 9512
rect 31852 9472 31892 9512
rect 32236 9472 32276 9512
rect 32620 9472 32660 9512
rect 33004 9472 33044 9512
rect 33388 9472 33428 9512
rect 33772 9472 33812 9512
rect 34156 9472 34196 9512
rect 34483 9472 34523 9512
rect 34684 9472 34724 9512
rect 34972 9472 35012 9512
rect 35308 9472 35348 9512
rect 35692 9472 35732 9512
rect 36076 9472 36116 9512
rect 36460 9472 36500 9512
rect 41836 9472 41876 9512
rect 42220 9472 42260 9512
rect 42604 9472 42644 9512
rect 42988 9472 43028 9512
rect 43372 9472 43412 9512
rect 43756 9472 43796 9512
rect 44140 9472 44180 9512
rect 44908 9472 44948 9512
rect 44620 9388 44660 9428
rect 2236 9304 2276 9344
rect 3388 9304 3428 9344
rect 11548 9304 11588 9344
rect 11932 9304 11972 9344
rect 14236 9304 14276 9344
rect 14620 9304 14660 9344
rect 16540 9304 16580 9344
rect 19996 9304 20036 9344
rect 20860 9304 20900 9344
rect 22012 9304 22052 9344
rect 23548 9304 23588 9344
rect 24220 9304 24260 9344
rect 24604 9304 24644 9344
rect 25084 9304 25124 9344
rect 25756 9304 25796 9344
rect 29596 9304 29636 9344
rect 33148 9304 33188 9344
rect 35068 9304 35108 9344
rect 42460 9304 42500 9344
rect 44380 9304 44420 9344
rect 1468 9220 1508 9260
rect 2620 9220 2660 9260
rect 10780 9220 10820 9260
rect 12316 9220 12356 9260
rect 15388 9220 15428 9260
rect 15772 9220 15812 9260
rect 20332 9220 20372 9260
rect 21628 9220 21668 9260
rect 22780 9220 22820 9260
rect 23164 9220 23204 9260
rect 24700 9220 24740 9260
rect 26236 9220 26276 9260
rect 27004 9220 27044 9260
rect 28156 9220 28196 9260
rect 30460 9220 30500 9260
rect 33916 9220 33956 9260
rect 34300 9220 34340 9260
rect 40483 9220 40523 9260
rect 40675 9220 40715 9260
rect 40963 9220 41003 9260
rect 41251 9220 41291 9260
rect 41539 9220 41579 9260
rect 42076 9220 42116 9260
rect 45148 9220 45188 9260
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 1468 8884 1508 8924
rect 3196 8884 3236 8924
rect 10300 8884 10340 8924
rect 11068 8884 11108 8924
rect 12604 8884 12644 8924
rect 14140 8884 14180 8924
rect 15148 8884 15188 8924
rect 15868 8884 15908 8924
rect 16252 8884 16292 8924
rect 18460 8884 18500 8924
rect 18844 8884 18884 8924
rect 19228 8884 19268 8924
rect 19612 8884 19652 8924
rect 19996 8884 20036 8924
rect 20380 8884 20420 8924
rect 20764 8884 20804 8924
rect 21436 8884 21476 8924
rect 29596 8884 29636 8924
rect 32188 8884 32228 8924
rect 32572 8884 32612 8924
rect 32956 8884 32996 8924
rect 33340 8884 33380 8924
rect 33724 8884 33764 8924
rect 34108 8884 34148 8924
rect 35740 8884 35780 8924
rect 43036 8884 43076 8924
rect 43420 8884 43460 8924
rect 1852 8800 1892 8840
rect 3580 8800 3620 8840
rect 11452 8800 11492 8840
rect 12220 8800 12260 8840
rect 12988 8800 13028 8840
rect 17980 8800 18020 8840
rect 23164 8800 23204 8840
rect 25276 8800 25316 8840
rect 25948 8800 25988 8840
rect 34492 8800 34532 8840
rect 35356 8800 35396 8840
rect 38092 8800 38132 8840
rect 38524 8800 38564 8840
rect 44380 8800 44420 8840
rect 15052 8716 15092 8756
rect 15235 8716 15275 8756
rect 17644 8716 17684 8756
rect 17836 8716 17876 8756
rect 41260 8716 41300 8756
rect 41644 8716 41684 8756
rect 41932 8716 41972 8756
rect 42220 8716 42260 8756
rect 42508 8716 42548 8756
rect 1228 8632 1268 8672
rect 1612 8632 1652 8672
rect 1996 8632 2036 8672
rect 2380 8632 2420 8672
rect 2620 8632 2660 8672
rect 2956 8632 2996 8672
rect 3340 8632 3380 8672
rect 10060 8632 10100 8672
rect 10444 8632 10484 8672
rect 10828 8632 10868 8672
rect 11212 8632 11252 8672
rect 11596 8632 11636 8672
rect 11980 8632 12020 8672
rect 12364 8632 12404 8672
rect 12748 8632 12788 8672
rect 13132 8632 13172 8672
rect 13516 8632 13556 8672
rect 13756 8632 13796 8672
rect 13900 8632 13940 8672
rect 14284 8632 14324 8672
rect 14524 8632 14564 8672
rect 14668 8632 14708 8672
rect 15628 8632 15668 8672
rect 16012 8632 16052 8672
rect 16396 8632 16436 8672
rect 16636 8632 16676 8672
rect 17260 8632 17300 8672
rect 18220 8632 18260 8672
rect 18700 8632 18740 8672
rect 19084 8632 19124 8672
rect 19468 8632 19508 8672
rect 19852 8632 19892 8672
rect 20236 8632 20276 8672
rect 20620 8632 20660 8672
rect 21004 8632 21044 8672
rect 21196 8632 21236 8672
rect 21868 8632 21908 8672
rect 22060 8632 22100 8672
rect 22300 8632 22340 8672
rect 22780 8632 22820 8672
rect 23020 8632 23060 8672
rect 23404 8632 23444 8672
rect 23548 8632 23588 8672
rect 23788 8632 23828 8672
rect 25516 8632 25556 8672
rect 25708 8632 25748 8672
rect 26284 8632 26324 8672
rect 26476 8632 26516 8672
rect 26716 8632 26756 8672
rect 29356 8632 29396 8672
rect 29836 8632 29876 8672
rect 32428 8632 32468 8672
rect 32812 8632 32852 8672
rect 33196 8632 33236 8672
rect 33580 8632 33620 8672
rect 33964 8632 34004 8672
rect 34348 8632 34388 8672
rect 34732 8632 34772 8672
rect 35116 8632 35156 8672
rect 35539 8632 35579 8672
rect 38092 8632 38132 8672
rect 38284 8632 38324 8672
rect 38764 8632 38804 8672
rect 39052 8632 39092 8672
rect 39340 8632 39380 8672
rect 39628 8632 39668 8672
rect 39916 8632 39956 8672
rect 40204 8632 40244 8672
rect 40492 8632 40532 8672
rect 40780 8632 40820 8672
rect 40972 8632 41012 8672
rect 42652 8632 42692 8672
rect 42892 8632 42932 8672
rect 43276 8632 43316 8672
rect 43660 8632 43700 8672
rect 43948 8632 43988 8672
rect 44140 8632 44180 8672
rect 44524 8632 44564 8672
rect 44908 8632 44948 8672
rect 2236 8548 2276 8588
rect 10684 8548 10724 8588
rect 13372 8548 13412 8588
rect 14908 8548 14948 8588
rect 17020 8548 17060 8588
rect 21628 8548 21668 8588
rect 44764 8548 44804 8588
rect 11836 8464 11876 8504
rect 17644 8464 17684 8504
rect 26044 8464 26084 8504
rect 29116 8464 29156 8504
rect 45148 8464 45188 8504
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 11164 8128 11204 8168
rect 14236 8128 14276 8168
rect 18604 8128 18644 8168
rect 28540 8128 28580 8168
rect 28924 8128 28964 8168
rect 31228 8128 31268 8168
rect 31996 8128 32036 8168
rect 34876 8128 34916 8168
rect 35356 8128 35396 8168
rect 43228 8128 43268 8168
rect 15340 8044 15380 8084
rect 19900 8044 19940 8084
rect 29836 8044 29876 8084
rect 31612 8044 31652 8084
rect 34972 8044 35012 8084
rect 43612 8044 43652 8084
rect 1228 7960 1268 8000
rect 1612 7960 1652 8000
rect 10924 7960 10964 8000
rect 11308 7960 11348 8000
rect 11788 7960 11828 8000
rect 13900 7960 13940 8000
rect 14476 7960 14516 8000
rect 15715 7960 15755 8000
rect 16195 7960 16235 8000
rect 17164 7960 17204 8000
rect 19660 7960 19700 8000
rect 25996 7960 26036 8000
rect 28780 7960 28820 8000
rect 29164 7960 29204 8000
rect 29443 7960 29483 8000
rect 31468 7960 31508 8000
rect 31852 7960 31892 8000
rect 32236 7960 32276 8000
rect 34636 7960 34676 8000
rect 35212 7960 35252 8000
rect 35596 7960 35636 8000
rect 38380 7960 38420 8000
rect 38956 7960 38996 8000
rect 39820 7960 39860 8000
rect 40156 7960 40196 8000
rect 40396 7960 40436 8000
rect 42316 7960 42356 8000
rect 42700 7960 42740 8000
rect 43084 7960 43124 8000
rect 43468 7960 43508 8000
rect 43852 7960 43892 8000
rect 44236 7960 44276 8000
rect 44620 7960 44660 8000
rect 44908 7960 44948 8000
rect 12172 7876 12212 7916
rect 13420 7876 13460 7916
rect 14659 7876 14699 7916
rect 14956 7876 14996 7916
rect 15134 7876 15174 7916
rect 15244 7876 15284 7916
rect 15437 7876 15477 7916
rect 15575 7876 15615 7916
rect 15820 7876 15860 7916
rect 16060 7876 16100 7916
rect 16300 7876 16340 7916
rect 16675 7894 16715 7934
rect 16780 7876 16820 7916
rect 17260 7876 17300 7916
rect 17740 7876 17780 7916
rect 18228 7876 18268 7916
rect 18604 7876 18644 7916
rect 18796 7876 18836 7916
rect 20236 7876 20276 7916
rect 21484 7876 21524 7916
rect 29308 7876 29348 7916
rect 29548 7876 29588 7916
rect 29836 7876 29876 7916
rect 29951 7876 29991 7916
rect 30124 7876 30164 7916
rect 30316 7876 30356 7916
rect 30508 7876 30548 7916
rect 12028 7792 12068 7832
rect 14140 7792 14180 7832
rect 14860 7792 14900 7832
rect 16387 7792 16427 7832
rect 37228 7792 37268 7832
rect 37516 7792 37556 7832
rect 37804 7792 37844 7832
rect 38092 7792 38132 7832
rect 40060 7792 40100 7832
rect 42844 7792 42884 7832
rect 43996 7792 44036 7832
rect 1468 7708 1508 7748
rect 1852 7708 1892 7748
rect 11548 7708 11588 7748
rect 13612 7708 13652 7748
rect 15907 7708 15947 7748
rect 18412 7708 18452 7748
rect 20044 7708 20084 7748
rect 26236 7708 26276 7748
rect 29635 7708 29675 7748
rect 30412 7708 30452 7748
rect 38620 7708 38660 7748
rect 39196 7708 39236 7748
rect 42076 7708 42116 7748
rect 42460 7708 42500 7748
rect 44380 7708 44420 7748
rect 45148 7708 45188 7748
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 16963 7372 17003 7412
rect 42787 7372 42827 7412
rect 44227 7372 44267 7412
rect 13036 7288 13076 7328
rect 16108 7288 16148 7328
rect 27340 7288 27380 7328
rect 29068 7288 29108 7328
rect 11596 7204 11636 7244
rect 12844 7195 12884 7235
rect 15907 7204 15947 7244
rect 16204 7204 16244 7244
rect 16631 7204 16671 7244
rect 16876 7204 16916 7244
rect 25900 7204 25940 7244
rect 27148 7195 27188 7235
rect 28492 7204 28532 7244
rect 28675 7204 28715 7244
rect 28855 7204 28895 7244
rect 29164 7204 29204 7244
rect 29355 7204 29395 7244
rect 29644 7204 29684 7244
rect 29931 7204 29971 7244
rect 30169 7204 30209 7244
rect 30499 7204 30539 7244
rect 30988 7195 31028 7235
rect 31468 7204 31508 7244
rect 31948 7204 31988 7244
rect 32066 7204 32106 7244
rect 3436 7120 3476 7160
rect 3820 7120 3860 7160
rect 4060 7120 4100 7160
rect 15052 7120 15092 7160
rect 15484 7120 15524 7160
rect 15724 7120 15764 7160
rect 16771 7120 16811 7160
rect 17500 7120 17540 7160
rect 17740 7120 17780 7160
rect 18124 7120 18164 7160
rect 21868 7120 21908 7160
rect 22156 7120 22196 7160
rect 25516 7120 25556 7160
rect 29836 7120 29876 7160
rect 30067 7111 30107 7151
rect 31564 7120 31604 7160
rect 35692 7120 35732 7160
rect 38092 7120 38132 7160
rect 38380 7120 38420 7160
rect 38668 7120 38708 7160
rect 39004 7120 39044 7160
rect 39436 7120 39476 7160
rect 39724 7120 39764 7160
rect 40012 7120 40052 7160
rect 40636 7120 40676 7160
rect 40876 7120 40916 7160
rect 42940 7120 42980 7160
rect 43180 7120 43220 7160
rect 43564 7120 43604 7160
rect 43948 7120 43988 7160
rect 44524 7120 44564 7160
rect 44908 7120 44948 7160
rect 15292 7036 15332 7076
rect 25756 7036 25796 7076
rect 35452 7036 35492 7076
rect 43324 7036 43364 7076
rect 3676 6952 3716 6992
rect 17884 6952 17924 6992
rect 21628 6952 21668 6992
rect 22396 6952 22436 6992
rect 28675 6952 28715 6992
rect 29356 6952 29396 6992
rect 30268 6952 30308 6992
rect 39292 6952 39332 6992
rect 43708 6952 43748 6992
rect 44764 6952 44804 6992
rect 45148 6952 45188 6992
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 27628 6616 27668 6656
rect 30019 6616 30059 6656
rect 29011 6439 29051 6479
rect 29404 6448 29444 6488
rect 29644 6448 29684 6488
rect 31180 6448 31220 6488
rect 34636 6448 34676 6488
rect 34876 6448 34916 6488
rect 35308 6448 35348 6488
rect 35692 6448 35732 6488
rect 37036 6448 37076 6488
rect 41644 6448 41684 6488
rect 44524 6448 44564 6488
rect 44908 6448 44948 6488
rect 26188 6364 26228 6404
rect 27436 6364 27476 6404
rect 28876 6364 28916 6404
rect 29113 6364 29153 6404
rect 29843 6364 29883 6404
rect 30019 6364 30059 6404
rect 41884 6280 41924 6320
rect 45148 6280 45188 6320
rect 28780 6196 28820 6236
rect 30940 6196 30980 6236
rect 35548 6196 35588 6236
rect 35932 6196 35972 6236
rect 37276 6196 37316 6236
rect 43555 6196 43595 6236
rect 43843 6196 43883 6236
rect 44131 6196 44171 6236
rect 44764 6196 44804 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 34636 5608 34676 5648
rect 34876 5608 34916 5648
rect 43132 5608 43172 5648
rect 43372 5608 43412 5648
rect 43564 5608 43604 5648
rect 43852 5608 43892 5648
rect 44140 5608 44180 5648
rect 44524 5608 44564 5648
rect 44908 5608 44948 5648
rect 45148 5608 45188 5648
rect 44764 5440 44804 5480
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 29068 5104 29108 5144
rect 20812 4936 20852 4976
rect 34732 4936 34772 4976
rect 35020 4936 35060 4976
rect 35308 4936 35348 4976
rect 35500 4936 35540 4976
rect 44524 4936 44564 4976
rect 44908 4936 44948 4976
rect 45148 4936 45188 4976
rect 12844 4852 12884 4892
rect 13027 4852 13067 4892
rect 21196 4852 21236 4892
rect 22444 4852 22484 4892
rect 23308 4852 23348 4892
rect 23491 4852 23531 4892
rect 27628 4852 27668 4892
rect 28876 4852 28916 4892
rect 12940 4684 12980 4724
rect 21052 4684 21092 4724
rect 22636 4684 22676 4724
rect 23404 4684 23444 4724
rect 44764 4684 44804 4724
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 12124 4348 12164 4388
rect 12844 4264 12884 4304
rect 17596 4264 17636 4304
rect 19276 4264 19316 4304
rect 23491 4264 23531 4304
rect 23692 4264 23732 4304
rect 45148 4264 45188 4304
rect 12643 4180 12683 4220
rect 12940 4180 12980 4220
rect 13130 4180 13170 4220
rect 13247 4180 13287 4220
rect 13420 4180 13460 4220
rect 15095 4180 15135 4220
rect 15340 4180 15380 4220
rect 17836 4180 17876 4220
rect 19084 4171 19124 4211
rect 22243 4180 22283 4220
rect 22540 4180 22580 4220
rect 22723 4180 22763 4220
rect 22999 4180 23039 4220
rect 23164 4180 23204 4220
rect 23404 4180 23444 4220
rect 23788 4180 23828 4220
rect 11884 4096 11924 4136
rect 12268 4096 12308 4136
rect 12508 4096 12548 4136
rect 13612 4096 13652 4136
rect 15235 4096 15275 4136
rect 15436 4096 15476 4136
rect 17356 4096 17396 4136
rect 23299 4096 23339 4136
rect 23907 4096 23947 4136
rect 24028 4138 24068 4178
rect 24172 4180 24212 4220
rect 24355 4180 24395 4220
rect 24571 4180 24611 4220
rect 24748 4180 24788 4220
rect 27724 4096 27764 4136
rect 33292 4096 33332 4136
rect 33532 4096 33572 4136
rect 38572 4096 38612 4136
rect 40492 4096 40532 4136
rect 40876 4096 40916 4136
rect 41260 4096 41300 4136
rect 42124 4096 42164 4136
rect 44524 4096 44564 4136
rect 44908 4096 44948 4136
rect 13324 4012 13364 4052
rect 22540 4012 22580 4052
rect 24355 4012 24395 4052
rect 40252 4012 40292 4052
rect 40636 4012 40676 4052
rect 41020 4012 41060 4052
rect 44764 4012 44804 4052
rect 13852 3928 13892 3968
rect 23020 3928 23060 3968
rect 24556 3928 24596 3968
rect 27964 3928 28004 3968
rect 38332 3928 38372 3968
rect 42364 3928 42404 3968
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 8956 3592 8996 3632
rect 11548 3592 11588 3632
rect 24076 3592 24116 3632
rect 24892 3592 24932 3632
rect 38716 3592 38756 3632
rect 40540 3592 40580 3632
rect 45148 3592 45188 3632
rect 16204 3508 16244 3548
rect 25852 3508 25892 3548
rect 42364 3508 42404 3548
rect 8716 3424 8756 3464
rect 9388 3424 9428 3464
rect 11788 3424 11828 3464
rect 12556 3424 12596 3464
rect 14755 3424 14795 3464
rect 14956 3424 14996 3464
rect 15820 3424 15860 3464
rect 21244 3424 21284 3464
rect 21484 3424 21524 3464
rect 21868 3424 21908 3464
rect 22636 3424 22676 3464
rect 24748 3424 24788 3464
rect 25132 3424 25172 3464
rect 25612 3424 25652 3464
rect 25987 3424 26027 3464
rect 37852 3424 37892 3464
rect 38092 3424 38132 3464
rect 38476 3424 38516 3464
rect 38956 3424 38996 3464
rect 39436 3424 39476 3464
rect 39724 3424 39764 3464
rect 40012 3424 40052 3464
rect 40300 3424 40340 3464
rect 40876 3424 40916 3464
rect 41356 3424 41396 3464
rect 41740 3424 41780 3464
rect 42124 3424 42164 3464
rect 42508 3424 42548 3464
rect 42892 3424 42932 3464
rect 44524 3424 44564 3464
rect 44908 3424 44948 3464
rect 9772 3340 9812 3380
rect 11020 3340 11060 3380
rect 12067 3340 12107 3380
rect 12172 3340 12212 3380
rect 12652 3340 12692 3380
rect 13132 3340 13172 3380
rect 13620 3340 13660 3380
rect 13987 3340 14027 3380
rect 14284 3340 14324 3380
rect 14615 3340 14655 3380
rect 14860 3340 14900 3380
rect 15244 3340 15284 3380
rect 15427 3340 15467 3380
rect 16396 3340 16436 3380
rect 17604 3340 17644 3380
rect 22126 3340 22166 3380
rect 22252 3340 22292 3380
rect 22732 3340 22772 3380
rect 23212 3340 23252 3380
rect 23700 3340 23740 3380
rect 24076 3340 24116 3380
rect 24191 3340 24231 3380
rect 24364 3340 24404 3380
rect 26188 3340 26228 3380
rect 27436 3340 27476 3380
rect 11212 3256 11252 3296
rect 14188 3256 14228 3296
rect 16060 3256 16100 3296
rect 24508 3256 24548 3296
rect 40636 3256 40676 3296
rect 41980 3256 42020 3296
rect 42748 3256 42788 3296
rect 44764 3256 44804 3296
rect 9628 3172 9668 3212
rect 13804 3172 13844 3212
rect 15340 3172 15380 3212
rect 21628 3172 21668 3212
rect 23884 3172 23924 3212
rect 38236 3172 38276 3212
rect 41596 3172 41636 3212
rect 43132 3172 43172 3212
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 38908 2836 38948 2876
rect 40099 2836 40139 2876
rect 40300 2836 40340 2876
rect 40588 2836 40628 2876
rect 40876 2836 40916 2876
rect 41164 2836 41204 2876
rect 41452 2836 41492 2876
rect 41731 2836 41771 2876
rect 45148 2836 45188 2876
rect 10540 2752 10580 2792
rect 12028 2752 12068 2792
rect 12892 2752 12932 2792
rect 13795 2752 13835 2792
rect 15052 2752 15092 2792
rect 22684 2752 22724 2792
rect 23395 2752 23435 2792
rect 39292 2752 39332 2792
rect 42748 2752 42788 2792
rect 9100 2668 9140 2708
rect 10348 2659 10388 2699
rect 13483 2668 13523 2708
rect 13708 2668 13748 2708
rect 14956 2668 14996 2708
rect 15148 2668 15188 2708
rect 23063 2668 23103 2708
rect 23309 2668 23349 2708
rect 12268 2584 12308 2624
rect 12652 2584 12692 2624
rect 13603 2584 13643 2624
rect 14188 2584 14228 2624
rect 14476 2584 14516 2624
rect 14716 2584 14756 2624
rect 22540 2584 22580 2624
rect 22924 2584 22964 2624
rect 23203 2584 23243 2624
rect 23788 2584 23828 2624
rect 24172 2584 24212 2624
rect 39148 2584 39188 2624
rect 39532 2584 39572 2624
rect 42124 2584 42164 2624
rect 42508 2584 42548 2624
rect 44140 2584 44180 2624
rect 44524 2584 44564 2624
rect 44908 2584 44948 2624
rect 42364 2500 42404 2540
rect 44764 2500 44804 2540
rect 13948 2416 13988 2456
rect 22300 2416 22340 2456
rect 23548 2416 23588 2456
rect 23932 2416 23972 2456
rect 44380 2416 44420 2456
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 1756 2080 1796 2120
rect 45148 2080 45188 2120
rect 1516 1912 1556 1952
rect 3436 1912 3476 1952
rect 5164 1912 5204 1952
rect 6892 1912 6932 1952
rect 8620 1912 8660 1952
rect 43372 1912 43412 1952
rect 43756 1912 43796 1952
rect 44140 1912 44180 1952
rect 44524 1912 44564 1952
rect 44908 1912 44948 1952
rect 43996 1744 44036 1784
rect 3196 1660 3236 1700
rect 4924 1660 4964 1700
rect 6652 1660 6692 1700
rect 8380 1660 8420 1700
rect 43612 1660 43652 1700
rect 44380 1660 44420 1700
rect 44764 1660 44804 1700
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal2 >>
rect 0 11024 90 11044
rect 46278 11024 46368 11044
rect 0 10984 1420 11024
rect 1460 10984 1469 11024
rect 44227 10984 44236 11024
rect 44276 10984 46368 11024
rect 0 10964 90 10984
rect 46278 10964 46368 10984
rect 0 10688 90 10708
rect 46278 10688 46368 10708
rect 0 10648 1132 10688
rect 1172 10648 1181 10688
rect 43747 10648 43756 10688
rect 43796 10648 46368 10688
rect 0 10628 90 10648
rect 46278 10628 46368 10648
rect 0 10352 90 10372
rect 46278 10352 46368 10372
rect 0 10312 1036 10352
rect 1076 10312 1085 10352
rect 43267 10312 43276 10352
rect 43316 10312 46368 10352
rect 0 10292 90 10312
rect 46278 10292 46368 10312
rect 16099 10228 16108 10268
rect 16148 10228 23060 10268
rect 14092 10144 16876 10184
rect 16916 10144 16925 10184
rect 14092 10100 14132 10144
rect 23020 10100 23060 10228
rect 2947 10060 2956 10100
rect 2996 10060 10060 10100
rect 10100 10060 10109 10100
rect 10243 10060 10252 10100
rect 10292 10060 11212 10100
rect 11252 10060 11261 10100
rect 12876 10060 12940 10100
rect 12980 10060 13036 10100
rect 13076 10060 13085 10100
rect 13708 10060 14132 10100
rect 14179 10060 14188 10100
rect 14228 10060 16396 10100
rect 16436 10060 16445 10100
rect 16492 10060 22252 10100
rect 22292 10060 22301 10100
rect 23020 10060 27764 10100
rect 27907 10060 27916 10100
rect 27956 10060 42892 10100
rect 42932 10060 42941 10100
rect 0 10016 90 10036
rect 13708 10016 13748 10060
rect 0 9976 500 10016
rect 1411 9976 1420 10016
rect 1460 9976 2764 10016
rect 2804 9976 2813 10016
rect 9379 9976 9388 10016
rect 9428 9976 13748 10016
rect 13987 9976 13996 10016
rect 14036 9976 16012 10016
rect 16052 9976 16061 10016
rect 0 9956 90 9976
rect 460 9848 500 9976
rect 1123 9892 1132 9932
rect 1172 9892 1748 9932
rect 12451 9892 12460 9932
rect 12500 9892 15916 9932
rect 15956 9892 15965 9932
rect 460 9808 1652 9848
rect 0 9680 90 9700
rect 0 9640 980 9680
rect 0 9620 90 9640
rect 0 9344 90 9364
rect 940 9344 980 9640
rect 1612 9512 1652 9808
rect 1708 9596 1748 9892
rect 16492 9848 16532 10060
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 10051 9808 10060 9848
rect 10100 9808 12652 9848
rect 12692 9808 12701 9848
rect 13612 9808 15052 9848
rect 15092 9808 15101 9848
rect 15331 9808 15340 9848
rect 15380 9808 16532 9848
rect 16780 9976 22828 10016
rect 22868 9976 22877 10016
rect 23395 9976 23404 10016
rect 23444 9976 26956 10016
rect 26996 9976 27005 10016
rect 13612 9764 13652 9808
rect 16780 9764 16820 9976
rect 27724 9932 27764 10060
rect 46278 10016 46368 10036
rect 27811 9976 27820 10016
rect 27860 9976 31468 10016
rect 31508 9976 31517 10016
rect 33571 9976 33580 10016
rect 33620 9976 40492 10016
rect 40532 9976 40541 10016
rect 43852 9976 46368 10016
rect 23587 9892 23596 9932
rect 23636 9892 26284 9932
rect 26324 9892 26333 9932
rect 27724 9892 30068 9932
rect 33379 9892 33388 9932
rect 33428 9892 39244 9932
rect 39284 9892 39293 9932
rect 9484 9724 11308 9764
rect 11348 9724 11357 9764
rect 11404 9724 12844 9764
rect 12884 9724 12893 9764
rect 13516 9724 13652 9764
rect 13708 9724 14900 9764
rect 14947 9724 14956 9764
rect 14996 9724 15628 9764
rect 15668 9724 15677 9764
rect 16012 9724 16820 9764
rect 16876 9808 18548 9848
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 23779 9808 23788 9848
rect 23828 9808 28972 9848
rect 29012 9808 29021 9848
rect 29443 9808 29452 9848
rect 29492 9808 29740 9848
rect 29780 9808 29789 9848
rect 9484 9680 9524 9724
rect 11404 9680 11444 9724
rect 1843 9640 1852 9680
rect 1892 9640 2900 9680
rect 2995 9640 3004 9680
rect 3044 9640 9524 9680
rect 9619 9640 9628 9680
rect 9668 9640 10252 9680
rect 10292 9640 10301 9680
rect 11155 9640 11164 9680
rect 11204 9640 11444 9680
rect 11500 9640 11788 9680
rect 11828 9640 11837 9680
rect 12691 9640 12700 9680
rect 12740 9640 13420 9680
rect 13460 9640 13469 9680
rect 2860 9596 2900 9640
rect 11500 9596 11540 9640
rect 13516 9596 13556 9724
rect 1708 9556 2420 9596
rect 2860 9556 9292 9596
rect 9332 9556 9341 9596
rect 10003 9556 10012 9596
rect 10052 9556 11540 9596
rect 11788 9556 12940 9596
rect 12980 9556 12989 9596
rect 13075 9556 13084 9596
rect 13124 9556 13556 9596
rect 2380 9512 2420 9556
rect 1097 9472 1228 9512
rect 1268 9472 1277 9512
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 1987 9472 1996 9512
rect 2036 9472 2045 9512
rect 2371 9472 2380 9512
rect 2420 9472 2429 9512
rect 2633 9472 2764 9512
rect 2804 9472 2813 9512
rect 2860 9472 3148 9512
rect 3188 9472 3197 9512
rect 9257 9472 9388 9512
rect 9428 9472 9437 9512
rect 9763 9472 9772 9512
rect 9812 9472 9821 9512
rect 10025 9472 10156 9512
rect 10196 9472 10205 9512
rect 10387 9472 10396 9512
rect 10436 9472 10484 9512
rect 10531 9472 10540 9512
rect 10580 9472 10711 9512
rect 10793 9472 10924 9512
rect 10964 9472 10973 9512
rect 11299 9472 11308 9512
rect 11348 9472 11357 9512
rect 11561 9472 11692 9512
rect 11732 9472 11741 9512
rect 1996 9428 2036 9472
rect 2860 9428 2900 9472
rect 9772 9428 9812 9472
rect 1027 9388 1036 9428
rect 1076 9388 2036 9428
rect 2092 9388 2900 9428
rect 4099 9388 4108 9428
rect 4148 9388 9812 9428
rect 10444 9428 10484 9472
rect 11308 9428 11348 9472
rect 10444 9388 10828 9428
rect 10868 9388 10877 9428
rect 11308 9388 11500 9428
rect 11540 9388 11549 9428
rect 2092 9344 2132 9388
rect 11788 9344 11828 9556
rect 13708 9512 13748 9724
rect 14860 9680 14900 9724
rect 16012 9680 16052 9724
rect 16876 9680 16916 9808
rect 18508 9764 18548 9808
rect 13843 9640 13852 9680
rect 13892 9640 13996 9680
rect 14036 9640 14045 9680
rect 14860 9640 16052 9680
rect 16147 9640 16156 9680
rect 16196 9640 16300 9680
rect 16340 9640 16349 9680
rect 16786 9640 16916 9680
rect 17020 9724 17932 9764
rect 17972 9724 17981 9764
rect 18403 9724 18412 9764
rect 18452 9724 18461 9764
rect 18508 9724 22060 9764
rect 22100 9724 22109 9764
rect 22252 9724 23116 9764
rect 23156 9724 23165 9764
rect 24748 9724 25132 9764
rect 25172 9724 25181 9764
rect 25411 9724 25420 9764
rect 25460 9724 25652 9764
rect 25795 9724 25804 9764
rect 25844 9724 26900 9764
rect 28867 9724 28876 9764
rect 28916 9724 29932 9764
rect 29972 9724 29981 9764
rect 16786 9596 16826 9640
rect 17020 9596 17060 9724
rect 18412 9680 18452 9724
rect 22252 9680 22292 9724
rect 24748 9680 24788 9724
rect 17299 9640 17308 9680
rect 17348 9640 17452 9680
rect 17492 9640 17501 9680
rect 17683 9640 17692 9680
rect 17732 9640 18316 9680
rect 18356 9640 18365 9680
rect 18412 9640 18460 9680
rect 18500 9640 18509 9680
rect 18835 9640 18844 9680
rect 18884 9640 19468 9680
rect 19508 9640 19517 9680
rect 19603 9640 19612 9680
rect 19652 9640 20236 9680
rect 20276 9640 20285 9680
rect 20524 9640 21196 9680
rect 21236 9640 21245 9680
rect 21523 9640 21532 9680
rect 21572 9640 22292 9680
rect 22675 9640 22684 9680
rect 22724 9640 24788 9680
rect 24835 9640 24844 9680
rect 24884 9640 25556 9680
rect 13795 9556 13804 9596
rect 13844 9556 14804 9596
rect 14764 9512 14804 9556
rect 16300 9556 16826 9596
rect 16972 9556 17060 9596
rect 18067 9556 18076 9596
rect 18116 9556 18604 9596
rect 18644 9556 18653 9596
rect 19219 9556 19228 9596
rect 19268 9556 19852 9596
rect 19892 9556 19901 9596
rect 16300 9512 16340 9556
rect 16972 9512 17012 9556
rect 20524 9512 20564 9640
rect 21100 9556 21388 9596
rect 21428 9556 21437 9596
rect 21763 9556 21772 9596
rect 21812 9556 21821 9596
rect 22147 9556 22156 9596
rect 22196 9556 22205 9596
rect 22252 9556 22348 9596
rect 22388 9556 22397 9596
rect 23020 9556 23500 9596
rect 23540 9556 23549 9596
rect 23683 9556 23692 9596
rect 23732 9556 23741 9596
rect 23875 9556 23884 9596
rect 23924 9556 23933 9596
rect 24451 9556 24460 9596
rect 24500 9556 24509 9596
rect 24643 9556 24652 9596
rect 24692 9556 25364 9596
rect 21100 9512 21140 9556
rect 21772 9512 21812 9556
rect 22156 9512 22196 9556
rect 22252 9512 22292 9556
rect 23020 9512 23060 9556
rect 23692 9512 23732 9556
rect 23884 9512 23924 9556
rect 24460 9512 24500 9556
rect 25324 9512 25364 9556
rect 25516 9512 25556 9640
rect 25612 9596 25652 9724
rect 26275 9640 26284 9680
rect 26324 9640 26620 9680
rect 26660 9640 26669 9680
rect 25612 9556 26516 9596
rect 26476 9512 26516 9556
rect 26860 9512 26900 9724
rect 30028 9680 30068 9892
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 34348 9808 37364 9848
rect 37411 9808 37420 9848
rect 37460 9808 41644 9848
rect 41684 9808 41693 9848
rect 31939 9724 31948 9764
rect 31988 9724 32372 9764
rect 32707 9724 32716 9764
rect 32756 9724 33524 9764
rect 32332 9680 32372 9724
rect 33484 9680 33524 9724
rect 28483 9640 28492 9680
rect 28532 9640 29204 9680
rect 30028 9640 30076 9680
rect 30116 9640 30125 9680
rect 31171 9640 31180 9680
rect 31220 9640 31228 9680
rect 31268 9640 31351 9680
rect 31555 9640 31564 9680
rect 31604 9640 31996 9680
rect 32036 9640 32045 9680
rect 32332 9640 32764 9680
rect 32804 9640 32813 9680
rect 33484 9640 33532 9680
rect 33572 9640 33581 9680
rect 28291 9556 28300 9596
rect 28340 9556 28820 9596
rect 28915 9556 28924 9596
rect 28964 9556 28972 9596
rect 29012 9556 29095 9596
rect 28780 9512 28820 9556
rect 29164 9512 29204 9640
rect 29251 9556 29260 9596
rect 29300 9556 30356 9596
rect 31363 9556 31372 9596
rect 31412 9556 31612 9596
rect 31652 9556 31661 9596
rect 31747 9556 31756 9596
rect 31796 9556 32380 9596
rect 32420 9556 32429 9596
rect 33091 9556 33100 9596
rect 33140 9556 33428 9596
rect 30316 9512 30356 9556
rect 33388 9512 33428 9556
rect 34348 9512 34388 9808
rect 37324 9764 37364 9808
rect 37324 9724 40588 9764
rect 40628 9724 40637 9764
rect 42988 9724 43756 9764
rect 43796 9724 43805 9764
rect 42988 9680 43028 9724
rect 43852 9680 43892 9976
rect 46278 9956 46368 9976
rect 46278 9680 46368 9700
rect 35395 9640 35404 9680
rect 35444 9640 35452 9680
rect 35492 9640 35575 9680
rect 36163 9640 36172 9680
rect 36212 9640 36220 9680
rect 36260 9640 36343 9680
rect 36451 9640 36460 9680
rect 36500 9640 40780 9680
rect 40820 9640 40829 9680
rect 42835 9640 42844 9680
rect 42884 9640 43028 9680
rect 43219 9640 43228 9680
rect 43268 9640 43276 9680
rect 43316 9640 43399 9680
rect 43603 9640 43612 9680
rect 43652 9640 43892 9680
rect 43987 9640 43996 9680
rect 44036 9640 46368 9680
rect 46278 9620 46368 9640
rect 34819 9556 34828 9596
rect 34868 9556 35836 9596
rect 35876 9556 35885 9596
rect 36355 9556 36364 9596
rect 36404 9556 43028 9596
rect 42988 9512 43028 9556
rect 11945 9472 12076 9512
rect 12116 9472 12125 9512
rect 12451 9472 12460 9512
rect 12500 9472 12509 9512
rect 12713 9472 12844 9512
rect 12884 9472 12893 9512
rect 13097 9472 13228 9512
rect 13268 9472 13277 9512
rect 13459 9472 13468 9512
rect 13508 9472 13556 9512
rect 13603 9472 13612 9512
rect 13652 9472 13748 9512
rect 13987 9472 13996 9512
rect 14036 9472 14167 9512
rect 14249 9472 14380 9512
rect 14420 9472 14429 9512
rect 14755 9472 14764 9512
rect 14804 9472 14813 9512
rect 14995 9472 15004 9512
rect 15044 9472 15092 9512
rect 15139 9472 15148 9512
rect 15188 9472 15319 9512
rect 15401 9472 15532 9512
rect 15572 9472 15581 9512
rect 15785 9472 15916 9512
rect 15956 9472 15965 9512
rect 16291 9472 16300 9512
rect 16340 9472 16349 9512
rect 16553 9472 16684 9512
rect 16724 9472 16733 9512
rect 16915 9472 16924 9512
rect 16964 9472 17012 9512
rect 17059 9472 17068 9512
rect 17108 9472 17117 9512
rect 17321 9472 17452 9512
rect 17492 9472 17501 9512
rect 17705 9472 17836 9512
rect 17876 9472 17885 9512
rect 18211 9472 18220 9512
rect 18260 9472 18412 9512
rect 18452 9472 18461 9512
rect 18595 9472 18604 9512
rect 18644 9472 18796 9512
rect 18836 9472 18845 9512
rect 18979 9472 18988 9512
rect 19028 9472 19037 9512
rect 19241 9472 19372 9512
rect 19412 9472 19421 9512
rect 19625 9472 19756 9512
rect 19796 9472 19805 9512
rect 20515 9472 20524 9512
rect 20564 9472 20573 9512
rect 20707 9472 20716 9512
rect 20756 9472 20764 9512
rect 20804 9472 20887 9512
rect 21091 9472 21100 9512
rect 21140 9472 21149 9512
rect 21283 9472 21292 9512
rect 21332 9472 21812 9512
rect 21859 9472 21868 9512
rect 21908 9472 22196 9512
rect 22243 9472 22252 9512
rect 22292 9472 22301 9512
rect 22435 9472 22444 9512
rect 22484 9472 22540 9512
rect 22580 9472 22615 9512
rect 23011 9472 23020 9512
rect 23060 9472 23069 9512
rect 23395 9472 23404 9512
rect 23444 9472 23732 9512
rect 23779 9472 23788 9512
rect 23828 9472 23924 9512
rect 23971 9472 23980 9512
rect 24020 9472 24076 9512
rect 24116 9472 24151 9512
rect 24233 9472 24268 9512
rect 24308 9472 24364 9512
rect 24404 9472 24413 9512
rect 24460 9472 24940 9512
rect 24980 9472 24989 9512
rect 25315 9472 25324 9512
rect 25364 9472 25373 9512
rect 25507 9472 25516 9512
rect 25556 9472 25565 9512
rect 25699 9472 25708 9512
rect 25748 9472 25852 9512
rect 25892 9472 25901 9512
rect 26083 9472 26092 9512
rect 26132 9472 26141 9512
rect 26467 9472 26476 9512
rect 26516 9472 26525 9512
rect 26851 9472 26860 9512
rect 26900 9472 26909 9512
rect 27235 9472 27244 9512
rect 27284 9472 27293 9512
rect 28099 9472 28108 9512
rect 28148 9472 28396 9512
rect 28436 9472 28445 9512
rect 28492 9472 28540 9512
rect 28580 9472 28589 9512
rect 28771 9472 28780 9512
rect 28820 9472 28829 9512
rect 29155 9472 29164 9512
rect 29204 9472 29213 9512
rect 29347 9472 29356 9512
rect 29396 9472 29405 9512
rect 29452 9472 29692 9512
rect 29732 9472 29741 9512
rect 29923 9472 29932 9512
rect 29972 9472 30103 9512
rect 30307 9472 30316 9512
rect 30356 9472 30365 9512
rect 30691 9472 30700 9512
rect 30740 9472 30749 9512
rect 31459 9472 31468 9512
rect 31508 9472 31796 9512
rect 31843 9472 31852 9512
rect 31892 9472 31901 9512
rect 32227 9472 32236 9512
rect 32276 9472 32285 9512
rect 32611 9472 32620 9512
rect 32660 9472 32716 9512
rect 32756 9472 32791 9512
rect 32873 9472 33004 9512
rect 33044 9472 33053 9512
rect 33379 9472 33388 9512
rect 33428 9472 33437 9512
rect 33571 9472 33580 9512
rect 33620 9472 33772 9512
rect 33812 9472 33821 9512
rect 34147 9472 34156 9512
rect 34196 9472 34205 9512
rect 34348 9472 34483 9512
rect 34523 9472 34532 9512
rect 34627 9472 34636 9512
rect 34676 9472 34684 9512
rect 34724 9472 34807 9512
rect 34963 9472 34972 9512
rect 35012 9472 35020 9512
rect 35060 9472 35143 9512
rect 35299 9472 35308 9512
rect 35348 9472 35636 9512
rect 35683 9472 35692 9512
rect 35732 9472 35863 9512
rect 35932 9472 36076 9512
rect 36116 9472 36125 9512
rect 36259 9472 36268 9512
rect 36308 9472 36460 9512
rect 36500 9472 36509 9512
rect 37708 9472 40012 9512
rect 40052 9472 40061 9512
rect 41705 9472 41836 9512
rect 41876 9472 41885 9512
rect 42019 9472 42028 9512
rect 42068 9472 42220 9512
rect 42260 9472 42269 9512
rect 42316 9472 42604 9512
rect 42644 9472 42653 9512
rect 42979 9472 42988 9512
rect 43028 9472 43037 9512
rect 43241 9472 43276 9512
rect 43316 9472 43372 9512
rect 43412 9472 43421 9512
rect 43625 9472 43660 9512
rect 43700 9472 43756 9512
rect 43796 9472 43805 9512
rect 44009 9472 44140 9512
rect 44180 9472 44189 9512
rect 44899 9472 44908 9512
rect 44948 9472 44957 9512
rect 12460 9428 12500 9472
rect 13516 9428 13556 9472
rect 15052 9428 15092 9472
rect 17068 9428 17108 9472
rect 18988 9428 19028 9472
rect 26092 9428 26132 9472
rect 27244 9428 27284 9472
rect 28492 9428 28532 9472
rect 29356 9428 29396 9472
rect 12460 9388 13420 9428
rect 13460 9388 13469 9428
rect 13516 9388 14956 9428
rect 14996 9388 15005 9428
rect 15052 9388 16780 9428
rect 16820 9388 16829 9428
rect 17068 9388 17260 9428
rect 17300 9388 17309 9428
rect 18115 9388 18124 9428
rect 18164 9388 19028 9428
rect 19075 9388 19084 9428
rect 19124 9388 21140 9428
rect 21859 9388 21868 9428
rect 21908 9388 24788 9428
rect 25027 9388 25036 9428
rect 25076 9388 26132 9428
rect 26179 9388 26188 9428
rect 26228 9388 27284 9428
rect 27331 9388 27340 9428
rect 27380 9388 28532 9428
rect 28675 9388 28684 9428
rect 28724 9388 29396 9428
rect 21100 9344 21140 9388
rect 24748 9344 24788 9388
rect 29452 9344 29492 9472
rect 30700 9428 30740 9472
rect 31756 9428 31796 9472
rect 29731 9388 29740 9428
rect 29780 9388 30740 9428
rect 31747 9388 31756 9428
rect 31796 9388 31805 9428
rect 0 9304 212 9344
rect 940 9304 2132 9344
rect 2227 9304 2236 9344
rect 2276 9304 3284 9344
rect 3379 9304 3388 9344
rect 3428 9304 10676 9344
rect 11539 9304 11548 9344
rect 11588 9304 11828 9344
rect 11923 9304 11932 9344
rect 11972 9304 13708 9344
rect 13748 9304 13757 9344
rect 14179 9304 14188 9344
rect 14228 9304 14236 9344
rect 14276 9304 14359 9344
rect 14611 9304 14620 9344
rect 14660 9304 16396 9344
rect 16436 9304 16445 9344
rect 16531 9304 16540 9344
rect 16580 9304 17740 9344
rect 17780 9304 17789 9344
rect 17923 9304 17932 9344
rect 17972 9304 19852 9344
rect 19892 9304 19901 9344
rect 19987 9304 19996 9344
rect 20036 9304 20620 9344
rect 20660 9304 20669 9344
rect 20851 9304 20860 9344
rect 20900 9304 20908 9344
rect 20948 9304 21031 9344
rect 21100 9304 22012 9344
rect 22052 9304 22061 9344
rect 22339 9304 22348 9344
rect 22388 9304 23548 9344
rect 23588 9304 23597 9344
rect 24211 9304 24220 9344
rect 24260 9304 24364 9344
rect 24404 9304 24413 9344
rect 24521 9304 24604 9344
rect 24644 9304 24652 9344
rect 24692 9304 24701 9344
rect 24748 9304 25084 9344
rect 25124 9304 25133 9344
rect 25747 9304 25756 9344
rect 25796 9304 25900 9344
rect 25940 9304 25949 9344
rect 27907 9304 27916 9344
rect 27956 9304 29492 9344
rect 29587 9304 29596 9344
rect 29636 9304 30028 9344
rect 30068 9304 30077 9344
rect 30124 9304 30892 9344
rect 30932 9304 30941 9344
rect 0 9284 90 9304
rect 172 9092 212 9304
rect 3244 9260 3284 9304
rect 1459 9220 1468 9260
rect 1508 9220 1748 9260
rect 1891 9220 1900 9260
rect 1940 9220 2228 9260
rect 2611 9220 2620 9260
rect 2660 9220 2764 9260
rect 2804 9220 2813 9260
rect 3244 9220 8852 9260
rect 1708 9176 1748 9220
rect 2188 9176 2228 9220
rect 1708 9136 2092 9176
rect 2132 9136 2141 9176
rect 2188 9136 8716 9176
rect 8756 9136 8765 9176
rect 8812 9092 8852 9220
rect 10636 9176 10676 9304
rect 30124 9260 30164 9304
rect 10771 9220 10780 9260
rect 10820 9220 11308 9260
rect 11348 9220 11357 9260
rect 11875 9220 11884 9260
rect 11924 9220 12172 9260
rect 12212 9220 12221 9260
rect 12307 9220 12316 9260
rect 12356 9220 12596 9260
rect 13411 9220 13420 9260
rect 13460 9220 14572 9260
rect 14612 9220 14621 9260
rect 15379 9220 15388 9260
rect 15428 9220 15668 9260
rect 15763 9220 15772 9260
rect 15812 9220 17356 9260
rect 17396 9220 17405 9260
rect 18211 9220 18220 9260
rect 18260 9220 19084 9260
rect 19124 9220 19133 9260
rect 20323 9220 20332 9260
rect 20372 9220 21004 9260
rect 21044 9220 21053 9260
rect 21619 9220 21628 9260
rect 21668 9220 21676 9260
rect 21716 9220 21799 9260
rect 22649 9220 22732 9260
rect 22772 9220 22780 9260
rect 22820 9220 22829 9260
rect 23020 9220 23164 9260
rect 23204 9220 23213 9260
rect 23404 9220 24700 9260
rect 24740 9220 24749 9260
rect 24835 9220 24844 9260
rect 24884 9220 26236 9260
rect 26276 9220 26285 9260
rect 26467 9220 26476 9260
rect 26516 9220 27004 9260
rect 27044 9220 27053 9260
rect 27715 9220 27724 9260
rect 27764 9220 28156 9260
rect 28196 9220 28205 9260
rect 29068 9220 30164 9260
rect 30220 9220 30460 9260
rect 30500 9220 30509 9260
rect 12556 9176 12596 9220
rect 15628 9176 15668 9220
rect 23020 9176 23060 9220
rect 10636 9136 11788 9176
rect 11828 9136 11837 9176
rect 12556 9136 12788 9176
rect 12748 9092 12788 9136
rect 12940 9136 14092 9176
rect 14132 9136 14141 9176
rect 14755 9136 14764 9176
rect 14804 9136 15340 9176
rect 15380 9136 15389 9176
rect 15628 9136 17164 9176
rect 17204 9136 17213 9176
rect 17731 9136 17740 9176
rect 17780 9136 19852 9176
rect 19892 9136 19901 9176
rect 19948 9136 20660 9176
rect 21283 9136 21292 9176
rect 21332 9136 23060 9176
rect 12940 9092 12980 9136
rect 19948 9092 19988 9136
rect 172 9052 2380 9092
rect 2420 9052 2429 9092
rect 2860 9052 4780 9092
rect 4820 9052 4829 9092
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 8812 9052 12268 9092
rect 12308 9052 12317 9092
rect 12748 9052 12980 9092
rect 14179 9052 14188 9092
rect 14228 9052 19988 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 0 9008 90 9028
rect 0 8968 1228 9008
rect 1268 8968 1277 9008
rect 0 8948 90 8968
rect 2860 8924 2900 9052
rect 20620 9008 20660 9136
rect 23404 9092 23444 9220
rect 29068 9176 29108 9220
rect 30220 9176 30260 9220
rect 23491 9136 23500 9176
rect 23540 9136 25804 9176
rect 25844 9136 25853 9176
rect 26851 9136 26860 9176
rect 26900 9136 29108 9176
rect 29155 9136 29164 9176
rect 29204 9136 30260 9176
rect 31852 9092 31892 9472
rect 32236 9428 32276 9472
rect 34156 9428 34196 9472
rect 35596 9428 35636 9472
rect 35932 9428 35972 9472
rect 37708 9428 37748 9472
rect 32236 9388 34060 9428
rect 34100 9388 34109 9428
rect 34156 9388 35404 9428
rect 35444 9388 35453 9428
rect 35587 9388 35596 9428
rect 35636 9388 35645 9428
rect 35779 9388 35788 9428
rect 35828 9388 35972 9428
rect 36163 9388 36172 9428
rect 36212 9388 37748 9428
rect 37891 9388 37900 9428
rect 37940 9388 42220 9428
rect 42260 9388 42269 9428
rect 42316 9344 42356 9472
rect 44908 9428 44948 9472
rect 43171 9388 43180 9428
rect 43220 9388 43468 9428
rect 43508 9388 44620 9428
rect 44660 9388 44948 9428
rect 46278 9344 46368 9364
rect 32323 9304 32332 9344
rect 32372 9304 33148 9344
rect 33188 9304 33197 9344
rect 33475 9304 33484 9344
rect 33524 9304 34484 9344
rect 34531 9304 34540 9344
rect 34580 9304 35068 9344
rect 35108 9304 35117 9344
rect 37411 9304 37420 9344
rect 37460 9304 42356 9344
rect 42451 9304 42460 9344
rect 42500 9304 44236 9344
rect 44276 9304 44285 9344
rect 44371 9304 44380 9344
rect 44420 9304 46368 9344
rect 34444 9260 34484 9304
rect 46278 9284 46368 9304
rect 33187 9220 33196 9260
rect 33236 9220 33916 9260
rect 33956 9220 33965 9260
rect 34169 9220 34252 9260
rect 34292 9220 34300 9260
rect 34340 9220 34349 9260
rect 34444 9220 35500 9260
rect 35540 9220 35549 9260
rect 35596 9220 36364 9260
rect 36404 9220 36413 9260
rect 40474 9220 40483 9260
rect 40523 9220 40675 9260
rect 40724 9220 40963 9260
rect 41003 9220 41251 9260
rect 41291 9220 41539 9260
rect 41579 9220 41740 9260
rect 41780 9220 41789 9260
rect 42067 9220 42076 9260
rect 42116 9220 42644 9260
rect 45139 9220 45148 9260
rect 45188 9220 45868 9260
rect 45908 9220 45917 9260
rect 35596 9176 35636 9220
rect 42604 9176 42644 9220
rect 20707 9052 20716 9092
rect 20756 9052 21484 9092
rect 21524 9052 21533 9092
rect 21763 9052 21772 9092
rect 21812 9052 23444 9092
rect 26179 9052 26188 9092
rect 26228 9052 31892 9092
rect 32332 9136 35636 9176
rect 35971 9136 35980 9176
rect 36020 9136 41164 9176
rect 41204 9136 41213 9176
rect 42604 9136 44804 9176
rect 32332 9008 32372 9136
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 38851 9052 38860 9092
rect 38900 9052 43700 9092
rect 3331 8968 3340 9008
rect 3380 8968 10060 9008
rect 10100 8968 10109 9008
rect 10636 8968 11020 9008
rect 11060 8968 11069 9008
rect 11875 8968 11884 9008
rect 11924 8968 12556 9008
rect 12596 8968 12605 9008
rect 12988 8968 13516 9008
rect 13556 8968 13565 9008
rect 13891 8968 13900 9008
rect 13940 8968 13949 9008
rect 16108 8968 16972 9008
rect 17012 8968 17021 9008
rect 17155 8968 17164 9008
rect 17204 8968 20276 9008
rect 20620 8968 20948 9008
rect 27331 8968 27340 9008
rect 27380 8968 32372 9008
rect 32428 8968 33484 9008
rect 33524 8968 33533 9008
rect 38947 8968 38956 9008
rect 38996 8968 43316 9008
rect 10636 8924 10676 8968
rect 12988 8924 13028 8968
rect 13900 8924 13940 8968
rect 16108 8924 16148 8968
rect 1459 8884 1468 8924
rect 1508 8884 2900 8924
rect 3187 8884 3196 8924
rect 3236 8884 10156 8924
rect 10196 8884 10205 8924
rect 10291 8884 10300 8924
rect 10340 8884 10676 8924
rect 11059 8884 11068 8924
rect 11108 8884 11980 8924
rect 12020 8884 12029 8924
rect 12076 8884 12364 8924
rect 12404 8884 12413 8924
rect 12595 8884 12604 8924
rect 12644 8884 13028 8924
rect 13324 8884 13940 8924
rect 14131 8884 14140 8924
rect 14180 8884 14956 8924
rect 14996 8884 15005 8924
rect 15139 8884 15148 8924
rect 15188 8884 15319 8924
rect 15859 8884 15868 8924
rect 15908 8884 16148 8924
rect 16243 8884 16252 8924
rect 16292 8884 18260 8924
rect 18377 8884 18460 8924
rect 18500 8884 18508 8924
rect 18548 8884 18557 8924
rect 18691 8884 18700 8924
rect 18740 8884 18844 8924
rect 18884 8884 18893 8924
rect 19145 8884 19228 8924
rect 19268 8884 19276 8924
rect 19316 8884 19325 8924
rect 19529 8884 19612 8924
rect 19652 8884 19660 8924
rect 19700 8884 19709 8924
rect 19939 8884 19948 8924
rect 19988 8884 19996 8924
rect 20036 8884 20119 8924
rect 12076 8840 12116 8884
rect 13324 8840 13364 8884
rect 18220 8840 18260 8884
rect 20236 8840 20276 8968
rect 20371 8884 20380 8924
rect 20420 8884 20524 8924
rect 20564 8884 20573 8924
rect 20681 8884 20764 8924
rect 20804 8884 20812 8924
rect 20852 8884 20861 8924
rect 20908 8840 20948 8968
rect 21427 8884 21436 8924
rect 21476 8884 23732 8924
rect 1769 8800 1852 8840
rect 1892 8800 1900 8840
rect 1940 8800 1949 8840
rect 3571 8800 3580 8840
rect 3620 8800 11116 8840
rect 11156 8800 11165 8840
rect 11443 8800 11452 8840
rect 11492 8800 12116 8840
rect 12172 8800 12220 8840
rect 12260 8800 12269 8840
rect 12979 8800 12988 8840
rect 13028 8800 13364 8840
rect 13411 8800 13420 8840
rect 13460 8800 17980 8840
rect 18020 8800 18029 8840
rect 18220 8800 19604 8840
rect 20236 8800 20756 8840
rect 20908 8800 23164 8840
rect 23204 8800 23213 8840
rect 12172 8756 12212 8800
rect 556 8716 2036 8756
rect 0 8672 90 8692
rect 556 8672 596 8716
rect 1996 8672 2036 8716
rect 2860 8716 10156 8756
rect 10196 8716 10205 8756
rect 10444 8716 11020 8756
rect 11060 8716 11069 8756
rect 11308 8716 11596 8756
rect 11636 8716 11645 8756
rect 11971 8716 11980 8756
rect 12020 8716 12212 8756
rect 13756 8716 14092 8756
rect 14132 8716 14141 8756
rect 14659 8716 14668 8756
rect 14708 8716 14717 8756
rect 14921 8716 15052 8756
rect 15092 8716 15101 8756
rect 15226 8716 15235 8756
rect 15275 8716 15628 8756
rect 15668 8716 15677 8756
rect 15916 8716 16204 8756
rect 16244 8716 16253 8756
rect 16387 8716 16396 8756
rect 16436 8716 17644 8756
rect 17684 8716 17693 8756
rect 17827 8716 17836 8756
rect 17876 8716 18604 8756
rect 18644 8716 18653 8756
rect 2860 8672 2900 8716
rect 10444 8672 10484 8716
rect 0 8632 596 8672
rect 643 8632 652 8672
rect 692 8632 1228 8672
rect 1268 8632 1277 8672
rect 1603 8632 1612 8672
rect 1652 8632 1661 8672
rect 1987 8632 1996 8672
rect 2036 8632 2045 8672
rect 2249 8632 2380 8672
rect 2420 8632 2429 8672
rect 2611 8632 2620 8672
rect 2660 8632 2900 8672
rect 2947 8632 2956 8672
rect 2996 8632 3127 8672
rect 3209 8632 3340 8672
rect 3380 8632 3389 8672
rect 3436 8632 9388 8672
rect 9428 8632 9437 8672
rect 10051 8632 10060 8672
rect 10100 8632 10252 8672
rect 10292 8632 10301 8672
rect 10435 8632 10444 8672
rect 10484 8632 10493 8672
rect 10697 8632 10828 8672
rect 10868 8632 10877 8672
rect 11081 8632 11212 8672
rect 11252 8632 11261 8672
rect 0 8612 90 8632
rect 0 8336 90 8356
rect 1612 8336 1652 8632
rect 3436 8588 3476 8632
rect 11308 8588 11348 8716
rect 13756 8672 13796 8716
rect 14668 8672 14708 8716
rect 15244 8672 15284 8716
rect 11587 8632 11596 8672
rect 11636 8632 11645 8672
rect 11971 8632 11980 8672
rect 12020 8632 12308 8672
rect 12355 8632 12364 8672
rect 12404 8632 12535 8672
rect 12739 8632 12748 8672
rect 12788 8632 12844 8672
rect 12884 8632 12919 8672
rect 13123 8632 13132 8672
rect 13172 8632 13181 8672
rect 13507 8632 13516 8672
rect 13556 8632 13687 8672
rect 13747 8632 13756 8672
rect 13796 8632 13805 8672
rect 13891 8632 13900 8672
rect 13940 8632 13949 8672
rect 14153 8632 14188 8672
rect 14228 8632 14284 8672
rect 14324 8632 14333 8672
rect 14515 8632 14524 8672
rect 14564 8632 14612 8672
rect 14659 8632 14668 8672
rect 14708 8632 14755 8672
rect 15235 8632 15244 8672
rect 15284 8632 15360 8672
rect 15619 8632 15628 8672
rect 15668 8632 15724 8672
rect 15764 8632 15799 8672
rect 2227 8548 2236 8588
rect 2276 8548 3476 8588
rect 10675 8548 10684 8588
rect 10724 8548 11348 8588
rect 11596 8588 11636 8632
rect 12268 8588 12308 8632
rect 13132 8588 13172 8632
rect 13900 8588 13940 8632
rect 14572 8588 14612 8632
rect 15916 8588 15956 8716
rect 19564 8672 19604 8800
rect 20236 8716 20620 8756
rect 20660 8716 20669 8756
rect 20236 8672 20276 8716
rect 20716 8672 20756 8800
rect 21955 8716 21964 8756
rect 22004 8716 22013 8756
rect 22243 8716 22252 8756
rect 22292 8716 22772 8756
rect 22819 8716 22828 8756
rect 22868 8716 22964 8756
rect 21964 8672 22004 8716
rect 22732 8672 22772 8716
rect 16003 8632 16012 8672
rect 16052 8632 16183 8672
rect 16291 8632 16300 8672
rect 16340 8632 16396 8672
rect 16436 8632 16492 8672
rect 16532 8632 16541 8672
rect 16627 8632 16636 8672
rect 16676 8632 17068 8672
rect 17108 8632 17117 8672
rect 17251 8632 17260 8672
rect 17300 8632 17309 8672
rect 17539 8632 17548 8672
rect 17588 8632 18220 8672
rect 18260 8632 18269 8672
rect 18569 8632 18700 8672
rect 18740 8632 18749 8672
rect 18953 8632 19084 8672
rect 19124 8632 19133 8672
rect 19337 8632 19468 8672
rect 19508 8632 19517 8672
rect 19564 8632 19852 8672
rect 19892 8632 19901 8672
rect 20227 8632 20236 8672
rect 20276 8632 20285 8672
rect 20611 8632 20620 8672
rect 20660 8632 20756 8672
rect 20873 8632 21004 8672
rect 21044 8632 21053 8672
rect 21187 8632 21196 8672
rect 21236 8632 21367 8672
rect 21571 8632 21580 8672
rect 21620 8632 21868 8672
rect 21908 8632 21917 8672
rect 21964 8632 22060 8672
rect 22100 8632 22109 8672
rect 22291 8632 22300 8672
rect 22340 8632 22636 8672
rect 22676 8632 22685 8672
rect 22732 8632 22780 8672
rect 22820 8632 22829 8672
rect 17260 8588 17300 8632
rect 22924 8588 22964 8716
rect 23020 8716 23500 8756
rect 23540 8716 23549 8756
rect 23020 8672 23060 8716
rect 23011 8632 23020 8672
rect 23060 8632 23069 8672
rect 23273 8632 23404 8672
rect 23444 8632 23453 8672
rect 23500 8632 23548 8672
rect 23588 8632 23597 8672
rect 23500 8588 23540 8632
rect 11596 8548 12020 8588
rect 12268 8548 12940 8588
rect 12980 8548 12989 8588
rect 13123 8548 13132 8588
rect 13172 8548 13219 8588
rect 13363 8548 13372 8588
rect 13412 8548 13612 8588
rect 13652 8548 13661 8588
rect 13891 8548 13900 8588
rect 13940 8548 13987 8588
rect 14572 8548 14764 8588
rect 14804 8548 14813 8588
rect 14899 8548 14908 8588
rect 14948 8548 15956 8588
rect 16867 8548 16876 8588
rect 16916 8548 17020 8588
rect 17060 8548 17069 8588
rect 17155 8548 17164 8588
rect 17204 8548 21628 8588
rect 21668 8548 21677 8588
rect 22924 8548 23540 8588
rect 23692 8588 23732 8884
rect 23788 8884 26764 8924
rect 26804 8884 26813 8924
rect 26947 8884 26956 8924
rect 26996 8884 29596 8924
rect 29636 8884 29645 8924
rect 32131 8884 32140 8924
rect 32180 8884 32188 8924
rect 32228 8884 32311 8924
rect 23788 8672 23828 8884
rect 24451 8800 24460 8840
rect 24500 8800 25276 8840
rect 25316 8800 25325 8840
rect 25420 8800 25748 8840
rect 25939 8800 25948 8840
rect 25988 8800 28396 8840
rect 28436 8800 28780 8840
rect 28820 8800 28829 8840
rect 25420 8756 25460 8800
rect 25708 8756 25748 8800
rect 23884 8716 25460 8756
rect 25603 8716 25612 8756
rect 25652 8716 25661 8756
rect 25708 8716 26188 8756
rect 26228 8716 26237 8756
rect 26371 8716 26380 8756
rect 26420 8716 26429 8756
rect 26563 8716 26572 8756
rect 26612 8716 29356 8756
rect 29396 8716 29405 8756
rect 23779 8632 23788 8672
rect 23828 8632 23837 8672
rect 23884 8588 23924 8716
rect 25612 8672 25652 8716
rect 26380 8672 26420 8716
rect 32428 8672 32468 8968
rect 32515 8884 32524 8924
rect 32564 8884 32572 8924
rect 32612 8884 32695 8924
rect 32899 8884 32908 8924
rect 32948 8884 32956 8924
rect 32996 8884 33079 8924
rect 33283 8884 33292 8924
rect 33332 8884 33340 8924
rect 33380 8884 33463 8924
rect 33667 8884 33676 8924
rect 33716 8884 33724 8924
rect 33764 8884 33847 8924
rect 34099 8884 34108 8924
rect 34148 8884 34348 8924
rect 34388 8884 34397 8924
rect 35657 8884 35740 8924
rect 35780 8884 35788 8924
rect 35828 8884 35837 8924
rect 37315 8884 37324 8924
rect 37364 8884 43036 8924
rect 43076 8884 43085 8924
rect 34435 8800 34444 8840
rect 34484 8800 34492 8840
rect 34532 8800 34615 8840
rect 35347 8800 35356 8840
rect 35396 8800 35692 8840
rect 35732 8800 35741 8840
rect 37795 8800 37804 8840
rect 37844 8800 38092 8840
rect 38132 8800 38141 8840
rect 38515 8800 38524 8840
rect 38564 8800 41068 8840
rect 41108 8800 41117 8840
rect 42211 8800 42220 8840
rect 42260 8800 42796 8840
rect 42836 8800 42845 8840
rect 33100 8716 33524 8756
rect 33100 8672 33140 8716
rect 25219 8632 25228 8672
rect 25268 8632 25516 8672
rect 25556 8632 25565 8672
rect 25612 8632 25708 8672
rect 25748 8632 25757 8672
rect 25987 8632 25996 8672
rect 26036 8632 26284 8672
rect 26324 8632 26333 8672
rect 26380 8632 26476 8672
rect 26516 8632 26525 8672
rect 26707 8632 26716 8672
rect 26756 8632 28780 8672
rect 28820 8632 28829 8672
rect 29059 8632 29068 8672
rect 29108 8632 29356 8672
rect 29396 8632 29405 8672
rect 29635 8632 29644 8672
rect 29684 8632 29836 8672
rect 29876 8632 29885 8672
rect 32419 8632 32428 8672
rect 32468 8632 32477 8672
rect 32803 8632 32812 8672
rect 32852 8632 33140 8672
rect 33187 8632 33196 8672
rect 33236 8632 33388 8672
rect 33428 8632 33437 8672
rect 33484 8588 33524 8716
rect 33964 8716 38860 8756
rect 38900 8716 38909 8756
rect 40675 8716 40684 8756
rect 40724 8716 41260 8756
rect 41300 8716 41309 8756
rect 41635 8716 41644 8756
rect 41684 8716 41932 8756
rect 41972 8716 42220 8756
rect 42260 8716 42508 8756
rect 42548 8716 43180 8756
rect 43220 8716 43229 8756
rect 33964 8672 34004 8716
rect 43276 8672 43316 8968
rect 43363 8884 43372 8924
rect 43412 8884 43420 8924
rect 43460 8884 43543 8924
rect 43660 8672 43700 9052
rect 44764 9008 44804 9136
rect 46278 9008 46368 9028
rect 44764 8968 46368 9008
rect 46278 8948 46368 8968
rect 44371 8800 44380 8840
rect 44420 8800 46196 8840
rect 46156 8672 46196 8800
rect 46278 8672 46368 8692
rect 33571 8632 33580 8672
rect 33620 8632 33772 8672
rect 33812 8632 33821 8672
rect 33955 8632 33964 8672
rect 34004 8632 34013 8672
rect 34339 8632 34348 8672
rect 34388 8632 34540 8672
rect 34580 8632 34589 8672
rect 34723 8632 34732 8672
rect 34772 8632 34781 8672
rect 35107 8632 35116 8672
rect 35156 8632 35404 8672
rect 35444 8632 35453 8672
rect 35530 8632 35539 8672
rect 35579 8632 37900 8672
rect 37940 8632 37949 8672
rect 38083 8632 38092 8672
rect 38132 8632 38284 8672
rect 38324 8632 38764 8672
rect 38804 8632 39052 8672
rect 39092 8632 39340 8672
rect 39380 8632 39628 8672
rect 39668 8632 39916 8672
rect 39956 8632 40204 8672
rect 40244 8632 40492 8672
rect 40532 8632 40780 8672
rect 40820 8632 40972 8672
rect 41012 8632 41021 8672
rect 41731 8632 41740 8672
rect 41780 8632 42652 8672
rect 42692 8632 42701 8672
rect 42761 8632 42892 8672
rect 42932 8632 42941 8672
rect 43075 8632 43084 8672
rect 43124 8632 43220 8672
rect 43267 8632 43276 8672
rect 43316 8632 43325 8672
rect 43651 8632 43660 8672
rect 43700 8632 43709 8672
rect 43843 8632 43852 8672
rect 43892 8632 43948 8672
rect 43988 8632 44140 8672
rect 44180 8632 44189 8672
rect 44323 8632 44332 8672
rect 44372 8632 44524 8672
rect 44564 8632 44573 8672
rect 44899 8632 44908 8672
rect 44948 8632 45004 8672
rect 45044 8632 45079 8672
rect 46156 8632 46368 8672
rect 34732 8588 34772 8632
rect 43180 8588 43220 8632
rect 46278 8612 46368 8632
rect 23692 8548 23924 8588
rect 25132 8548 25844 8588
rect 27523 8548 27532 8588
rect 27572 8548 31948 8588
rect 31988 8548 31997 8588
rect 33484 8548 34636 8588
rect 34676 8548 34685 8588
rect 34732 8548 35308 8588
rect 35348 8548 35357 8588
rect 35404 8548 43124 8588
rect 43180 8548 44660 8588
rect 44755 8548 44764 8588
rect 44804 8548 45772 8588
rect 45812 8548 45821 8588
rect 11980 8504 12020 8548
rect 25132 8504 25172 8548
rect 11753 8464 11836 8504
rect 11876 8464 11884 8504
rect 11924 8464 11933 8504
rect 11980 8464 13420 8504
rect 13460 8464 13469 8504
rect 13987 8464 13996 8504
rect 14036 8464 16972 8504
rect 17012 8464 17021 8504
rect 17443 8464 17452 8504
rect 17492 8464 17644 8504
rect 17684 8464 17693 8504
rect 18691 8464 18700 8504
rect 18740 8464 19756 8504
rect 19796 8464 19805 8504
rect 19939 8464 19948 8504
rect 19988 8464 19997 8504
rect 20131 8464 20140 8504
rect 20180 8464 20189 8504
rect 20812 8464 25172 8504
rect 25804 8504 25844 8548
rect 35404 8504 35444 8548
rect 43084 8504 43124 8548
rect 25804 8464 25940 8504
rect 26035 8464 26044 8504
rect 26084 8464 26092 8504
rect 26132 8464 26215 8504
rect 27619 8464 27628 8504
rect 27668 8464 28684 8504
rect 28724 8464 28733 8504
rect 29107 8464 29116 8504
rect 29156 8464 29260 8504
rect 29300 8464 29309 8504
rect 29827 8464 29836 8504
rect 29876 8464 35444 8504
rect 35491 8464 35500 8504
rect 35540 8464 38380 8504
rect 38420 8464 38429 8504
rect 38851 8464 38860 8504
rect 38900 8464 40108 8504
rect 40148 8464 40157 8504
rect 40291 8464 40300 8504
rect 40340 8464 43028 8504
rect 43084 8464 43372 8504
rect 43412 8464 43421 8504
rect 12067 8380 12076 8420
rect 12116 8380 19852 8420
rect 19892 8380 19901 8420
rect 19948 8336 19988 8464
rect 20140 8420 20180 8464
rect 20812 8420 20852 8464
rect 20140 8380 20852 8420
rect 20899 8380 20908 8420
rect 20948 8380 25844 8420
rect 0 8296 1652 8336
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19948 8296 25612 8336
rect 25652 8296 25661 8336
rect 0 8276 90 8296
rect 15340 8212 15916 8252
rect 15956 8212 15965 8252
rect 19843 8212 19852 8252
rect 19892 8212 19901 8252
rect 20131 8212 20140 8252
rect 20180 8212 25708 8252
rect 25748 8212 25757 8252
rect 11155 8128 11164 8168
rect 11204 8128 11404 8168
rect 11444 8128 11453 8168
rect 14227 8128 14236 8168
rect 14276 8128 14380 8168
rect 14420 8128 14429 8168
rect 15340 8084 15380 8212
rect 19852 8168 19892 8212
rect 25804 8168 25844 8380
rect 25900 8252 25940 8464
rect 42988 8420 43028 8464
rect 25987 8380 25996 8420
rect 26036 8380 29740 8420
rect 29780 8380 29789 8420
rect 30211 8380 30220 8420
rect 30260 8380 36692 8420
rect 36739 8380 36748 8420
rect 36788 8380 42892 8420
rect 42932 8380 42941 8420
rect 42988 8380 43220 8420
rect 36652 8336 36692 8380
rect 27427 8296 27436 8336
rect 27476 8296 28492 8336
rect 28532 8296 28541 8336
rect 28675 8296 28684 8336
rect 28724 8296 31564 8336
rect 31604 8296 31613 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 36652 8296 43084 8336
rect 43124 8296 43133 8336
rect 43180 8252 43220 8380
rect 25900 8212 28724 8252
rect 30115 8212 30124 8252
rect 30164 8212 32620 8252
rect 32660 8212 32669 8252
rect 35683 8212 35692 8252
rect 35732 8212 43124 8252
rect 43180 8212 44276 8252
rect 28684 8168 28724 8212
rect 15532 8128 16724 8168
rect 18473 8128 18604 8168
rect 18644 8128 18653 8168
rect 19651 8128 19660 8168
rect 19700 8128 19796 8168
rect 19852 8128 25748 8168
rect 25804 8128 28540 8168
rect 28580 8128 28589 8168
rect 28684 8128 28924 8168
rect 28964 8128 28973 8168
rect 29731 8128 29740 8168
rect 29780 8128 31228 8168
rect 31268 8128 31277 8168
rect 31939 8128 31948 8168
rect 31988 8128 31996 8168
rect 32036 8128 32119 8168
rect 34867 8128 34876 8168
rect 34916 8128 35020 8168
rect 35060 8128 35069 8168
rect 35225 8128 35308 8168
rect 35348 8128 35356 8168
rect 35396 8128 35405 8168
rect 37699 8128 37708 8168
rect 37748 8128 42356 8168
rect 10147 8044 10156 8084
rect 10196 8044 11348 8084
rect 12835 8044 12844 8084
rect 12884 8044 13940 8084
rect 15043 8044 15052 8084
rect 15092 8044 15284 8084
rect 15331 8044 15340 8084
rect 15380 8044 15389 8084
rect 0 8000 90 8020
rect 11308 8000 11348 8044
rect 13900 8000 13940 8044
rect 15244 8000 15284 8044
rect 15532 8000 15572 8128
rect 15724 8044 16300 8084
rect 16340 8044 16349 8084
rect 15724 8000 15764 8044
rect 0 7960 652 8000
rect 692 7960 701 8000
rect 1097 7960 1228 8000
rect 1268 7960 1277 8000
rect 1603 7960 1612 8000
rect 1652 7960 1661 8000
rect 10915 7960 10924 8000
rect 10964 7960 10973 8000
rect 11177 7960 11308 8000
rect 11348 7960 11357 8000
rect 11657 7960 11788 8000
rect 11828 7960 12212 8000
rect 13891 7960 13900 8000
rect 13940 7960 13949 8000
rect 14467 7960 14476 8000
rect 14516 7960 14996 8000
rect 15139 7960 15148 8000
rect 15188 7960 15197 8000
rect 15244 7960 15340 8000
rect 15380 7960 15572 8000
rect 15706 7960 15715 8000
rect 15755 7960 15764 8000
rect 15907 7960 15916 8000
rect 15956 7960 16100 8000
rect 16186 7960 16195 8000
rect 16244 7960 16375 8000
rect 0 7940 90 7960
rect 1612 7832 1652 7960
rect 10924 7916 10964 7960
rect 12172 7916 12212 7960
rect 13420 7916 13460 7925
rect 14956 7916 14996 7960
rect 15148 7916 15188 7960
rect 15532 7916 15572 7960
rect 16060 7916 16100 7960
rect 16684 7943 16724 8128
rect 19756 8084 19796 8128
rect 25708 8084 25748 8128
rect 16771 8044 16780 8084
rect 16820 8044 18740 8084
rect 19756 8044 19900 8084
rect 19940 8044 19949 8084
rect 20131 8044 20140 8084
rect 20180 8044 23060 8084
rect 25708 8044 28684 8084
rect 28724 8044 28733 8084
rect 28780 8044 29068 8084
rect 29108 8044 29356 8084
rect 29396 8044 29405 8084
rect 29635 8044 29644 8084
rect 29684 8044 29836 8084
rect 29876 8044 29885 8084
rect 31555 8044 31564 8084
rect 31604 8044 31612 8084
rect 31652 8044 31735 8084
rect 34531 8044 34540 8084
rect 34580 8044 34972 8084
rect 35012 8044 35021 8084
rect 35875 8044 35884 8084
rect 35924 8044 42124 8084
rect 42164 8044 42173 8084
rect 18700 8000 18740 8044
rect 17155 7960 17164 8000
rect 17204 7960 17548 8000
rect 17588 7960 17597 8000
rect 18700 7960 19660 8000
rect 19700 7960 20180 8000
rect 16666 7934 16724 7943
rect 10924 7876 11980 7916
rect 12020 7876 12029 7916
rect 12163 7876 12172 7916
rect 12212 7876 12221 7916
rect 13289 7876 13420 7916
rect 13460 7876 13469 7916
rect 14537 7876 14659 7916
rect 14708 7876 14717 7916
rect 14825 7876 14956 7916
rect 14996 7876 15005 7916
rect 15101 7876 15134 7916
rect 15174 7876 15188 7916
rect 15235 7876 15244 7916
rect 15284 7876 15293 7916
rect 15388 7876 15437 7916
rect 15477 7876 15486 7916
rect 15532 7876 15575 7916
rect 15615 7876 15624 7916
rect 15811 7876 15820 7916
rect 15860 7876 15869 7916
rect 16051 7876 16060 7916
rect 16100 7876 16109 7916
rect 16291 7876 16300 7916
rect 16340 7876 16471 7916
rect 16666 7894 16675 7934
rect 16715 7894 16724 7934
rect 17740 7916 17780 7925
rect 16666 7893 16724 7894
rect 16771 7876 16780 7916
rect 16820 7876 17068 7916
rect 17108 7876 17117 7916
rect 17251 7876 17260 7916
rect 17300 7876 17492 7916
rect 17609 7876 17740 7916
rect 17780 7876 17789 7916
rect 18219 7876 18228 7916
rect 18268 7876 18277 7916
rect 13420 7867 13460 7876
rect 15244 7832 15284 7876
rect 15388 7832 15428 7876
rect 15820 7832 15860 7876
rect 17452 7832 17492 7876
rect 17740 7867 17780 7876
rect 844 7792 1652 7832
rect 12019 7792 12028 7832
rect 12068 7792 12940 7832
rect 12980 7792 12989 7832
rect 14131 7792 14140 7832
rect 14180 7792 14476 7832
rect 14516 7792 14525 7832
rect 14851 7792 14860 7832
rect 14900 7792 15284 7832
rect 15361 7792 16052 7832
rect 16265 7792 16387 7832
rect 16436 7792 16445 7832
rect 17452 7792 17548 7832
rect 17588 7792 17597 7832
rect 0 7664 90 7684
rect 844 7664 884 7792
rect 15388 7748 15428 7792
rect 16012 7748 16052 7792
rect 18237 7748 18277 7876
rect 18412 7876 18604 7916
rect 18644 7876 18653 7916
rect 18787 7876 18796 7916
rect 18836 7876 18967 7916
rect 18412 7748 18452 7876
rect 20140 7748 20180 7960
rect 20236 7916 20276 7925
rect 23020 7916 23060 8044
rect 28780 8000 28820 8044
rect 42316 8000 42356 8128
rect 43084 8000 43124 8212
rect 43219 8128 43228 8168
rect 43268 8128 43276 8168
rect 43316 8128 43399 8168
rect 43555 8044 43564 8084
rect 43604 8044 43612 8084
rect 43652 8044 43735 8084
rect 44236 8000 44276 8212
rect 44620 8000 44660 8548
rect 45139 8464 45148 8504
rect 45188 8464 45676 8504
rect 45716 8464 45725 8504
rect 46278 8336 46368 8356
rect 45859 8296 45868 8336
rect 45908 8296 46368 8336
rect 46278 8276 46368 8296
rect 46278 8000 46368 8020
rect 25603 7960 25612 8000
rect 25652 7960 25996 8000
rect 26036 7960 26188 8000
rect 26228 7960 26237 8000
rect 28771 7960 28780 8000
rect 28820 7960 28829 8000
rect 28963 7960 28972 8000
rect 29012 7960 29164 8000
rect 29204 7960 29213 8000
rect 29434 7960 29443 8000
rect 29483 7960 29836 8000
rect 29876 7960 29885 8000
rect 31459 7960 31468 8000
rect 31508 7960 31639 8000
rect 31747 7960 31756 8000
rect 31796 7960 31852 8000
rect 31892 7960 31927 8000
rect 32105 7960 32236 8000
rect 32276 7960 32285 8000
rect 34339 7960 34348 8000
rect 34388 7960 34636 8000
rect 34676 7960 34685 8000
rect 35203 7960 35212 8000
rect 35252 7960 35261 8000
rect 35587 7960 35596 8000
rect 35636 7960 38188 8000
rect 38228 7960 38237 8000
rect 38371 7960 38380 8000
rect 38420 7960 38429 8000
rect 38825 7960 38860 8000
rect 38900 7960 38956 8000
rect 38996 7960 39005 8000
rect 39689 7960 39820 8000
rect 39860 7960 39869 8000
rect 40025 7960 40108 8000
rect 40148 7960 40156 8000
rect 40196 7960 40205 8000
rect 40265 7960 40396 8000
rect 40436 7960 40445 8000
rect 42307 7960 42316 8000
rect 42356 7960 42365 8000
rect 42691 7960 42700 8000
rect 42740 7960 42749 8000
rect 43075 7960 43084 8000
rect 43124 7960 43133 8000
rect 43337 7960 43372 8000
rect 43412 7960 43468 8000
rect 43508 7960 43517 8000
rect 43721 7960 43756 8000
rect 43796 7960 43852 8000
rect 43892 7960 43901 8000
rect 44227 7960 44236 8000
rect 44276 7960 44285 8000
rect 44611 7960 44620 8000
rect 44660 7960 44669 8000
rect 44777 7960 44908 8000
rect 44948 7960 44957 8000
rect 45763 7960 45772 8000
rect 45812 7960 46368 8000
rect 35212 7916 35252 7960
rect 20276 7876 20716 7916
rect 20756 7876 21196 7916
rect 21236 7876 21245 7916
rect 21475 7876 21484 7916
rect 21524 7876 21533 7916
rect 23020 7876 27532 7916
rect 27572 7876 27581 7916
rect 29059 7876 29068 7916
rect 29108 7876 29308 7916
rect 29348 7876 29357 7916
rect 29452 7876 29548 7916
rect 29588 7876 29597 7916
rect 29705 7876 29740 7916
rect 29780 7876 29836 7916
rect 29876 7876 29885 7916
rect 29942 7876 29951 7916
rect 29991 7876 30000 7916
rect 30115 7876 30124 7916
rect 30164 7876 30211 7916
rect 30307 7876 30316 7916
rect 30356 7876 30365 7916
rect 30499 7876 30508 7916
rect 30548 7876 30679 7916
rect 35212 7876 35980 7916
rect 36020 7876 36029 7916
rect 36844 7876 38284 7916
rect 38324 7876 38333 7916
rect 20236 7867 20276 7876
rect 21484 7748 21524 7876
rect 29452 7832 29492 7876
rect 29951 7832 29991 7876
rect 30124 7832 30164 7876
rect 30316 7832 30356 7876
rect 36844 7832 36884 7876
rect 38380 7832 38420 7960
rect 42700 7916 42740 7960
rect 46278 7940 46368 7960
rect 38467 7876 38476 7916
rect 38516 7876 42740 7916
rect 28291 7792 28300 7832
rect 28340 7792 29492 7832
rect 29904 7792 29932 7832
rect 29972 7792 29991 7832
rect 30115 7792 30124 7832
rect 30164 7792 30173 7832
rect 30307 7792 30316 7832
rect 30356 7792 30403 7832
rect 30787 7792 30796 7832
rect 30836 7792 36884 7832
rect 37027 7792 37036 7832
rect 37076 7792 37228 7832
rect 37268 7792 37516 7832
rect 37556 7792 37804 7832
rect 37844 7792 38092 7832
rect 38132 7792 38420 7832
rect 40051 7792 40060 7832
rect 40100 7792 41684 7832
rect 41827 7792 41836 7832
rect 41876 7792 42844 7832
rect 42884 7792 42893 7832
rect 42979 7792 42988 7832
rect 43028 7792 43996 7832
rect 44036 7792 44045 7832
rect 1459 7708 1468 7748
rect 1508 7708 1748 7748
rect 1843 7708 1852 7748
rect 1892 7708 10060 7748
rect 10100 7708 10109 7748
rect 11539 7708 11548 7748
rect 11588 7708 11884 7748
rect 11924 7708 11933 7748
rect 13603 7708 13612 7748
rect 13652 7708 15428 7748
rect 15785 7708 15907 7748
rect 15956 7708 15965 7748
rect 16012 7708 18277 7748
rect 18403 7708 18412 7748
rect 18452 7708 18461 7748
rect 18787 7708 18796 7748
rect 18836 7708 20044 7748
rect 20084 7708 20093 7748
rect 20140 7708 21524 7748
rect 26227 7708 26236 7748
rect 26276 7708 27340 7748
rect 27380 7708 27389 7748
rect 28780 7708 29108 7748
rect 29155 7708 29164 7748
rect 29204 7708 29635 7748
rect 29675 7708 29684 7748
rect 30403 7708 30412 7748
rect 30452 7708 30700 7748
rect 30740 7708 30749 7748
rect 30883 7708 30892 7748
rect 30932 7708 32236 7748
rect 32276 7708 32285 7748
rect 32419 7708 32428 7748
rect 32468 7708 37708 7748
rect 37748 7708 37757 7748
rect 38611 7708 38620 7748
rect 38660 7708 39052 7748
rect 39092 7708 39101 7748
rect 39187 7708 39196 7748
rect 39236 7708 39916 7748
rect 39956 7708 39965 7748
rect 0 7624 884 7664
rect 0 7604 90 7624
rect 1708 7412 1748 7708
rect 28780 7664 28820 7708
rect 12163 7624 12172 7664
rect 12212 7624 16916 7664
rect 17251 7624 17260 7664
rect 17300 7624 25420 7664
rect 25460 7624 25469 7664
rect 28195 7624 28204 7664
rect 28244 7624 28628 7664
rect 28675 7624 28684 7664
rect 28724 7624 28820 7664
rect 29068 7664 29108 7708
rect 41644 7664 41684 7792
rect 41731 7708 41740 7748
rect 41780 7708 42076 7748
rect 42116 7708 42125 7748
rect 42211 7708 42220 7748
rect 42260 7708 42460 7748
rect 42500 7708 42509 7748
rect 43747 7708 43756 7748
rect 43796 7708 44380 7748
rect 44420 7708 44429 7748
rect 45139 7708 45148 7748
rect 45188 7708 45868 7748
rect 45908 7708 45917 7748
rect 46278 7664 46368 7684
rect 29068 7624 32564 7664
rect 38563 7624 38572 7664
rect 38612 7624 40396 7664
rect 40436 7624 40445 7664
rect 41644 7624 44908 7664
rect 44948 7624 44957 7664
rect 45667 7624 45676 7664
rect 45716 7624 46368 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 9283 7540 9292 7580
rect 9332 7540 16780 7580
rect 16820 7540 16829 7580
rect 16876 7496 16916 7624
rect 28588 7580 28628 7624
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 20515 7540 20524 7580
rect 20564 7540 24940 7580
rect 24980 7540 24989 7580
rect 25324 7540 28492 7580
rect 28532 7540 28541 7580
rect 28588 7540 28780 7580
rect 28820 7540 28829 7580
rect 32419 7540 32428 7580
rect 32468 7540 32477 7580
rect 25324 7496 25364 7540
rect 32428 7496 32468 7540
rect 16876 7456 17108 7496
rect 19651 7456 19660 7496
rect 19700 7456 25364 7496
rect 25411 7456 25420 7496
rect 25460 7456 28532 7496
rect 28963 7456 28972 7496
rect 29012 7456 29204 7496
rect 17068 7412 17108 7456
rect 28492 7412 28532 7456
rect 1708 7372 16012 7412
rect 16052 7372 16061 7412
rect 16195 7372 16204 7412
rect 16244 7372 16963 7412
rect 17003 7372 17012 7412
rect 17068 7372 25516 7412
rect 25556 7372 25565 7412
rect 28492 7372 28876 7412
rect 28916 7372 28925 7412
rect 0 7328 90 7348
rect 0 7288 1228 7328
rect 1268 7288 1277 7328
rect 13027 7288 13036 7328
rect 13076 7288 14668 7328
rect 14708 7288 15340 7328
rect 15380 7288 15956 7328
rect 16099 7288 16108 7328
rect 16148 7288 16436 7328
rect 27331 7288 27340 7328
rect 27380 7288 28300 7328
rect 28340 7288 28349 7328
rect 28540 7288 28820 7328
rect 28937 7288 29068 7328
rect 29108 7288 29117 7328
rect 0 7268 90 7288
rect 15916 7244 15956 7288
rect 16396 7244 16436 7288
rect 28540 7244 28580 7288
rect 28780 7244 28820 7288
rect 29164 7244 29204 7456
rect 29644 7456 30548 7496
rect 30595 7456 30604 7496
rect 30644 7456 32468 7496
rect 29308 7372 29356 7412
rect 29396 7372 29405 7412
rect 29308 7244 29348 7372
rect 29644 7244 29684 7456
rect 29951 7288 30124 7328
rect 30164 7288 30173 7328
rect 29951 7251 29991 7288
rect 29941 7244 29991 7251
rect 30220 7244 30260 7456
rect 30508 7412 30548 7456
rect 32524 7412 32564 7624
rect 46278 7604 46368 7624
rect 32611 7540 32620 7580
rect 32660 7540 35020 7580
rect 35060 7540 35069 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 35779 7540 35788 7580
rect 35828 7540 42988 7580
rect 43028 7540 43037 7580
rect 39043 7456 39052 7496
rect 39092 7456 44620 7496
rect 44660 7456 44669 7496
rect 30508 7372 32140 7412
rect 32180 7372 32189 7412
rect 32524 7372 41740 7412
rect 41780 7372 41789 7412
rect 42778 7372 42787 7412
rect 42827 7372 43468 7412
rect 43508 7372 44227 7412
rect 44267 7372 44276 7412
rect 46278 7328 46368 7348
rect 30787 7288 30796 7328
rect 30836 7288 42220 7328
rect 42260 7288 42269 7328
rect 45859 7288 45868 7328
rect 45908 7288 46368 7328
rect 46278 7268 46368 7288
rect 11299 7204 11308 7244
rect 11348 7204 11596 7244
rect 11636 7204 11645 7244
rect 12809 7235 12940 7244
rect 12809 7204 12844 7235
rect 12884 7204 12940 7235
rect 12980 7204 13420 7244
rect 13460 7204 13469 7244
rect 15898 7204 15907 7244
rect 15947 7204 15956 7244
rect 16099 7204 16108 7244
rect 16148 7204 16204 7244
rect 16244 7204 16279 7244
rect 16396 7204 16631 7244
rect 16671 7204 16680 7244
rect 16867 7204 16876 7244
rect 16916 7204 18796 7244
rect 18836 7204 18845 7244
rect 25516 7204 25900 7244
rect 25940 7204 25949 7244
rect 27017 7204 27148 7244
rect 27188 7204 27197 7244
rect 28483 7204 28492 7244
rect 28532 7204 28580 7244
rect 28666 7204 28675 7244
rect 28715 7204 28724 7244
rect 12844 7186 12884 7195
rect 25516 7160 25556 7204
rect 27148 7186 27188 7195
rect 28684 7160 28724 7204
rect 28780 7204 28855 7244
rect 28895 7204 28904 7244
rect 29155 7204 29164 7244
rect 29204 7204 29213 7244
rect 29308 7204 29355 7244
rect 29395 7204 29404 7244
rect 29596 7204 29644 7244
rect 29684 7204 29693 7244
rect 29922 7204 29931 7244
rect 29971 7211 29991 7244
rect 29971 7204 29981 7211
rect 30160 7204 30169 7244
rect 30209 7204 30260 7244
rect 30473 7204 30499 7244
rect 30539 7204 30604 7244
rect 30644 7204 30653 7244
rect 30883 7204 30892 7244
rect 30932 7235 31063 7244
rect 30932 7204 30988 7235
rect 28780 7160 28820 7204
rect 29596 7202 29636 7204
rect 29548 7162 29636 7202
rect 31028 7204 31063 7235
rect 31433 7204 31468 7244
rect 31508 7204 31564 7244
rect 31604 7204 31613 7244
rect 31747 7204 31756 7244
rect 31796 7204 31948 7244
rect 31988 7204 31997 7244
rect 32057 7204 32066 7244
rect 32106 7204 32140 7244
rect 32180 7204 32246 7244
rect 38179 7204 38188 7244
rect 38228 7204 39436 7244
rect 39476 7204 39485 7244
rect 39907 7204 39916 7244
rect 39956 7204 41836 7244
rect 41876 7204 41885 7244
rect 30988 7186 31028 7195
rect 29548 7160 29588 7162
rect 3427 7120 3436 7160
rect 3476 7120 3485 7160
rect 3811 7120 3820 7160
rect 3860 7120 3869 7160
rect 3977 7120 4060 7160
rect 4100 7120 4108 7160
rect 4148 7120 4157 7160
rect 15043 7120 15052 7160
rect 15092 7120 15244 7160
rect 15284 7120 15293 7160
rect 15427 7120 15436 7160
rect 15476 7120 15484 7160
rect 15524 7120 15607 7160
rect 15715 7120 15724 7160
rect 15764 7120 15860 7160
rect 15907 7120 15916 7160
rect 15956 7120 16771 7160
rect 16811 7120 16820 7160
rect 17347 7120 17356 7160
rect 17396 7120 17500 7160
rect 17540 7120 17549 7160
rect 17644 7120 17740 7160
rect 17780 7120 17932 7160
rect 17972 7120 17981 7160
rect 18115 7120 18124 7160
rect 18164 7120 18173 7160
rect 18691 7120 18700 7160
rect 18740 7120 21868 7160
rect 21908 7120 22156 7160
rect 22196 7120 22205 7160
rect 25385 7120 25516 7160
rect 25556 7120 25565 7160
rect 28483 7120 28492 7160
rect 28532 7120 28724 7160
rect 28771 7120 28780 7160
rect 28820 7120 29588 7160
rect 29705 7120 29836 7160
rect 29876 7120 29885 7160
rect 30051 7151 30116 7160
rect 0 6992 90 7012
rect 0 6952 748 6992
rect 788 6952 797 6992
rect 0 6932 90 6952
rect 0 6656 90 6676
rect 3436 6656 3476 7120
rect 3820 7076 3860 7120
rect 15820 7076 15860 7120
rect 17644 7076 17684 7120
rect 18124 7076 18164 7120
rect 30051 7111 30067 7151
rect 30107 7111 30116 7151
rect 31459 7120 31468 7160
rect 31508 7120 31564 7160
rect 31604 7120 31639 7160
rect 35683 7120 35692 7160
rect 35732 7120 37708 7160
rect 37748 7120 37757 7160
rect 37961 7120 38092 7160
rect 38132 7120 38380 7160
rect 38420 7120 38668 7160
rect 38708 7120 38717 7160
rect 38873 7120 38956 7160
rect 38996 7120 39004 7160
rect 39044 7120 39053 7160
rect 39331 7120 39340 7160
rect 39380 7120 39436 7160
rect 39476 7120 39724 7160
rect 39764 7120 40012 7160
rect 40052 7120 40061 7160
rect 40505 7120 40588 7160
rect 40628 7120 40636 7160
rect 40676 7120 40685 7160
rect 40745 7120 40876 7160
rect 40916 7120 40925 7160
rect 41251 7120 41260 7160
rect 41300 7120 42940 7160
rect 42980 7120 42989 7160
rect 43049 7120 43084 7160
rect 43124 7120 43180 7160
rect 43220 7120 43284 7160
rect 43433 7120 43564 7160
rect 43604 7120 43613 7160
rect 43939 7120 43948 7160
rect 43988 7120 43997 7160
rect 44393 7120 44524 7160
rect 44564 7120 44573 7160
rect 44899 7120 44908 7160
rect 44948 7120 44957 7160
rect 30051 7110 30116 7111
rect 30051 7076 30091 7110
rect 3820 7036 8428 7076
rect 8468 7036 8477 7076
rect 15283 7036 15292 7076
rect 15332 7036 15532 7076
rect 15572 7036 15581 7076
rect 15811 7036 15820 7076
rect 15860 7036 15869 7076
rect 17539 7036 17548 7076
rect 17588 7036 17684 7076
rect 17731 7036 17740 7076
rect 17780 7036 18164 7076
rect 18220 7036 23692 7076
rect 23732 7036 23741 7076
rect 25747 7036 25756 7076
rect 25796 7036 28396 7076
rect 28436 7036 28445 7076
rect 30019 7036 30028 7076
rect 30068 7036 30091 7076
rect 35443 7036 35452 7076
rect 35492 7036 35596 7076
rect 35636 7036 35645 7076
rect 39139 7036 39148 7076
rect 39188 7036 43324 7076
rect 43364 7036 43373 7076
rect 3667 6952 3676 6992
rect 3716 6952 10828 6992
rect 10868 6952 10877 6992
rect 17644 6952 17884 6992
rect 17924 6952 17933 6992
rect 17644 6908 17684 6952
rect 18220 6908 18260 7036
rect 20707 6952 20716 6992
rect 20756 6952 21628 6992
rect 21668 6952 21677 6992
rect 22313 6952 22396 6992
rect 22436 6952 22444 6992
rect 22484 6952 23060 6992
rect 28195 6952 28204 6992
rect 28244 6952 28675 6992
rect 28715 6952 28724 6992
rect 29059 6952 29068 6992
rect 29108 6952 29356 6992
rect 29396 6952 29405 6992
rect 30259 6952 30268 6992
rect 30308 6952 30316 6992
rect 30356 6952 30439 6992
rect 33004 6952 35156 6992
rect 35779 6952 35788 6992
rect 35828 6952 38668 6992
rect 38708 6952 38717 6992
rect 39283 6952 39292 6992
rect 39332 6952 39341 6992
rect 41347 6952 41356 6992
rect 41396 6952 41972 6992
rect 12355 6868 12364 6908
rect 12404 6868 17684 6908
rect 17836 6868 18260 6908
rect 23020 6908 23060 6952
rect 33004 6908 33044 6952
rect 23020 6868 27148 6908
rect 27188 6868 27197 6908
rect 28675 6868 28684 6908
rect 28724 6868 29356 6908
rect 29396 6868 29405 6908
rect 29539 6868 29548 6908
rect 29588 6868 33044 6908
rect 33100 6868 35020 6908
rect 35060 6868 35069 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 11875 6784 11884 6824
rect 11924 6784 17740 6824
rect 17780 6784 17789 6824
rect 17836 6740 17876 6868
rect 33100 6824 33140 6868
rect 17923 6784 17932 6824
rect 17972 6784 18700 6824
rect 18740 6784 18749 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 24163 6784 24172 6824
rect 24212 6784 27284 6824
rect 27331 6784 27340 6824
rect 27380 6784 33140 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 27244 6740 27284 6784
rect 35116 6740 35156 6952
rect 35299 6868 35308 6908
rect 35348 6868 37996 6908
rect 38036 6868 38045 6908
rect 39292 6824 39332 6952
rect 41932 6824 41972 6952
rect 43180 6952 43708 6992
rect 43748 6952 43757 6992
rect 43180 6824 43220 6952
rect 39292 6784 41740 6824
rect 41780 6784 41789 6824
rect 41932 6784 43220 6824
rect 13219 6700 13228 6740
rect 13268 6700 17876 6740
rect 17932 6700 25612 6740
rect 25652 6700 25661 6740
rect 27244 6700 29356 6740
rect 29396 6700 29405 6740
rect 29539 6700 29548 6740
rect 29588 6700 35020 6740
rect 35060 6700 35069 6740
rect 35116 6700 43084 6740
rect 43124 6700 43133 6740
rect 0 6616 844 6656
rect 884 6616 893 6656
rect 3436 6616 17836 6656
rect 17876 6616 17885 6656
rect 0 6596 90 6616
rect 17932 6572 17972 6700
rect 18019 6616 18028 6656
rect 18068 6616 23212 6656
rect 23252 6616 23261 6656
rect 27244 6616 27340 6656
rect 27380 6616 27389 6656
rect 27497 6616 27628 6656
rect 27668 6616 27677 6656
rect 28291 6616 28300 6656
rect 28340 6616 29836 6656
rect 29876 6616 29885 6656
rect 30010 6616 30019 6656
rect 30059 6616 30508 6656
rect 30548 6616 30557 6656
rect 40291 6616 40300 6656
rect 40340 6616 41780 6656
rect 27244 6572 27284 6616
rect 10051 6532 10060 6572
rect 10100 6532 17972 6572
rect 19459 6532 19468 6572
rect 19508 6532 27284 6572
rect 27340 6532 35116 6572
rect 35156 6532 35165 6572
rect 35299 6532 35308 6572
rect 35348 6532 41684 6572
rect 27340 6488 27380 6532
rect 41644 6488 41684 6532
rect 41740 6488 41780 6616
rect 43948 6572 43988 7120
rect 44908 7076 44948 7120
rect 41932 6532 43988 6572
rect 44044 7036 44948 7076
rect 41932 6488 41972 6532
rect 44044 6488 44084 7036
rect 46278 6992 46368 7012
rect 44755 6952 44764 6992
rect 44804 6952 44813 6992
rect 45139 6952 45148 6992
rect 45188 6952 46368 6992
rect 44764 6824 44804 6952
rect 46278 6932 46368 6952
rect 44764 6784 46252 6824
rect 46292 6784 46301 6824
rect 46278 6656 46368 6676
rect 46243 6616 46252 6656
rect 46292 6616 46368 6656
rect 46278 6596 46368 6616
rect 1219 6448 1228 6488
rect 1268 6448 27380 6488
rect 27811 6448 27820 6488
rect 27860 6448 28780 6488
rect 28820 6448 28829 6488
rect 29002 6479 29164 6488
rect 29002 6439 29011 6479
rect 29051 6448 29164 6479
rect 29204 6448 29213 6488
rect 29347 6448 29356 6488
rect 29396 6448 29404 6488
rect 29444 6448 29527 6488
rect 29635 6448 29644 6488
rect 29684 6448 29780 6488
rect 29827 6448 29836 6488
rect 29876 6448 29885 6488
rect 30403 6448 30412 6488
rect 30452 6448 31180 6488
rect 31220 6448 31660 6488
rect 31700 6448 31709 6488
rect 34505 6448 34636 6488
rect 34676 6448 34685 6488
rect 34793 6448 34876 6488
rect 34916 6448 34924 6488
rect 34964 6448 34973 6488
rect 35299 6448 35308 6488
rect 35348 6448 35357 6488
rect 35561 6448 35692 6488
rect 35732 6448 35741 6488
rect 36451 6448 36460 6488
rect 36500 6448 37036 6488
rect 37076 6448 37085 6488
rect 37987 6448 37996 6488
rect 38036 6448 41260 6488
rect 41300 6448 41309 6488
rect 41635 6448 41644 6488
rect 41684 6448 41693 6488
rect 41740 6448 41972 6488
rect 43171 6448 43180 6488
rect 43220 6448 44084 6488
rect 44140 6532 44812 6572
rect 44852 6532 44861 6572
rect 29051 6439 29060 6448
rect 29002 6438 29060 6439
rect 27436 6404 27476 6413
rect 8419 6364 8428 6404
rect 8468 6364 23308 6404
rect 23348 6364 23357 6404
rect 26057 6364 26188 6404
rect 26228 6364 26237 6404
rect 27523 6364 27532 6404
rect 27572 6364 28876 6404
rect 28916 6364 28925 6404
rect 29104 6364 29113 6404
rect 29153 6364 29548 6404
rect 29588 6364 29597 6404
rect 0 6320 90 6340
rect 27436 6320 27476 6364
rect 29740 6320 29780 6448
rect 29836 6404 29876 6448
rect 29834 6364 29843 6404
rect 29883 6364 29923 6404
rect 30010 6364 30019 6404
rect 30059 6364 30316 6404
rect 30356 6364 30365 6404
rect 0 6280 23060 6320
rect 27139 6280 27148 6320
rect 27188 6280 27476 6320
rect 27532 6280 29684 6320
rect 29740 6280 30028 6320
rect 30068 6280 30077 6320
rect 31363 6280 31372 6320
rect 31412 6280 34924 6320
rect 34964 6280 34973 6320
rect 0 6260 90 6280
rect 23020 6236 23060 6280
rect 27532 6236 27572 6280
rect 23020 6196 27572 6236
rect 28771 6196 28780 6236
rect 28820 6196 28876 6236
rect 28916 6196 28951 6236
rect 29644 6152 29684 6280
rect 29731 6196 29740 6236
rect 29780 6196 30940 6236
rect 30980 6196 30989 6236
rect 35308 6152 35348 6448
rect 35875 6364 35884 6404
rect 35924 6364 43564 6404
rect 43604 6364 43613 6404
rect 44140 6320 44180 6532
rect 44515 6448 44524 6488
rect 44564 6448 44573 6488
rect 44620 6448 44908 6488
rect 44948 6448 44957 6488
rect 37123 6280 37132 6320
rect 37172 6280 40876 6320
rect 40916 6280 40925 6320
rect 41875 6280 41884 6320
rect 41924 6280 44180 6320
rect 35539 6196 35548 6236
rect 35588 6196 35597 6236
rect 35923 6196 35932 6236
rect 35972 6196 37172 6236
rect 37267 6196 37276 6236
rect 37316 6196 40204 6236
rect 40244 6196 40253 6236
rect 40387 6196 40396 6236
rect 40436 6196 43084 6236
rect 43124 6196 43133 6236
rect 43459 6196 43468 6236
rect 43508 6196 43555 6236
rect 43595 6196 43639 6236
rect 43721 6196 43843 6236
rect 43892 6196 44131 6236
rect 44171 6196 44180 6236
rect 1315 6112 1324 6152
rect 1364 6112 17836 6152
rect 17876 6112 17885 6152
rect 18019 6112 18028 6152
rect 18068 6112 20524 6152
rect 20564 6112 20573 6152
rect 29644 6112 31084 6152
rect 31124 6112 31133 6152
rect 31267 6112 31276 6152
rect 31316 6112 35348 6152
rect 35548 6152 35588 6196
rect 37132 6152 37172 6196
rect 44524 6152 44564 6448
rect 35548 6112 37076 6152
rect 37132 6112 44564 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 27811 6028 27820 6068
rect 27860 6028 30988 6068
rect 31028 6028 31037 6068
rect 31459 6028 31468 6068
rect 31508 6028 35020 6068
rect 35060 6028 35069 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 0 5984 90 6004
rect 37036 5984 37076 6112
rect 38851 6028 38860 6068
rect 38900 6028 44524 6068
rect 44564 6028 44573 6068
rect 44620 5984 44660 6448
rect 46278 6320 46368 6340
rect 45139 6280 45148 6320
rect 45188 6280 46368 6320
rect 46278 6260 46368 6280
rect 44755 6196 44764 6236
rect 44804 6196 44813 6236
rect 44764 6152 44804 6196
rect 44764 6112 46252 6152
rect 46292 6112 46301 6152
rect 46278 5984 46368 6004
rect 0 5944 23692 5984
rect 23732 5944 23741 5984
rect 28003 5944 28012 5984
rect 28052 5944 30220 5984
rect 30260 5944 30269 5984
rect 37036 5944 44660 5984
rect 46243 5944 46252 5984
rect 46292 5944 46368 5984
rect 0 5924 90 5944
rect 46278 5924 46368 5944
rect 1411 5860 1420 5900
rect 1460 5860 18700 5900
rect 18740 5860 18749 5900
rect 25795 5860 25804 5900
rect 25844 5860 32908 5900
rect 32948 5860 32957 5900
rect 35500 5860 39148 5900
rect 39188 5860 39197 5900
rect 40108 5860 43084 5900
rect 43124 5860 43133 5900
rect 43267 5860 43276 5900
rect 43316 5860 44716 5900
rect 44756 5860 44765 5900
rect 12739 5776 12748 5816
rect 12788 5776 34580 5816
rect 34627 5776 34636 5816
rect 34676 5776 35404 5816
rect 35444 5776 35453 5816
rect 34540 5732 34580 5776
rect 35500 5732 35540 5860
rect 40108 5816 40148 5860
rect 35587 5776 35596 5816
rect 35636 5776 40148 5816
rect 40195 5776 40204 5816
rect 40244 5776 44948 5816
rect 23020 5692 34444 5732
rect 34484 5692 34493 5732
rect 34540 5692 35540 5732
rect 41731 5692 41740 5732
rect 41780 5692 44564 5732
rect 0 5648 90 5668
rect 0 5608 1324 5648
rect 1364 5608 1373 5648
rect 0 5588 90 5608
rect 23020 5564 23060 5692
rect 44524 5648 44564 5692
rect 44908 5648 44948 5776
rect 46278 5648 46368 5668
rect 16963 5524 16972 5564
rect 17012 5524 23060 5564
rect 33100 5608 34636 5648
rect 34676 5608 34685 5648
rect 34867 5608 34876 5648
rect 34916 5608 38860 5648
rect 38900 5608 38909 5648
rect 41635 5608 41644 5648
rect 41684 5608 43132 5648
rect 43172 5608 43181 5648
rect 43363 5608 43372 5648
rect 43412 5608 43421 5648
rect 43555 5608 43564 5648
rect 43604 5608 43852 5648
rect 43892 5608 44140 5648
rect 44180 5608 44189 5648
rect 44515 5608 44524 5648
rect 44564 5608 44573 5648
rect 44899 5608 44908 5648
rect 44948 5608 44957 5648
rect 45139 5608 45148 5648
rect 45188 5608 46368 5648
rect 33100 5396 33140 5608
rect 835 5356 844 5396
rect 884 5356 33140 5396
rect 0 5312 90 5332
rect 0 5272 1420 5312
rect 1460 5272 1469 5312
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 0 5252 90 5272
rect 2755 5188 2764 5228
rect 2804 5188 27628 5228
rect 27668 5188 27677 5228
rect 16387 5104 16396 5144
rect 16436 5104 24460 5144
rect 24500 5104 24509 5144
rect 29059 5104 29068 5144
rect 29108 5104 30604 5144
rect 30644 5104 30653 5144
rect 4771 5020 4780 5060
rect 4820 5020 20852 5060
rect 0 4976 90 4996
rect 20812 4976 20852 5020
rect 21292 5020 33140 5060
rect 0 4936 2900 4976
rect 12259 4936 12268 4976
rect 12308 4936 13076 4976
rect 20803 4936 20812 4976
rect 20852 4936 20861 4976
rect 0 4916 90 4936
rect 2860 4808 2900 4936
rect 13036 4892 13076 4936
rect 20812 4892 20852 4936
rect 12643 4852 12652 4892
rect 12692 4852 12844 4892
rect 12884 4852 12893 4892
rect 13018 4852 13027 4892
rect 13067 4852 16396 4892
rect 16436 4852 16445 4892
rect 20812 4852 21196 4892
rect 21236 4852 21245 4892
rect 21292 4808 21332 5020
rect 27139 4936 27148 4976
rect 27188 4936 28916 4976
rect 22444 4892 22484 4901
rect 28876 4892 28916 4936
rect 22313 4852 22444 4892
rect 22484 4852 22493 4892
rect 23011 4852 23020 4892
rect 23060 4852 23308 4892
rect 23348 4852 23357 4892
rect 23482 4852 23491 4892
rect 23531 4852 24844 4892
rect 24884 4852 25324 4892
rect 25364 4852 25373 4892
rect 27497 4852 27628 4892
rect 27668 4852 27677 4892
rect 33100 4892 33140 5020
rect 34540 4976 34580 5608
rect 43372 5564 43412 5608
rect 46278 5588 46368 5608
rect 34627 5524 34636 5564
rect 34676 5524 43412 5564
rect 44755 5440 44764 5480
rect 44804 5440 46252 5480
rect 46292 5440 46301 5480
rect 46278 5312 46368 5332
rect 46243 5272 46252 5312
rect 46292 5272 46368 5312
rect 46278 5252 46368 5272
rect 46278 4976 46368 4996
rect 34540 4936 34732 4976
rect 34772 4936 35020 4976
rect 35060 4936 35308 4976
rect 35348 4936 35500 4976
rect 35540 4936 35549 4976
rect 41827 4936 41836 4976
rect 41876 4936 44524 4976
rect 44564 4936 44573 4976
rect 44777 4936 44908 4976
rect 44948 4936 44957 4976
rect 45139 4936 45148 4976
rect 45188 4936 46368 4976
rect 46278 4916 46368 4936
rect 33100 4852 39820 4892
rect 39860 4852 39869 4892
rect 22444 4843 22484 4852
rect 28876 4843 28916 4852
rect 2860 4768 21332 4808
rect 22540 4768 28052 4808
rect 22540 4724 22580 4768
rect 28012 4724 28052 4768
rect 28972 4768 44332 4808
rect 44372 4768 44381 4808
rect 28972 4724 29012 4768
rect 12931 4684 12940 4724
rect 12980 4684 13132 4724
rect 13172 4684 13181 4724
rect 21043 4684 21052 4724
rect 21092 4684 22580 4724
rect 22627 4684 22636 4724
rect 22676 4684 23212 4724
rect 23252 4684 23261 4724
rect 23395 4684 23404 4724
rect 23444 4684 24076 4724
rect 24116 4684 24125 4724
rect 28012 4684 29012 4724
rect 44755 4684 44764 4724
rect 44804 4684 44813 4724
rect 0 4640 90 4660
rect 44764 4640 44804 4684
rect 46278 4640 46368 4660
rect 0 4600 38956 4640
rect 38996 4600 39005 4640
rect 44764 4600 46368 4640
rect 0 4580 90 4600
rect 46278 4580 46368 4600
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 20524 4516 23788 4556
rect 23828 4516 23837 4556
rect 23971 4516 23980 4556
rect 24020 4516 24692 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 20524 4388 20564 4516
rect 12115 4348 12124 4388
rect 12164 4348 13804 4388
rect 13844 4348 13853 4388
rect 17356 4348 17780 4388
rect 0 4304 90 4324
rect 17356 4304 17396 4348
rect 17740 4304 17780 4348
rect 18700 4348 20564 4388
rect 22732 4348 23020 4388
rect 23060 4348 23069 4388
rect 23299 4348 23308 4388
rect 23348 4348 24212 4388
rect 18700 4304 18740 4348
rect 22732 4304 22772 4348
rect 0 4264 1420 4304
rect 1460 4264 1469 4304
rect 12835 4264 12844 4304
rect 12884 4264 13268 4304
rect 13507 4264 13516 4304
rect 13556 4264 15148 4304
rect 15188 4264 15197 4304
rect 15340 4264 15532 4304
rect 15572 4264 15820 4304
rect 15860 4264 17396 4304
rect 17513 4264 17596 4304
rect 17636 4264 17644 4304
rect 17684 4264 17693 4304
rect 17740 4264 18740 4304
rect 19267 4264 19276 4304
rect 19316 4264 19325 4304
rect 22252 4264 22772 4304
rect 23203 4264 23212 4304
rect 23252 4264 23491 4304
rect 23531 4264 23540 4304
rect 23683 4264 23692 4304
rect 23732 4264 23980 4304
rect 24020 4264 24029 4304
rect 0 4244 90 4264
rect 13228 4220 13268 4264
rect 15340 4220 15380 4264
rect 19276 4220 19316 4264
rect 22252 4220 22292 4264
rect 22732 4220 22772 4264
rect 24172 4220 24212 4348
rect 24652 4220 24692 4516
rect 46278 4304 46368 4324
rect 25027 4264 25036 4304
rect 25076 4264 40916 4304
rect 45139 4264 45148 4304
rect 45188 4264 46368 4304
rect 11779 4180 11788 4220
rect 11828 4180 12643 4220
rect 12692 4180 12701 4220
rect 12931 4180 12940 4220
rect 12980 4180 12989 4220
rect 13121 4180 13130 4220
rect 13170 4180 13179 4220
rect 13228 4180 13247 4220
rect 13287 4180 13296 4220
rect 13411 4180 13420 4220
rect 13460 4180 13591 4220
rect 14092 4180 15095 4220
rect 15135 4180 15144 4220
rect 15331 4180 15340 4220
rect 15380 4180 15389 4220
rect 17356 4180 17836 4220
rect 17876 4180 17885 4220
rect 18953 4180 19084 4220
rect 19124 4180 19133 4220
rect 19276 4180 22156 4220
rect 22196 4180 22243 4220
rect 22283 4180 22292 4220
rect 22409 4180 22540 4220
rect 22580 4180 22589 4220
rect 22714 4180 22723 4220
rect 22763 4180 22772 4220
rect 22868 4180 22924 4220
rect 22964 4180 22999 4220
rect 23039 4180 23048 4220
rect 23155 4180 23164 4220
rect 23204 4180 23213 4220
rect 23369 4180 23404 4220
rect 23444 4180 23500 4220
rect 23540 4180 23549 4220
rect 23657 4180 23788 4220
rect 23828 4180 23837 4220
rect 24163 4180 24172 4220
rect 24212 4180 24221 4220
rect 24268 4180 24355 4220
rect 24395 4180 24404 4220
rect 24562 4180 24571 4220
rect 24611 4180 24692 4220
rect 24739 4180 24748 4220
rect 24788 4180 24797 4220
rect 35875 4180 35884 4220
rect 35924 4180 38284 4220
rect 38324 4180 38333 4220
rect 38380 4180 40300 4220
rect 40340 4180 40349 4220
rect 11875 4096 11884 4136
rect 11924 4096 11933 4136
rect 12137 4096 12268 4136
rect 12308 4096 12317 4136
rect 12451 4096 12460 4136
rect 12500 4096 12508 4136
rect 12548 4096 12631 4136
rect 11884 4052 11924 4096
rect 12940 4052 12980 4180
rect 13132 4136 13172 4180
rect 13123 4096 13132 4136
rect 13172 4096 13217 4136
rect 13481 4096 13612 4136
rect 13652 4096 13661 4136
rect 14092 4052 14132 4180
rect 17356 4136 17396 4180
rect 19084 4162 19124 4171
rect 23164 4136 23204 4180
rect 24019 4138 24028 4178
rect 24068 4138 24077 4178
rect 14947 4096 14956 4136
rect 14996 4096 15235 4136
rect 15275 4096 15284 4136
rect 15427 4096 15436 4136
rect 15476 4096 15607 4136
rect 16003 4096 16012 4136
rect 16052 4096 17356 4136
rect 17396 4096 17405 4136
rect 23116 4096 23204 4136
rect 23290 4096 23299 4136
rect 23339 4096 23348 4136
rect 23395 4096 23404 4136
rect 23444 4096 23907 4136
rect 23947 4096 23956 4136
rect 23116 4052 23156 4096
rect 23308 4052 23348 4096
rect 24028 4052 24068 4138
rect 24268 4136 24308 4180
rect 24748 4136 24788 4180
rect 38380 4136 38420 4180
rect 40876 4136 40916 4264
rect 46278 4244 46368 4264
rect 41059 4180 41068 4220
rect 41108 4180 43220 4220
rect 44611 4180 44620 4220
rect 44660 4180 44948 4220
rect 43180 4136 43220 4180
rect 44908 4136 44948 4180
rect 24259 4096 24268 4136
rect 24308 4096 24317 4136
rect 24460 4096 24788 4136
rect 27619 4096 27628 4136
rect 27668 4096 27724 4136
rect 27764 4096 27799 4136
rect 33161 4096 33292 4136
rect 33332 4096 33341 4136
rect 33523 4096 33532 4136
rect 33572 4096 38420 4136
rect 38563 4096 38572 4136
rect 38612 4096 38621 4136
rect 38755 4096 38764 4136
rect 38804 4096 40492 4136
rect 40532 4096 40541 4136
rect 40867 4096 40876 4136
rect 40916 4096 40925 4136
rect 41129 4096 41260 4136
rect 41300 4096 41309 4136
rect 41993 4096 42124 4136
rect 42164 4096 42173 4136
rect 43180 4096 44524 4136
rect 44564 4096 44573 4136
rect 44899 4096 44908 4136
rect 44948 4096 44957 4136
rect 24460 4052 24500 4096
rect 38572 4052 38612 4096
rect 11884 4012 12980 4052
rect 13315 4012 13324 4052
rect 13364 4012 14132 4052
rect 14755 4012 14764 4052
rect 14804 4012 21196 4052
rect 21236 4012 21245 4052
rect 22531 4012 22540 4052
rect 22580 4012 22924 4052
rect 22964 4012 22973 4052
rect 23107 4012 23116 4052
rect 23156 4012 23165 4052
rect 23308 4012 23788 4052
rect 23828 4012 23837 4052
rect 23971 4012 23980 4052
rect 24020 4012 24068 4052
rect 24346 4012 24355 4052
rect 24395 4012 24500 4052
rect 27331 4012 27340 4052
rect 27380 4012 38612 4052
rect 40003 4012 40012 4052
rect 40052 4012 40252 4052
rect 40292 4012 40301 4052
rect 40483 4012 40492 4052
rect 40532 4012 40636 4052
rect 40676 4012 40685 4052
rect 40771 4012 40780 4052
rect 40820 4012 41020 4052
rect 41060 4012 41069 4052
rect 44755 4012 44764 4052
rect 44804 4012 45620 4052
rect 0 3968 90 3988
rect 12940 3968 12980 4012
rect 45580 3968 45620 4012
rect 46278 3968 46368 3988
rect 0 3928 1420 3968
rect 1460 3928 1469 3968
rect 12940 3928 13708 3968
rect 13748 3928 13757 3968
rect 13843 3928 13852 3968
rect 13892 3928 16588 3968
rect 16628 3928 16637 3968
rect 20131 3928 20140 3968
rect 20180 3928 21292 3968
rect 21332 3928 21341 3968
rect 23011 3928 23020 3968
rect 23060 3928 23596 3968
rect 23636 3928 23645 3968
rect 24547 3928 24556 3968
rect 24596 3928 25132 3968
rect 25172 3928 25181 3968
rect 25891 3928 25900 3968
rect 25940 3928 27244 3968
rect 27284 3928 27293 3968
rect 27955 3928 27964 3968
rect 28004 3928 36020 3968
rect 36067 3928 36076 3968
rect 36116 3928 38332 3968
rect 38372 3928 38381 3968
rect 38467 3928 38476 3968
rect 38516 3928 40684 3968
rect 40724 3928 40733 3968
rect 42355 3928 42364 3968
rect 42404 3928 44908 3968
rect 44948 3928 44957 3968
rect 45580 3928 46368 3968
rect 0 3908 90 3928
rect 9772 3844 35884 3884
rect 35924 3844 35933 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 0 3632 90 3652
rect 9772 3632 9812 3844
rect 35980 3800 36020 3928
rect 46278 3908 46368 3928
rect 36163 3844 36172 3884
rect 36212 3844 38668 3884
rect 38708 3844 38717 3884
rect 12163 3760 12172 3800
rect 12212 3760 14188 3800
rect 14228 3760 14237 3800
rect 14371 3760 14380 3800
rect 14420 3760 16396 3800
rect 16436 3760 16445 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 19276 3760 33140 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 35980 3760 37420 3800
rect 37460 3760 37469 3800
rect 39436 3760 45004 3800
rect 45044 3760 45053 3800
rect 19276 3716 19316 3760
rect 33100 3716 33140 3760
rect 0 3592 1228 3632
rect 1268 3592 1277 3632
rect 8947 3592 8956 3632
rect 8996 3592 9812 3632
rect 9868 3676 19316 3716
rect 23369 3676 23500 3716
rect 23540 3676 24500 3716
rect 25027 3676 25036 3716
rect 25076 3676 29260 3716
rect 29300 3676 29309 3716
rect 33100 3676 39340 3716
rect 39380 3676 39389 3716
rect 0 3572 90 3592
rect 9868 3548 9908 3676
rect 10915 3592 10924 3632
rect 10964 3592 11548 3632
rect 11588 3592 11597 3632
rect 12940 3592 13516 3632
rect 13556 3592 13565 3632
rect 13699 3592 13708 3632
rect 13748 3592 23020 3632
rect 23060 3592 23069 3632
rect 2860 3508 9908 3548
rect 2860 3464 2900 3508
rect 12940 3464 12980 3592
rect 14860 3508 15148 3548
rect 15188 3508 16204 3548
rect 16244 3508 16253 3548
rect 16387 3508 16396 3548
rect 16436 3508 23116 3548
rect 23156 3508 23165 3548
rect 172 3424 2900 3464
rect 8585 3424 8716 3464
rect 8756 3424 8765 3464
rect 9257 3424 9388 3464
rect 9428 3424 9437 3464
rect 11779 3424 11788 3464
rect 11828 3424 12556 3464
rect 12596 3424 12980 3464
rect 13132 3424 14092 3464
rect 14132 3424 14141 3464
rect 14284 3424 14380 3464
rect 14420 3424 14429 3464
rect 14633 3424 14755 3464
rect 14804 3424 14813 3464
rect 0 3296 90 3316
rect 172 3296 212 3424
rect 9388 3380 9428 3424
rect 11020 3380 11060 3389
rect 13132 3380 13172 3424
rect 14284 3380 14324 3424
rect 14860 3380 14900 3508
rect 14947 3424 14956 3464
rect 14996 3424 15127 3464
rect 15811 3424 15820 3464
rect 15860 3424 15869 3464
rect 16396 3424 19276 3464
rect 19316 3424 19325 3464
rect 21187 3424 21196 3464
rect 21236 3424 21244 3464
rect 21284 3424 21367 3464
rect 21475 3424 21484 3464
rect 21524 3424 21655 3464
rect 21833 3424 21868 3464
rect 21908 3424 21964 3464
rect 22004 3424 22013 3464
rect 22060 3424 22156 3464
rect 22196 3424 22205 3464
rect 22505 3424 22636 3464
rect 22676 3424 22685 3464
rect 9388 3340 9772 3380
rect 9812 3340 9821 3380
rect 10889 3340 11020 3380
rect 11060 3340 11069 3380
rect 11779 3340 11788 3380
rect 11828 3340 12067 3380
rect 12107 3340 12116 3380
rect 12163 3340 12172 3380
rect 12212 3340 12343 3380
rect 12521 3340 12652 3380
rect 12692 3340 12701 3380
rect 13411 3340 13420 3380
rect 13460 3340 13620 3380
rect 13660 3340 13669 3380
rect 13978 3340 13987 3380
rect 14027 3340 14036 3380
rect 14275 3340 14284 3380
rect 14324 3340 14333 3380
rect 14380 3340 14615 3380
rect 14655 3340 14664 3380
rect 14851 3340 14860 3380
rect 14900 3340 14909 3380
rect 15043 3340 15052 3380
rect 15092 3340 15244 3380
rect 15284 3340 15293 3380
rect 15418 3340 15427 3380
rect 15476 3340 15607 3380
rect 11020 3331 11060 3340
rect 13132 3331 13172 3340
rect 13996 3296 14036 3340
rect 14380 3296 14420 3340
rect 15820 3296 15860 3424
rect 16396 3380 16436 3424
rect 22060 3380 22100 3424
rect 23212 3380 23252 3389
rect 16265 3340 16396 3380
rect 16436 3340 16445 3380
rect 17548 3340 17604 3380
rect 17644 3340 17653 3380
rect 17731 3340 17740 3380
rect 17780 3340 20812 3380
rect 20852 3340 20861 3380
rect 20908 3340 21772 3380
rect 21812 3340 21821 3380
rect 22060 3340 22126 3380
rect 22166 3340 22175 3380
rect 22243 3340 22252 3380
rect 22292 3340 22301 3380
rect 22601 3340 22732 3380
rect 22772 3340 22781 3380
rect 23500 3380 23540 3676
rect 23971 3592 23980 3632
rect 24020 3592 24076 3632
rect 24116 3592 24151 3632
rect 23587 3424 23596 3464
rect 23636 3424 24212 3464
rect 24172 3380 24212 3424
rect 24460 3380 24500 3676
rect 24809 3592 24892 3632
rect 24932 3592 24940 3632
rect 24980 3592 24989 3632
rect 25603 3592 25612 3632
rect 25652 3592 27436 3632
rect 27476 3592 27485 3632
rect 29059 3592 29068 3632
rect 29108 3592 37996 3632
rect 38036 3592 38045 3632
rect 38659 3592 38668 3632
rect 38708 3592 38716 3632
rect 38756 3592 38839 3632
rect 39436 3548 39476 3760
rect 46278 3632 46368 3652
rect 40531 3592 40540 3632
rect 40580 3592 44564 3632
rect 45139 3592 45148 3632
rect 45188 3592 46368 3632
rect 24739 3508 24748 3548
rect 24788 3508 25172 3548
rect 25843 3508 25852 3548
rect 25892 3508 39476 3548
rect 42355 3508 42364 3548
rect 42404 3508 44140 3548
rect 44180 3508 44189 3548
rect 25132 3464 25172 3508
rect 44524 3464 44564 3592
rect 46278 3572 46368 3592
rect 24713 3424 24748 3464
rect 24788 3424 24844 3464
rect 24884 3424 24893 3464
rect 25123 3424 25132 3464
rect 25172 3424 25181 3464
rect 25481 3424 25612 3464
rect 25652 3424 25661 3464
rect 25978 3424 25987 3464
rect 26027 3424 26036 3464
rect 36355 3424 36364 3464
rect 36404 3424 37852 3464
rect 37892 3424 37901 3464
rect 37987 3424 37996 3464
rect 38036 3424 38092 3464
rect 38132 3424 38167 3464
rect 38345 3424 38476 3464
rect 38516 3424 38525 3464
rect 38947 3424 38956 3464
rect 38996 3424 39005 3464
rect 39331 3424 39340 3464
rect 39380 3424 39436 3464
rect 39476 3424 39724 3464
rect 39764 3424 40012 3464
rect 40052 3424 40300 3464
rect 40340 3424 40349 3464
rect 40745 3424 40876 3464
rect 40916 3424 40925 3464
rect 41347 3424 41356 3464
rect 41396 3424 41405 3464
rect 41609 3424 41740 3464
rect 41780 3424 41789 3464
rect 41993 3424 42124 3464
rect 42164 3424 42173 3464
rect 42377 3424 42508 3464
rect 42548 3424 42557 3464
rect 42691 3424 42700 3464
rect 42740 3424 42892 3464
rect 42932 3424 42941 3464
rect 44515 3424 44524 3464
rect 44564 3424 44573 3464
rect 44777 3424 44812 3464
rect 44852 3424 44908 3464
rect 44948 3424 44957 3464
rect 25996 3380 26036 3424
rect 23500 3340 23700 3380
rect 23740 3340 23749 3380
rect 23945 3340 24076 3380
rect 24116 3340 24125 3380
rect 24172 3340 24191 3380
rect 24231 3340 24240 3380
rect 24355 3340 24364 3380
rect 24404 3340 26036 3380
rect 26188 3380 26228 3389
rect 38956 3380 38996 3424
rect 26228 3340 27148 3380
rect 27188 3340 27197 3380
rect 27305 3340 27436 3380
rect 27476 3340 27485 3380
rect 28012 3340 38996 3380
rect 16396 3331 16436 3340
rect 0 3256 212 3296
rect 2083 3256 2092 3296
rect 2132 3256 2900 3296
rect 11203 3256 11212 3296
rect 11252 3256 12116 3296
rect 13507 3256 13516 3296
rect 13556 3256 14036 3296
rect 14179 3256 14188 3296
rect 14228 3256 14420 3296
rect 15244 3256 15860 3296
rect 16051 3256 16060 3296
rect 16100 3256 16300 3296
rect 16340 3256 16349 3296
rect 0 3236 90 3256
rect 2860 3128 2900 3256
rect 12076 3212 12116 3256
rect 9619 3172 9628 3212
rect 9668 3172 10060 3212
rect 10100 3172 10109 3212
rect 12076 3172 13420 3212
rect 13460 3172 13469 3212
rect 13795 3172 13804 3212
rect 13844 3172 14956 3212
rect 14996 3172 15005 3212
rect 15244 3128 15284 3256
rect 15820 3212 15860 3256
rect 17548 3212 17588 3340
rect 20908 3296 20948 3340
rect 22252 3296 22292 3340
rect 23212 3296 23252 3340
rect 26188 3331 26228 3340
rect 17923 3256 17932 3296
rect 17972 3256 20948 3296
rect 21475 3256 21484 3296
rect 21524 3256 22292 3296
rect 22348 3256 22964 3296
rect 23212 3256 23788 3296
rect 23828 3256 23837 3296
rect 24355 3256 24364 3296
rect 24404 3256 24508 3296
rect 24548 3256 24557 3296
rect 15331 3172 15340 3212
rect 15380 3172 15628 3212
rect 15668 3172 15677 3212
rect 15820 3172 17588 3212
rect 17644 3172 21628 3212
rect 21668 3172 21677 3212
rect 2860 3088 15284 3128
rect 15427 3088 15436 3128
rect 15476 3088 17548 3128
rect 17588 3088 17597 3128
rect 17644 3044 17684 3172
rect 22348 3128 22388 3256
rect 17731 3088 17740 3128
rect 17780 3088 22388 3128
rect 22924 3128 22964 3256
rect 23875 3172 23884 3212
rect 23924 3172 24268 3212
rect 24308 3172 24317 3212
rect 28012 3128 28052 3340
rect 31843 3256 31852 3296
rect 31892 3256 40636 3296
rect 40676 3256 40685 3296
rect 33091 3172 33100 3212
rect 33140 3172 38236 3212
rect 38276 3172 38285 3212
rect 22924 3088 28052 3128
rect 33100 3088 38476 3128
rect 38516 3088 38525 3128
rect 33100 3044 33140 3088
rect 41356 3044 41396 3424
rect 42604 3340 44428 3380
rect 44468 3340 44477 3380
rect 42604 3296 42644 3340
rect 46278 3296 46368 3316
rect 41971 3256 41980 3296
rect 42020 3256 42644 3296
rect 42739 3256 42748 3296
rect 42788 3256 43756 3296
rect 43796 3256 43805 3296
rect 44755 3256 44764 3296
rect 44804 3256 46368 3296
rect 46278 3236 46368 3256
rect 41587 3172 41596 3212
rect 41636 3172 41876 3212
rect 43123 3172 43132 3212
rect 43172 3172 43372 3212
rect 43412 3172 43421 3212
rect 41836 3128 41876 3172
rect 41836 3088 44524 3128
rect 44564 3088 44573 3128
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 12643 3004 12652 3044
rect 12692 3004 13804 3044
rect 13844 3004 13853 3044
rect 15619 3004 15628 3044
rect 15668 3004 17684 3044
rect 17827 3004 17836 3044
rect 17876 3004 19948 3044
rect 19988 3004 19997 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 24739 3004 24748 3044
rect 24788 3004 33140 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 35788 3004 41396 3044
rect 0 2960 90 2980
rect 35788 2960 35828 3004
rect 46278 2960 46368 2980
rect 0 2920 1460 2960
rect 15811 2920 15820 2960
rect 15860 2920 22732 2960
rect 22772 2920 22781 2960
rect 24451 2920 24460 2960
rect 24500 2920 35828 2960
rect 40108 2920 40300 2960
rect 40340 2920 40349 2960
rect 45484 2920 46368 2960
rect 0 2900 90 2920
rect 1420 2876 1460 2920
rect 40108 2876 40148 2920
rect 45484 2876 45524 2920
rect 46278 2900 46368 2920
rect 1420 2836 33140 2876
rect 38899 2836 38908 2876
rect 38948 2836 39148 2876
rect 39188 2836 39197 2876
rect 40090 2836 40099 2876
rect 40139 2836 40300 2876
rect 40340 2836 40588 2876
rect 40628 2836 40876 2876
rect 40916 2836 41164 2876
rect 41204 2836 41452 2876
rect 41492 2836 41731 2876
rect 41771 2836 41780 2876
rect 45139 2836 45148 2876
rect 45188 2836 45524 2876
rect 10531 2752 10540 2792
rect 10580 2752 11788 2792
rect 11828 2752 11837 2792
rect 11971 2752 11980 2792
rect 12020 2752 12028 2792
rect 12068 2752 12151 2792
rect 12761 2752 12844 2792
rect 12884 2752 12892 2792
rect 12932 2752 12941 2792
rect 13411 2752 13420 2792
rect 13460 2752 13652 2792
rect 13786 2752 13795 2792
rect 13835 2752 14764 2792
rect 14804 2752 14813 2792
rect 14921 2752 15052 2792
rect 15092 2752 15101 2792
rect 20611 2752 20620 2792
rect 20660 2752 22684 2792
rect 22724 2752 22733 2792
rect 23273 2752 23395 2792
rect 23444 2752 23453 2792
rect 11788 2708 11828 2752
rect 13612 2708 13652 2752
rect 33100 2708 33140 2836
rect 34819 2752 34828 2792
rect 34868 2752 39292 2792
rect 39332 2752 39341 2792
rect 42739 2752 42748 2792
rect 42788 2752 44948 2792
rect 8707 2668 8716 2708
rect 8756 2668 9100 2708
rect 9140 2668 9149 2708
rect 10348 2699 11020 2708
rect 10388 2668 11020 2699
rect 11060 2668 11069 2708
rect 11788 2668 13483 2708
rect 13556 2668 13565 2708
rect 13612 2668 13708 2708
rect 13748 2668 13757 2708
rect 14825 2668 14956 2708
rect 14996 2668 15005 2708
rect 15139 2668 15148 2708
rect 15188 2668 15319 2708
rect 15715 2668 15724 2708
rect 15764 2668 22540 2708
rect 22580 2668 22589 2708
rect 23011 2668 23020 2708
rect 23060 2668 23063 2708
rect 23103 2668 23191 2708
rect 23299 2668 23308 2708
rect 23349 2668 23479 2708
rect 23683 2668 23692 2708
rect 23732 2668 24212 2708
rect 33100 2668 42548 2708
rect 10348 2650 10388 2659
rect 0 2624 90 2644
rect 24172 2624 24212 2668
rect 42508 2624 42548 2668
rect 44908 2624 44948 2752
rect 46278 2624 46368 2644
rect 0 2584 8908 2624
rect 8948 2584 8957 2624
rect 12137 2584 12172 2624
rect 12212 2584 12268 2624
rect 12308 2584 12317 2624
rect 12521 2584 12652 2624
rect 12692 2584 12701 2624
rect 13481 2584 13603 2624
rect 13652 2584 13661 2624
rect 14057 2584 14092 2624
rect 14132 2584 14188 2624
rect 14228 2584 14237 2624
rect 14345 2584 14476 2624
rect 14516 2584 14525 2624
rect 14707 2584 14716 2624
rect 14756 2584 18124 2624
rect 18164 2584 18173 2624
rect 22531 2584 22540 2624
rect 22580 2584 22636 2624
rect 22676 2584 22711 2624
rect 22819 2584 22828 2624
rect 22868 2584 22924 2624
rect 22964 2584 22999 2624
rect 23165 2584 23203 2624
rect 23243 2584 23252 2624
rect 23779 2584 23788 2624
rect 23828 2584 23837 2624
rect 24163 2584 24172 2624
rect 24212 2584 24221 2624
rect 39139 2584 39148 2624
rect 39188 2584 39244 2624
rect 39284 2584 39319 2624
rect 39523 2584 39532 2624
rect 39572 2584 39581 2624
rect 42115 2584 42124 2624
rect 42164 2584 42173 2624
rect 42499 2584 42508 2624
rect 42548 2584 42557 2624
rect 44131 2584 44140 2624
rect 44180 2584 44189 2624
rect 44393 2584 44524 2624
rect 44564 2584 44573 2624
rect 44899 2584 44908 2624
rect 44948 2584 44957 2624
rect 45772 2584 46368 2624
rect 0 2564 90 2584
rect 13612 2540 13652 2584
rect 23212 2540 23252 2584
rect 23788 2540 23828 2584
rect 39532 2540 39572 2584
rect 13612 2500 15820 2540
rect 15860 2500 15869 2540
rect 20995 2500 21004 2540
rect 21044 2500 22484 2540
rect 22531 2500 22540 2540
rect 22580 2500 23156 2540
rect 23203 2500 23212 2540
rect 23252 2500 23261 2540
rect 23788 2500 24172 2540
rect 24212 2500 24221 2540
rect 39139 2500 39148 2540
rect 39188 2500 39572 2540
rect 22444 2456 22484 2500
rect 2860 2416 8812 2456
rect 8852 2416 8861 2456
rect 11683 2416 11692 2456
rect 11732 2416 13948 2456
rect 13988 2416 13997 2456
rect 17740 2416 22300 2456
rect 22340 2416 22349 2456
rect 22444 2416 23020 2456
rect 23060 2416 23069 2456
rect 0 2288 90 2308
rect 2860 2288 2900 2416
rect 4108 2332 15436 2372
rect 15476 2332 15485 2372
rect 0 2248 2900 2288
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 0 2228 90 2248
rect 4108 2120 4148 2332
rect 17740 2288 17780 2416
rect 23116 2372 23156 2500
rect 23299 2416 23308 2456
rect 23348 2416 23548 2456
rect 23588 2416 23597 2456
rect 23692 2416 23932 2456
rect 23972 2416 23981 2456
rect 28012 2416 38956 2456
rect 38996 2416 39005 2456
rect 23692 2372 23732 2416
rect 23116 2332 23732 2372
rect 1747 2080 1756 2120
rect 1796 2080 4148 2120
rect 5164 2248 12556 2288
rect 12596 2248 12605 2288
rect 13219 2248 13228 2288
rect 13268 2248 17780 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 0 1952 90 1972
rect 5164 1952 5204 2248
rect 28012 2204 28052 2416
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 6892 2164 17452 2204
rect 17492 2164 17501 2204
rect 22147 2164 22156 2204
rect 22196 2164 28052 2204
rect 6892 1952 6932 2164
rect 8236 2080 25132 2120
rect 25172 2080 25181 2120
rect 25603 2080 25612 2120
rect 25652 2080 39244 2120
rect 39284 2080 39293 2120
rect 0 1912 212 1952
rect 1385 1912 1420 1952
rect 1460 1912 1516 1952
rect 1556 1912 1565 1952
rect 3427 1912 3436 1952
rect 3476 1912 3485 1952
rect 5155 1912 5164 1952
rect 5204 1912 5213 1952
rect 6883 1912 6892 1952
rect 6932 1912 6941 1952
rect 0 1892 90 1912
rect 172 1784 212 1912
rect 3436 1868 3476 1912
rect 8236 1868 8276 2080
rect 8620 1996 30700 2036
rect 30740 1996 30749 2036
rect 8620 1952 8660 1996
rect 42124 1952 42164 2584
rect 44140 2540 44180 2584
rect 45772 2540 45812 2584
rect 46278 2564 46368 2584
rect 42355 2500 42364 2540
rect 42404 2500 44180 2540
rect 44755 2500 44764 2540
rect 44804 2500 45812 2540
rect 44371 2416 44380 2456
rect 44420 2416 45044 2456
rect 45004 1952 45044 2416
rect 46278 2288 46368 2308
rect 45580 2248 46368 2288
rect 45580 2120 45620 2248
rect 46278 2228 46368 2248
rect 45139 2080 45148 2120
rect 45188 2080 45620 2120
rect 46278 1952 46368 1972
rect 8611 1912 8620 1952
rect 8660 1912 8669 1952
rect 8716 1912 42164 1952
rect 43241 1912 43372 1952
rect 43412 1912 43421 1952
rect 43625 1912 43756 1952
rect 43796 1912 43805 1952
rect 44009 1912 44140 1952
rect 44180 1912 44189 1952
rect 44419 1912 44428 1952
rect 44468 1912 44524 1952
rect 44564 1912 44599 1952
rect 44777 1912 44908 1952
rect 44948 1912 44957 1952
rect 45004 1912 46368 1952
rect 3436 1828 8276 1868
rect 8716 1784 8756 1912
rect 46278 1892 46368 1912
rect 8899 1828 8908 1868
rect 8948 1828 24460 1868
rect 24500 1828 24509 1868
rect 172 1744 8756 1784
rect 8803 1744 8812 1784
rect 8852 1744 24652 1784
rect 24692 1744 24701 1784
rect 43987 1744 43996 1784
rect 44036 1744 45580 1784
rect 45620 1744 45629 1784
rect 3065 1660 3148 1700
rect 3188 1660 3196 1700
rect 3236 1660 3245 1700
rect 4771 1660 4780 1700
rect 4820 1660 4924 1700
rect 4964 1660 4973 1700
rect 6521 1660 6604 1700
rect 6644 1660 6652 1700
rect 6692 1660 6701 1700
rect 8249 1660 8332 1700
rect 8372 1660 8380 1700
rect 8420 1660 8429 1700
rect 43603 1660 43612 1700
rect 43652 1660 44276 1700
rect 44371 1660 44380 1700
rect 44420 1660 44620 1700
rect 44660 1660 44669 1700
rect 44755 1660 44764 1700
rect 44804 1660 45044 1700
rect 0 1616 90 1636
rect 0 1576 41740 1616
rect 41780 1576 41789 1616
rect 0 1556 90 1576
rect 44236 1532 44276 1660
rect 45004 1616 45044 1660
rect 46278 1616 46368 1636
rect 45004 1576 46368 1616
rect 46278 1556 46368 1576
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 44236 1492 46196 1532
rect 46156 1448 46196 1492
rect 46156 1408 46252 1448
rect 46292 1408 46301 1448
rect 0 1280 90 1300
rect 46278 1280 46368 1300
rect 0 1240 42700 1280
rect 42740 1240 42749 1280
rect 46243 1240 46252 1280
rect 46292 1240 46368 1280
rect 0 1220 90 1240
rect 46278 1220 46368 1240
rect 0 944 90 964
rect 46278 944 46368 964
rect 0 904 42508 944
rect 42548 904 42557 944
rect 45571 904 45580 944
rect 45620 904 46368 944
rect 0 884 90 904
rect 46278 884 46368 904
rect 0 608 90 628
rect 46278 608 46368 628
rect 0 568 42124 608
rect 42164 568 42173 608
rect 44611 568 44620 608
rect 44660 568 46368 608
rect 0 548 90 568
rect 46278 548 46368 568
rect 13507 148 13516 188
rect 13556 148 41260 188
rect 41300 148 41309 188
rect 10051 64 10060 104
rect 10100 64 40876 104
rect 40916 64 40925 104
<< via2 >>
rect 1420 10984 1460 11024
rect 44236 10984 44276 11024
rect 1132 10648 1172 10688
rect 43756 10648 43796 10688
rect 1036 10312 1076 10352
rect 43276 10312 43316 10352
rect 16108 10228 16148 10268
rect 16876 10144 16916 10184
rect 2956 10060 2996 10100
rect 10060 10060 10100 10100
rect 10252 10060 10292 10100
rect 11212 10060 11252 10100
rect 12940 10060 12980 10100
rect 13036 10060 13076 10100
rect 14188 10060 14228 10100
rect 16396 10060 16436 10100
rect 22252 10060 22292 10100
rect 27916 10060 27956 10100
rect 42892 10060 42932 10100
rect 1420 9976 1460 10016
rect 2764 9976 2804 10016
rect 9388 9976 9428 10016
rect 13996 9976 14036 10016
rect 16012 9976 16052 10016
rect 1132 9892 1172 9932
rect 12460 9892 12500 9932
rect 15916 9892 15956 9932
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 10060 9808 10100 9848
rect 12652 9808 12692 9848
rect 15052 9808 15092 9848
rect 15340 9808 15380 9848
rect 22828 9976 22868 10016
rect 23404 9976 23444 10016
rect 26956 9976 26996 10016
rect 27820 9976 27860 10016
rect 31468 9976 31508 10016
rect 33580 9976 33620 10016
rect 40492 9976 40532 10016
rect 23596 9892 23636 9932
rect 26284 9892 26324 9932
rect 33388 9892 33428 9932
rect 39244 9892 39284 9932
rect 11308 9724 11348 9764
rect 12844 9724 12884 9764
rect 14956 9724 14996 9764
rect 15628 9724 15668 9764
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 23788 9808 23828 9848
rect 28972 9808 29012 9848
rect 29452 9808 29492 9848
rect 29740 9808 29780 9848
rect 10252 9640 10292 9680
rect 11788 9640 11828 9680
rect 13420 9640 13460 9680
rect 9292 9556 9332 9596
rect 12940 9556 12980 9596
rect 1228 9472 1268 9512
rect 2764 9472 2804 9512
rect 9388 9472 9428 9512
rect 10156 9472 10196 9512
rect 10540 9472 10580 9512
rect 10924 9472 10964 9512
rect 11692 9472 11732 9512
rect 1036 9388 1076 9428
rect 4108 9388 4148 9428
rect 10828 9388 10868 9428
rect 11500 9388 11540 9428
rect 13996 9640 14036 9680
rect 16300 9640 16340 9680
rect 17932 9724 17972 9764
rect 18412 9724 18452 9764
rect 22060 9724 22100 9764
rect 23116 9724 23156 9764
rect 25132 9724 25172 9764
rect 25420 9724 25460 9764
rect 25804 9724 25844 9764
rect 28876 9724 28916 9764
rect 29932 9724 29972 9764
rect 17452 9640 17492 9680
rect 18316 9640 18356 9680
rect 19468 9640 19508 9680
rect 20236 9640 20276 9680
rect 21196 9640 21236 9680
rect 24844 9640 24884 9680
rect 13804 9556 13844 9596
rect 18604 9556 18644 9596
rect 19852 9556 19892 9596
rect 21388 9556 21428 9596
rect 21772 9556 21812 9596
rect 22156 9556 22196 9596
rect 22348 9556 22388 9596
rect 23500 9556 23540 9596
rect 23692 9556 23732 9596
rect 23884 9556 23924 9596
rect 24460 9556 24500 9596
rect 24652 9556 24692 9596
rect 26284 9640 26324 9680
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 37420 9808 37460 9848
rect 41644 9808 41684 9848
rect 31948 9724 31988 9764
rect 32716 9724 32756 9764
rect 28492 9640 28532 9680
rect 31180 9640 31220 9680
rect 31564 9640 31604 9680
rect 28300 9556 28340 9596
rect 28972 9556 29012 9596
rect 29260 9556 29300 9596
rect 31372 9556 31412 9596
rect 31756 9556 31796 9596
rect 33100 9556 33140 9596
rect 40588 9724 40628 9764
rect 43756 9724 43796 9764
rect 35404 9640 35444 9680
rect 36172 9640 36212 9680
rect 36460 9640 36500 9680
rect 40780 9640 40820 9680
rect 43276 9640 43316 9680
rect 34828 9556 34868 9596
rect 36364 9556 36404 9596
rect 12076 9472 12116 9512
rect 12844 9472 12884 9512
rect 13228 9472 13268 9512
rect 13996 9472 14036 9512
rect 14380 9472 14420 9512
rect 15148 9472 15188 9512
rect 15532 9472 15572 9512
rect 15916 9472 15956 9512
rect 16684 9472 16724 9512
rect 17452 9472 17492 9512
rect 17836 9472 17876 9512
rect 18412 9472 18452 9512
rect 18796 9472 18836 9512
rect 19372 9472 19412 9512
rect 19756 9472 19796 9512
rect 20716 9472 20756 9512
rect 22540 9472 22580 9512
rect 24076 9472 24116 9512
rect 24268 9472 24308 9512
rect 25708 9472 25748 9512
rect 28108 9472 28148 9512
rect 29932 9472 29972 9512
rect 32716 9472 32756 9512
rect 33004 9472 33044 9512
rect 33580 9472 33620 9512
rect 34636 9472 34676 9512
rect 35020 9472 35060 9512
rect 35692 9472 35732 9512
rect 36268 9472 36308 9512
rect 40012 9472 40052 9512
rect 41836 9472 41876 9512
rect 42028 9472 42068 9512
rect 43276 9472 43316 9512
rect 43660 9472 43700 9512
rect 44140 9472 44180 9512
rect 13420 9388 13460 9428
rect 14956 9388 14996 9428
rect 16780 9388 16820 9428
rect 17260 9388 17300 9428
rect 18124 9388 18164 9428
rect 19084 9388 19124 9428
rect 21868 9388 21908 9428
rect 25036 9388 25076 9428
rect 26188 9388 26228 9428
rect 27340 9388 27380 9428
rect 28684 9388 28724 9428
rect 29740 9388 29780 9428
rect 31756 9388 31796 9428
rect 13708 9304 13748 9344
rect 14188 9304 14228 9344
rect 16396 9304 16436 9344
rect 17740 9304 17780 9344
rect 17932 9304 17972 9344
rect 19852 9304 19892 9344
rect 20620 9304 20660 9344
rect 20908 9304 20948 9344
rect 22348 9304 22388 9344
rect 24364 9304 24404 9344
rect 24652 9304 24692 9344
rect 25900 9304 25940 9344
rect 27916 9304 27956 9344
rect 30028 9304 30068 9344
rect 30892 9304 30932 9344
rect 1900 9220 1940 9260
rect 2764 9220 2804 9260
rect 2092 9136 2132 9176
rect 8716 9136 8756 9176
rect 11308 9220 11348 9260
rect 11884 9220 11924 9260
rect 12172 9220 12212 9260
rect 13420 9220 13460 9260
rect 14572 9220 14612 9260
rect 17356 9220 17396 9260
rect 18220 9220 18260 9260
rect 19084 9220 19124 9260
rect 21004 9220 21044 9260
rect 21676 9220 21716 9260
rect 22732 9220 22772 9260
rect 24844 9220 24884 9260
rect 26476 9220 26516 9260
rect 27724 9220 27764 9260
rect 11788 9136 11828 9176
rect 14092 9136 14132 9176
rect 14764 9136 14804 9176
rect 15340 9136 15380 9176
rect 17164 9136 17204 9176
rect 17740 9136 17780 9176
rect 19852 9136 19892 9176
rect 21292 9136 21332 9176
rect 2380 9052 2420 9092
rect 4780 9052 4820 9092
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 12268 9052 12308 9092
rect 14188 9052 14228 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 1228 8968 1268 9008
rect 23500 9136 23540 9176
rect 25804 9136 25844 9176
rect 26860 9136 26900 9176
rect 29164 9136 29204 9176
rect 34060 9388 34100 9428
rect 35404 9388 35444 9428
rect 35596 9388 35636 9428
rect 35788 9388 35828 9428
rect 36172 9388 36212 9428
rect 37900 9388 37940 9428
rect 42220 9388 42260 9428
rect 43180 9388 43220 9428
rect 43468 9388 43508 9428
rect 32332 9304 32372 9344
rect 33484 9304 33524 9344
rect 34540 9304 34580 9344
rect 37420 9304 37460 9344
rect 44236 9304 44276 9344
rect 33196 9220 33236 9260
rect 34252 9220 34292 9260
rect 35500 9220 35540 9260
rect 36364 9220 36404 9260
rect 40684 9220 40715 9260
rect 40715 9220 40724 9260
rect 41740 9220 41780 9260
rect 45868 9220 45908 9260
rect 20716 9052 20756 9092
rect 21484 9052 21524 9092
rect 21772 9052 21812 9092
rect 26188 9052 26228 9092
rect 35980 9136 36020 9176
rect 41164 9136 41204 9176
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 38860 9052 38900 9092
rect 3340 8968 3380 9008
rect 10060 8968 10100 9008
rect 11020 8968 11060 9008
rect 11884 8968 11924 9008
rect 12556 8968 12596 9008
rect 13516 8968 13556 9008
rect 13900 8968 13940 9008
rect 16972 8968 17012 9008
rect 17164 8968 17204 9008
rect 27340 8968 27380 9008
rect 33484 8968 33524 9008
rect 38956 8968 38996 9008
rect 10156 8884 10196 8924
rect 11980 8884 12020 8924
rect 12364 8884 12404 8924
rect 14956 8884 14996 8924
rect 15148 8884 15188 8924
rect 18508 8884 18548 8924
rect 18700 8884 18740 8924
rect 19276 8884 19316 8924
rect 19660 8884 19700 8924
rect 19948 8884 19988 8924
rect 20524 8884 20564 8924
rect 20812 8884 20852 8924
rect 1900 8800 1940 8840
rect 11116 8800 11156 8840
rect 13420 8800 13460 8840
rect 10156 8716 10196 8756
rect 11020 8716 11060 8756
rect 11596 8716 11636 8756
rect 11980 8716 12020 8756
rect 14092 8716 14132 8756
rect 14668 8716 14708 8756
rect 15052 8716 15092 8756
rect 15628 8716 15668 8756
rect 16204 8716 16244 8756
rect 16396 8716 16436 8756
rect 18604 8716 18644 8756
rect 652 8632 692 8672
rect 2380 8632 2420 8672
rect 2956 8632 2996 8672
rect 3340 8632 3380 8672
rect 9388 8632 9428 8672
rect 10252 8632 10292 8672
rect 10828 8632 10868 8672
rect 11212 8632 11252 8672
rect 12364 8632 12404 8672
rect 12844 8632 12884 8672
rect 13516 8632 13556 8672
rect 14188 8632 14228 8672
rect 15244 8632 15284 8672
rect 15724 8632 15764 8672
rect 20620 8716 20660 8756
rect 21964 8716 22004 8756
rect 22252 8716 22292 8756
rect 22828 8716 22868 8756
rect 16012 8632 16052 8672
rect 16300 8632 16340 8672
rect 16492 8632 16532 8672
rect 17068 8632 17108 8672
rect 17548 8632 17588 8672
rect 18220 8632 18260 8672
rect 18700 8632 18740 8672
rect 19084 8632 19124 8672
rect 19468 8632 19508 8672
rect 21004 8632 21044 8672
rect 21196 8632 21236 8672
rect 21580 8632 21620 8672
rect 22636 8632 22676 8672
rect 23500 8716 23540 8756
rect 23404 8632 23444 8672
rect 12940 8548 12980 8588
rect 13132 8548 13172 8588
rect 13612 8548 13652 8588
rect 13900 8548 13940 8588
rect 14764 8548 14804 8588
rect 16876 8548 16916 8588
rect 17164 8548 17204 8588
rect 26764 8884 26804 8924
rect 26956 8884 26996 8924
rect 32140 8884 32180 8924
rect 24460 8800 24500 8840
rect 28396 8800 28436 8840
rect 28780 8800 28820 8840
rect 25612 8716 25652 8756
rect 26188 8716 26228 8756
rect 26380 8716 26420 8756
rect 26572 8716 26612 8756
rect 29356 8716 29396 8756
rect 32524 8884 32564 8924
rect 32908 8884 32948 8924
rect 33292 8884 33332 8924
rect 33676 8884 33716 8924
rect 34348 8884 34388 8924
rect 35788 8884 35828 8924
rect 37324 8884 37364 8924
rect 34444 8800 34484 8840
rect 35692 8800 35732 8840
rect 37804 8800 37844 8840
rect 41068 8800 41108 8840
rect 42220 8800 42260 8840
rect 42796 8800 42836 8840
rect 25228 8632 25268 8672
rect 25996 8632 26036 8672
rect 28780 8632 28820 8672
rect 29068 8632 29108 8672
rect 29644 8632 29684 8672
rect 33388 8632 33428 8672
rect 38860 8716 38900 8756
rect 40684 8716 40724 8756
rect 43180 8716 43220 8756
rect 43372 8884 43412 8924
rect 33772 8632 33812 8672
rect 34540 8632 34580 8672
rect 35404 8632 35444 8672
rect 37900 8632 37940 8672
rect 41740 8632 41780 8672
rect 42892 8632 42932 8672
rect 43084 8632 43124 8672
rect 43852 8632 43892 8672
rect 44332 8632 44372 8672
rect 45004 8632 45044 8672
rect 27532 8548 27572 8588
rect 31948 8548 31988 8588
rect 34636 8548 34676 8588
rect 35308 8548 35348 8588
rect 45772 8548 45812 8588
rect 11884 8464 11924 8504
rect 13420 8464 13460 8504
rect 13996 8464 14036 8504
rect 16972 8464 17012 8504
rect 17452 8464 17492 8504
rect 18700 8464 18740 8504
rect 19756 8464 19796 8504
rect 19948 8464 19988 8504
rect 20140 8464 20180 8504
rect 26092 8464 26132 8504
rect 27628 8464 27668 8504
rect 28684 8464 28724 8504
rect 29260 8464 29300 8504
rect 29836 8464 29876 8504
rect 35500 8464 35540 8504
rect 38380 8464 38420 8504
rect 38860 8464 38900 8504
rect 40108 8464 40148 8504
rect 40300 8464 40340 8504
rect 43372 8464 43412 8504
rect 12076 8380 12116 8420
rect 19852 8380 19892 8420
rect 20908 8380 20948 8420
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 25612 8296 25652 8336
rect 15916 8212 15956 8252
rect 19852 8212 19892 8252
rect 20140 8212 20180 8252
rect 25708 8212 25748 8252
rect 11404 8128 11444 8168
rect 14380 8128 14420 8168
rect 25996 8380 26036 8420
rect 29740 8380 29780 8420
rect 30220 8380 30260 8420
rect 36748 8380 36788 8420
rect 42892 8380 42932 8420
rect 27436 8296 27476 8336
rect 28492 8296 28532 8336
rect 28684 8296 28724 8336
rect 31564 8296 31604 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 43084 8296 43124 8336
rect 30124 8212 30164 8252
rect 32620 8212 32660 8252
rect 35692 8212 35732 8252
rect 18604 8128 18644 8168
rect 19660 8128 19700 8168
rect 29740 8128 29780 8168
rect 31948 8128 31988 8168
rect 35020 8128 35060 8168
rect 35308 8128 35348 8168
rect 37708 8128 37748 8168
rect 10156 8044 10196 8084
rect 12844 8044 12884 8084
rect 15052 8044 15092 8084
rect 16300 8044 16340 8084
rect 652 7960 692 8000
rect 1228 7960 1268 8000
rect 11308 7960 11348 8000
rect 11788 7960 11828 8000
rect 15148 7960 15188 8000
rect 15340 7960 15380 8000
rect 15916 7960 15956 8000
rect 16204 7960 16235 8000
rect 16235 7960 16244 8000
rect 16780 8044 16820 8084
rect 20140 8044 20180 8084
rect 28684 8044 28724 8084
rect 29068 8044 29108 8084
rect 29356 8044 29396 8084
rect 29644 8044 29684 8084
rect 31564 8044 31604 8084
rect 34540 8044 34580 8084
rect 35884 8044 35924 8084
rect 42124 8044 42164 8084
rect 17548 7960 17588 8000
rect 11980 7876 12020 7916
rect 13420 7876 13460 7916
rect 14668 7876 14699 7916
rect 14699 7876 14708 7916
rect 14956 7876 14996 7916
rect 16300 7876 16340 7916
rect 17068 7876 17108 7916
rect 17740 7876 17780 7916
rect 12940 7792 12980 7832
rect 14476 7792 14516 7832
rect 16396 7792 16427 7832
rect 16427 7792 16436 7832
rect 17548 7792 17588 7832
rect 18796 7876 18836 7916
rect 43276 8128 43316 8168
rect 43564 8044 43604 8084
rect 45676 8464 45716 8504
rect 45868 8296 45908 8336
rect 25612 7960 25652 8000
rect 26188 7960 26228 8000
rect 28972 7960 29012 8000
rect 29164 7960 29204 8000
rect 29836 7960 29876 8000
rect 31468 7960 31508 8000
rect 31756 7960 31796 8000
rect 32236 7960 32276 8000
rect 34348 7960 34388 8000
rect 38188 7960 38228 8000
rect 38860 7960 38900 8000
rect 39820 7960 39860 8000
rect 40108 7960 40148 8000
rect 40396 7960 40436 8000
rect 43372 7960 43412 8000
rect 43756 7960 43796 8000
rect 44908 7960 44948 8000
rect 45772 7960 45812 8000
rect 20716 7876 20756 7916
rect 21196 7876 21236 7916
rect 27532 7876 27572 7916
rect 29068 7876 29108 7916
rect 29740 7876 29780 7916
rect 30508 7876 30548 7916
rect 35980 7876 36020 7916
rect 38284 7876 38324 7916
rect 38476 7876 38516 7916
rect 28300 7792 28340 7832
rect 29932 7792 29972 7832
rect 30124 7792 30164 7832
rect 30316 7792 30356 7832
rect 30796 7792 30836 7832
rect 37036 7792 37076 7832
rect 38092 7792 38132 7832
rect 41836 7792 41876 7832
rect 42988 7792 43028 7832
rect 10060 7708 10100 7748
rect 11884 7708 11924 7748
rect 15916 7708 15947 7748
rect 15947 7708 15956 7748
rect 18796 7708 18836 7748
rect 27340 7708 27380 7748
rect 29164 7708 29204 7748
rect 30700 7708 30740 7748
rect 30892 7708 30932 7748
rect 32236 7708 32276 7748
rect 32428 7708 32468 7748
rect 37708 7708 37748 7748
rect 39052 7708 39092 7748
rect 39916 7708 39956 7748
rect 12172 7624 12212 7664
rect 17260 7624 17300 7664
rect 25420 7624 25460 7664
rect 28204 7624 28244 7664
rect 28684 7624 28724 7664
rect 41740 7708 41780 7748
rect 42220 7708 42260 7748
rect 43756 7708 43796 7748
rect 45868 7708 45908 7748
rect 38572 7624 38612 7664
rect 40396 7624 40436 7664
rect 44908 7624 44948 7664
rect 45676 7624 45716 7664
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 9292 7540 9332 7580
rect 16780 7540 16820 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20524 7540 20564 7580
rect 24940 7540 24980 7580
rect 28492 7540 28532 7580
rect 28780 7540 28820 7580
rect 32428 7540 32468 7580
rect 19660 7456 19700 7496
rect 25420 7456 25460 7496
rect 28972 7456 29012 7496
rect 16012 7372 16052 7412
rect 16204 7372 16244 7412
rect 25516 7372 25556 7412
rect 28876 7372 28916 7412
rect 1228 7288 1268 7328
rect 14668 7288 14708 7328
rect 15340 7288 15380 7328
rect 28300 7288 28340 7328
rect 29068 7288 29108 7328
rect 30604 7456 30644 7496
rect 29356 7372 29396 7412
rect 30124 7288 30164 7328
rect 32620 7540 32660 7580
rect 35020 7540 35060 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 35788 7540 35828 7580
rect 42988 7540 43028 7580
rect 39052 7456 39092 7496
rect 44620 7456 44660 7496
rect 32140 7372 32180 7412
rect 41740 7372 41780 7412
rect 43468 7372 43508 7412
rect 30796 7288 30836 7328
rect 42220 7288 42260 7328
rect 45868 7288 45908 7328
rect 11308 7204 11348 7244
rect 12940 7204 12980 7244
rect 13420 7204 13460 7244
rect 16108 7204 16148 7244
rect 18796 7204 18836 7244
rect 27148 7235 27188 7244
rect 27148 7204 27188 7235
rect 30604 7204 30644 7244
rect 30892 7204 30932 7244
rect 31564 7204 31604 7244
rect 31756 7204 31796 7244
rect 32140 7204 32180 7244
rect 38188 7204 38228 7244
rect 39436 7204 39476 7244
rect 39916 7204 39956 7244
rect 41836 7204 41876 7244
rect 4108 7120 4148 7160
rect 15244 7120 15284 7160
rect 15436 7120 15476 7160
rect 15916 7120 15956 7160
rect 17356 7120 17396 7160
rect 17932 7120 17972 7160
rect 18700 7120 18740 7160
rect 25516 7120 25556 7160
rect 28492 7120 28532 7160
rect 28780 7120 28820 7160
rect 29836 7120 29876 7160
rect 748 6952 788 6992
rect 31468 7120 31508 7160
rect 37708 7120 37748 7160
rect 38092 7120 38132 7160
rect 38668 7120 38708 7160
rect 38956 7120 38996 7160
rect 39340 7120 39380 7160
rect 40588 7120 40628 7160
rect 40876 7120 40916 7160
rect 41260 7120 41300 7160
rect 43084 7120 43124 7160
rect 43564 7120 43604 7160
rect 44524 7120 44564 7160
rect 8428 7036 8468 7076
rect 15532 7036 15572 7076
rect 15820 7036 15860 7076
rect 17548 7036 17588 7076
rect 17740 7036 17780 7076
rect 23692 7036 23732 7076
rect 28396 7036 28436 7076
rect 30028 7036 30068 7076
rect 35596 7036 35636 7076
rect 39148 7036 39188 7076
rect 10828 6952 10868 6992
rect 20716 6952 20756 6992
rect 22444 6952 22484 6992
rect 28204 6952 28244 6992
rect 29068 6952 29108 6992
rect 30316 6952 30356 6992
rect 35788 6952 35828 6992
rect 38668 6952 38708 6992
rect 41356 6952 41396 6992
rect 12364 6868 12404 6908
rect 27148 6868 27188 6908
rect 28684 6868 28724 6908
rect 29356 6868 29396 6908
rect 29548 6868 29588 6908
rect 35020 6868 35060 6908
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 11884 6784 11924 6824
rect 17740 6784 17780 6824
rect 17932 6784 17972 6824
rect 18700 6784 18740 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 24172 6784 24212 6824
rect 27340 6784 27380 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 35308 6868 35348 6908
rect 37996 6868 38036 6908
rect 41740 6784 41780 6824
rect 13228 6700 13268 6740
rect 25612 6700 25652 6740
rect 29356 6700 29396 6740
rect 29548 6700 29588 6740
rect 35020 6700 35060 6740
rect 43084 6700 43124 6740
rect 844 6616 884 6656
rect 17836 6616 17876 6656
rect 18028 6616 18068 6656
rect 23212 6616 23252 6656
rect 27340 6616 27380 6656
rect 27628 6616 27668 6656
rect 28300 6616 28340 6656
rect 29836 6616 29876 6656
rect 30508 6616 30548 6656
rect 40300 6616 40340 6656
rect 10060 6532 10100 6572
rect 19468 6532 19508 6572
rect 35116 6532 35156 6572
rect 35308 6532 35348 6572
rect 46252 6784 46292 6824
rect 46252 6616 46292 6656
rect 1228 6448 1268 6488
rect 27820 6448 27860 6488
rect 28780 6448 28820 6488
rect 29164 6448 29204 6488
rect 29356 6448 29396 6488
rect 29836 6448 29876 6488
rect 30412 6448 30452 6488
rect 31660 6448 31700 6488
rect 34636 6448 34676 6488
rect 34924 6448 34964 6488
rect 35692 6448 35732 6488
rect 36460 6448 36500 6488
rect 37996 6448 38036 6488
rect 41260 6448 41300 6488
rect 43180 6448 43220 6488
rect 44812 6532 44852 6572
rect 8428 6364 8468 6404
rect 23308 6364 23348 6404
rect 26188 6364 26228 6404
rect 27532 6364 27572 6404
rect 29548 6364 29588 6404
rect 30316 6364 30356 6404
rect 27148 6280 27188 6320
rect 30028 6280 30068 6320
rect 31372 6280 31412 6320
rect 34924 6280 34964 6320
rect 28876 6196 28916 6236
rect 29740 6196 29780 6236
rect 35884 6364 35924 6404
rect 43564 6364 43604 6404
rect 37132 6280 37172 6320
rect 40876 6280 40916 6320
rect 40204 6196 40244 6236
rect 40396 6196 40436 6236
rect 43084 6196 43124 6236
rect 43468 6196 43508 6236
rect 43852 6196 43883 6236
rect 43883 6196 43892 6236
rect 1324 6112 1364 6152
rect 17836 6112 17876 6152
rect 18028 6112 18068 6152
rect 20524 6112 20564 6152
rect 31084 6112 31124 6152
rect 31276 6112 31316 6152
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 27820 6028 27860 6068
rect 30988 6028 31028 6068
rect 31468 6028 31508 6068
rect 35020 6028 35060 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 38860 6028 38900 6068
rect 44524 6028 44564 6068
rect 46252 6112 46292 6152
rect 23692 5944 23732 5984
rect 28012 5944 28052 5984
rect 30220 5944 30260 5984
rect 46252 5944 46292 5984
rect 1420 5860 1460 5900
rect 18700 5860 18740 5900
rect 25804 5860 25844 5900
rect 32908 5860 32948 5900
rect 39148 5860 39188 5900
rect 43084 5860 43124 5900
rect 43276 5860 43316 5900
rect 44716 5860 44756 5900
rect 12748 5776 12788 5816
rect 34636 5776 34676 5816
rect 35404 5776 35444 5816
rect 35596 5776 35636 5816
rect 40204 5776 40244 5816
rect 34444 5692 34484 5732
rect 41740 5692 41780 5732
rect 1324 5608 1364 5648
rect 16972 5524 17012 5564
rect 38860 5608 38900 5648
rect 41644 5608 41684 5648
rect 43564 5608 43604 5648
rect 43852 5608 43892 5648
rect 844 5356 884 5396
rect 1420 5272 1460 5312
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 2764 5188 2804 5228
rect 27628 5188 27668 5228
rect 16396 5104 16436 5144
rect 24460 5104 24500 5144
rect 30604 5104 30644 5144
rect 4780 5020 4820 5060
rect 12268 4936 12308 4976
rect 12652 4852 12692 4892
rect 16396 4852 16436 4892
rect 27148 4936 27188 4976
rect 22444 4852 22484 4892
rect 23020 4852 23060 4892
rect 24844 4852 24884 4892
rect 25324 4852 25364 4892
rect 27628 4852 27668 4892
rect 34636 5524 34676 5564
rect 46252 5440 46292 5480
rect 46252 5272 46292 5312
rect 41836 4936 41876 4976
rect 44908 4936 44948 4976
rect 39820 4852 39860 4892
rect 44332 4768 44372 4808
rect 13132 4684 13172 4724
rect 23212 4684 23252 4724
rect 24076 4684 24116 4724
rect 38956 4600 38996 4640
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 23788 4516 23828 4556
rect 23980 4516 24020 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 13804 4348 13844 4388
rect 23020 4348 23060 4388
rect 23308 4348 23348 4388
rect 1420 4264 1460 4304
rect 13516 4264 13556 4304
rect 15148 4264 15188 4304
rect 15532 4264 15572 4304
rect 15820 4264 15860 4304
rect 17644 4264 17684 4304
rect 23212 4264 23252 4304
rect 23980 4264 24020 4304
rect 25036 4264 25076 4304
rect 11788 4180 11828 4220
rect 12652 4180 12683 4220
rect 12683 4180 12692 4220
rect 13420 4180 13460 4220
rect 19084 4211 19124 4220
rect 19084 4180 19124 4211
rect 22156 4180 22196 4220
rect 22540 4180 22580 4220
rect 22924 4180 22964 4220
rect 23500 4180 23540 4220
rect 23788 4180 23828 4220
rect 35884 4180 35924 4220
rect 38284 4180 38324 4220
rect 40300 4180 40340 4220
rect 12268 4096 12308 4136
rect 12460 4096 12500 4136
rect 13132 4096 13172 4136
rect 13612 4096 13652 4136
rect 14956 4096 14996 4136
rect 15436 4096 15476 4136
rect 16012 4096 16052 4136
rect 23404 4096 23444 4136
rect 41068 4180 41108 4220
rect 44620 4180 44660 4220
rect 24268 4096 24308 4136
rect 27628 4096 27668 4136
rect 33292 4096 33332 4136
rect 38764 4096 38804 4136
rect 41260 4096 41300 4136
rect 42124 4096 42164 4136
rect 14764 4012 14804 4052
rect 21196 4012 21236 4052
rect 22924 4012 22964 4052
rect 23116 4012 23156 4052
rect 23788 4012 23828 4052
rect 23980 4012 24020 4052
rect 27340 4012 27380 4052
rect 40012 4012 40052 4052
rect 40492 4012 40532 4052
rect 40780 4012 40820 4052
rect 1420 3928 1460 3968
rect 13708 3928 13748 3968
rect 16588 3928 16628 3968
rect 20140 3928 20180 3968
rect 21292 3928 21332 3968
rect 23596 3928 23636 3968
rect 25132 3928 25172 3968
rect 25900 3928 25940 3968
rect 27244 3928 27284 3968
rect 36076 3928 36116 3968
rect 38476 3928 38516 3968
rect 40684 3928 40724 3968
rect 44908 3928 44948 3968
rect 35884 3844 35924 3884
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 36172 3844 36212 3884
rect 38668 3844 38708 3884
rect 12172 3760 12212 3800
rect 14188 3760 14228 3800
rect 14380 3760 14420 3800
rect 16396 3760 16436 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 37420 3760 37460 3800
rect 45004 3760 45044 3800
rect 1228 3592 1268 3632
rect 23500 3676 23540 3716
rect 25036 3676 25076 3716
rect 29260 3676 29300 3716
rect 39340 3676 39380 3716
rect 10924 3592 10964 3632
rect 13516 3592 13556 3632
rect 13708 3592 13748 3632
rect 23020 3592 23060 3632
rect 15148 3508 15188 3548
rect 16396 3508 16436 3548
rect 23116 3508 23156 3548
rect 8716 3424 8756 3464
rect 9388 3424 9428 3464
rect 14092 3424 14132 3464
rect 14380 3424 14420 3464
rect 14764 3424 14795 3464
rect 14795 3424 14804 3464
rect 14956 3424 14996 3464
rect 19276 3424 19316 3464
rect 21196 3424 21236 3464
rect 21484 3424 21524 3464
rect 21964 3424 22004 3464
rect 22156 3424 22196 3464
rect 22636 3424 22676 3464
rect 11020 3340 11060 3380
rect 11788 3340 11828 3380
rect 12172 3340 12212 3380
rect 12652 3340 12692 3380
rect 13420 3340 13460 3380
rect 15052 3340 15092 3380
rect 15436 3340 15467 3380
rect 15467 3340 15476 3380
rect 16396 3340 16436 3380
rect 17740 3340 17780 3380
rect 20812 3340 20852 3380
rect 21772 3340 21812 3380
rect 22732 3340 22772 3380
rect 23980 3592 24020 3632
rect 23596 3424 23636 3464
rect 24940 3592 24980 3632
rect 25612 3592 25652 3632
rect 27436 3592 27476 3632
rect 29068 3592 29108 3632
rect 37996 3592 38036 3632
rect 38668 3592 38708 3632
rect 24748 3508 24788 3548
rect 44140 3508 44180 3548
rect 24844 3424 24884 3464
rect 25612 3424 25652 3464
rect 36364 3424 36404 3464
rect 37996 3424 38036 3464
rect 38476 3424 38516 3464
rect 39340 3424 39380 3464
rect 40300 3424 40340 3464
rect 40876 3424 40916 3464
rect 41740 3424 41780 3464
rect 42124 3424 42164 3464
rect 42508 3424 42548 3464
rect 42700 3424 42740 3464
rect 44812 3424 44852 3464
rect 24076 3340 24116 3380
rect 27148 3340 27188 3380
rect 27436 3340 27476 3380
rect 2092 3256 2132 3296
rect 13516 3256 13556 3296
rect 16300 3256 16340 3296
rect 10060 3172 10100 3212
rect 13420 3172 13460 3212
rect 14956 3172 14996 3212
rect 17932 3256 17972 3296
rect 21484 3256 21524 3296
rect 23788 3256 23828 3296
rect 24364 3256 24404 3296
rect 15628 3172 15668 3212
rect 15436 3088 15476 3128
rect 17548 3088 17588 3128
rect 17740 3088 17780 3128
rect 24268 3172 24308 3212
rect 31852 3256 31892 3296
rect 33100 3172 33140 3212
rect 38476 3088 38516 3128
rect 44428 3340 44468 3380
rect 43756 3256 43796 3296
rect 43372 3172 43412 3212
rect 44524 3088 44564 3128
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 12652 3004 12692 3044
rect 13804 3004 13844 3044
rect 15628 3004 15668 3044
rect 17836 3004 17876 3044
rect 19948 3004 19988 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 24748 3004 24788 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 15820 2920 15860 2960
rect 22732 2920 22772 2960
rect 24460 2920 24500 2960
rect 40300 2920 40340 2960
rect 39148 2836 39188 2876
rect 11788 2752 11828 2792
rect 11980 2752 12020 2792
rect 12844 2752 12884 2792
rect 13420 2752 13460 2792
rect 14764 2752 14804 2792
rect 15052 2752 15092 2792
rect 20620 2752 20660 2792
rect 23404 2752 23435 2792
rect 23435 2752 23444 2792
rect 34828 2752 34868 2792
rect 8716 2668 8756 2708
rect 11020 2668 11060 2708
rect 13516 2668 13523 2708
rect 13523 2668 13556 2708
rect 14956 2668 14996 2708
rect 15148 2668 15188 2708
rect 15724 2668 15764 2708
rect 22540 2668 22580 2708
rect 23020 2668 23060 2708
rect 23308 2668 23309 2708
rect 23309 2668 23348 2708
rect 23692 2668 23732 2708
rect 8908 2584 8948 2624
rect 12172 2584 12212 2624
rect 12652 2584 12692 2624
rect 13612 2584 13643 2624
rect 13643 2584 13652 2624
rect 14092 2584 14132 2624
rect 14476 2584 14516 2624
rect 18124 2584 18164 2624
rect 22636 2584 22676 2624
rect 22828 2584 22868 2624
rect 39244 2584 39284 2624
rect 44524 2584 44564 2624
rect 15820 2500 15860 2540
rect 21004 2500 21044 2540
rect 22540 2500 22580 2540
rect 23212 2500 23252 2540
rect 24172 2500 24212 2540
rect 39148 2500 39188 2540
rect 8812 2416 8852 2456
rect 11692 2416 11732 2456
rect 23020 2416 23060 2456
rect 15436 2332 15476 2372
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 23308 2416 23348 2456
rect 38956 2416 38996 2456
rect 12556 2248 12596 2288
rect 13228 2248 13268 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 17452 2164 17492 2204
rect 22156 2164 22196 2204
rect 25132 2080 25172 2120
rect 25612 2080 25652 2120
rect 39244 2080 39284 2120
rect 1420 1912 1460 1952
rect 30700 1996 30740 2036
rect 43372 1912 43412 1952
rect 43756 1912 43796 1952
rect 44140 1912 44180 1952
rect 44428 1912 44468 1952
rect 44908 1912 44948 1952
rect 8908 1828 8948 1868
rect 24460 1828 24500 1868
rect 8812 1744 8852 1784
rect 24652 1744 24692 1784
rect 45580 1744 45620 1784
rect 3148 1660 3188 1700
rect 4780 1660 4820 1700
rect 6604 1660 6644 1700
rect 8332 1660 8372 1700
rect 44620 1660 44660 1700
rect 41740 1576 41780 1616
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 46252 1408 46292 1448
rect 42700 1240 42740 1280
rect 46252 1240 46292 1280
rect 42508 904 42548 944
rect 45580 904 45620 944
rect 42124 568 42164 608
rect 44620 568 44660 608
rect 13516 148 13556 188
rect 41260 148 41300 188
rect 10060 64 10100 104
rect 40876 64 40916 104
<< metal3 >>
rect 11000 11764 11080 11844
rect 11192 11764 11272 11844
rect 11384 11764 11464 11844
rect 11576 11764 11656 11844
rect 11768 11764 11848 11844
rect 11960 11764 12040 11844
rect 12152 11764 12232 11844
rect 12344 11764 12424 11844
rect 12536 11764 12616 11844
rect 12728 11764 12808 11844
rect 12920 11764 13000 11844
rect 13112 11764 13192 11844
rect 13304 11764 13384 11844
rect 13496 11764 13576 11844
rect 13688 11764 13768 11844
rect 13880 11764 13960 11844
rect 14072 11764 14152 11844
rect 14264 11764 14344 11844
rect 14456 11764 14536 11844
rect 14648 11764 14728 11844
rect 14840 11764 14920 11844
rect 15032 11764 15112 11844
rect 15224 11764 15304 11844
rect 15416 11764 15496 11844
rect 15608 11764 15688 11844
rect 15800 11764 15880 11844
rect 15992 11764 16072 11844
rect 16184 11764 16264 11844
rect 16376 11764 16456 11844
rect 16568 11764 16648 11844
rect 16760 11764 16840 11844
rect 16952 11764 17032 11844
rect 17144 11764 17224 11844
rect 17336 11764 17416 11844
rect 17528 11764 17608 11844
rect 17720 11764 17800 11844
rect 17912 11764 17992 11844
rect 18104 11764 18184 11844
rect 18296 11764 18376 11844
rect 18488 11764 18568 11844
rect 18680 11764 18760 11844
rect 18872 11764 18952 11844
rect 19064 11764 19144 11844
rect 19256 11764 19336 11844
rect 19448 11764 19528 11844
rect 19640 11764 19720 11844
rect 19832 11764 19912 11844
rect 20024 11764 20104 11844
rect 20216 11764 20296 11844
rect 20408 11764 20488 11844
rect 20600 11764 20680 11844
rect 20792 11764 20872 11844
rect 20984 11764 21064 11844
rect 21176 11764 21256 11844
rect 21368 11764 21448 11844
rect 21560 11764 21640 11844
rect 21752 11764 21832 11844
rect 21944 11764 22024 11844
rect 22136 11764 22216 11844
rect 22328 11764 22408 11844
rect 22520 11764 22600 11844
rect 22712 11764 22792 11844
rect 22904 11764 22984 11844
rect 23096 11764 23176 11844
rect 23288 11764 23368 11844
rect 23480 11764 23560 11844
rect 23672 11764 23752 11844
rect 23864 11764 23944 11844
rect 24056 11764 24136 11844
rect 24248 11764 24328 11844
rect 24440 11764 24520 11844
rect 24632 11764 24712 11844
rect 24824 11764 24904 11844
rect 25016 11764 25096 11844
rect 25208 11764 25288 11844
rect 25400 11764 25480 11844
rect 25592 11764 25672 11844
rect 25784 11764 25864 11844
rect 25976 11764 26056 11844
rect 26168 11764 26248 11844
rect 26360 11764 26440 11844
rect 26552 11764 26632 11844
rect 26744 11764 26824 11844
rect 26936 11764 27016 11844
rect 27128 11764 27208 11844
rect 27320 11764 27400 11844
rect 27512 11764 27592 11844
rect 27704 11764 27784 11844
rect 27896 11764 27976 11844
rect 28088 11764 28168 11844
rect 28280 11764 28360 11844
rect 28472 11764 28552 11844
rect 28664 11764 28744 11844
rect 28856 11764 28936 11844
rect 29048 11764 29128 11844
rect 29240 11764 29320 11844
rect 29432 11764 29512 11844
rect 29624 11764 29704 11844
rect 29816 11764 29896 11844
rect 30008 11764 30088 11844
rect 30200 11764 30280 11844
rect 30392 11764 30472 11844
rect 30584 11764 30664 11844
rect 30776 11764 30856 11844
rect 30968 11764 31048 11844
rect 31160 11764 31240 11844
rect 31352 11764 31432 11844
rect 31544 11764 31624 11844
rect 31736 11764 31816 11844
rect 31928 11764 32008 11844
rect 32120 11764 32200 11844
rect 32312 11764 32392 11844
rect 32504 11764 32584 11844
rect 32696 11764 32776 11844
rect 32888 11764 32968 11844
rect 33080 11764 33160 11844
rect 33272 11764 33352 11844
rect 33464 11764 33544 11844
rect 33656 11764 33736 11844
rect 33848 11764 33928 11844
rect 34040 11764 34120 11844
rect 34232 11764 34312 11844
rect 34424 11764 34504 11844
rect 34616 11764 34696 11844
rect 34808 11764 34888 11844
rect 35000 11764 35080 11844
rect 1420 11024 1460 11033
rect 1132 10688 1172 10697
rect 1036 10352 1076 10361
rect 1036 9428 1076 10312
rect 1132 9932 1172 10648
rect 1420 10016 1460 10984
rect 2956 10100 2996 10109
rect 1420 9967 1460 9976
rect 2764 10016 2804 10025
rect 1132 9883 1172 9892
rect 1036 9379 1076 9388
rect 1228 9512 1268 9521
rect 1228 9008 1268 9472
rect 2764 9512 2804 9976
rect 2764 9463 2804 9472
rect 1228 8959 1268 8968
rect 1900 9260 1940 9269
rect 1900 8840 1940 9220
rect 2764 9260 2804 9269
rect 1900 8791 1940 8800
rect 2092 9176 2132 9185
rect 652 8672 692 8681
rect 652 8000 692 8632
rect 652 7951 692 7960
rect 1228 8000 1268 8009
rect 1228 7328 1268 7960
rect 1228 7279 1268 7288
rect 748 6992 788 7001
rect 748 4136 788 6952
rect 844 6656 884 6665
rect 844 5396 884 6616
rect 844 5347 884 5356
rect 1228 6488 1268 6497
rect 748 4087 788 4096
rect 1228 3632 1268 6448
rect 1324 6152 1364 6161
rect 1324 5648 1364 6112
rect 1324 5599 1364 5608
rect 1420 5900 1460 5909
rect 1420 5312 1460 5860
rect 1420 5263 1460 5272
rect 1420 4304 1460 4313
rect 1420 4169 1460 4264
rect 1420 3968 1460 3977
rect 1420 3833 1460 3928
rect 1228 3583 1268 3592
rect 2092 3296 2132 9136
rect 2380 9092 2420 9101
rect 2380 8672 2420 9052
rect 2380 8623 2420 8632
rect 2764 5228 2804 9220
rect 2956 8672 2996 10060
rect 10060 10100 10100 10109
rect 10252 10100 10292 10109
rect 10100 10060 10196 10100
rect 10060 10051 10100 10060
rect 9388 10016 9428 10025
rect 3688 9848 4056 9857
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 3688 9799 4056 9808
rect 9292 9596 9332 9605
rect 4108 9428 4148 9437
rect 2956 8623 2996 8632
rect 3340 9008 3380 9017
rect 3340 8672 3380 8968
rect 3340 8623 3380 8632
rect 3688 8336 4056 8345
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 3688 8287 4056 8296
rect 4108 7160 4148 9388
rect 8716 9176 8756 9185
rect 4108 7111 4148 7120
rect 4780 9092 4820 9101
rect 3688 6824 4056 6833
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 3688 6775 4056 6784
rect 3688 5312 4056 5321
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 3688 5263 4056 5272
rect 2764 5179 2804 5188
rect 4780 5060 4820 9052
rect 4928 9092 5296 9101
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 4928 9043 5296 9052
rect 4928 7580 5296 7589
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 4928 7531 5296 7540
rect 8428 7076 8468 7085
rect 8428 6404 8468 7036
rect 8428 6355 8468 6364
rect 4928 6068 5296 6077
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 4928 6019 5296 6028
rect 4780 5011 4820 5020
rect 4928 4556 5296 4565
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 4928 4507 5296 4516
rect 3688 3800 4056 3809
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 3688 3751 4056 3760
rect 2092 3247 2132 3256
rect 8716 3464 8756 9136
rect 9292 7580 9332 9556
rect 9388 9512 9428 9976
rect 10156 9932 10196 10060
rect 10156 9883 10196 9892
rect 9388 9463 9428 9472
rect 10060 9848 10100 9857
rect 10060 9008 10100 9808
rect 10252 9680 10292 10060
rect 10252 9631 10292 9640
rect 10060 8959 10100 8968
rect 10156 9512 10196 9521
rect 10156 8924 10196 9472
rect 10156 8875 10196 8884
rect 10540 9512 10580 9521
rect 10156 8756 10196 8765
rect 9292 7531 9332 7540
rect 9388 8672 9428 8681
rect 4928 3044 5296 3053
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 4928 2995 5296 3004
rect 8716 2708 8756 3424
rect 9388 3464 9428 8632
rect 10156 8084 10196 8716
rect 10156 8035 10196 8044
rect 10252 8672 10292 8681
rect 10060 7748 10100 7757
rect 10060 6572 10100 7708
rect 10060 6523 10100 6532
rect 10252 6236 10292 8632
rect 10540 8420 10580 9472
rect 10828 9512 10868 9521
rect 10828 9428 10868 9472
rect 10828 9377 10868 9388
rect 10924 9512 10964 9521
rect 10540 8371 10580 8380
rect 10828 8672 10868 8681
rect 10828 6992 10868 8632
rect 10828 6943 10868 6952
rect 10252 6187 10292 6196
rect 10924 3632 10964 9472
rect 11020 9008 11060 11764
rect 11212 10100 11252 11764
rect 11212 10051 11252 10060
rect 11308 9764 11348 9773
rect 11308 9629 11348 9724
rect 11308 9428 11348 9437
rect 11308 9260 11348 9388
rect 11308 9211 11348 9220
rect 11020 8959 11060 8968
rect 11116 8840 11156 8849
rect 11020 8756 11060 8765
rect 11020 8336 11060 8716
rect 11116 8672 11156 8800
rect 11212 8672 11252 8681
rect 11116 8632 11212 8672
rect 11212 8623 11252 8632
rect 11020 8287 11060 8296
rect 11404 8168 11444 11764
rect 11500 9428 11540 9437
rect 11500 9260 11540 9388
rect 11500 9211 11540 9220
rect 11596 8756 11636 11764
rect 11788 9680 11828 11764
rect 11788 9631 11828 9640
rect 11884 9764 11924 9773
rect 11596 8707 11636 8716
rect 11692 9512 11732 9521
rect 11404 8119 11444 8128
rect 11308 8000 11348 8009
rect 11308 7244 11348 7960
rect 11308 7195 11348 7204
rect 10924 3583 10964 3592
rect 9388 3415 9428 3424
rect 11020 3380 11060 3389
rect 10060 3212 10100 3221
rect 10060 3077 10100 3172
rect 8716 2659 8756 2668
rect 11020 2708 11060 3340
rect 11020 2659 11060 2668
rect 8908 2624 8948 2633
rect 8812 2456 8852 2465
rect 3688 2288 4056 2297
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 3688 2239 4056 2248
rect 1420 1952 1460 1961
rect 1420 80 1460 1912
rect 8812 1784 8852 2416
rect 8908 1868 8948 2584
rect 11692 2456 11732 9472
rect 11884 9260 11924 9724
rect 11884 9211 11924 9220
rect 11788 9176 11828 9185
rect 11788 8000 11828 9136
rect 11884 9008 11924 9017
rect 11884 8504 11924 8968
rect 11980 8924 12020 11764
rect 11980 8875 12020 8884
rect 12076 9512 12116 9521
rect 11980 8756 12020 8765
rect 11980 8621 12020 8716
rect 11884 8455 11924 8464
rect 12076 8420 12116 9472
rect 12172 9512 12212 11764
rect 12172 9463 12212 9472
rect 12076 8371 12116 8380
rect 12172 9260 12212 9269
rect 11788 7951 11828 7960
rect 11980 7916 12020 7925
rect 11884 7748 11924 7757
rect 11884 7613 11924 7708
rect 11884 6824 11924 6833
rect 11788 4220 11828 4229
rect 11788 3380 11828 4180
rect 11788 2792 11828 3340
rect 11788 2743 11828 2752
rect 11692 2407 11732 2416
rect 8908 1819 8948 1828
rect 8812 1735 8852 1744
rect 3148 1700 3188 1709
rect 3148 80 3188 1660
rect 4780 1700 4820 1709
rect 4780 860 4820 1660
rect 6604 1700 6644 1709
rect 4928 1532 5296 1541
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 4928 1483 5296 1492
rect 4780 820 4916 860
rect 4876 80 4916 820
rect 6604 80 6644 1660
rect 8332 1700 8372 1709
rect 8332 80 8372 1660
rect 11884 1448 11924 6784
rect 11980 2792 12020 7876
rect 12172 7664 12212 9220
rect 12268 9176 12308 9185
rect 12268 9092 12308 9136
rect 12268 9041 12308 9052
rect 12364 8924 12404 11764
rect 12364 8875 12404 8884
rect 12460 9932 12500 9941
rect 12172 7615 12212 7624
rect 12364 8672 12404 8681
rect 12364 6908 12404 8632
rect 12364 6859 12404 6868
rect 12268 4976 12308 4985
rect 12268 4136 12308 4936
rect 12268 4087 12308 4096
rect 12460 4136 12500 9892
rect 12556 9428 12596 11764
rect 12652 9848 12692 9857
rect 12652 9596 12692 9808
rect 12652 9547 12692 9556
rect 12556 9379 12596 9388
rect 12748 9260 12788 11764
rect 12940 11444 12980 11764
rect 12940 11404 13076 11444
rect 12940 10100 12980 10109
rect 12844 10060 12940 10100
rect 12844 9764 12884 10060
rect 12940 10051 12980 10060
rect 13036 10100 13076 11404
rect 13036 10051 13076 10060
rect 12844 9715 12884 9724
rect 12940 9680 12980 9689
rect 12940 9596 12980 9640
rect 12940 9545 12980 9556
rect 12556 9220 12788 9260
rect 12844 9512 12884 9521
rect 12556 9008 12596 9220
rect 12844 9092 12884 9472
rect 12844 9043 12884 9052
rect 12556 8959 12596 8968
rect 13132 8924 13172 11764
rect 13324 9680 13364 11764
rect 13324 9631 13364 9640
rect 13420 9764 13460 9775
rect 13420 9680 13460 9724
rect 13420 9631 13460 9640
rect 13132 8875 13172 8884
rect 13228 9512 13268 9521
rect 12748 8840 12788 8849
rect 12748 5816 12788 8800
rect 12844 8672 12884 8681
rect 12844 8252 12884 8632
rect 12940 8588 12980 8597
rect 13132 8588 13172 8597
rect 12980 8548 13076 8588
rect 12940 8520 12980 8548
rect 12844 8203 12884 8212
rect 12748 5767 12788 5776
rect 12844 8084 12884 8093
rect 12652 4892 12692 4901
rect 12652 4220 12692 4852
rect 12652 4171 12692 4180
rect 12460 4087 12500 4096
rect 11980 2743 12020 2752
rect 12172 3800 12212 3809
rect 12172 3380 12212 3760
rect 12172 2624 12212 3340
rect 12652 3380 12692 3389
rect 12172 2575 12212 2584
rect 12556 3296 12596 3305
rect 12556 2288 12596 3256
rect 12652 3044 12692 3340
rect 12652 2624 12692 3004
rect 12844 2792 12884 8044
rect 12940 7832 12980 7841
rect 12940 7697 12980 7792
rect 12940 7244 12980 7253
rect 12940 3380 12980 7204
rect 12940 3331 12980 3340
rect 13036 2900 13076 8548
rect 13132 8504 13172 8548
rect 13132 8453 13172 8464
rect 13228 6740 13268 9472
rect 13420 9428 13460 9437
rect 13420 9260 13460 9388
rect 13420 9211 13460 9220
rect 13516 9008 13556 11764
rect 13708 9344 13748 11764
rect 13708 9295 13748 9304
rect 13804 9596 13844 9605
rect 13516 8959 13556 8968
rect 13420 8840 13460 8849
rect 13420 8504 13460 8800
rect 13516 8672 13556 8681
rect 13516 8537 13556 8632
rect 13612 8588 13652 8597
rect 13420 8455 13460 8464
rect 13612 8453 13652 8548
rect 13420 7916 13460 7925
rect 13420 7244 13460 7876
rect 13420 7195 13460 7204
rect 13228 6691 13268 6700
rect 13132 4724 13172 4733
rect 13132 4136 13172 4684
rect 13804 4388 13844 9556
rect 13900 9008 13940 11764
rect 13996 10016 14036 10025
rect 13996 9680 14036 9976
rect 13996 9631 14036 9640
rect 13900 8959 13940 8968
rect 13996 9512 14036 9521
rect 13900 8588 13940 8597
rect 13900 7916 13940 8548
rect 13996 8504 14036 9472
rect 14092 9176 14132 11764
rect 14188 10100 14228 10109
rect 14188 9344 14228 10060
rect 14188 9295 14228 9304
rect 14092 9127 14132 9136
rect 14188 9092 14228 9101
rect 14092 8756 14132 8765
rect 14092 8621 14132 8716
rect 14188 8672 14228 9052
rect 14188 8623 14228 8632
rect 14284 8588 14324 11764
rect 14284 8539 14324 8548
rect 14380 9512 14420 9521
rect 13996 8455 14036 8464
rect 14380 8168 14420 9472
rect 14380 8119 14420 8128
rect 13900 7867 13940 7876
rect 14476 7832 14516 11764
rect 14668 9764 14708 11764
rect 14668 9715 14708 9724
rect 14476 7783 14516 7792
rect 14572 9260 14612 9269
rect 13804 4339 13844 4348
rect 13516 4304 13556 4313
rect 13132 4087 13172 4096
rect 13420 4220 13460 4229
rect 13420 3380 13460 4180
rect 13516 3632 13556 4264
rect 13516 3583 13556 3592
rect 13612 4136 13652 4145
rect 13420 3212 13460 3340
rect 13036 2860 13268 2900
rect 12844 2743 12884 2752
rect 12652 2575 12692 2584
rect 12556 2239 12596 2248
rect 13228 2288 13268 2860
rect 13420 2792 13460 3172
rect 13420 2743 13460 2752
rect 13516 3296 13556 3305
rect 13516 2708 13556 3256
rect 13516 2659 13556 2668
rect 13612 2624 13652 4096
rect 13708 3968 13748 3977
rect 13708 3632 13748 3928
rect 14188 3800 14228 3809
rect 14188 3665 14228 3760
rect 14380 3800 14420 3809
rect 13708 3583 13748 3592
rect 14092 3464 14132 3473
rect 14092 3128 14132 3424
rect 13804 3044 13844 3055
rect 13804 2960 13844 3004
rect 13804 2911 13844 2920
rect 13612 2575 13652 2584
rect 14092 2624 14132 3088
rect 14380 3464 14420 3760
rect 14380 2900 14420 3424
rect 14572 3044 14612 9220
rect 14764 9176 14804 9185
rect 14764 8840 14804 9136
rect 14668 8800 14804 8840
rect 14668 8756 14708 8800
rect 14668 8707 14708 8716
rect 14860 8756 14900 11764
rect 15052 9848 15092 11764
rect 15052 9799 15092 9808
rect 14956 9764 14996 9773
rect 14956 9428 14996 9724
rect 15148 9596 15188 9607
rect 15148 9512 15188 9556
rect 15148 9463 15188 9472
rect 14956 9379 14996 9388
rect 15244 9176 15284 11764
rect 14956 9136 15284 9176
rect 15340 9848 15380 9857
rect 15340 9176 15380 9808
rect 14956 8924 14996 9136
rect 15340 9127 15380 9136
rect 14956 8875 14996 8884
rect 15148 8924 15188 8933
rect 14860 8707 14900 8716
rect 15052 8756 15092 8765
rect 14764 8588 14804 8683
rect 14764 8539 14804 8548
rect 14764 8336 14804 8345
rect 14668 7916 14708 7925
rect 14668 7328 14708 7876
rect 14668 7279 14708 7288
rect 14764 4052 14804 8296
rect 15052 8084 15092 8716
rect 15052 8035 15092 8044
rect 15148 8000 15188 8884
rect 15148 7951 15188 7960
rect 15244 8672 15284 8681
rect 14956 7916 14996 7925
rect 14956 7580 14996 7876
rect 14956 7531 14996 7540
rect 15148 7244 15188 7253
rect 15148 4304 15188 7204
rect 15244 7160 15284 8632
rect 15340 8000 15380 8009
rect 15340 7328 15380 7960
rect 15340 7279 15380 7288
rect 15244 7111 15284 7120
rect 15436 7160 15476 11764
rect 15628 9764 15668 11764
rect 15628 9715 15668 9724
rect 15436 7111 15476 7120
rect 15532 9512 15572 9521
rect 15532 7076 15572 9472
rect 15628 8756 15668 8765
rect 15628 8621 15668 8716
rect 15724 8672 15764 8681
rect 15532 7027 15572 7036
rect 15148 4255 15188 4264
rect 15532 4304 15572 4313
rect 14764 4003 14804 4012
rect 14956 4136 14996 4145
rect 14572 2995 14612 3004
rect 14764 3464 14804 3473
rect 14380 2860 14516 2900
rect 14092 2575 14132 2584
rect 14476 2624 14516 2860
rect 14764 2792 14804 3424
rect 14956 3464 14996 4096
rect 15436 4136 15476 4145
rect 14956 3415 14996 3424
rect 15148 3548 15188 3557
rect 15052 3380 15092 3389
rect 14764 2743 14804 2752
rect 14956 3212 14996 3221
rect 14956 2708 14996 3172
rect 15052 2792 15092 3340
rect 15052 2743 15092 2752
rect 14956 2659 14996 2668
rect 15148 2708 15188 3508
rect 15436 3380 15476 4096
rect 15436 3331 15476 3340
rect 15436 3128 15476 3137
rect 15148 2659 15188 2668
rect 15244 3088 15436 3128
rect 14476 2575 14516 2584
rect 13228 2239 13268 2248
rect 11788 1408 11924 1448
rect 10060 104 10100 113
rect 1400 0 1480 80
rect 3128 0 3208 80
rect 4856 0 4936 80
rect 6584 0 6664 80
rect 8312 0 8392 80
rect 10040 64 10060 80
rect 11788 80 11828 1408
rect 13516 188 13556 197
rect 13516 80 13556 148
rect 15244 80 15284 3088
rect 15436 3079 15476 3088
rect 15532 2900 15572 4264
rect 15628 3296 15668 3307
rect 15628 3212 15668 3256
rect 15628 3163 15668 3172
rect 15628 3044 15668 3053
rect 15628 2909 15668 3004
rect 15436 2860 15572 2900
rect 15436 2372 15476 2860
rect 15724 2708 15764 8632
rect 15820 8588 15860 11764
rect 16012 10016 16052 11764
rect 16012 9967 16052 9976
rect 16108 10268 16148 10277
rect 15916 9932 15956 9941
rect 15916 9512 15956 9892
rect 15916 9463 15956 9472
rect 16108 8756 16148 10228
rect 15820 8539 15860 8548
rect 16012 8716 16148 8756
rect 16204 8756 16244 11764
rect 16396 10100 16436 11764
rect 16396 10051 16436 10060
rect 16300 9848 16340 9857
rect 16300 9680 16340 9808
rect 16300 9631 16340 9640
rect 16588 9596 16628 11764
rect 16492 9556 16628 9596
rect 16396 9344 16436 9353
rect 16492 9344 16532 9556
rect 16436 9304 16532 9344
rect 16684 9512 16724 9521
rect 16396 9295 16436 9304
rect 16492 9176 16532 9185
rect 16012 8672 16052 8716
rect 16204 8707 16244 8716
rect 16396 8756 16436 8765
rect 15916 8252 15956 8261
rect 15916 8000 15956 8212
rect 15916 7951 15956 7960
rect 15916 7748 15956 7757
rect 15820 7664 15860 7673
rect 15820 7076 15860 7624
rect 15916 7160 15956 7708
rect 16012 7580 16052 8632
rect 16300 8672 16340 8681
rect 16300 8084 16340 8632
rect 16300 8035 16340 8044
rect 16204 8000 16244 8009
rect 16012 7540 16148 7580
rect 15916 7111 15956 7120
rect 16012 7412 16052 7421
rect 15820 7027 15860 7036
rect 15820 6908 15860 6917
rect 15820 4304 15860 6868
rect 15820 4255 15860 4264
rect 16012 4136 16052 7372
rect 16108 7244 16148 7540
rect 16204 7412 16244 7960
rect 16204 7363 16244 7372
rect 16300 7916 16340 7925
rect 16108 7195 16148 7204
rect 16300 6908 16340 7876
rect 16396 7832 16436 8716
rect 16492 8672 16532 9136
rect 16492 8623 16532 8632
rect 16588 8840 16628 8849
rect 16396 7783 16436 7792
rect 16492 8252 16532 8261
rect 16492 7496 16532 8212
rect 16492 7447 16532 7456
rect 16300 6859 16340 6868
rect 16396 5144 16436 5153
rect 16396 4892 16436 5104
rect 16396 4843 16436 4852
rect 16012 4087 16052 4096
rect 16588 3968 16628 8800
rect 16684 8084 16724 9472
rect 16780 9428 16820 11764
rect 16780 9379 16820 9388
rect 16876 10184 16916 10193
rect 16876 8588 16916 10144
rect 16972 9008 17012 11764
rect 17164 9176 17204 11764
rect 17164 9127 17204 9136
rect 17260 9428 17300 9437
rect 17164 9008 17204 9017
rect 16972 8959 17012 8968
rect 17068 8968 17164 9008
rect 17068 8672 17108 8968
rect 17164 8959 17204 8968
rect 17068 8623 17108 8632
rect 16876 8539 16916 8548
rect 16972 8588 17012 8599
rect 16972 8504 17012 8548
rect 16972 8455 17012 8464
rect 17164 8588 17204 8597
rect 16684 8035 16724 8044
rect 16780 8084 16820 8093
rect 16780 7580 16820 8044
rect 17068 7916 17108 7925
rect 17164 7916 17204 8548
rect 17108 7876 17204 7916
rect 17068 7867 17108 7876
rect 17260 7664 17300 9388
rect 17356 9260 17396 11764
rect 17548 9848 17588 11764
rect 17548 9799 17588 9808
rect 17452 9764 17492 9775
rect 17452 9680 17492 9724
rect 17452 9631 17492 9640
rect 17452 9512 17492 9521
rect 17452 9428 17492 9472
rect 17452 9377 17492 9388
rect 17740 9344 17780 11764
rect 17932 9764 17972 11764
rect 17932 9715 17972 9724
rect 18124 9764 18164 11764
rect 18124 9715 18164 9724
rect 18316 9680 18356 11764
rect 18412 10016 18452 10025
rect 18412 9764 18452 9976
rect 18412 9715 18452 9724
rect 18316 9631 18356 9640
rect 17836 9512 17876 9521
rect 17836 9377 17876 9472
rect 18412 9512 18452 9521
rect 18124 9428 18164 9437
rect 17740 9295 17780 9304
rect 17932 9344 17972 9353
rect 17356 9211 17396 9220
rect 17740 9176 17780 9185
rect 17548 8672 17588 8681
rect 17260 7615 17300 7624
rect 17356 8504 17396 8513
rect 16780 7531 16820 7540
rect 17356 7160 17396 8464
rect 17356 7111 17396 7120
rect 17452 8504 17492 8513
rect 16588 3919 16628 3928
rect 16972 5564 17012 5573
rect 16396 3800 16436 3809
rect 16396 3548 16436 3760
rect 16396 3499 16436 3508
rect 16396 3380 16436 3389
rect 16300 3296 16340 3305
rect 16300 3161 16340 3256
rect 16396 3245 16436 3340
rect 15724 2659 15764 2668
rect 15820 2960 15860 2969
rect 15820 2540 15860 2920
rect 15820 2491 15860 2500
rect 15436 2323 15476 2332
rect 16972 80 17012 5524
rect 17452 2204 17492 8464
rect 17548 8000 17588 8632
rect 17548 7951 17588 7960
rect 17644 8000 17684 8009
rect 17548 7832 17588 7841
rect 17548 7076 17588 7792
rect 17548 7027 17588 7036
rect 17644 4304 17684 7960
rect 17740 7916 17780 9136
rect 17740 7076 17780 7876
rect 17932 7160 17972 9304
rect 17932 7111 17972 7120
rect 17740 7027 17780 7036
rect 17740 6824 17780 6833
rect 17932 6824 17972 6833
rect 17780 6784 17932 6824
rect 17740 6775 17780 6784
rect 17932 6775 17972 6784
rect 17836 6656 17876 6665
rect 18028 6656 18068 6665
rect 17876 6616 18028 6656
rect 17836 6607 17876 6616
rect 18028 6607 18068 6616
rect 17836 6152 17876 6161
rect 18028 6152 18068 6161
rect 17876 6112 18028 6152
rect 17836 6103 17876 6112
rect 18028 6103 18068 6112
rect 17644 4255 17684 4264
rect 17740 3800 17780 3809
rect 17740 3380 17780 3760
rect 17740 3331 17780 3340
rect 17932 3296 17972 3305
rect 17548 3128 17588 3137
rect 17740 3128 17780 3137
rect 17588 3088 17740 3128
rect 17548 3079 17588 3088
rect 17740 3079 17780 3088
rect 17932 3128 17972 3256
rect 17932 3079 17972 3088
rect 17836 3044 17876 3053
rect 17836 2960 17876 3004
rect 17836 2909 17876 2920
rect 18124 2624 18164 9388
rect 18220 9260 18260 9269
rect 18220 8672 18260 9220
rect 18220 8623 18260 8632
rect 18412 8252 18452 9472
rect 18508 8924 18548 11764
rect 18700 10268 18740 11764
rect 18604 10228 18740 10268
rect 18604 9596 18644 10228
rect 18892 10184 18932 11764
rect 18604 9547 18644 9556
rect 18700 10144 18932 10184
rect 18508 8875 18548 8884
rect 18700 8924 18740 10144
rect 19084 10016 19124 11764
rect 19084 9967 19124 9976
rect 18808 9848 19176 9857
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 18808 9799 19176 9808
rect 18700 8875 18740 8884
rect 18796 9512 18836 9521
rect 18412 8203 18452 8212
rect 18604 8756 18644 8765
rect 18604 8168 18644 8716
rect 18700 8672 18740 8681
rect 18700 8504 18740 8632
rect 18700 8455 18740 8464
rect 18796 8504 18836 9472
rect 19084 9428 19124 9437
rect 19084 9260 19124 9388
rect 19084 9211 19124 9220
rect 19276 8924 19316 11764
rect 19468 9680 19508 11764
rect 19468 9631 19508 9640
rect 19276 8875 19316 8884
rect 19372 9512 19412 9521
rect 19372 8924 19412 9472
rect 19372 8875 19412 8884
rect 19564 9260 19604 9269
rect 19084 8672 19124 8681
rect 19468 8672 19508 8681
rect 19124 8632 19316 8660
rect 19084 8620 19316 8632
rect 18796 8455 18836 8464
rect 18808 8336 19176 8345
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 18808 8287 19176 8296
rect 18604 8119 18644 8128
rect 19276 8168 19316 8620
rect 19276 8119 19316 8128
rect 18796 7916 18836 7925
rect 18796 7748 18836 7876
rect 18796 7244 18836 7708
rect 18796 7195 18836 7204
rect 18700 7160 18740 7169
rect 18700 6824 18740 7120
rect 18700 6775 18740 6784
rect 18808 6824 19176 6833
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 18808 6775 19176 6784
rect 19468 6572 19508 8632
rect 19564 8336 19604 9220
rect 19660 8924 19700 11764
rect 19852 9596 19892 11764
rect 20044 10100 20084 11764
rect 19852 9547 19892 9556
rect 19948 10060 20084 10100
rect 19660 8875 19700 8884
rect 19756 9512 19796 9521
rect 19756 8840 19796 9472
rect 19852 9344 19892 9439
rect 19852 9295 19892 9304
rect 19852 9176 19892 9185
rect 19852 9041 19892 9136
rect 19948 8924 19988 10060
rect 20236 9680 20276 11764
rect 20236 9631 20276 9640
rect 20428 9260 20468 11764
rect 20620 9344 20660 11764
rect 20620 9295 20660 9304
rect 20716 9512 20756 9521
rect 20428 9220 20564 9260
rect 20048 9092 20416 9101
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20048 9043 20416 9052
rect 19948 8875 19988 8884
rect 20044 8924 20084 8933
rect 19756 8791 19796 8800
rect 20044 8660 20084 8884
rect 20524 8924 20564 9220
rect 20716 9092 20756 9472
rect 20716 9043 20756 9052
rect 20524 8875 20564 8884
rect 20812 8924 20852 11764
rect 20812 8875 20852 8884
rect 20908 9344 20948 9353
rect 19948 8620 20084 8660
rect 20620 8756 20660 8765
rect 20908 8756 20948 9304
rect 21004 9260 21044 11764
rect 21196 9680 21236 11764
rect 21196 9631 21236 9640
rect 21388 9596 21428 11764
rect 21388 9547 21428 9556
rect 21004 9211 21044 9220
rect 19564 8287 19604 8296
rect 19756 8504 19796 8513
rect 19660 8168 19700 8177
rect 19660 7496 19700 8128
rect 19660 7447 19700 7456
rect 19756 7328 19796 8464
rect 19948 8504 19988 8620
rect 19948 8455 19988 8464
rect 20140 8504 20180 8599
rect 20140 8455 20180 8464
rect 19852 8420 19892 8429
rect 19852 8252 19892 8380
rect 20044 8420 20084 8429
rect 19852 8203 19892 8212
rect 19948 8336 19988 8345
rect 19948 8084 19988 8296
rect 20044 8252 20084 8380
rect 20140 8252 20180 8261
rect 20044 8212 20140 8252
rect 20140 8203 20180 8212
rect 20140 8084 20180 8093
rect 19948 8044 20140 8084
rect 20140 8035 20180 8044
rect 19948 7580 19988 7589
rect 19948 7412 19988 7540
rect 20048 7580 20416 7589
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20048 7531 20416 7540
rect 20524 7580 20564 7589
rect 20524 7496 20564 7540
rect 20524 7445 20564 7456
rect 19948 7363 19988 7372
rect 19756 7279 19796 7288
rect 19468 6523 19508 6532
rect 20524 6152 20564 6161
rect 20048 6068 20416 6077
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20048 6019 20416 6028
rect 20524 5984 20564 6112
rect 20524 5935 20564 5944
rect 18700 5900 18740 5909
rect 18700 5765 18740 5860
rect 18808 5312 19176 5321
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 18808 5263 19176 5272
rect 20048 4556 20416 4565
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20048 4507 20416 4516
rect 19084 4220 19124 4229
rect 19276 4220 19316 4229
rect 19124 4180 19276 4220
rect 19084 4171 19124 4180
rect 18808 3800 19176 3809
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 18808 3751 19176 3760
rect 19276 3464 19316 4180
rect 19276 3415 19316 3424
rect 20140 3968 20180 3977
rect 20140 3212 20180 3928
rect 19948 3172 20180 3212
rect 19948 3044 19988 3172
rect 19948 2995 19988 3004
rect 20048 3044 20416 3053
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20048 2995 20416 3004
rect 18124 2575 18164 2584
rect 18700 2960 18740 2969
rect 17452 2155 17492 2164
rect 18700 80 18740 2920
rect 20620 2792 20660 8716
rect 20812 8716 20948 8756
rect 21292 9176 21332 9185
rect 20716 7916 20756 7925
rect 20716 6992 20756 7876
rect 20716 4220 20756 6952
rect 20716 4171 20756 4180
rect 20812 3380 20852 8716
rect 21004 8672 21044 8681
rect 20908 8588 20948 8597
rect 20908 8420 20948 8548
rect 20908 8371 20948 8380
rect 20812 3331 20852 3340
rect 20620 2743 20660 2752
rect 21004 2540 21044 8632
rect 21196 8672 21236 8681
rect 21196 7916 21236 8632
rect 21196 7867 21236 7876
rect 21196 4052 21236 4061
rect 21196 3464 21236 4012
rect 21292 3968 21332 9136
rect 21292 3919 21332 3928
rect 21484 9092 21524 9101
rect 21196 3415 21236 3424
rect 21484 3464 21524 9052
rect 21580 8672 21620 11764
rect 21772 9596 21812 11764
rect 21772 9547 21812 9556
rect 21868 9428 21908 9437
rect 21580 8623 21620 8632
rect 21676 9260 21716 9269
rect 21676 7244 21716 9220
rect 21868 9176 21908 9388
rect 21868 9127 21908 9136
rect 21676 7195 21716 7204
rect 21772 9092 21812 9101
rect 21484 3296 21524 3424
rect 21772 3380 21812 9052
rect 21964 8756 22004 11764
rect 21964 8707 22004 8716
rect 22060 9764 22100 9773
rect 22060 4388 22100 9724
rect 22156 9596 22196 11764
rect 22156 9547 22196 9556
rect 22252 10100 22292 10109
rect 22252 8756 22292 10060
rect 22348 9596 22388 11764
rect 22348 9547 22388 9556
rect 22540 9512 22580 11764
rect 22732 9680 22772 11764
rect 22732 9631 22772 9640
rect 22828 10016 22868 10025
rect 22540 9463 22580 9472
rect 22348 9344 22388 9353
rect 22348 9209 22388 9304
rect 22732 9260 22772 9269
rect 22252 8707 22292 8716
rect 22636 8672 22676 8681
rect 22444 6992 22484 7001
rect 22444 4892 22484 6952
rect 22444 4843 22484 4852
rect 22060 4339 22100 4348
rect 22540 4472 22580 4481
rect 22156 4220 22196 4229
rect 21772 3331 21812 3340
rect 21964 3464 22004 3473
rect 21964 3329 22004 3424
rect 22156 3464 22196 4180
rect 22540 4220 22580 4432
rect 22540 4171 22580 4180
rect 22156 3415 22196 3424
rect 22636 3464 22676 8632
rect 21484 3247 21524 3256
rect 21004 2491 21044 2500
rect 22540 2708 22580 2717
rect 22540 2540 22580 2668
rect 22636 2624 22676 3424
rect 22732 3464 22772 9220
rect 22828 8756 22868 9976
rect 22924 10016 22964 11764
rect 23116 10100 23156 11764
rect 23116 10060 23252 10100
rect 22924 9967 22964 9976
rect 23020 9932 23060 9941
rect 23020 9848 23060 9892
rect 22828 8707 22868 8716
rect 22924 9808 23060 9848
rect 22732 3380 22772 3424
rect 22732 3329 22772 3340
rect 22828 4472 22868 4481
rect 22732 3128 22772 3137
rect 22732 2960 22772 3088
rect 22732 2911 22772 2920
rect 22636 2575 22676 2584
rect 22828 2624 22868 4432
rect 22924 4220 22964 9808
rect 23116 9764 23156 9773
rect 23116 9680 23156 9724
rect 23116 9629 23156 9640
rect 23212 6656 23252 10060
rect 23212 6607 23252 6616
rect 23308 6404 23348 11764
rect 23404 10016 23444 10025
rect 23404 8672 23444 9976
rect 23500 9596 23540 11764
rect 23596 9932 23636 9941
rect 23596 9797 23636 9892
rect 23500 9547 23540 9556
rect 23692 9596 23732 11764
rect 23692 9547 23732 9556
rect 23788 9848 23828 9857
rect 23788 9260 23828 9808
rect 23884 9596 23924 11764
rect 23884 9547 23924 9556
rect 24076 9512 24116 11764
rect 24076 9463 24116 9472
rect 24268 9512 24308 11764
rect 24460 9596 24500 11764
rect 24460 9547 24500 9556
rect 24652 9596 24692 11764
rect 24844 9680 24884 11764
rect 24844 9631 24884 9640
rect 24652 9547 24692 9556
rect 24268 9463 24308 9472
rect 25036 9428 25076 11764
rect 25132 9764 25172 9773
rect 25132 9629 25172 9724
rect 25036 9379 25076 9388
rect 23788 9211 23828 9220
rect 24364 9344 24404 9353
rect 23500 9176 23540 9185
rect 23500 8756 23540 9136
rect 23500 8707 23540 8716
rect 24172 8840 24212 8849
rect 23404 8623 23444 8632
rect 23692 7076 23732 7087
rect 23692 6992 23732 7036
rect 23692 6943 23732 6952
rect 24172 6824 24212 8800
rect 24364 8756 24404 9304
rect 24652 9344 24692 9353
rect 24692 9304 24788 9344
rect 24652 9295 24692 9304
rect 24364 8707 24404 8716
rect 24460 8840 24500 8849
rect 24172 6775 24212 6784
rect 23308 6355 23348 6364
rect 23788 6404 23828 6413
rect 23692 6068 23732 6077
rect 23692 5984 23732 6028
rect 23692 5933 23732 5944
rect 23020 4892 23060 4901
rect 23020 4388 23060 4852
rect 23212 4724 23252 4733
rect 23252 4684 23348 4724
rect 23212 4675 23252 4684
rect 23308 4388 23348 4684
rect 23060 4348 23156 4388
rect 23020 4339 23060 4348
rect 22924 4171 22964 4180
rect 22924 4052 22964 4061
rect 22924 3044 22964 4012
rect 23116 4052 23156 4348
rect 23116 4003 23156 4012
rect 23212 4304 23252 4313
rect 23020 3632 23060 3641
rect 23020 3497 23060 3592
rect 23116 3548 23156 3557
rect 23116 3413 23156 3508
rect 22924 3004 23060 3044
rect 23020 2708 23060 3004
rect 23020 2659 23060 2668
rect 22828 2575 22868 2584
rect 22540 2491 22580 2500
rect 23212 2540 23252 4264
rect 23308 2708 23348 4348
rect 23788 4556 23828 6364
rect 24460 5144 24500 8800
rect 24460 5095 24500 5104
rect 24076 4724 24116 4733
rect 23500 4220 23540 4229
rect 23404 4136 23444 4145
rect 23404 2792 23444 4096
rect 23500 3716 23540 4180
rect 23692 4220 23732 4229
rect 23500 3667 23540 3676
rect 23596 3968 23636 3977
rect 23596 3464 23636 3928
rect 23596 3415 23636 3424
rect 23404 2743 23444 2752
rect 23308 2659 23348 2668
rect 23692 2708 23732 4180
rect 23788 4220 23828 4516
rect 23980 4556 24020 4565
rect 23980 4304 24020 4516
rect 23980 4255 24020 4264
rect 23788 4171 23828 4180
rect 23884 4220 23924 4229
rect 23788 4052 23828 4061
rect 23884 4052 23924 4180
rect 23828 4012 23924 4052
rect 23980 4052 24020 4061
rect 23788 4003 23828 4012
rect 23884 3884 23924 3893
rect 23788 3380 23828 3389
rect 23788 3296 23828 3340
rect 23788 3245 23828 3256
rect 23692 2659 23732 2668
rect 23212 2491 23252 2500
rect 23020 2456 23060 2465
rect 23308 2456 23348 2465
rect 23060 2416 23156 2456
rect 23020 2407 23060 2416
rect 23116 2372 23156 2416
rect 23308 2372 23348 2416
rect 23116 2332 23348 2372
rect 18808 2288 19176 2297
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 18808 2239 19176 2248
rect 22156 2204 22196 2213
rect 20048 1532 20416 1541
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20048 1483 20416 1492
rect 20428 860 20468 869
rect 20428 80 20468 820
rect 22156 80 22196 2164
rect 23884 80 23924 3844
rect 23980 3632 24020 4012
rect 23980 3583 24020 3592
rect 24076 3380 24116 4684
rect 24364 4388 24404 4397
rect 24076 3331 24116 3340
rect 24172 4220 24212 4229
rect 24172 2540 24212 4180
rect 24268 4136 24308 4145
rect 24268 3212 24308 4096
rect 24364 3296 24404 4348
rect 24556 4052 24596 4061
rect 24596 4012 24692 4052
rect 24556 4003 24596 4012
rect 24364 3247 24404 3256
rect 24268 3163 24308 3172
rect 24172 2491 24212 2500
rect 24460 2960 24500 2969
rect 24460 1868 24500 2920
rect 24460 1819 24500 1828
rect 24652 1784 24692 4012
rect 24748 3548 24788 9304
rect 24844 9260 24884 9269
rect 24844 8840 24884 9220
rect 24844 8791 24884 8800
rect 25228 8672 25268 11764
rect 25420 9764 25460 11764
rect 25420 9715 25460 9724
rect 25612 8756 25652 11764
rect 25804 9764 25844 11764
rect 25804 9715 25844 9724
rect 25612 8707 25652 8716
rect 25708 9512 25748 9521
rect 25228 8623 25268 8632
rect 25708 8504 25748 9472
rect 25900 9344 25940 9353
rect 25804 9260 25844 9269
rect 25804 9176 25844 9220
rect 25804 9125 25844 9136
rect 25900 9176 25940 9304
rect 25900 9127 25940 9136
rect 25996 8672 26036 11764
rect 26188 9428 26228 11764
rect 26284 9932 26324 9941
rect 26284 9680 26324 9892
rect 26284 9631 26324 9640
rect 26188 9379 26228 9388
rect 26188 9092 26228 9101
rect 26188 8756 26228 9052
rect 26188 8707 26228 8716
rect 26380 8756 26420 11764
rect 26380 8707 26420 8716
rect 26476 9260 26516 9269
rect 25996 8623 26036 8632
rect 25324 8464 25748 8504
rect 26092 8504 26132 8513
rect 24940 7580 24980 7589
rect 24748 3380 24788 3508
rect 24844 4892 24884 4901
rect 24844 3464 24884 4852
rect 24940 3632 24980 7540
rect 25324 4892 25364 8464
rect 25996 8420 26036 8429
rect 25708 8380 25996 8420
rect 25612 8336 25652 8345
rect 25612 8000 25652 8296
rect 25708 8252 25748 8380
rect 25996 8371 26036 8380
rect 25708 8203 25748 8212
rect 25612 7951 25652 7960
rect 25420 7664 25460 7673
rect 25420 7496 25460 7624
rect 25420 7447 25460 7456
rect 25516 7412 25556 7421
rect 25516 7160 25556 7372
rect 25516 7111 25556 7120
rect 25324 4843 25364 4852
rect 25612 6740 25652 6749
rect 25036 4304 25076 4313
rect 25036 3884 25076 4264
rect 25036 3835 25076 3844
rect 25132 3968 25172 3977
rect 24940 3583 24980 3592
rect 25036 3716 25076 3725
rect 25036 3548 25076 3676
rect 25036 3499 25076 3508
rect 24844 3415 24884 3424
rect 24748 3331 24788 3340
rect 24652 1735 24692 1744
rect 24748 3044 24788 3053
rect 24748 860 24788 3004
rect 25132 2120 25172 3928
rect 25612 3632 25652 6700
rect 25804 6068 25844 6077
rect 25804 5900 25844 6028
rect 25804 5851 25844 5860
rect 25612 3464 25652 3592
rect 25612 3415 25652 3424
rect 25900 3968 25940 3977
rect 25900 3044 25940 3928
rect 26092 3632 26132 8464
rect 26188 8000 26228 8009
rect 26188 6404 26228 7960
rect 26476 7412 26516 9220
rect 26572 9260 26612 11764
rect 26572 9211 26612 9220
rect 26764 8924 26804 11764
rect 26956 10016 26996 11764
rect 26956 9967 26996 9976
rect 26956 9596 26996 9605
rect 26860 9176 26900 9185
rect 26860 9041 26900 9136
rect 26764 8875 26804 8884
rect 26956 8924 26996 9556
rect 27148 9260 27188 11764
rect 27340 10100 27380 11764
rect 27532 10184 27572 11764
rect 27532 10144 27668 10184
rect 27340 10060 27476 10100
rect 27340 9428 27380 9437
rect 26956 8875 26996 8884
rect 27052 9220 27188 9260
rect 27244 9388 27340 9428
rect 26572 8756 26612 8851
rect 26572 8707 26612 8716
rect 26476 7363 26516 7372
rect 27052 6656 27092 9220
rect 27052 6607 27092 6616
rect 27148 7244 27188 7253
rect 27148 6908 27188 7204
rect 26188 6355 26228 6364
rect 26092 3583 26132 3592
rect 27148 6320 27188 6868
rect 27148 4976 27188 6280
rect 27148 3380 27188 4936
rect 27244 3968 27284 9388
rect 27340 9379 27380 9388
rect 27340 9008 27380 9017
rect 27340 7748 27380 8968
rect 27436 8336 27476 10060
rect 27436 8287 27476 8296
rect 27532 8588 27572 8597
rect 27532 7916 27572 8548
rect 27628 8504 27668 10144
rect 27724 9428 27764 11764
rect 27916 10100 27956 11764
rect 27916 10051 27956 10060
rect 27820 10016 27860 10025
rect 27820 9764 27860 9976
rect 27820 9715 27860 9724
rect 28108 9512 28148 11764
rect 28300 9596 28340 11764
rect 28492 9680 28532 11764
rect 28492 9631 28532 9640
rect 28300 9547 28340 9556
rect 28108 9463 28148 9472
rect 28684 9428 28724 11764
rect 28876 9764 28916 11764
rect 28876 9715 28916 9724
rect 28972 9848 29012 9857
rect 28972 9596 29012 9808
rect 28972 9547 29012 9556
rect 27724 9388 27860 9428
rect 27628 8455 27668 8464
rect 27724 9260 27764 9269
rect 27532 7867 27572 7876
rect 27340 7699 27380 7708
rect 27628 7160 27668 7169
rect 27340 6824 27380 6833
rect 27340 6656 27380 6784
rect 27340 6607 27380 6616
rect 27628 6656 27668 7120
rect 27628 6607 27668 6616
rect 27532 6404 27572 6413
rect 27532 6269 27572 6364
rect 27628 5228 27668 5237
rect 27628 4892 27668 5188
rect 27628 4136 27668 4852
rect 27724 4220 27764 9220
rect 27820 6488 27860 9388
rect 28684 9379 28724 9388
rect 27820 6439 27860 6448
rect 27916 9344 27956 9353
rect 27820 6068 27860 6077
rect 27820 5900 27860 6028
rect 27820 5851 27860 5860
rect 27916 4472 27956 9304
rect 28396 8840 28436 8849
rect 28300 7832 28340 7841
rect 28204 7664 28244 7673
rect 28204 6992 28244 7624
rect 28204 6943 28244 6952
rect 28300 7328 28340 7792
rect 28300 6656 28340 7288
rect 28396 7244 28436 8800
rect 28780 8840 28820 8935
rect 28780 8791 28820 8800
rect 28780 8672 28820 8681
rect 29068 8672 29108 11764
rect 29260 9596 29300 11764
rect 29452 9848 29492 11764
rect 29452 9799 29492 9808
rect 29260 9547 29300 9556
rect 29644 9428 29684 11764
rect 29548 9388 29684 9428
rect 29740 9848 29780 9857
rect 29740 9428 29780 9808
rect 28820 8632 29012 8660
rect 28780 8620 29012 8632
rect 29068 8623 29108 8632
rect 29164 9176 29204 9185
rect 28684 8504 28724 8599
rect 28972 8504 29012 8620
rect 28972 8464 29108 8504
rect 28684 8455 28724 8464
rect 28492 8420 28532 8429
rect 28492 8336 28532 8380
rect 28492 8285 28532 8296
rect 28684 8336 28724 8345
rect 28588 8168 28628 8177
rect 28588 7832 28628 8128
rect 28684 8084 28724 8296
rect 28684 8035 28724 8044
rect 28876 8168 28916 8177
rect 28876 7832 28916 8128
rect 29068 8084 29108 8464
rect 29068 8035 29108 8044
rect 28588 7792 28916 7832
rect 28972 8000 29012 8009
rect 28684 7664 28724 7673
rect 28492 7580 28532 7589
rect 28492 7445 28532 7540
rect 28684 7328 28724 7624
rect 28780 7580 28820 7591
rect 28780 7496 28820 7540
rect 28780 7447 28820 7456
rect 28972 7496 29012 7960
rect 29164 8000 29204 9136
rect 29356 8756 29396 8851
rect 29356 8707 29396 8716
rect 29164 7951 29204 7960
rect 29260 8504 29300 8513
rect 28972 7447 29012 7456
rect 29068 7916 29108 7925
rect 28684 7279 28724 7288
rect 28876 7412 28916 7421
rect 28876 7277 28916 7372
rect 29068 7328 29108 7876
rect 29068 7279 29108 7288
rect 29164 7748 29204 7757
rect 28396 7204 28532 7244
rect 28492 7160 28532 7204
rect 28492 7111 28532 7120
rect 28780 7160 28820 7169
rect 28396 7076 28436 7085
rect 28396 6992 28436 7036
rect 28780 7025 28820 7120
rect 29068 6992 29108 7001
rect 28396 6952 28628 6992
rect 28588 6908 28628 6952
rect 28684 6908 28724 6917
rect 28588 6868 28684 6908
rect 28684 6859 28724 6868
rect 29068 6857 29108 6952
rect 28300 6607 28340 6616
rect 28780 6488 28820 6497
rect 28780 6068 28820 6448
rect 29164 6488 29204 7708
rect 29164 6439 29204 6448
rect 28876 6236 28916 6245
rect 28876 6101 28916 6196
rect 28780 6019 28820 6028
rect 28012 5984 28052 5993
rect 28012 5849 28052 5944
rect 27916 4423 27956 4432
rect 27724 4171 27764 4180
rect 27628 4087 27668 4096
rect 27244 3919 27284 3928
rect 27340 4052 27380 4061
rect 27148 3331 27188 3340
rect 25900 2995 25940 3004
rect 25132 2071 25172 2080
rect 25612 2120 25652 2129
rect 24748 811 24788 820
rect 25612 80 25652 2080
rect 27340 80 27380 4012
rect 29260 3716 29300 8464
rect 29356 8084 29396 8093
rect 29356 7412 29396 8044
rect 29356 7363 29396 7372
rect 29356 6908 29396 6917
rect 29548 6908 29588 9388
rect 29740 9379 29780 9388
rect 29644 8840 29684 8849
rect 29644 8672 29684 8800
rect 29644 8623 29684 8632
rect 29836 8504 29876 11764
rect 29932 9764 29972 9773
rect 29932 9512 29972 9724
rect 30028 9680 30068 11764
rect 30220 11444 30260 11764
rect 30220 11395 30260 11404
rect 30412 9764 30452 11764
rect 30604 11192 30644 11764
rect 30604 11143 30644 11152
rect 30412 9724 30644 9764
rect 30316 9680 30356 9689
rect 30028 9640 30164 9680
rect 29932 9463 29972 9472
rect 29836 8455 29876 8464
rect 30028 9344 30068 9353
rect 29740 8420 29780 8429
rect 29740 8168 29780 8380
rect 29740 8119 29780 8128
rect 29396 6868 29492 6908
rect 29356 6859 29396 6868
rect 29356 6740 29396 6749
rect 29452 6740 29492 6868
rect 29548 6859 29588 6868
rect 29644 8084 29684 8093
rect 29548 6740 29588 6749
rect 29452 6700 29548 6740
rect 29356 6488 29396 6700
rect 29548 6691 29588 6700
rect 29356 6439 29396 6448
rect 29548 6404 29588 6413
rect 29644 6404 29684 8044
rect 29836 8000 29876 8009
rect 29740 7916 29780 7925
rect 29740 7496 29780 7876
rect 29740 7447 29780 7456
rect 29836 7160 29876 7960
rect 29836 7111 29876 7120
rect 29932 7832 29972 7841
rect 29932 6992 29972 7792
rect 29932 6943 29972 6952
rect 30028 7076 30068 9304
rect 30124 8252 30164 9640
rect 30356 9640 30452 9680
rect 30316 9631 30356 9640
rect 30220 8420 30260 8429
rect 30220 8285 30260 8380
rect 30124 8203 30164 8212
rect 30124 7832 30164 7841
rect 30124 7328 30164 7792
rect 30316 7832 30356 7841
rect 30316 7496 30356 7792
rect 30316 7447 30356 7456
rect 30124 7193 30164 7288
rect 29836 6656 29876 6665
rect 29836 6488 29876 6616
rect 29836 6439 29876 6448
rect 29588 6364 29684 6404
rect 29548 6355 29588 6364
rect 30028 6320 30068 7036
rect 30316 6992 30356 7001
rect 30316 6404 30356 6952
rect 30412 6488 30452 9640
rect 30508 7916 30548 7925
rect 30508 6656 30548 7876
rect 30604 7496 30644 9724
rect 30796 7832 30836 11764
rect 30796 7783 30836 7792
rect 30892 9344 30932 9353
rect 30604 7447 30644 7456
rect 30700 7748 30740 7757
rect 30508 6607 30548 6616
rect 30604 7328 30644 7368
rect 30604 7244 30644 7288
rect 30412 6439 30452 6448
rect 30316 6355 30356 6364
rect 30028 6271 30068 6280
rect 29740 6236 29780 6245
rect 29740 6152 29780 6196
rect 29740 6101 29780 6112
rect 30220 5984 30260 5993
rect 30220 5849 30260 5944
rect 30604 5144 30644 7204
rect 30604 5095 30644 5104
rect 29260 3667 29300 3676
rect 27436 3632 27476 3641
rect 27436 3380 27476 3592
rect 27436 3331 27476 3340
rect 29068 3632 29108 3641
rect 29068 80 29108 3592
rect 30700 2036 30740 7708
rect 30892 7748 30932 9304
rect 30988 9176 31028 11764
rect 31180 9680 31220 11764
rect 31180 9631 31220 9640
rect 31372 9596 31412 11764
rect 31372 9547 31412 9556
rect 31468 10016 31508 10025
rect 30988 9127 31028 9136
rect 30796 7412 30836 7423
rect 30796 7328 30836 7372
rect 30796 7279 30836 7288
rect 30892 7244 30932 7708
rect 30892 7195 30932 7204
rect 31468 8000 31508 9976
rect 31564 9680 31604 11764
rect 31564 9631 31604 9640
rect 31756 9596 31796 11764
rect 31948 9764 31988 11764
rect 31948 9715 31988 9724
rect 31756 9547 31796 9556
rect 31756 9428 31796 9437
rect 31796 9388 31892 9428
rect 31756 9379 31796 9388
rect 31660 8756 31700 8765
rect 31564 8336 31604 8345
rect 31564 8084 31604 8296
rect 31564 8035 31604 8044
rect 31468 7160 31508 7960
rect 31660 8000 31700 8716
rect 31756 8000 31796 8009
rect 31660 7960 31756 8000
rect 31564 7244 31604 7253
rect 31660 7244 31700 7960
rect 31756 7951 31796 7960
rect 31604 7204 31700 7244
rect 31756 7244 31796 7253
rect 31564 7195 31604 7204
rect 31756 7160 31796 7204
rect 31468 7111 31508 7120
rect 31660 7120 31796 7160
rect 30988 6572 31028 6581
rect 30988 6068 31028 6532
rect 31660 6488 31700 7120
rect 31660 6439 31700 6448
rect 31372 6320 31412 6329
rect 31084 6152 31124 6161
rect 31276 6152 31316 6161
rect 31124 6112 31276 6152
rect 31084 6103 31124 6112
rect 31276 6103 31316 6112
rect 30988 6019 31028 6028
rect 31372 2900 31412 6280
rect 31468 6068 31508 6077
rect 31468 5933 31508 6028
rect 31852 3296 31892 9388
rect 32140 8924 32180 11764
rect 32332 9344 32372 11764
rect 32332 9295 32372 9304
rect 32140 8875 32180 8884
rect 32524 8924 32564 11764
rect 32716 9764 32756 11764
rect 32716 9715 32756 9724
rect 32716 9512 32756 9521
rect 32716 9008 32756 9472
rect 32716 8959 32756 8968
rect 32524 8875 32564 8884
rect 32908 8924 32948 11764
rect 33100 11444 33140 11764
rect 33100 11404 33236 11444
rect 33004 9932 33044 9941
rect 33004 9512 33044 9892
rect 33004 9463 33044 9472
rect 33100 9596 33140 9605
rect 32908 8875 32948 8884
rect 31948 8588 31988 8597
rect 31948 8168 31988 8548
rect 31948 8119 31988 8128
rect 32620 8252 32660 8261
rect 32236 8000 32276 8009
rect 32236 7748 32276 7960
rect 32236 7699 32276 7708
rect 32428 7748 32468 7757
rect 32428 7580 32468 7708
rect 32428 7531 32468 7540
rect 32620 7580 32660 8212
rect 32620 7531 32660 7540
rect 32140 7412 32180 7421
rect 32140 7244 32180 7372
rect 32140 7195 32180 7204
rect 32908 5900 32948 5909
rect 32908 5765 32948 5860
rect 31852 3247 31892 3256
rect 33100 3212 33140 9556
rect 33196 9260 33236 11404
rect 33196 9211 33236 9220
rect 33292 8924 33332 11764
rect 33292 8875 33332 8884
rect 33388 9932 33428 9941
rect 33388 8672 33428 9892
rect 33484 9680 33524 11764
rect 33484 9631 33524 9640
rect 33580 10016 33620 10025
rect 33580 9512 33620 9976
rect 33580 9463 33620 9472
rect 33484 9344 33524 9353
rect 33484 9008 33524 9304
rect 33484 8959 33524 8968
rect 33676 8924 33716 11764
rect 33868 10016 33908 11764
rect 34060 10184 34100 11764
rect 34252 10352 34292 11764
rect 34252 10303 34292 10312
rect 34060 10144 34388 10184
rect 33868 9967 33908 9976
rect 33928 9848 34296 9857
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 33928 9799 34296 9808
rect 34252 9680 34292 9689
rect 34060 9596 34100 9605
rect 34060 9428 34100 9556
rect 34060 9379 34100 9388
rect 34252 9260 34292 9640
rect 34252 9211 34292 9220
rect 33676 8875 33716 8884
rect 34348 8924 34388 10144
rect 34348 8875 34388 8884
rect 34444 8840 34484 11764
rect 34540 10352 34580 10361
rect 34540 9344 34580 10312
rect 34636 9764 34676 11764
rect 34636 9715 34676 9724
rect 34732 10016 34772 10025
rect 34636 9512 34676 9521
rect 34732 9512 34772 9976
rect 34828 9596 34868 11764
rect 35020 9680 35060 11764
rect 38860 11444 38900 11453
rect 37420 9932 37460 9941
rect 37420 9848 37460 9892
rect 37420 9797 37460 9808
rect 35020 9631 35060 9640
rect 35404 9764 35444 9773
rect 35404 9680 35444 9724
rect 35404 9629 35444 9640
rect 36172 9680 36212 9689
rect 34828 9547 34868 9556
rect 36172 9545 36212 9640
rect 36460 9680 36500 9691
rect 36364 9596 36404 9605
rect 34676 9472 34772 9512
rect 35020 9512 35060 9521
rect 34636 9463 34676 9472
rect 34540 9295 34580 9304
rect 34444 8791 34484 8800
rect 33388 8623 33428 8632
rect 33772 8672 33812 8681
rect 33772 8588 33812 8632
rect 33772 8537 33812 8548
rect 34540 8672 34580 8681
rect 33928 8336 34296 8345
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 33928 8287 34296 8296
rect 34540 8084 34580 8632
rect 34636 8588 34676 8597
rect 34676 8548 34772 8588
rect 34636 8539 34676 8548
rect 34540 8035 34580 8044
rect 34348 8000 34388 8009
rect 33928 6824 34296 6833
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 33928 6775 34296 6784
rect 33928 5312 34296 5321
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 33928 5263 34296 5272
rect 33292 4136 33332 4145
rect 33292 4001 33332 4096
rect 33928 3800 34296 3809
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 33928 3751 34296 3760
rect 33100 3163 33140 3172
rect 30700 1987 30740 1996
rect 31276 2860 31412 2900
rect 30796 148 31124 188
rect 30796 80 30836 148
rect 10100 64 10120 80
rect 10040 0 10120 64
rect 11768 0 11848 80
rect 13496 0 13576 80
rect 15224 0 15304 80
rect 16952 0 17032 80
rect 18680 0 18760 80
rect 20408 0 20488 80
rect 22136 0 22216 80
rect 23864 0 23944 80
rect 25592 0 25672 80
rect 27320 0 27400 80
rect 29048 0 29128 80
rect 30776 0 30856 80
rect 31084 60 31124 148
rect 31276 60 31316 2860
rect 33928 2288 34296 2297
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 33928 2239 34296 2248
rect 34348 1448 34388 7960
rect 34636 6488 34676 6497
rect 34636 5816 34676 6448
rect 34636 5767 34676 5776
rect 34444 5732 34484 5741
rect 34444 5564 34484 5692
rect 34636 5564 34676 5573
rect 34444 5524 34636 5564
rect 34636 5515 34676 5524
rect 34732 2900 34772 8548
rect 35020 8168 35060 9472
rect 35692 9512 35732 9521
rect 35404 9428 35444 9437
rect 35404 9293 35444 9388
rect 35596 9428 35636 9437
rect 35500 9260 35540 9355
rect 35500 9211 35540 9220
rect 35168 9092 35536 9101
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35168 9043 35536 9052
rect 35404 8924 35444 8933
rect 35404 8672 35444 8884
rect 35404 8623 35444 8632
rect 35020 8119 35060 8128
rect 35308 8588 35348 8597
rect 35308 8168 35348 8548
rect 35308 8119 35348 8128
rect 35500 8504 35540 8513
rect 35500 8000 35540 8464
rect 35020 7960 35540 8000
rect 35020 7580 35060 7960
rect 35020 7531 35060 7540
rect 35168 7580 35536 7589
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35168 7531 35536 7540
rect 35596 7076 35636 9388
rect 35692 8840 35732 9472
rect 36268 9512 36308 9521
rect 35788 9428 35828 9437
rect 35788 8924 35828 9388
rect 36076 9428 36116 9437
rect 35788 8875 35828 8884
rect 35884 9176 35924 9185
rect 35692 8791 35732 8800
rect 35692 8504 35732 8513
rect 35692 8252 35732 8464
rect 35692 8203 35732 8212
rect 35788 8168 35828 8177
rect 35788 7580 35828 8128
rect 35884 8084 35924 9136
rect 35980 9176 36020 9185
rect 35980 8924 36020 9136
rect 35980 8875 36020 8884
rect 35884 8035 35924 8044
rect 35788 7531 35828 7540
rect 35980 7916 36020 7925
rect 35596 7027 35636 7036
rect 35788 6992 35828 7001
rect 35020 6908 35060 6917
rect 35308 6908 35348 6917
rect 35060 6868 35308 6908
rect 35020 6859 35060 6868
rect 35308 6859 35348 6868
rect 35020 6740 35060 6749
rect 35020 6605 35060 6700
rect 35788 6740 35828 6952
rect 35788 6691 35828 6700
rect 34924 6488 34964 6583
rect 35116 6572 35156 6581
rect 35308 6572 35348 6581
rect 35156 6532 35308 6572
rect 35116 6523 35156 6532
rect 35308 6523 35348 6532
rect 34924 6439 34964 6448
rect 35692 6488 35732 6497
rect 35020 6404 35060 6413
rect 34924 6320 34964 6329
rect 34924 6185 34964 6280
rect 35020 6068 35060 6364
rect 35020 6019 35060 6028
rect 35168 6068 35536 6077
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35168 6019 35536 6028
rect 35692 5900 35732 6448
rect 35884 6404 35924 6413
rect 35884 6269 35924 6364
rect 35692 5851 35732 5860
rect 35404 5816 35444 5825
rect 35596 5816 35636 5825
rect 35444 5776 35596 5816
rect 35404 5767 35444 5776
rect 35596 5767 35636 5776
rect 35168 4556 35536 4565
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35168 4507 35536 4516
rect 35884 4220 35924 4229
rect 35884 3884 35924 4180
rect 35884 3835 35924 3844
rect 35168 3044 35536 3053
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35168 2995 35536 3004
rect 34732 2860 34868 2900
rect 34828 2792 34868 2860
rect 34828 2743 34868 2752
rect 35168 1532 35536 1541
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35168 1483 35536 1492
rect 34252 1408 34388 1448
rect 32524 860 32564 869
rect 32524 80 32564 820
rect 34252 80 34292 1408
rect 35980 80 36020 7876
rect 36076 3968 36116 9388
rect 36172 9428 36212 9437
rect 36172 9260 36212 9388
rect 36172 9211 36212 9220
rect 36076 3919 36116 3928
rect 36172 9008 36212 9017
rect 36172 3884 36212 8968
rect 36268 6488 36308 9472
rect 36364 9260 36404 9556
rect 36460 9596 36500 9640
rect 36460 9547 36500 9556
rect 37900 9428 37940 9437
rect 36364 9211 36404 9220
rect 37324 9344 37364 9353
rect 37324 8924 37364 9304
rect 37324 8875 37364 8884
rect 37420 9344 37460 9353
rect 36268 6439 36308 6448
rect 36364 8588 36404 8597
rect 36172 3835 36212 3844
rect 36364 3464 36404 8548
rect 36748 8420 36788 8429
rect 36748 7496 36788 8380
rect 36748 7447 36788 7456
rect 37036 7832 37076 7841
rect 36460 6488 36500 6497
rect 36460 5984 36500 6448
rect 36460 5935 36500 5944
rect 37036 4304 37076 7792
rect 37132 6320 37172 6329
rect 37132 6185 37172 6280
rect 37036 4255 37076 4264
rect 37420 3800 37460 9304
rect 37804 8840 37844 8849
rect 37708 8168 37748 8177
rect 37708 7748 37748 8128
rect 37708 7699 37748 7708
rect 37420 3751 37460 3760
rect 37708 7160 37748 7169
rect 36364 3415 36404 3424
rect 37708 80 37748 7120
rect 37804 3968 37844 8800
rect 37900 8672 37940 9388
rect 38860 9092 38900 11404
rect 38860 9043 38900 9052
rect 38956 11192 38996 11201
rect 38956 9008 38996 11152
rect 44236 11024 44276 11033
rect 43756 10688 43796 10697
rect 43276 10352 43316 10361
rect 42892 10100 42932 10109
rect 40492 10016 40532 10025
rect 38956 8959 38996 8968
rect 39244 9932 39284 9941
rect 37900 8623 37940 8632
rect 38860 8756 38900 8765
rect 38380 8504 38420 8513
rect 38380 8369 38420 8464
rect 38860 8504 38900 8716
rect 38860 8455 38900 8464
rect 38188 8000 38228 8009
rect 38092 7832 38132 7841
rect 38092 7160 38132 7792
rect 38188 7244 38228 7960
rect 38860 8000 38900 8009
rect 38284 7916 38324 7925
rect 38476 7916 38516 7925
rect 38324 7876 38476 7916
rect 38284 7867 38324 7876
rect 38476 7867 38516 7876
rect 38188 7195 38228 7204
rect 38572 7664 38612 7673
rect 38092 7111 38132 7120
rect 37996 6908 38036 6917
rect 37996 6488 38036 6868
rect 37996 6439 38036 6448
rect 38284 4220 38324 4229
rect 38284 3968 38324 4180
rect 38476 3968 38516 3977
rect 38284 3928 38476 3968
rect 37804 3919 37844 3928
rect 38476 3919 38516 3928
rect 37996 3632 38036 3641
rect 37996 3464 38036 3592
rect 37996 3415 38036 3424
rect 38476 3464 38516 3473
rect 38476 3128 38516 3424
rect 38476 3079 38516 3088
rect 38572 860 38612 7624
rect 38668 7160 38708 7255
rect 38668 7111 38708 7120
rect 38668 6992 38708 7001
rect 38668 6857 38708 6952
rect 38860 6236 38900 7960
rect 39052 7748 39092 7757
rect 39052 7496 39092 7708
rect 39052 7447 39092 7456
rect 38956 7160 38996 7169
rect 38956 6572 38996 7120
rect 38956 6523 38996 6532
rect 39148 7076 39188 7085
rect 38860 6196 38996 6236
rect 38860 6068 38900 6077
rect 38860 5648 38900 6028
rect 38860 5599 38900 5608
rect 38956 4640 38996 6196
rect 39148 5900 39188 7036
rect 39148 5851 39188 5860
rect 38956 4591 38996 4600
rect 38764 4136 38804 4145
rect 38668 3884 38708 3893
rect 38668 3632 38708 3844
rect 38668 3583 38708 3592
rect 38764 2960 38804 4096
rect 38764 2911 38804 2920
rect 39244 2900 39284 9892
rect 40012 9512 40052 9521
rect 39820 8000 39860 8009
rect 39436 7244 39476 7253
rect 39340 7160 39380 7169
rect 39340 7025 39380 7120
rect 39340 3716 39380 3725
rect 39340 3464 39380 3676
rect 39340 3415 39380 3424
rect 39148 2876 39284 2900
rect 39188 2860 39284 2876
rect 39148 2827 39188 2836
rect 39244 2624 39284 2633
rect 39148 2540 39188 2549
rect 38956 2456 38996 2465
rect 39148 2456 39188 2500
rect 38996 2416 39188 2456
rect 38956 2407 38996 2416
rect 39244 2120 39284 2584
rect 39244 2071 39284 2080
rect 38572 811 38612 820
rect 39436 80 39476 7204
rect 39820 4892 39860 7960
rect 39916 7748 39956 7757
rect 39916 7244 39956 7708
rect 39916 7195 39956 7204
rect 39820 4843 39860 4852
rect 40012 4052 40052 9472
rect 40108 8504 40148 8513
rect 40108 8000 40148 8464
rect 40300 8504 40340 8513
rect 40300 8369 40340 8464
rect 40108 7951 40148 7960
rect 40396 8000 40436 8009
rect 40396 7664 40436 7960
rect 40396 7615 40436 7624
rect 40300 6656 40340 6665
rect 40300 6521 40340 6616
rect 40204 6236 40244 6245
rect 40396 6236 40436 6245
rect 40204 5816 40244 6196
rect 40204 5767 40244 5776
rect 40300 6196 40396 6236
rect 40300 4220 40340 6196
rect 40396 6187 40436 6196
rect 40300 4171 40340 4180
rect 40012 4003 40052 4012
rect 40492 4052 40532 9976
rect 41644 9848 41684 9857
rect 40588 9764 40628 9773
rect 40588 7160 40628 9724
rect 40780 9680 40820 9689
rect 40588 7111 40628 7120
rect 40684 9260 40724 9269
rect 40684 8756 40724 9220
rect 40492 4003 40532 4012
rect 40684 3968 40724 8716
rect 40780 4052 40820 9640
rect 41164 9176 41204 9185
rect 41068 8840 41108 8849
rect 40876 7160 40916 7169
rect 40876 6320 40916 7120
rect 40876 6271 40916 6280
rect 41068 4220 41108 8800
rect 41068 4171 41108 4180
rect 40780 4003 40820 4012
rect 40684 3919 40724 3928
rect 40300 3464 40340 3473
rect 40300 2960 40340 3424
rect 40300 2911 40340 2920
rect 40876 3464 40916 3473
rect 40876 104 40916 3424
rect 31084 20 31316 60
rect 32504 0 32584 80
rect 34232 0 34312 80
rect 35960 0 36040 80
rect 37688 0 37768 80
rect 39416 0 39496 80
rect 41164 80 41204 9136
rect 41260 7160 41300 7169
rect 41260 6488 41300 7120
rect 41356 7076 41396 7087
rect 41356 6992 41396 7036
rect 41356 6943 41396 6952
rect 41260 6439 41300 6448
rect 41644 5648 41684 9808
rect 41836 9512 41876 9521
rect 42028 9512 42068 9521
rect 41876 9472 41972 9512
rect 41836 9463 41876 9472
rect 41740 9428 41780 9437
rect 41740 9260 41780 9388
rect 41740 9211 41780 9220
rect 41740 8672 41780 8681
rect 41740 8537 41780 8632
rect 41836 7916 41876 7927
rect 41836 7832 41876 7876
rect 41836 7783 41876 7792
rect 41740 7748 41780 7757
rect 41740 7412 41780 7708
rect 41740 7363 41780 7372
rect 41836 7244 41876 7253
rect 41740 6824 41780 6833
rect 41740 5732 41780 6784
rect 41740 5683 41780 5692
rect 41644 5599 41684 5608
rect 41836 4976 41876 7204
rect 41836 4927 41876 4936
rect 41260 4136 41300 4145
rect 41260 188 41300 4096
rect 41740 3464 41780 3473
rect 41740 1616 41780 3424
rect 41932 3296 41972 9472
rect 42028 6992 42068 9472
rect 42220 9428 42260 9437
rect 42220 8840 42260 9388
rect 42220 8791 42260 8800
rect 42796 8840 42836 8849
rect 42124 8168 42164 8177
rect 42124 8084 42164 8128
rect 42124 8033 42164 8044
rect 42220 7748 42260 7757
rect 42220 7328 42260 7708
rect 42220 7279 42260 7288
rect 42028 6943 42068 6952
rect 42124 4136 42164 4145
rect 42124 4052 42164 4096
rect 42124 4001 42164 4012
rect 41932 3247 41972 3256
rect 42124 3464 42164 3473
rect 41740 1567 41780 1576
rect 42124 608 42164 3424
rect 42508 3464 42548 3473
rect 42508 944 42548 3424
rect 42700 3464 42740 3473
rect 42700 1280 42740 3424
rect 42796 2900 42836 8800
rect 42892 8672 42932 10060
rect 43276 9680 43316 10312
rect 43756 9764 43796 10648
rect 43756 9715 43796 9724
rect 43276 9631 43316 9640
rect 43276 9512 43316 9521
rect 43180 9428 43220 9437
rect 43180 9293 43220 9388
rect 43180 8756 43220 8765
rect 42892 8623 42932 8632
rect 43084 8672 43124 8681
rect 42892 8420 42932 8429
rect 42892 8285 42932 8380
rect 43084 8336 43124 8632
rect 43180 8621 43220 8716
rect 43276 8420 43316 9472
rect 43372 9512 43412 9521
rect 43372 8924 43412 9472
rect 43660 9512 43700 9521
rect 43372 8875 43412 8884
rect 43468 9428 43508 9437
rect 43276 8371 43316 8380
rect 43372 8504 43412 8513
rect 43084 8287 43124 8296
rect 43276 8252 43316 8261
rect 43276 8168 43316 8212
rect 43276 8117 43316 8128
rect 43372 8000 43412 8464
rect 43372 7951 43412 7960
rect 42988 7832 43028 7841
rect 42988 7580 43028 7792
rect 42988 7531 43028 7540
rect 43468 7412 43508 9388
rect 43564 8084 43604 8093
rect 43564 7949 43604 8044
rect 43660 7832 43700 9472
rect 44140 9512 44180 9521
rect 43852 8756 43892 8796
rect 43852 8672 43892 8716
rect 43756 8168 43796 8177
rect 43756 8000 43796 8128
rect 43756 7951 43796 7960
rect 43660 7783 43700 7792
rect 43756 7748 43796 7757
rect 43756 7664 43796 7708
rect 43756 7613 43796 7624
rect 43084 7160 43124 7169
rect 43084 6740 43124 7120
rect 43084 6691 43124 6700
rect 43084 6532 43220 6572
rect 43084 6236 43124 6532
rect 43180 6488 43220 6532
rect 43180 6439 43220 6448
rect 43084 6187 43124 6196
rect 43468 6236 43508 7372
rect 43564 7160 43604 7169
rect 43564 6404 43604 7120
rect 43564 6355 43604 6364
rect 43468 6187 43508 6196
rect 43852 6236 43892 8632
rect 44140 7748 44180 9472
rect 44236 9344 44276 10984
rect 44236 9295 44276 9304
rect 45868 9260 45908 9269
rect 44140 7699 44180 7708
rect 44332 8672 44372 8681
rect 43084 5900 43124 5909
rect 43084 5816 43124 5860
rect 43084 5765 43124 5776
rect 43276 5900 43316 5909
rect 43276 5816 43316 5860
rect 43276 5765 43316 5776
rect 43564 5648 43604 5657
rect 43372 3212 43412 3221
rect 42796 2860 42932 2900
rect 42700 1231 42740 1240
rect 42508 895 42548 904
rect 42124 559 42164 568
rect 41260 139 41300 148
rect 42892 80 42932 2860
rect 43372 1952 43412 3172
rect 43564 3212 43604 5608
rect 43852 5648 43892 6196
rect 43852 5599 43892 5608
rect 44332 4808 44372 8632
rect 45004 8672 45044 8681
rect 44908 8000 44948 8009
rect 44908 7865 44948 7960
rect 44908 7664 44948 7673
rect 44620 7496 44660 7505
rect 44524 7160 44564 7169
rect 44524 6068 44564 7120
rect 44524 6019 44564 6028
rect 44332 4759 44372 4768
rect 44620 4220 44660 7456
rect 44812 6572 44852 6581
rect 44620 4171 44660 4180
rect 44716 5900 44756 5909
rect 44140 3548 44180 3557
rect 43564 3163 43604 3172
rect 43756 3296 43796 3305
rect 43372 1903 43412 1912
rect 43756 1952 43796 3256
rect 43756 1903 43796 1912
rect 44140 1952 44180 3508
rect 44140 1903 44180 1912
rect 44428 3380 44468 3389
rect 44428 1952 44468 3340
rect 44524 3128 44564 3137
rect 44524 2624 44564 3088
rect 44524 2575 44564 2584
rect 44428 1903 44468 1912
rect 44620 1700 44660 1709
rect 44620 608 44660 1660
rect 44620 559 44660 568
rect 44716 440 44756 5860
rect 44812 3464 44852 6532
rect 44908 4976 44948 7624
rect 44908 4927 44948 4936
rect 44812 3415 44852 3424
rect 44908 3968 44948 3977
rect 44908 1952 44948 3928
rect 45004 3800 45044 8632
rect 45772 8588 45812 8597
rect 45676 8504 45716 8513
rect 45676 7664 45716 8464
rect 45772 8000 45812 8548
rect 45868 8336 45908 9220
rect 45868 8287 45908 8296
rect 45772 7951 45812 7960
rect 45676 7615 45716 7624
rect 45868 7748 45908 7757
rect 45868 7328 45908 7708
rect 45868 7279 45908 7288
rect 46252 6824 46292 6833
rect 46252 6656 46292 6784
rect 46252 6607 46292 6616
rect 46252 6152 46292 6161
rect 46252 5984 46292 6112
rect 46252 5935 46292 5944
rect 46252 5480 46292 5489
rect 46252 5312 46292 5440
rect 46252 5263 46292 5272
rect 45004 3751 45044 3760
rect 44908 1903 44948 1912
rect 45580 1784 45620 1793
rect 45580 944 45620 1744
rect 46252 1448 46292 1457
rect 46252 1280 46292 1408
rect 46252 1231 46292 1240
rect 45580 895 45620 904
rect 44620 400 44756 440
rect 44620 80 44660 400
rect 40876 55 40916 64
rect 41144 0 41224 80
rect 42872 0 42952 80
rect 44600 0 44680 80
<< via3 >>
rect 748 4096 788 4136
rect 1420 4264 1460 4304
rect 1420 3928 1460 3968
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 10156 9892 10196 9932
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 10828 9472 10868 9512
rect 10540 8380 10580 8420
rect 10252 6196 10292 6236
rect 11308 9724 11348 9764
rect 11308 9388 11348 9428
rect 11020 8296 11060 8336
rect 11500 9220 11540 9260
rect 11884 9724 11924 9764
rect 11020 3340 11060 3380
rect 10060 3172 10100 3212
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 11980 8716 12020 8756
rect 12172 9472 12212 9512
rect 11884 7708 11924 7748
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 12268 9136 12308 9176
rect 12652 9556 12692 9596
rect 12556 9388 12596 9428
rect 12940 9640 12980 9680
rect 12844 9052 12884 9092
rect 13324 9640 13364 9680
rect 13420 9724 13460 9764
rect 13132 8884 13172 8924
rect 12748 8800 12788 8840
rect 12844 8212 12884 8252
rect 12556 3256 12596 3296
rect 12940 7792 12980 7832
rect 12940 3340 12980 3380
rect 13132 8464 13172 8504
rect 13516 8632 13556 8672
rect 13612 8548 13652 8588
rect 14092 8716 14132 8756
rect 14284 8548 14324 8588
rect 13900 7876 13940 7916
rect 14668 9724 14708 9764
rect 14188 3760 14228 3800
rect 14092 3088 14132 3128
rect 13804 2920 13844 2960
rect 15148 9556 15188 9596
rect 14860 8716 14900 8756
rect 14764 8548 14804 8588
rect 14764 8296 14804 8336
rect 14956 7540 14996 7580
rect 15148 7204 15188 7244
rect 15628 8716 15668 8756
rect 14572 3004 14612 3044
rect 15628 3256 15668 3296
rect 15628 3004 15668 3044
rect 15820 8548 15860 8588
rect 16300 9808 16340 9848
rect 16492 9136 16532 9176
rect 15820 7624 15860 7664
rect 15820 6868 15860 6908
rect 16588 8800 16628 8840
rect 16492 8212 16532 8252
rect 16492 7456 16532 7496
rect 16300 6868 16340 6908
rect 16972 8548 17012 8588
rect 16684 8044 16724 8084
rect 17548 9808 17588 9848
rect 17452 9724 17492 9764
rect 17452 9388 17492 9428
rect 18124 9724 18164 9764
rect 18412 9976 18452 10016
rect 17836 9472 17876 9512
rect 17356 8464 17396 8504
rect 16396 3340 16436 3380
rect 16300 3256 16340 3296
rect 17644 7960 17684 8000
rect 17740 3760 17780 3800
rect 17932 3088 17972 3128
rect 17836 2920 17876 2960
rect 19084 9976 19124 10016
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 18412 8212 18452 8252
rect 19372 8884 19412 8924
rect 19564 9220 19604 9260
rect 18796 8464 18836 8504
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 19276 8128 19316 8168
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 19852 9304 19892 9344
rect 19852 9136 19892 9176
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 20044 8884 20084 8924
rect 19756 8800 19796 8840
rect 19564 8296 19604 8336
rect 20140 8464 20180 8504
rect 20044 8380 20084 8420
rect 19948 8296 19988 8336
rect 19948 7540 19988 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 20524 7456 20564 7496
rect 19948 7372 19988 7412
rect 19756 7288 19796 7328
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 20524 5944 20564 5984
rect 18700 5860 18740 5900
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 19276 4180 19316 4220
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 18700 2920 18740 2960
rect 20716 4180 20756 4220
rect 20908 8548 20948 8588
rect 21868 9136 21908 9176
rect 21676 7204 21716 7244
rect 22732 9640 22772 9680
rect 22348 9304 22388 9344
rect 22060 4348 22100 4388
rect 22540 4432 22580 4472
rect 21964 3424 22004 3464
rect 22924 9976 22964 10016
rect 23020 9892 23060 9932
rect 22732 3424 22772 3464
rect 22828 4432 22868 4472
rect 22732 3088 22772 3128
rect 23116 9640 23156 9680
rect 23596 9892 23636 9932
rect 25132 9724 25172 9764
rect 23788 9220 23828 9260
rect 24172 8800 24212 8840
rect 23692 6952 23732 6992
rect 24364 8716 24404 8756
rect 23788 6364 23828 6404
rect 23692 6028 23732 6068
rect 22924 4180 22964 4220
rect 23020 3592 23060 3632
rect 23116 3508 23156 3548
rect 23692 4180 23732 4220
rect 23884 4180 23924 4220
rect 23884 3844 23924 3884
rect 23788 3340 23828 3380
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 20428 820 20468 860
rect 24364 4348 24404 4388
rect 24172 4180 24212 4220
rect 24556 4012 24596 4052
rect 24844 8800 24884 8840
rect 25804 9220 25844 9260
rect 25900 9136 25940 9176
rect 25036 3844 25076 3884
rect 25036 3508 25076 3548
rect 24748 3340 24788 3380
rect 25804 6028 25844 6068
rect 26572 9220 26612 9260
rect 26956 9556 26996 9596
rect 26860 9136 26900 9176
rect 26572 8716 26612 8756
rect 26476 7372 26516 7412
rect 27052 6616 27092 6656
rect 26092 3592 26132 3632
rect 27820 9724 27860 9764
rect 27628 7120 27668 7160
rect 27532 6364 27572 6404
rect 27820 5860 27860 5900
rect 28780 8800 28820 8840
rect 28684 8464 28724 8504
rect 28492 8380 28532 8420
rect 28588 8128 28628 8168
rect 28876 8128 28916 8168
rect 28492 7540 28532 7580
rect 28780 7456 28820 7496
rect 29356 8716 29396 8756
rect 28684 7288 28724 7328
rect 28876 7372 28916 7412
rect 28780 7120 28820 7160
rect 29068 6952 29108 6992
rect 28876 6196 28916 6236
rect 28780 6028 28820 6068
rect 28012 5944 28052 5984
rect 27916 4432 27956 4472
rect 27724 4180 27764 4220
rect 25900 3004 25940 3044
rect 24748 820 24788 860
rect 29644 8800 29684 8840
rect 30220 11404 30260 11444
rect 30604 11152 30644 11192
rect 29740 7456 29780 7496
rect 29932 6952 29972 6992
rect 30316 9640 30356 9680
rect 30220 8380 30260 8420
rect 30316 7456 30356 7496
rect 30124 7288 30164 7328
rect 30604 7288 30644 7328
rect 29740 6112 29780 6152
rect 30220 5944 30260 5984
rect 30988 9136 31028 9176
rect 30796 7372 30836 7412
rect 31660 8716 31700 8756
rect 30988 6532 31028 6572
rect 31468 6028 31508 6068
rect 32716 8968 32756 9008
rect 33004 9892 33044 9932
rect 32908 5860 32948 5900
rect 33484 9640 33524 9680
rect 34252 10312 34292 10352
rect 33868 9976 33908 10016
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 34252 9640 34292 9680
rect 34060 9556 34100 9596
rect 34540 10312 34580 10352
rect 34636 9724 34676 9764
rect 34732 9976 34772 10016
rect 38860 11404 38900 11444
rect 37420 9892 37460 9932
rect 35020 9640 35060 9680
rect 35404 9724 35444 9764
rect 36172 9640 36212 9680
rect 33772 8548 33812 8588
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 33292 4096 33332 4136
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 35404 9388 35444 9428
rect 35500 9220 35540 9260
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 35404 8884 35444 8924
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 36076 9388 36116 9428
rect 35884 9136 35924 9176
rect 35692 8464 35732 8504
rect 35788 8128 35828 8168
rect 35980 8884 36020 8924
rect 35020 6700 35060 6740
rect 35788 6700 35828 6740
rect 34924 6448 34964 6488
rect 35020 6364 35060 6404
rect 34924 6280 34964 6320
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 35884 6364 35924 6404
rect 35692 5860 35732 5900
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
rect 32524 820 32564 860
rect 36172 9220 36212 9260
rect 36172 8968 36212 9008
rect 36460 9556 36500 9596
rect 37324 9304 37364 9344
rect 36268 6448 36308 6488
rect 36364 8548 36404 8588
rect 36748 7456 36788 7496
rect 36460 5944 36500 5984
rect 37132 6280 37172 6320
rect 37036 4264 37076 4304
rect 38956 11152 38996 11192
rect 38380 8464 38420 8504
rect 37804 3928 37844 3968
rect 38668 7120 38708 7160
rect 38668 6952 38708 6992
rect 38956 6532 38996 6572
rect 38764 2920 38804 2960
rect 39340 7120 39380 7160
rect 38572 820 38612 860
rect 40300 8464 40340 8504
rect 40300 6616 40340 6656
rect 41356 7036 41396 7076
rect 41740 9388 41780 9428
rect 41740 8632 41780 8672
rect 41836 7876 41876 7916
rect 42124 8128 42164 8168
rect 42028 6952 42068 6992
rect 42124 4012 42164 4052
rect 41932 3256 41972 3296
rect 43180 9388 43220 9428
rect 43180 8716 43220 8756
rect 42892 8380 42932 8420
rect 43372 9472 43412 9512
rect 43276 8380 43316 8420
rect 43276 8212 43316 8252
rect 43564 8044 43604 8084
rect 43852 8716 43892 8756
rect 43756 8128 43796 8168
rect 43660 7792 43700 7832
rect 43756 7624 43796 7664
rect 44140 7708 44180 7748
rect 43084 5776 43124 5816
rect 43276 5776 43316 5816
rect 44908 7960 44948 8000
rect 43564 3172 43604 3212
<< metal4 >>
rect 30211 11404 30220 11444
rect 30260 11404 38860 11444
rect 38900 11404 38909 11444
rect 30595 11152 30604 11192
rect 30644 11152 38956 11192
rect 38996 11152 39005 11192
rect 34243 10312 34252 10352
rect 34292 10312 34540 10352
rect 34580 10312 34589 10352
rect 18403 9976 18412 10016
rect 18452 9976 19084 10016
rect 19124 9976 19133 10016
rect 20140 9976 22924 10016
rect 22964 9976 22973 10016
rect 33859 9976 33868 10016
rect 33908 9976 34732 10016
rect 34772 9976 34781 10016
rect 10147 9892 10156 9932
rect 10196 9892 18260 9932
rect 3679 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4065 9848
rect 16291 9808 16300 9848
rect 16340 9808 17548 9848
rect 17588 9808 17597 9848
rect 18220 9764 18260 9892
rect 18799 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19185 9848
rect 20140 9764 20180 9976
rect 23011 9892 23020 9932
rect 23060 9892 23596 9932
rect 23636 9892 23645 9932
rect 32995 9892 33004 9932
rect 33044 9892 37420 9932
rect 37460 9892 37469 9932
rect 33919 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34305 9848
rect 11299 9724 11308 9764
rect 11348 9724 11884 9764
rect 11924 9724 11933 9764
rect 13411 9724 13420 9764
rect 13460 9724 14668 9764
rect 14708 9724 14717 9764
rect 17443 9724 17452 9764
rect 17492 9724 18124 9764
rect 18164 9724 18173 9764
rect 18220 9724 20180 9764
rect 25123 9724 25132 9764
rect 25172 9724 27820 9764
rect 27860 9724 27869 9764
rect 34627 9724 34636 9764
rect 34676 9724 35404 9764
rect 35444 9724 35453 9764
rect 12931 9640 12940 9680
rect 12980 9640 13324 9680
rect 13364 9640 13373 9680
rect 15052 9640 22732 9680
rect 22772 9640 22781 9680
rect 23107 9640 23116 9680
rect 23156 9640 30316 9680
rect 30356 9640 30365 9680
rect 33475 9640 33484 9680
rect 33524 9640 34252 9680
rect 34292 9640 34301 9680
rect 35011 9640 35020 9680
rect 35060 9640 36172 9680
rect 36212 9640 36221 9680
rect 15052 9596 15092 9640
rect 12643 9556 12652 9596
rect 12692 9556 15092 9596
rect 15139 9556 15148 9596
rect 15188 9556 26956 9596
rect 26996 9556 27005 9596
rect 34051 9556 34060 9596
rect 34100 9556 36460 9596
rect 36500 9556 36509 9596
rect 10819 9472 10828 9512
rect 10868 9472 12172 9512
rect 12212 9472 12221 9512
rect 17827 9472 17836 9512
rect 17876 9472 43372 9512
rect 43412 9472 43421 9512
rect 11299 9388 11308 9428
rect 11348 9388 12556 9428
rect 12596 9388 12605 9428
rect 17443 9388 17452 9428
rect 17492 9388 23060 9428
rect 35395 9388 35404 9428
rect 35444 9388 36076 9428
rect 36116 9388 36125 9428
rect 41731 9388 41740 9428
rect 41780 9388 43180 9428
rect 43220 9388 43229 9428
rect 23020 9344 23060 9388
rect 19843 9304 19852 9344
rect 19892 9304 22348 9344
rect 22388 9304 22397 9344
rect 23020 9304 37324 9344
rect 37364 9304 37373 9344
rect 11491 9220 11500 9260
rect 11540 9220 19564 9260
rect 19604 9220 19613 9260
rect 19756 9220 23788 9260
rect 23828 9220 23837 9260
rect 25795 9220 25804 9260
rect 25844 9220 26572 9260
rect 26612 9220 26621 9260
rect 35491 9220 35500 9260
rect 35540 9220 36172 9260
rect 36212 9220 36221 9260
rect 19756 9176 19796 9220
rect 12259 9136 12268 9176
rect 12308 9136 12980 9176
rect 16483 9136 16492 9176
rect 16532 9136 19796 9176
rect 19843 9136 19852 9176
rect 19892 9136 21868 9176
rect 21908 9136 21917 9176
rect 25891 9136 25900 9176
rect 25940 9136 26860 9176
rect 26900 9136 26909 9176
rect 30979 9136 30988 9176
rect 31028 9136 35884 9176
rect 35924 9136 35933 9176
rect 12940 9092 12980 9136
rect 4919 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5305 9092
rect 12748 9052 12844 9092
rect 12884 9052 12893 9092
rect 12940 9052 18740 9092
rect 20039 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20425 9092
rect 35159 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35545 9092
rect 12748 8840 12788 9052
rect 18700 9008 18740 9052
rect 18700 8968 20084 9008
rect 32707 8968 32716 9008
rect 32756 8968 36172 9008
rect 36212 8968 36221 9008
rect 20044 8924 20084 8968
rect 12940 8884 13132 8924
rect 13172 8884 13181 8924
rect 19363 8884 19372 8924
rect 19412 8884 19892 8924
rect 20035 8884 20044 8924
rect 20084 8884 20093 8924
rect 35395 8884 35404 8924
rect 35444 8884 35980 8924
rect 36020 8884 36029 8924
rect 12739 8800 12748 8840
rect 12788 8800 12797 8840
rect 12940 8756 12980 8884
rect 19852 8840 19892 8884
rect 16579 8800 16588 8840
rect 16628 8800 19756 8840
rect 19796 8800 19805 8840
rect 19852 8800 24172 8840
rect 24212 8800 24221 8840
rect 24268 8800 24844 8840
rect 24884 8800 24893 8840
rect 28771 8800 28780 8840
rect 28820 8800 29644 8840
rect 29684 8800 29693 8840
rect 24268 8756 24308 8800
rect 11971 8716 11980 8756
rect 12020 8716 12980 8756
rect 14083 8716 14092 8756
rect 14132 8716 14860 8756
rect 14900 8716 14909 8756
rect 15619 8716 15628 8756
rect 15668 8716 24308 8756
rect 24355 8716 24364 8756
rect 24404 8716 26572 8756
rect 26612 8716 26621 8756
rect 29347 8716 29356 8756
rect 29396 8716 31660 8756
rect 31700 8716 31709 8756
rect 43171 8716 43180 8756
rect 43220 8716 43852 8756
rect 43892 8716 43901 8756
rect 13507 8632 13516 8672
rect 13556 8632 41740 8672
rect 41780 8632 41789 8672
rect 13603 8548 13612 8588
rect 13652 8548 14284 8588
rect 14324 8548 14333 8588
rect 14755 8548 14764 8588
rect 14804 8548 15820 8588
rect 15860 8548 15869 8588
rect 16963 8548 16972 8588
rect 17012 8548 20908 8588
rect 20948 8548 20957 8588
rect 33763 8548 33772 8588
rect 33812 8548 36364 8588
rect 36404 8548 36413 8588
rect 13123 8464 13132 8504
rect 13172 8464 17356 8504
rect 17396 8464 17405 8504
rect 18787 8464 18796 8504
rect 18836 8464 20140 8504
rect 20180 8464 20189 8504
rect 28675 8464 28684 8504
rect 28724 8464 35692 8504
rect 35732 8464 35741 8504
rect 38371 8464 38380 8504
rect 38420 8464 40300 8504
rect 40340 8464 40349 8504
rect 10531 8380 10540 8420
rect 10580 8380 20044 8420
rect 20084 8380 20093 8420
rect 28483 8380 28492 8420
rect 28532 8380 30220 8420
rect 30260 8380 30269 8420
rect 42883 8380 42892 8420
rect 42932 8380 43276 8420
rect 43316 8380 43325 8420
rect 3679 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4065 8336
rect 11011 8296 11020 8336
rect 11060 8296 14764 8336
rect 14804 8296 14813 8336
rect 18799 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19185 8336
rect 19555 8296 19564 8336
rect 19604 8296 19948 8336
rect 19988 8296 19997 8336
rect 33919 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34305 8336
rect 12835 8212 12844 8252
rect 12884 8212 16492 8252
rect 16532 8212 16541 8252
rect 18403 8212 18412 8252
rect 18452 8212 43276 8252
rect 43316 8212 43325 8252
rect 19267 8128 19276 8168
rect 19316 8128 28588 8168
rect 28628 8128 28637 8168
rect 28867 8128 28876 8168
rect 28916 8128 35788 8168
rect 35828 8128 35837 8168
rect 42115 8128 42124 8168
rect 42164 8128 43756 8168
rect 43796 8128 43805 8168
rect 16675 8044 16684 8084
rect 16724 8044 43564 8084
rect 43604 8044 43613 8084
rect 17635 7960 17644 8000
rect 17684 7960 44908 8000
rect 44948 7960 44957 8000
rect 13891 7876 13900 7916
rect 13940 7876 41836 7916
rect 41876 7876 41885 7916
rect 12931 7792 12940 7832
rect 12980 7792 43660 7832
rect 43700 7792 43709 7832
rect 11875 7708 11884 7748
rect 11924 7708 44140 7748
rect 44180 7708 44189 7748
rect 15811 7624 15820 7664
rect 15860 7624 43756 7664
rect 43796 7624 43805 7664
rect 4919 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5305 7580
rect 14947 7540 14956 7580
rect 14996 7540 19948 7580
rect 19988 7540 19997 7580
rect 20039 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20425 7580
rect 28483 7540 28492 7580
rect 28532 7540 33812 7580
rect 35159 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35545 7580
rect 33772 7496 33812 7540
rect 16483 7456 16492 7496
rect 16532 7456 20524 7496
rect 20564 7456 20573 7496
rect 28771 7456 28780 7496
rect 28820 7456 29740 7496
rect 29780 7456 29789 7496
rect 30221 7456 30316 7496
rect 30356 7456 30365 7496
rect 33772 7456 36748 7496
rect 36788 7456 36797 7496
rect 19939 7372 19948 7412
rect 19988 7372 26476 7412
rect 26516 7372 26525 7412
rect 28867 7372 28876 7412
rect 28916 7372 30796 7412
rect 30836 7372 30845 7412
rect 19747 7288 19756 7328
rect 19796 7288 28684 7328
rect 28724 7288 28733 7328
rect 30115 7288 30124 7328
rect 30164 7288 30604 7328
rect 30644 7288 30653 7328
rect 15139 7204 15148 7244
rect 15188 7204 21676 7244
rect 21716 7204 21725 7244
rect 27619 7120 27628 7160
rect 27668 7120 28780 7160
rect 28820 7120 28829 7160
rect 38659 7120 38668 7160
rect 38708 7120 39340 7160
rect 39380 7120 39389 7160
rect 28780 7036 41356 7076
rect 41396 7036 41405 7076
rect 28780 6992 28820 7036
rect 23683 6952 23692 6992
rect 23732 6952 28820 6992
rect 29059 6952 29068 6992
rect 29108 6952 29932 6992
rect 29972 6952 29981 6992
rect 38659 6952 38668 6992
rect 38708 6952 42028 6992
rect 42068 6952 42077 6992
rect 15811 6868 15820 6908
rect 15860 6868 16300 6908
rect 16340 6868 16349 6908
rect 3679 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4065 6824
rect 18799 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19185 6824
rect 33919 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34305 6824
rect 35011 6700 35020 6740
rect 35060 6700 35788 6740
rect 35828 6700 35837 6740
rect 27043 6616 27052 6656
rect 27092 6616 40300 6656
rect 40340 6616 40349 6656
rect 30979 6532 30988 6572
rect 31028 6532 38956 6572
rect 38996 6532 39005 6572
rect 34915 6448 34924 6488
rect 34964 6448 36268 6488
rect 36308 6448 36317 6488
rect 23779 6364 23788 6404
rect 23828 6364 27532 6404
rect 27572 6364 27581 6404
rect 35011 6364 35020 6404
rect 35060 6364 35884 6404
rect 35924 6364 35933 6404
rect 34915 6280 34924 6320
rect 34964 6280 37132 6320
rect 37172 6280 37181 6320
rect 10243 6196 10252 6236
rect 10292 6196 18740 6236
rect 28867 6196 28876 6236
rect 28916 6196 30316 6236
rect 30356 6196 30365 6236
rect 18700 6152 18740 6196
rect 18700 6112 29740 6152
rect 29780 6112 29789 6152
rect 4919 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5305 6068
rect 20039 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20425 6068
rect 23683 6028 23692 6068
rect 23732 6028 25804 6068
rect 25844 6028 25853 6068
rect 28771 6028 28780 6068
rect 28820 6028 31468 6068
rect 31508 6028 31517 6068
rect 35159 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35545 6068
rect 20515 5944 20524 5984
rect 20564 5944 28012 5984
rect 28052 5944 28061 5984
rect 30211 5944 30220 5984
rect 30260 5944 36460 5984
rect 36500 5944 36509 5984
rect 18691 5860 18700 5900
rect 18740 5860 27820 5900
rect 27860 5860 27869 5900
rect 32899 5860 32908 5900
rect 32948 5860 35692 5900
rect 35732 5860 35741 5900
rect 43075 5776 43084 5816
rect 43124 5776 43276 5816
rect 43316 5776 43325 5816
rect 3679 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4065 5312
rect 18799 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19185 5312
rect 33919 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34305 5312
rect 4919 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5305 4556
rect 20039 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20425 4556
rect 35159 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35545 4556
rect 22531 4432 22540 4472
rect 22580 4432 22828 4472
rect 22868 4432 27916 4472
rect 27956 4432 27965 4472
rect 22051 4348 22060 4388
rect 22100 4348 24364 4388
rect 24404 4348 24413 4388
rect 1411 4264 1420 4304
rect 1460 4264 37036 4304
rect 37076 4264 37085 4304
rect 19267 4180 19276 4220
rect 19316 4180 20716 4220
rect 20756 4180 20765 4220
rect 22915 4180 22924 4220
rect 22964 4180 23692 4220
rect 23732 4180 23741 4220
rect 23875 4180 23884 4220
rect 23924 4180 24172 4220
rect 24212 4180 27724 4220
rect 27764 4180 27773 4220
rect 739 4096 748 4136
rect 788 4096 33292 4136
rect 33332 4096 33341 4136
rect 24547 4012 24556 4052
rect 24596 4012 42124 4052
rect 42164 4012 42173 4052
rect 1411 3928 1420 3968
rect 1460 3928 37804 3968
rect 37844 3928 37853 3968
rect 23875 3844 23884 3884
rect 23924 3844 25036 3884
rect 25076 3844 25085 3884
rect 3679 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4065 3800
rect 14179 3760 14188 3800
rect 14228 3760 17740 3800
rect 17780 3760 17789 3800
rect 18799 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19185 3800
rect 33919 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34305 3800
rect 23011 3592 23020 3632
rect 23060 3592 26092 3632
rect 26132 3592 26141 3632
rect 23107 3508 23116 3548
rect 23156 3508 25036 3548
rect 25076 3508 25085 3548
rect 21955 3424 21964 3464
rect 22004 3424 22732 3464
rect 22772 3424 22781 3464
rect 11011 3340 11020 3380
rect 11060 3340 12940 3380
rect 12980 3340 16396 3380
rect 16436 3340 16445 3380
rect 23779 3340 23788 3380
rect 23828 3340 24748 3380
rect 24788 3340 24797 3380
rect 12547 3256 12556 3296
rect 12596 3256 15628 3296
rect 15668 3256 15677 3296
rect 16291 3256 16300 3296
rect 16340 3256 41932 3296
rect 41972 3256 41981 3296
rect 10051 3172 10060 3212
rect 10100 3172 43564 3212
rect 43604 3172 43613 3212
rect 14083 3088 14092 3128
rect 14132 3088 17932 3128
rect 17972 3088 17981 3128
rect 22723 3088 22732 3128
rect 22772 3088 23060 3128
rect 23020 3044 23060 3088
rect 4919 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5305 3044
rect 14563 3004 14572 3044
rect 14612 3004 15628 3044
rect 15668 3004 15677 3044
rect 20039 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20425 3044
rect 23020 3004 25900 3044
rect 25940 3004 25949 3044
rect 35159 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35545 3044
rect 13795 2920 13804 2960
rect 13844 2920 17836 2960
rect 17876 2920 17885 2960
rect 18691 2920 18700 2960
rect 18740 2920 38764 2960
rect 38804 2920 38813 2960
rect 3679 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4065 2288
rect 18799 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19185 2288
rect 33919 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34305 2288
rect 4919 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5305 1532
rect 20039 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20425 1532
rect 35159 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35545 1532
rect 20419 820 20428 860
rect 20468 820 24748 860
rect 24788 820 24797 860
rect 32515 820 32524 860
rect 32564 820 38572 860
rect 38612 820 38621 860
<< via4 >>
rect 3688 9808 3728 9848
rect 3770 9808 3810 9848
rect 3852 9808 3892 9848
rect 3934 9808 3974 9848
rect 4016 9808 4056 9848
rect 18808 9808 18848 9848
rect 18890 9808 18930 9848
rect 18972 9808 19012 9848
rect 19054 9808 19094 9848
rect 19136 9808 19176 9848
rect 33928 9808 33968 9848
rect 34010 9808 34050 9848
rect 34092 9808 34132 9848
rect 34174 9808 34214 9848
rect 34256 9808 34296 9848
rect 4928 9052 4968 9092
rect 5010 9052 5050 9092
rect 5092 9052 5132 9092
rect 5174 9052 5214 9092
rect 5256 9052 5296 9092
rect 20048 9052 20088 9092
rect 20130 9052 20170 9092
rect 20212 9052 20252 9092
rect 20294 9052 20334 9092
rect 20376 9052 20416 9092
rect 35168 9052 35208 9092
rect 35250 9052 35290 9092
rect 35332 9052 35372 9092
rect 35414 9052 35454 9092
rect 35496 9052 35536 9092
rect 3688 8296 3728 8336
rect 3770 8296 3810 8336
rect 3852 8296 3892 8336
rect 3934 8296 3974 8336
rect 4016 8296 4056 8336
rect 18808 8296 18848 8336
rect 18890 8296 18930 8336
rect 18972 8296 19012 8336
rect 19054 8296 19094 8336
rect 19136 8296 19176 8336
rect 33928 8296 33968 8336
rect 34010 8296 34050 8336
rect 34092 8296 34132 8336
rect 34174 8296 34214 8336
rect 34256 8296 34296 8336
rect 4928 7540 4968 7580
rect 5010 7540 5050 7580
rect 5092 7540 5132 7580
rect 5174 7540 5214 7580
rect 5256 7540 5296 7580
rect 20048 7540 20088 7580
rect 20130 7540 20170 7580
rect 20212 7540 20252 7580
rect 20294 7540 20334 7580
rect 20376 7540 20416 7580
rect 35168 7540 35208 7580
rect 35250 7540 35290 7580
rect 35332 7540 35372 7580
rect 35414 7540 35454 7580
rect 35496 7540 35536 7580
rect 30316 7456 30356 7496
rect 3688 6784 3728 6824
rect 3770 6784 3810 6824
rect 3852 6784 3892 6824
rect 3934 6784 3974 6824
rect 4016 6784 4056 6824
rect 18808 6784 18848 6824
rect 18890 6784 18930 6824
rect 18972 6784 19012 6824
rect 19054 6784 19094 6824
rect 19136 6784 19176 6824
rect 33928 6784 33968 6824
rect 34010 6784 34050 6824
rect 34092 6784 34132 6824
rect 34174 6784 34214 6824
rect 34256 6784 34296 6824
rect 30316 6196 30356 6236
rect 4928 6028 4968 6068
rect 5010 6028 5050 6068
rect 5092 6028 5132 6068
rect 5174 6028 5214 6068
rect 5256 6028 5296 6068
rect 20048 6028 20088 6068
rect 20130 6028 20170 6068
rect 20212 6028 20252 6068
rect 20294 6028 20334 6068
rect 20376 6028 20416 6068
rect 35168 6028 35208 6068
rect 35250 6028 35290 6068
rect 35332 6028 35372 6068
rect 35414 6028 35454 6068
rect 35496 6028 35536 6068
rect 3688 5272 3728 5312
rect 3770 5272 3810 5312
rect 3852 5272 3892 5312
rect 3934 5272 3974 5312
rect 4016 5272 4056 5312
rect 18808 5272 18848 5312
rect 18890 5272 18930 5312
rect 18972 5272 19012 5312
rect 19054 5272 19094 5312
rect 19136 5272 19176 5312
rect 33928 5272 33968 5312
rect 34010 5272 34050 5312
rect 34092 5272 34132 5312
rect 34174 5272 34214 5312
rect 34256 5272 34296 5312
rect 4928 4516 4968 4556
rect 5010 4516 5050 4556
rect 5092 4516 5132 4556
rect 5174 4516 5214 4556
rect 5256 4516 5296 4556
rect 20048 4516 20088 4556
rect 20130 4516 20170 4556
rect 20212 4516 20252 4556
rect 20294 4516 20334 4556
rect 20376 4516 20416 4556
rect 35168 4516 35208 4556
rect 35250 4516 35290 4556
rect 35332 4516 35372 4556
rect 35414 4516 35454 4556
rect 35496 4516 35536 4556
rect 3688 3760 3728 3800
rect 3770 3760 3810 3800
rect 3852 3760 3892 3800
rect 3934 3760 3974 3800
rect 4016 3760 4056 3800
rect 18808 3760 18848 3800
rect 18890 3760 18930 3800
rect 18972 3760 19012 3800
rect 19054 3760 19094 3800
rect 19136 3760 19176 3800
rect 33928 3760 33968 3800
rect 34010 3760 34050 3800
rect 34092 3760 34132 3800
rect 34174 3760 34214 3800
rect 34256 3760 34296 3800
rect 4928 3004 4968 3044
rect 5010 3004 5050 3044
rect 5092 3004 5132 3044
rect 5174 3004 5214 3044
rect 5256 3004 5296 3044
rect 20048 3004 20088 3044
rect 20130 3004 20170 3044
rect 20212 3004 20252 3044
rect 20294 3004 20334 3044
rect 20376 3004 20416 3044
rect 35168 3004 35208 3044
rect 35250 3004 35290 3044
rect 35332 3004 35372 3044
rect 35414 3004 35454 3044
rect 35496 3004 35536 3044
rect 3688 2248 3728 2288
rect 3770 2248 3810 2288
rect 3852 2248 3892 2288
rect 3934 2248 3974 2288
rect 4016 2248 4056 2288
rect 18808 2248 18848 2288
rect 18890 2248 18930 2288
rect 18972 2248 19012 2288
rect 19054 2248 19094 2288
rect 19136 2248 19176 2288
rect 33928 2248 33968 2288
rect 34010 2248 34050 2288
rect 34092 2248 34132 2288
rect 34174 2248 34214 2288
rect 34256 2248 34296 2288
rect 4928 1492 4968 1532
rect 5010 1492 5050 1532
rect 5092 1492 5132 1532
rect 5174 1492 5214 1532
rect 5256 1492 5296 1532
rect 20048 1492 20088 1532
rect 20130 1492 20170 1532
rect 20212 1492 20252 1532
rect 20294 1492 20334 1532
rect 20376 1492 20416 1532
rect 35168 1492 35208 1532
rect 35250 1492 35290 1532
rect 35332 1492 35372 1532
rect 35414 1492 35454 1532
rect 35496 1492 35536 1532
<< metal5 >>
rect 3652 9848 4092 11844
rect 3652 9808 3688 9848
rect 3728 9808 3770 9848
rect 3810 9808 3852 9848
rect 3892 9808 3934 9848
rect 3974 9808 4016 9848
rect 4056 9808 4092 9848
rect 3652 8336 4092 9808
rect 3652 8296 3688 8336
rect 3728 8296 3770 8336
rect 3810 8296 3852 8336
rect 3892 8296 3934 8336
rect 3974 8296 4016 8336
rect 4056 8296 4092 8336
rect 3652 6824 4092 8296
rect 3652 6784 3688 6824
rect 3728 6784 3770 6824
rect 3810 6784 3852 6824
rect 3892 6784 3934 6824
rect 3974 6784 4016 6824
rect 4056 6784 4092 6824
rect 3652 5312 4092 6784
rect 3652 5272 3688 5312
rect 3728 5272 3770 5312
rect 3810 5272 3852 5312
rect 3892 5272 3934 5312
rect 3974 5272 4016 5312
rect 4056 5272 4092 5312
rect 3652 3800 4092 5272
rect 3652 3760 3688 3800
rect 3728 3760 3770 3800
rect 3810 3760 3852 3800
rect 3892 3760 3934 3800
rect 3974 3760 4016 3800
rect 4056 3760 4092 3800
rect 3652 2288 4092 3760
rect 3652 2248 3688 2288
rect 3728 2248 3770 2288
rect 3810 2248 3852 2288
rect 3892 2248 3934 2288
rect 3974 2248 4016 2288
rect 4056 2248 4092 2288
rect 3652 0 4092 2248
rect 4892 9092 5332 11844
rect 4892 9052 4928 9092
rect 4968 9052 5010 9092
rect 5050 9052 5092 9092
rect 5132 9052 5174 9092
rect 5214 9052 5256 9092
rect 5296 9052 5332 9092
rect 4892 7580 5332 9052
rect 4892 7540 4928 7580
rect 4968 7540 5010 7580
rect 5050 7540 5092 7580
rect 5132 7540 5174 7580
rect 5214 7540 5256 7580
rect 5296 7540 5332 7580
rect 4892 6068 5332 7540
rect 4892 6028 4928 6068
rect 4968 6028 5010 6068
rect 5050 6028 5092 6068
rect 5132 6028 5174 6068
rect 5214 6028 5256 6068
rect 5296 6028 5332 6068
rect 4892 4556 5332 6028
rect 4892 4516 4928 4556
rect 4968 4516 5010 4556
rect 5050 4516 5092 4556
rect 5132 4516 5174 4556
rect 5214 4516 5256 4556
rect 5296 4516 5332 4556
rect 4892 3044 5332 4516
rect 4892 3004 4928 3044
rect 4968 3004 5010 3044
rect 5050 3004 5092 3044
rect 5132 3004 5174 3044
rect 5214 3004 5256 3044
rect 5296 3004 5332 3044
rect 4892 1532 5332 3004
rect 4892 1492 4928 1532
rect 4968 1492 5010 1532
rect 5050 1492 5092 1532
rect 5132 1492 5174 1532
rect 5214 1492 5256 1532
rect 5296 1492 5332 1532
rect 4892 0 5332 1492
rect 18772 9848 19212 11844
rect 18772 9808 18808 9848
rect 18848 9808 18890 9848
rect 18930 9808 18972 9848
rect 19012 9808 19054 9848
rect 19094 9808 19136 9848
rect 19176 9808 19212 9848
rect 18772 8336 19212 9808
rect 18772 8296 18808 8336
rect 18848 8296 18890 8336
rect 18930 8296 18972 8336
rect 19012 8296 19054 8336
rect 19094 8296 19136 8336
rect 19176 8296 19212 8336
rect 18772 6824 19212 8296
rect 18772 6784 18808 6824
rect 18848 6784 18890 6824
rect 18930 6784 18972 6824
rect 19012 6784 19054 6824
rect 19094 6784 19136 6824
rect 19176 6784 19212 6824
rect 18772 5312 19212 6784
rect 18772 5272 18808 5312
rect 18848 5272 18890 5312
rect 18930 5272 18972 5312
rect 19012 5272 19054 5312
rect 19094 5272 19136 5312
rect 19176 5272 19212 5312
rect 18772 3800 19212 5272
rect 18772 3760 18808 3800
rect 18848 3760 18890 3800
rect 18930 3760 18972 3800
rect 19012 3760 19054 3800
rect 19094 3760 19136 3800
rect 19176 3760 19212 3800
rect 18772 2288 19212 3760
rect 18772 2248 18808 2288
rect 18848 2248 18890 2288
rect 18930 2248 18972 2288
rect 19012 2248 19054 2288
rect 19094 2248 19136 2288
rect 19176 2248 19212 2288
rect 18772 0 19212 2248
rect 20012 9092 20452 11844
rect 20012 9052 20048 9092
rect 20088 9052 20130 9092
rect 20170 9052 20212 9092
rect 20252 9052 20294 9092
rect 20334 9052 20376 9092
rect 20416 9052 20452 9092
rect 20012 7580 20452 9052
rect 20012 7540 20048 7580
rect 20088 7540 20130 7580
rect 20170 7540 20212 7580
rect 20252 7540 20294 7580
rect 20334 7540 20376 7580
rect 20416 7540 20452 7580
rect 20012 6068 20452 7540
rect 33892 9848 34332 11844
rect 33892 9808 33928 9848
rect 33968 9808 34010 9848
rect 34050 9808 34092 9848
rect 34132 9808 34174 9848
rect 34214 9808 34256 9848
rect 34296 9808 34332 9848
rect 33892 8336 34332 9808
rect 33892 8296 33928 8336
rect 33968 8296 34010 8336
rect 34050 8296 34092 8336
rect 34132 8296 34174 8336
rect 34214 8296 34256 8336
rect 34296 8296 34332 8336
rect 30316 7496 30356 7505
rect 30316 6236 30356 7456
rect 30316 6187 30356 6196
rect 33892 6824 34332 8296
rect 33892 6784 33928 6824
rect 33968 6784 34010 6824
rect 34050 6784 34092 6824
rect 34132 6784 34174 6824
rect 34214 6784 34256 6824
rect 34296 6784 34332 6824
rect 20012 6028 20048 6068
rect 20088 6028 20130 6068
rect 20170 6028 20212 6068
rect 20252 6028 20294 6068
rect 20334 6028 20376 6068
rect 20416 6028 20452 6068
rect 20012 4556 20452 6028
rect 20012 4516 20048 4556
rect 20088 4516 20130 4556
rect 20170 4516 20212 4556
rect 20252 4516 20294 4556
rect 20334 4516 20376 4556
rect 20416 4516 20452 4556
rect 20012 3044 20452 4516
rect 20012 3004 20048 3044
rect 20088 3004 20130 3044
rect 20170 3004 20212 3044
rect 20252 3004 20294 3044
rect 20334 3004 20376 3044
rect 20416 3004 20452 3044
rect 20012 1532 20452 3004
rect 20012 1492 20048 1532
rect 20088 1492 20130 1532
rect 20170 1492 20212 1532
rect 20252 1492 20294 1532
rect 20334 1492 20376 1532
rect 20416 1492 20452 1532
rect 20012 0 20452 1492
rect 33892 5312 34332 6784
rect 33892 5272 33928 5312
rect 33968 5272 34010 5312
rect 34050 5272 34092 5312
rect 34132 5272 34174 5312
rect 34214 5272 34256 5312
rect 34296 5272 34332 5312
rect 33892 3800 34332 5272
rect 33892 3760 33928 3800
rect 33968 3760 34010 3800
rect 34050 3760 34092 3800
rect 34132 3760 34174 3800
rect 34214 3760 34256 3800
rect 34296 3760 34332 3800
rect 33892 2288 34332 3760
rect 33892 2248 33928 2288
rect 33968 2248 34010 2288
rect 34050 2248 34092 2288
rect 34132 2248 34174 2288
rect 34214 2248 34256 2288
rect 34296 2248 34332 2288
rect 33892 0 34332 2248
rect 35132 9092 35572 11844
rect 35132 9052 35168 9092
rect 35208 9052 35250 9092
rect 35290 9052 35332 9092
rect 35372 9052 35414 9092
rect 35454 9052 35496 9092
rect 35536 9052 35572 9092
rect 35132 7580 35572 9052
rect 35132 7540 35168 7580
rect 35208 7540 35250 7580
rect 35290 7540 35332 7580
rect 35372 7540 35414 7580
rect 35454 7540 35496 7580
rect 35536 7540 35572 7580
rect 35132 6068 35572 7540
rect 35132 6028 35168 6068
rect 35208 6028 35250 6068
rect 35290 6028 35332 6068
rect 35372 6028 35414 6068
rect 35454 6028 35496 6068
rect 35536 6028 35572 6068
rect 35132 4556 35572 6028
rect 35132 4516 35168 4556
rect 35208 4516 35250 4556
rect 35290 4516 35332 4556
rect 35372 4516 35414 4556
rect 35454 4516 35496 4556
rect 35536 4516 35572 4556
rect 35132 3044 35572 4516
rect 35132 3004 35168 3044
rect 35208 3004 35250 3044
rect 35290 3004 35332 3044
rect 35372 3004 35414 3044
rect 35454 3004 35496 3044
rect 35536 3004 35572 3044
rect 35132 1532 35572 3004
rect 35132 1492 35168 1532
rect 35208 1492 35250 1532
rect 35290 1492 35332 1532
rect 35372 1492 35414 1532
rect 35454 1492 35496 1532
rect 35536 1492 35572 1532
rect 35132 0 35572 1492
use sg13g2_mux4_1  _036_
timestamp 1677257233
transform 1 0 21984 0 1 3024
box -48 -56 2064 834
use sg13g2_nor2_1  _037_
timestamp 1676627187
transform 1 0 24096 0 -1 4536
box -48 -56 432 834
use sg13g2_nor2b_1  _038_
timestamp 1685181386
transform 1 0 22656 0 -1 4536
box -54 -56 528 834
use sg13g2_nor2_1  _039_
timestamp 1676627187
transform 1 0 23232 0 1 4536
box -48 -56 432 834
use sg13g2_nor3_1  _040_
timestamp 1676639442
transform -1 0 24480 0 1 3024
box -48 -56 528 834
use sg13g2_nor2b_1  _041_
timestamp 1685181386
transform 1 0 22176 0 -1 4536
box -54 -56 528 834
use sg13g2_o21ai_1  _042_
timestamp 1685175443
transform 1 0 23136 0 -1 4536
box -48 -56 538 834
use sg13g2_o21ai_1  _043_
timestamp 1685175443
transform 1 0 23040 0 -1 3024
box -48 -56 538 834
use sg13g2_o21ai_1  _044_
timestamp 1685175443
transform -1 0 24096 0 -1 4536
box -48 -56 538 834
use sg13g2_nor2_1  _045_
timestamp 1676627187
transform -1 0 24864 0 -1 4536
box -48 -56 432 834
use sg13g2_mux4_1  _046_
timestamp 1677257233
transform 1 0 11904 0 1 3024
box -48 -56 2064 834
use sg13g2_nor2_1  _047_
timestamp 1676627187
transform -1 0 15264 0 -1 3024
box -48 -56 432 834
use sg13g2_nor2b_1  _048_
timestamp 1685181386
transform 1 0 12576 0 -1 4536
box -54 -56 528 834
use sg13g2_nor2_1  _049_
timestamp 1676627187
transform 1 0 12768 0 1 4536
box -48 -56 432 834
use sg13g2_nor3_1  _050_
timestamp 1676639442
transform -1 0 13536 0 -1 4536
box -48 -56 528 834
use sg13g2_nor2b_1  _051_
timestamp 1685181386
transform 1 0 13920 0 1 3024
box -54 -56 528 834
use sg13g2_o21ai_1  _052_
timestamp 1685175443
transform 1 0 13440 0 -1 3024
box -48 -56 538 834
use sg13g2_o21ai_1  _053_
timestamp 1685175443
transform 1 0 14592 0 1 3024
box -48 -56 538 834
use sg13g2_o21ai_1  _054_
timestamp 1685175443
transform 1 0 15072 0 -1 4536
box -48 -56 538 834
use sg13g2_nor2_1  _055_
timestamp 1676627187
transform 1 0 15168 0 1 3024
box -48 -56 432 834
use sg13g2_mux4_1  _056_
timestamp 1677257233
transform 1 0 16512 0 1 7560
box -48 -56 2064 834
use sg13g2_nor2_1  _057_
timestamp 1676627187
transform -1 0 18912 0 1 7560
box -48 -56 432 834
use sg13g2_nor2b_1  _058_
timestamp 1685181386
transform 1 0 14592 0 1 7560
box -54 -56 528 834
use sg13g2_nor2_1  _059_
timestamp 1676627187
transform 1 0 14976 0 -1 9072
box -48 -56 432 834
use sg13g2_nor3_1  _060_
timestamp 1676639442
transform -1 0 15552 0 1 7560
box -48 -56 528 834
use sg13g2_nor2b_1  _061_
timestamp 1685181386
transform 1 0 15840 0 -1 7560
box -54 -56 528 834
use sg13g2_o21ai_1  _062_
timestamp 1685175443
transform 1 0 15552 0 1 7560
box -48 -56 538 834
use sg13g2_o21ai_1  _063_
timestamp 1685175443
transform 1 0 16608 0 -1 7560
box -48 -56 538 834
use sg13g2_o21ai_1  _064_
timestamp 1685175443
transform 1 0 16032 0 1 7560
box -48 -56 538 834
use sg13g2_nor2_1  _065_
timestamp 1676627187
transform -1 0 17952 0 -1 9072
box -48 -56 432 834
use sg13g2_mux4_1  _066_
timestamp 1677257233
transform -1 0 32256 0 -1 7560
box -48 -56 2064 834
use sg13g2_nor2_1  _067_
timestamp 1676627187
transform 1 0 29760 0 1 6048
box -48 -56 432 834
use sg13g2_nor2b_1  _068_
timestamp 1685181386
transform -1 0 29760 0 -1 7560
box -54 -56 528 834
use sg13g2_nor2_1  _069_
timestamp 1676627187
transform 1 0 28416 0 -1 7560
box -48 -56 432 834
use sg13g2_nor3_1  _070_
timestamp 1676639442
transform -1 0 30240 0 1 7560
box -48 -56 528 834
use sg13g2_nor2b_1  _071_
timestamp 1685181386
transform 1 0 28800 0 -1 7560
box -54 -56 528 834
use sg13g2_o21ai_1  _072_
timestamp 1685175443
transform -1 0 30240 0 -1 7560
box -48 -56 538 834
use sg13g2_o21ai_1  _073_
timestamp 1685175443
transform 1 0 29280 0 1 7560
box -48 -56 538 834
use sg13g2_o21ai_1  _074_
timestamp 1685175443
transform -1 0 29184 0 1 6048
box -48 -56 538 834
use sg13g2_nor2_1  _075_
timestamp 1676627187
transform -1 0 30624 0 1 7560
box -48 -56 432 834
use sg13g2_dlhq_1  _076_
timestamp 1678805552
transform 1 0 17760 0 -1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _077_
timestamp 1678805552
transform -1 0 27552 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _078_
timestamp 1678805552
transform 1 0 21120 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _079_
timestamp 1678805552
transform 1 0 9024 0 -1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _080_
timestamp 1678805552
transform 1 0 9696 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _081_
timestamp 1678805552
transform -1 0 17760 0 1 3024
box -50 -56 1692 834
use sg13g2_dlhq_1  _082_
timestamp 1678805552
transform 1 0 11520 0 -1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _083_
timestamp 1678805552
transform 1 0 12096 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _084_
timestamp 1678805552
transform -1 0 21600 0 1 7560
box -50 -56 1692 834
use sg13g2_dlhq_1  _085_
timestamp 1678805552
transform 1 0 26112 0 1 6048
box -50 -56 1692 834
use sg13g2_dlhq_1  _086_
timestamp 1678805552
transform 1 0 27552 0 1 4536
box -50 -56 1692 834
use sg13g2_dlhq_1  _087_
timestamp 1678805552
transform 1 0 25824 0 -1 7560
box -50 -56 1692 834
use sg13g2_buf_1  _089_
timestamp 1676381911
transform 1 0 42048 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _090_
timestamp 1676381911
transform 1 0 42432 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _091_
timestamp 1676381911
transform 1 0 42816 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _092_
timestamp 1676381911
transform 1 0 41664 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _093_
timestamp 1676381911
transform 1 0 42048 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _094_
timestamp 1676381911
transform 1 0 42048 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _095_
timestamp 1676381911
transform 1 0 41280 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _096_
timestamp 1676381911
transform 1 0 42432 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _097_
timestamp 1676381911
transform 1 0 40224 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _098_
timestamp 1676381911
transform 1 0 41568 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _099_
timestamp 1676381911
transform 1 0 38208 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _100_
timestamp 1676381911
transform 1 0 38304 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _101_
timestamp 1676381911
transform 1 0 38880 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _102_
timestamp 1676381911
transform 1 0 39744 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _103_
timestamp 1676381911
transform 1 0 38976 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _104_
timestamp 1676381911
transform 1 0 36960 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _105_
timestamp 1676381911
transform 1 0 35616 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _106_
timestamp 1676381911
transform 1 0 35232 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _107_
timestamp 1676381911
transform 1 0 34560 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _108_
timestamp 1676381911
transform 1 0 33216 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _109_
timestamp 1676381911
transform 1 0 17280 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _110_
timestamp 1676381911
transform 1 0 25536 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _111_
timestamp 1676381911
transform 1 0 20736 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  _112_
timestamp 1676381911
transform 1 0 8640 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _113_
timestamp 1676381911
transform 1 0 9312 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _114_
timestamp 1676381911
transform 1 0 15744 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _115_
timestamp 1676381911
transform 1 0 11232 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _116_
timestamp 1676381911
transform 1 0 11712 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _117_
timestamp 1676381911
transform 1 0 19584 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _118_
timestamp 1676381911
transform 1 0 25920 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _119_
timestamp 1676381911
transform 1 0 27648 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _120_
timestamp 1676381911
transform 1 0 25440 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _121_
timestamp 1676381911
transform 1 0 21120 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _122_
timestamp 1676381911
transform -1 0 41376 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _123_
timestamp 1676381911
transform -1 0 39072 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _124_
timestamp 1676381911
transform -1 0 43488 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  _125_
timestamp 1676381911
transform -1 0 40608 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _126_
timestamp 1676381911
transform -1 0 38592 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _127_
timestamp 1676381911
transform -1 0 39648 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _128_
timestamp 1676381911
transform -1 0 40992 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _129_
timestamp 1676381911
transform -1 0 39264 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _130_
timestamp 1676381911
transform -1 0 38688 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _131_
timestamp 1676381911
transform -1 0 38208 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _132_
timestamp 1676381911
transform -1 0 40992 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _133_
timestamp 1676381911
transform -1 0 40512 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _134_
timestamp 1676381911
transform 1 0 34560 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _135_
timestamp 1676381911
transform -1 0 35328 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _136_
timestamp 1676381911
transform -1 0 35808 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _137_
timestamp 1676381911
transform -1 0 35712 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _138_
timestamp 1676381911
transform 1 0 35040 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _139_
timestamp 1676381911
transform 1 0 35424 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _140_
timestamp 1676381911
transform 1 0 34560 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _141_
timestamp 1676381911
transform -1 0 31296 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _142_
timestamp 1676381911
transform -1 0 17376 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _143_
timestamp 1676381911
transform -1 0 12384 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _144_
timestamp 1676381911
transform -1 0 21600 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _145_
timestamp 1676381911
transform 1 0 3744 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _146_
timestamp 1676381911
transform 1 0 3360 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _147_
timestamp 1676381911
transform 1 0 2880 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _148_
timestamp 1676381911
transform 1 0 3264 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _149_
timestamp 1676381911
transform -1 0 31584 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _150_
timestamp 1676381911
transform -1 0 18336 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _151_
timestamp 1676381911
transform -1 0 11904 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _152_
timestamp 1676381911
transform -1 0 22656 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _153_
timestamp 1676381911
transform -1 0 32352 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _154_
timestamp 1676381911
transform -1 0 18240 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _155_
timestamp 1676381911
transform -1 0 14304 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _156_
timestamp 1676381911
transform -1 0 25248 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _157_
timestamp 1676381911
transform -1 0 31968 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _158_
timestamp 1676381911
transform -1 0 17856 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _159_
timestamp 1676381911
transform 1 0 12576 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _160_
timestamp 1676381911
transform -1 0 21984 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _161_
timestamp 1676381911
transform -1 0 43008 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _162_
timestamp 1676381911
transform -1 0 43680 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _163_
timestamp 1676381911
transform -1 0 43200 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _164_
timestamp 1676381911
transform -1 0 44736 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _165_
timestamp 1676381911
transform -1 0 44064 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _166_
timestamp 1676381911
transform -1 0 23520 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _167_
timestamp 1676381911
transform -1 0 23904 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _168_
timestamp 1676381911
transform -1 0 23136 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _169_
timestamp 1676381911
transform -1 0 28896 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _170_
timestamp 1676381911
transform -1 0 14592 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _171_
timestamp 1676381911
transform 1 0 11808 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _172_
timestamp 1676381911
transform -1 0 24288 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _173_
timestamp 1676381911
transform -1 0 29952 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _174_
timestamp 1676381911
transform 1 0 14976 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _175_
timestamp 1676381911
transform 1 0 12192 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _176_
timestamp 1676381911
transform -1 0 24864 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  _177_
timestamp 1676381911
transform -1 0 43968 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _178_
timestamp 1676381911
transform -1 0 42816 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _179_
timestamp 1676381911
transform -1 0 43392 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _180_
timestamp 1676381911
transform -1 0 42432 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _181_
timestamp 1676381911
transform -1 0 43776 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _182_
timestamp 1676381911
transform -1 0 44352 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _183_
timestamp 1676381911
transform -1 0 43584 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _184_
timestamp 1676381911
transform -1 0 43296 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  _185_
timestamp 1676381911
transform -1 0 29280 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  _186_
timestamp 1676381911
transform 1 0 15936 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _187_
timestamp 1676381911
transform 1 0 14400 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _188_
timestamp 1676381911
transform -1 0 23040 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _189_
timestamp 1676381911
transform -1 0 29760 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  _190_
timestamp 1676381911
transform 1 0 16320 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  _191_
timestamp 1676381911
transform 1 0 13536 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  _192_
timestamp 1676381911
transform -1 0 23904 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  _193_
timestamp 1676381911
transform -1 0 40992 0 1 3024
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 40896 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 37728 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 35424 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 39648 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 44160 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform -1 0 42624 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform -1 0 40896 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform 1 0 37440 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform -1 0 35424 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 39360 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 41472 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform -1 0 42336 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform -1 0 40608 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 38016 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform -1 0 35136 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 41664 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 41184 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform -1 0 42048 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform -1 0 40320 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 37152 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform -1 0 34848 0 1 4536
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform -1 0 41664 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 40896 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 43776 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform -1 0 40032 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 39936 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform -1 0 41376 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 43488 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform -1 0 41760 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform -1 0 39744 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 39648 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform -1 0 41088 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 40608 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform 1 0 43776 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform -1 0 39456 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 39360 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform -1 0 40800 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 41184 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 43488 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform -1 0 39168 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 38592 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform -1 0 40512 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 42624 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 44064 0 -1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform -1 0 38880 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 38304 0 -1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform -1 0 40224 0 -1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 40320 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform 1 0 44064 0 1 6048
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform -1 0 38208 0 -1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 38016 0 1 7560
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform 1 0 39936 0 1 3024
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 44544 0 1 9072
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform -1 0 44064 0 -1 9072
box -48 -56 336 834
use sg13g2_buf_1  fanout5
timestamp 1676381911
transform -1 0 21984 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  fanout6
timestamp 1676381911
transform 1 0 22080 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_0_0
timestamp 1677580104
transform 1 0 1152 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_2
timestamp 1677579658
transform 1 0 1344 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 1824 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 2496 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_25
timestamp 1679581782
transform 1 0 3552 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_32
timestamp 1679581782
transform 1 0 4224 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_43
timestamp 1679581782
transform 1 0 5280 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_50
timestamp 1679581782
transform 1 0 5952 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_61
timestamp 1679581782
transform 1 0 7008 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_68
timestamp 1679581782
transform 1 0 7680 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_79
timestamp 1679581782
transform 1 0 8736 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_86
timestamp 1679581782
transform 1 0 9408 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_93
timestamp 1679581782
transform 1 0 10080 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_100
timestamp 1679581782
transform 1 0 10752 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_107
timestamp 1679581782
transform 1 0 11424 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_114
timestamp 1679581782
transform 1 0 12096 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_121
timestamp 1679581782
transform 1 0 12768 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_128
timestamp 1679581782
transform 1 0 13440 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_135
timestamp 1679581782
transform 1 0 14112 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_142
timestamp 1679581782
transform 1 0 14784 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_149
timestamp 1679581782
transform 1 0 15456 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_156
timestamp 1679581782
transform 1 0 16128 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_163
timestamp 1679581782
transform 1 0 16800 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_170
timestamp 1679581782
transform 1 0 17472 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_177
timestamp 1679581782
transform 1 0 18144 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_184
timestamp 1679581782
transform 1 0 18816 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_191
timestamp 1679581782
transform 1 0 19488 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_198
timestamp 1679581782
transform 1 0 20160 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_205
timestamp 1679581782
transform 1 0 20832 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_212
timestamp 1679581782
transform 1 0 21504 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_219
timestamp 1679581782
transform 1 0 22176 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_226
timestamp 1679581782
transform 1 0 22848 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_233
timestamp 1679581782
transform 1 0 23520 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_240
timestamp 1679581782
transform 1 0 24192 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_247
timestamp 1679581782
transform 1 0 24864 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_254
timestamp 1679581782
transform 1 0 25536 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_261
timestamp 1679581782
transform 1 0 26208 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_268
timestamp 1679581782
transform 1 0 26880 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_275
timestamp 1679581782
transform 1 0 27552 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_282
timestamp 1679581782
transform 1 0 28224 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_289
timestamp 1679581782
transform 1 0 28896 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_296
timestamp 1679581782
transform 1 0 29568 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_303
timestamp 1679581782
transform 1 0 30240 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_310
timestamp 1679581782
transform 1 0 30912 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_317
timestamp 1679581782
transform 1 0 31584 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_324
timestamp 1679581782
transform 1 0 32256 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_331
timestamp 1679581782
transform 1 0 32928 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_338
timestamp 1679581782
transform 1 0 33600 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_345
timestamp 1679581782
transform 1 0 34272 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_352
timestamp 1679581782
transform 1 0 34944 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_359
timestamp 1679581782
transform 1 0 35616 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_366
timestamp 1679581782
transform 1 0 36288 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_373
timestamp 1679581782
transform 1 0 36960 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_380
timestamp 1679581782
transform 1 0 37632 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_387
timestamp 1679581782
transform 1 0 38304 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_394
timestamp 1679581782
transform 1 0 38976 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_401
timestamp 1679581782
transform 1 0 39648 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_408
timestamp 1679581782
transform 1 0 40320 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_415
timestamp 1679581782
transform 1 0 40992 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_422
timestamp 1679581782
transform 1 0 41664 0 1 1512
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_429
timestamp 1679581782
transform 1 0 42336 0 1 1512
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_436
timestamp 1677580104
transform 1 0 43008 0 1 1512
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_438
timestamp 1677579658
transform 1 0 43200 0 1 1512
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 1152 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 1824 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 2496 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 3168 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 3840 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 4512 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 5184 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 5856 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 6528 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 7200 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 7872 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_77
timestamp 1679577901
transform 1 0 8544 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_81
timestamp 1677579658
transform 1 0 8928 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_99
timestamp 1679581782
transform 1 0 10656 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_106
timestamp 1679581782
transform 1 0 11328 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_117
timestamp 1677580104
transform 1 0 12384 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_123
timestamp 1679577901
transform 1 0 12960 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_127
timestamp 1677579658
transform 1 0 13344 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_137
timestamp 1677579658
transform 1 0 14304 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_142
timestamp 1677579658
transform 1 0 14784 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 15264 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 15936 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 16608 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 17280 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 17952 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 18624 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 19296 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19968 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 20640 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 21312 0 -1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_217
timestamp 1677580104
transform 1 0 21984 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_219
timestamp 1677579658
transform 1 0 22176 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_241
timestamp 1679581782
transform 1 0 24288 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_248
timestamp 1679581782
transform 1 0 24960 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_255
timestamp 1679581782
transform 1 0 25632 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_262
timestamp 1679581782
transform 1 0 26304 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_269
timestamp 1679581782
transform 1 0 26976 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_276
timestamp 1679581782
transform 1 0 27648 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_283
timestamp 1679581782
transform 1 0 28320 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_290
timestamp 1679581782
transform 1 0 28992 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_297
timestamp 1679581782
transform 1 0 29664 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_304
timestamp 1679581782
transform 1 0 30336 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_311
timestamp 1679581782
transform 1 0 31008 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_318
timestamp 1679581782
transform 1 0 31680 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_325
timestamp 1679581782
transform 1 0 32352 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_332
timestamp 1679581782
transform 1 0 33024 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_339
timestamp 1679581782
transform 1 0 33696 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_346
timestamp 1679581782
transform 1 0 34368 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_353
timestamp 1679581782
transform 1 0 35040 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_360
timestamp 1679581782
transform 1 0 35712 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_367
timestamp 1679581782
transform 1 0 36384 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_374
timestamp 1679581782
transform 1 0 37056 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_381
timestamp 1679581782
transform 1 0 37728 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_388
timestamp 1679577901
transform 1 0 38400 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_392
timestamp 1677579658
transform 1 0 38784 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_401
timestamp 1677580104
transform 1 0 39648 0 -1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_403
timestamp 1677579658
transform 1 0 39840 0 -1 3024
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_425
timestamp 1677579658
transform 1 0 41952 0 -1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 42816 0 -1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_1_441
timestamp 1679577901
transform 1 0 43488 0 -1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_1_445
timestamp 1677580104
transform 1 0 43872 0 -1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 1152 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 1824 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 2496 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 3168 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 3840 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 4512 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 5184 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 5856 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 6528 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 7200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 7872 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_77
timestamp 1677579658
transform 1 0 8544 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_82
timestamp 1677580104
transform 1 0 9024 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_84
timestamp 1677579658
transform 1 0 9216 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_106
timestamp 1677580104
transform 1 0 11328 0 1 3024
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_138
timestamp 1677580104
transform 1 0 14400 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_145
timestamp 1677579658
transform 1 0 15072 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_150
timestamp 1677580104
transform 1 0 15552 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_2_173
timestamp 1679581782
transform 1 0 17760 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_180
timestamp 1679581782
transform 1 0 18432 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_187
timestamp 1679581782
transform 1 0 19104 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_194
timestamp 1679581782
transform 1 0 19776 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_201
timestamp 1679581782
transform 1 0 20448 0 1 3024
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_208
timestamp 1677579658
transform 1 0 21120 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_251
timestamp 1677580104
transform 1 0 25248 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_253
timestamp 1677579658
transform 1 0 25440 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_275
timestamp 1679581782
transform 1 0 27552 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_282
timestamp 1679581782
transform 1 0 28224 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_289
timestamp 1679581782
transform 1 0 28896 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_296
timestamp 1679581782
transform 1 0 29568 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_303
timestamp 1679581782
transform 1 0 30240 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_310
timestamp 1679581782
transform 1 0 30912 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_317
timestamp 1679581782
transform 1 0 31584 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_324
timestamp 1679581782
transform 1 0 32256 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_331
timestamp 1679581782
transform 1 0 32928 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_338
timestamp 1679581782
transform 1 0 33600 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_345
timestamp 1679581782
transform 1 0 34272 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_352
timestamp 1679581782
transform 1 0 34944 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_359
timestamp 1679581782
transform 1 0 35616 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_366
timestamp 1679581782
transform 1 0 36288 0 1 3024
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_373
timestamp 1679581782
transform 1 0 36960 0 1 3024
box -48 -56 720 834
use sg13g2_fill_2  FILLER_2_380
timestamp 1677580104
transform 1 0 37632 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_390
timestamp 1677579658
transform 1 0 38592 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_395
timestamp 1677580104
transform 1 0 39072 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_397
timestamp 1677579658
transform 1 0 39264 0 1 3024
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_415
timestamp 1677580104
transform 1 0 40992 0 1 3024
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_417
timestamp 1677579658
transform 1 0 41184 0 1 3024
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_438
timestamp 1679581782
transform 1 0 43200 0 1 3024
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_445
timestamp 1679577901
transform 1 0 43872 0 1 3024
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_449
timestamp 1677580104
transform 1 0 44256 0 1 3024
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 1152 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 1824 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 2496 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 3168 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 3840 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 4512 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 5184 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 5856 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 6528 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 7200 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 7872 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 8544 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 9216 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 9888 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 10560 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_105
timestamp 1679577901
transform 1 0 11232 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_109
timestamp 1677580104
transform 1 0 11616 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 13920 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_140
timestamp 1679577901
transform 1 0 14592 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_144
timestamp 1677579658
transform 1 0 14976 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_150
timestamp 1679581782
transform 1 0 15552 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_157
timestamp 1679581782
transform 1 0 16224 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_164
timestamp 1679577901
transform 1 0 16896 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_172
timestamp 1677579658
transform 1 0 17664 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_190
timestamp 1679581782
transform 1 0 19392 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_197
timestamp 1679581782
transform 1 0 20064 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_204
timestamp 1679581782
transform 1 0 20736 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_211
timestamp 1679581782
transform 1 0 21408 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_218
timestamp 1677579658
transform 1 0 22080 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_247
timestamp 1679581782
transform 1 0 24864 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_254
timestamp 1679581782
transform 1 0 25536 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_261
timestamp 1679581782
transform 1 0 26208 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_268
timestamp 1679581782
transform 1 0 26880 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_275
timestamp 1677579658
transform 1 0 27552 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679581782
transform 1 0 28032 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679581782
transform 1 0 28704 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1679581782
transform 1 0 29376 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1679581782
transform 1 0 30048 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1679581782
transform 1 0 30720 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_315
timestamp 1679581782
transform 1 0 31392 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_322
timestamp 1679581782
transform 1 0 32064 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_3_329
timestamp 1679577901
transform 1 0 32736 0 -1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_333
timestamp 1677579658
transform 1 0 33120 0 -1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_338
timestamp 1679581782
transform 1 0 33600 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_345
timestamp 1679581782
transform 1 0 34272 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_352
timestamp 1679581782
transform 1 0 34944 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_359
timestamp 1679581782
transform 1 0 35616 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_366
timestamp 1679581782
transform 1 0 36288 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_373
timestamp 1679581782
transform 1 0 36960 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_380
timestamp 1679581782
transform 1 0 37632 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_391
timestamp 1679581782
transform 1 0 38688 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_398
timestamp 1679581782
transform 1 0 39360 0 -1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_405
timestamp 1677580104
transform 1 0 40032 0 -1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_419
timestamp 1679581782
transform 1 0 41376 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_430
timestamp 1679581782
transform 1 0 42432 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_437
timestamp 1679581782
transform 1 0 43104 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_444
timestamp 1679581782
transform 1 0 43776 0 -1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 1152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 1824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 2496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 3168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 3840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 4512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 5184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 5856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 6528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 7200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679581782
transform 1 0 7872 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 8544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 9216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 9888 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 10560 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679581782
transform 1 0 11232 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679581782
transform 1 0 11904 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_119
timestamp 1677580104
transform 1 0 12576 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_125
timestamp 1679581782
transform 1 0 13152 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_132
timestamp 1679581782
transform 1 0 13824 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_139
timestamp 1679581782
transform 1 0 14496 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_146
timestamp 1679581782
transform 1 0 15168 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_153
timestamp 1679581782
transform 1 0 15840 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_160
timestamp 1679581782
transform 1 0 16512 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_167
timestamp 1679581782
transform 1 0 17184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_174
timestamp 1679581782
transform 1 0 17856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_181
timestamp 1679581782
transform 1 0 18528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_188
timestamp 1679581782
transform 1 0 19200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_195
timestamp 1679581782
transform 1 0 19872 0 1 4536
box -48 -56 720 834
use sg13g2_fill_2  FILLER_4_202
timestamp 1677580104
transform 1 0 20544 0 1 4536
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_225
timestamp 1679577901
transform 1 0 22752 0 1 4536
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_229
timestamp 1677579658
transform 1 0 23136 0 1 4536
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_234
timestamp 1679581782
transform 1 0 23616 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_241
timestamp 1679581782
transform 1 0 24288 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_248
timestamp 1679581782
transform 1 0 24960 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_255
timestamp 1679581782
transform 1 0 25632 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_262
timestamp 1679581782
transform 1 0 26304 0 1 4536
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_269
timestamp 1679577901
transform 1 0 26976 0 1 4536
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_273
timestamp 1677580104
transform 1 0 27360 0 1 4536
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_292
timestamp 1679581782
transform 1 0 29184 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_299
timestamp 1679581782
transform 1 0 29856 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_306
timestamp 1679581782
transform 1 0 30528 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_313
timestamp 1679581782
transform 1 0 31200 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_320
timestamp 1679581782
transform 1 0 31872 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_327
timestamp 1679581782
transform 1 0 32544 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_334
timestamp 1679581782
transform 1 0 33216 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_341
timestamp 1679581782
transform 1 0 33888 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_360
timestamp 1679581782
transform 1 0 35712 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_367
timestamp 1679581782
transform 1 0 36384 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_374
timestamp 1679581782
transform 1 0 37056 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_381
timestamp 1679581782
transform 1 0 37728 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_388
timestamp 1679581782
transform 1 0 38400 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_395
timestamp 1679581782
transform 1 0 39072 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_402
timestamp 1679581782
transform 1 0 39744 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_409
timestamp 1679581782
transform 1 0 40416 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_416
timestamp 1679581782
transform 1 0 41088 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_423
timestamp 1679581782
transform 1 0 41760 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_430
timestamp 1679581782
transform 1 0 42432 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_437
timestamp 1679581782
transform 1 0 43104 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_444
timestamp 1679581782
transform 1 0 43776 0 1 4536
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 1152 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 1824 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 2496 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 3168 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 3840 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 4512 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 5184 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 5856 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 6528 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 7200 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 7872 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 8544 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_84
timestamp 1679581782
transform 1 0 9216 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_91
timestamp 1679581782
transform 1 0 9888 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_98
timestamp 1679581782
transform 1 0 10560 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679581782
transform 1 0 11232 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_112
timestamp 1679581782
transform 1 0 11904 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679581782
transform 1 0 12576 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_126
timestamp 1679581782
transform 1 0 13248 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_133
timestamp 1679581782
transform 1 0 13920 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679581782
transform 1 0 14592 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 15264 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 15936 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 16608 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 17280 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679581782
transform 1 0 17952 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679581782
transform 1 0 18624 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679581782
transform 1 0 19296 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679581782
transform 1 0 19968 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679581782
transform 1 0 20640 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679581782
transform 1 0 21312 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679581782
transform 1 0 21984 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_224
timestamp 1679581782
transform 1 0 22656 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_231
timestamp 1679581782
transform 1 0 23328 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_238
timestamp 1679581782
transform 1 0 24000 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_245
timestamp 1679581782
transform 1 0 24672 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_252
timestamp 1679581782
transform 1 0 25344 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_259
timestamp 1679581782
transform 1 0 26016 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_266
timestamp 1679581782
transform 1 0 26688 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_273
timestamp 1679581782
transform 1 0 27360 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_280
timestamp 1679581782
transform 1 0 28032 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_287
timestamp 1679581782
transform 1 0 28704 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_294
timestamp 1679581782
transform 1 0 29376 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_301
timestamp 1679581782
transform 1 0 30048 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_308
timestamp 1679581782
transform 1 0 30720 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_315
timestamp 1679581782
transform 1 0 31392 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_322
timestamp 1679581782
transform 1 0 32064 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_329
timestamp 1679581782
transform 1 0 32736 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_336
timestamp 1679581782
transform 1 0 33408 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_343
timestamp 1679577901
transform 1 0 34080 0 -1 6048
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_347
timestamp 1677579658
transform 1 0 34464 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_352
timestamp 1679581782
transform 1 0 34944 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_359
timestamp 1679581782
transform 1 0 35616 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_366
timestamp 1679581782
transform 1 0 36288 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_373
timestamp 1679581782
transform 1 0 36960 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_380
timestamp 1679581782
transform 1 0 37632 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_387
timestamp 1679581782
transform 1 0 38304 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_394
timestamp 1679581782
transform 1 0 38976 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_401
timestamp 1679581782
transform 1 0 39648 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_408
timestamp 1679581782
transform 1 0 40320 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_415
timestamp 1679581782
transform 1 0 40992 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_422
timestamp 1679581782
transform 1 0 41664 0 -1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_429
timestamp 1679581782
transform 1 0 42336 0 -1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_436
timestamp 1677579658
transform 1 0 43008 0 -1 6048
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_450
timestamp 1677579658
transform 1 0 44352 0 -1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 1152 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 1824 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 2496 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 3168 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 3840 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 4512 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 5184 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 5856 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 6528 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 7200 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 7872 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 8544 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 9216 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 9888 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 10560 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 11232 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 11904 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 12576 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 13248 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 13920 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 14592 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 15264 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 15936 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 16608 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 17280 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 17952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 18624 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 19296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 19968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 20640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 21312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 21984 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_224
timestamp 1679581782
transform 1 0 22656 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_231
timestamp 1679581782
transform 1 0 23328 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_238
timestamp 1679581782
transform 1 0 24000 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1679581782
transform 1 0 24672 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1679581782
transform 1 0 25344 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_259
timestamp 1677579658
transform 1 0 26016 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_277
timestamp 1679581782
transform 1 0 27744 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_284
timestamp 1677580104
transform 1 0 28416 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_286
timestamp 1677579658
transform 1 0 28608 0 1 6048
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_292
timestamp 1677580104
transform 1 0 29184 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_302
timestamp 1679581782
transform 1 0 30144 0 1 6048
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_309
timestamp 1677579658
transform 1 0 30816 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_314
timestamp 1679581782
transform 1 0 31296 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_321
timestamp 1679581782
transform 1 0 31968 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_328
timestamp 1679581782
transform 1 0 32640 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_335
timestamp 1679581782
transform 1 0 33312 0 1 6048
box -48 -56 720 834
use sg13g2_decap_4  FILLER_6_342
timestamp 1679577901
transform 1 0 33984 0 1 6048
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_346
timestamp 1677580104
transform 1 0 34368 0 1 6048
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_352
timestamp 1677580104
transform 1 0 34944 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_354
timestamp 1677579658
transform 1 0 35136 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_363
timestamp 1679581782
transform 1 0 36000 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_370
timestamp 1677580104
transform 1 0 36672 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_372
timestamp 1677579658
transform 1 0 36864 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_377
timestamp 1679581782
transform 1 0 37344 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_384
timestamp 1679581782
transform 1 0 38016 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_391
timestamp 1679581782
transform 1 0 38688 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_398
timestamp 1679581782
transform 1 0 39360 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_405
timestamp 1679581782
transform 1 0 40032 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_412
timestamp 1679581782
transform 1 0 40704 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_419
timestamp 1677580104
transform 1 0 41376 0 1 6048
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_425
timestamp 1679581782
transform 1 0 41952 0 1 6048
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_432
timestamp 1679581782
transform 1 0 42624 0 1 6048
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_439
timestamp 1677580104
transform 1 0 43296 0 1 6048
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_450
timestamp 1677579658
transform 1 0 44352 0 1 6048
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 1152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 1824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 2496 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_21
timestamp 1677580104
transform 1 0 3168 0 -1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_31
timestamp 1679581782
transform 1 0 4128 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_38
timestamp 1679581782
transform 1 0 4800 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_45
timestamp 1679581782
transform 1 0 5472 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_52
timestamp 1679581782
transform 1 0 6144 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_59
timestamp 1679581782
transform 1 0 6816 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_66
timestamp 1679581782
transform 1 0 7488 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_73
timestamp 1679581782
transform 1 0 8160 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_80
timestamp 1679581782
transform 1 0 8832 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_87
timestamp 1679581782
transform 1 0 9504 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_94
timestamp 1679581782
transform 1 0 10176 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_101
timestamp 1679581782
transform 1 0 10848 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_125
timestamp 1679581782
transform 1 0 13152 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_132
timestamp 1679581782
transform 1 0 13824 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_139
timestamp 1679577901
transform 1 0 14496 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_143
timestamp 1677579658
transform 1 0 14880 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_148
timestamp 1677579658
transform 1 0 15360 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_158
timestamp 1677580104
transform 1 0 16320 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_160
timestamp 1677579658
transform 1 0 16512 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_166
timestamp 1679577901
transform 1 0 17088 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_178
timestamp 1679581782
transform 1 0 18240 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_185
timestamp 1679581782
transform 1 0 18912 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_192
timestamp 1679581782
transform 1 0 19584 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_199
timestamp 1679581782
transform 1 0 20256 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_206
timestamp 1679581782
transform 1 0 20928 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_217
timestamp 1677579658
transform 1 0 21984 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_222
timestamp 1679581782
transform 1 0 22464 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_229
timestamp 1679581782
transform 1 0 23136 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_236
timestamp 1679581782
transform 1 0 23808 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_243
timestamp 1679581782
transform 1 0 24480 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_250
timestamp 1677580104
transform 1 0 25152 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_252
timestamp 1677579658
transform 1 0 25344 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_274
timestamp 1679581782
transform 1 0 27456 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_281
timestamp 1677580104
transform 1 0 28128 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_283
timestamp 1677579658
transform 1 0 28320 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_324
timestamp 1679581782
transform 1 0 32256 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_331
timestamp 1679581782
transform 1 0 32928 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_338
timestamp 1679581782
transform 1 0 33600 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_345
timestamp 1679581782
transform 1 0 34272 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_4  FILLER_7_352
timestamp 1679577901
transform 1 0 34944 0 -1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_356
timestamp 1677579658
transform 1 0 35328 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_361
timestamp 1679581782
transform 1 0 35808 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_368
timestamp 1679581782
transform 1 0 36480 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_375
timestamp 1679581782
transform 1 0 37152 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_382
timestamp 1677580104
transform 1 0 37824 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_393
timestamp 1677579658
transform 1 0 38880 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_4  FILLER_7_407
timestamp 1679577901
transform 1 0 40224 0 -1 7560
box -48 -56 432 834
use sg13g2_decap_8  FILLER_7_415
timestamp 1679581782
transform 1 0 40992 0 -1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_422
timestamp 1679581782
transform 1 0 41664 0 -1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_429
timestamp 1677580104
transform 1 0 42336 0 -1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_431
timestamp 1677579658
transform 1 0 42528 0 -1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_447
timestamp 1677579658
transform 1 0 44064 0 -1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_8
timestamp 1679581782
transform 1 0 1920 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_15
timestamp 1679581782
transform 1 0 2592 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_22
timestamp 1679581782
transform 1 0 3264 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_29
timestamp 1679581782
transform 1 0 3936 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_36
timestamp 1679581782
transform 1 0 4608 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_43
timestamp 1679581782
transform 1 0 5280 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_50
timestamp 1679581782
transform 1 0 5952 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_57
timestamp 1679581782
transform 1 0 6624 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_64
timestamp 1679581782
transform 1 0 7296 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_71
timestamp 1679581782
transform 1 0 7968 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_78
timestamp 1679581782
transform 1 0 8640 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_85
timestamp 1679581782
transform 1 0 9312 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_92
timestamp 1679581782
transform 1 0 9984 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_99
timestamp 1677580104
transform 1 0 10656 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_109
timestamp 1677579658
transform 1 0 11616 0 1 7560
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_131
timestamp 1677579658
transform 1 0 13728 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_185
timestamp 1679581782
transform 1 0 18912 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_213
timestamp 1679581782
transform 1 0 21600 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_220
timestamp 1679581782
transform 1 0 22272 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_227
timestamp 1679581782
transform 1 0 22944 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_234
timestamp 1679581782
transform 1 0 23616 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_241
timestamp 1679581782
transform 1 0 24288 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_248
timestamp 1679581782
transform 1 0 24960 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_255
timestamp 1677580104
transform 1 0 25632 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_257
timestamp 1677579658
transform 1 0 25824 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_262
timestamp 1679581782
transform 1 0 26304 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_269
timestamp 1679581782
transform 1 0 26976 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_276
timestamp 1679581782
transform 1 0 27648 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_283
timestamp 1677580104
transform 1 0 28320 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_307
timestamp 1679577901
transform 1 0 30624 0 1 7560
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_311
timestamp 1677580104
transform 1 0 31008 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_325
timestamp 1679581782
transform 1 0 32352 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_332
timestamp 1679581782
transform 1 0 33024 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_339
timestamp 1679581782
transform 1 0 33696 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_346
timestamp 1677580104
transform 1 0 34368 0 1 7560
box -48 -56 240 834
use sg13g2_decap_8  FILLER_8_360
timestamp 1679581782
transform 1 0 35712 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_367
timestamp 1679581782
transform 1 0 36384 0 1 7560
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_374
timestamp 1677579658
transform 1 0 37056 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_391
timestamp 1677580104
transform 1 0 38688 0 1 7560
box -48 -56 240 834
use sg13g2_decap_4  FILLER_8_397
timestamp 1679577901
transform 1 0 39264 0 1 7560
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_401
timestamp 1677579658
transform 1 0 39648 0 1 7560
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_410
timestamp 1679581782
transform 1 0 40512 0 1 7560
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_417
timestamp 1679581782
transform 1 0 41184 0 1 7560
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_424
timestamp 1677580104
transform 1 0 41856 0 1 7560
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_454
timestamp 1677579658
transform 1 0 44736 0 1 7560
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_16
timestamp 1677580104
transform 1 0 2688 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_26
timestamp 1679581782
transform 1 0 3648 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_33
timestamp 1679581782
transform 1 0 4320 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_40
timestamp 1679581782
transform 1 0 4992 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_47
timestamp 1679581782
transform 1 0 5664 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_54
timestamp 1679581782
transform 1 0 6336 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_61
timestamp 1679581782
transform 1 0 7008 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_68
timestamp 1679581782
transform 1 0 7680 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_75
timestamp 1679581782
transform 1 0 8352 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_82
timestamp 1679581782
transform 1 0 9024 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_89
timestamp 1677580104
transform 1 0 9696 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_91
timestamp 1677579658
transform 1 0 9888 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_148
timestamp 1677580104
transform 1 0 15360 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_162
timestamp 1677580104
transform 1 0 16704 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_164
timestamp 1677579658
transform 1 0 16896 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_169
timestamp 1677580104
transform 1 0 17376 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_179
timestamp 1677579658
transform 1 0 18336 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_212
timestamp 1677579658
transform 1 0 21504 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_221
timestamp 1679577901
transform 1 0 22368 0 -1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_9_237
timestamp 1679581782
transform 1 0 23904 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_244
timestamp 1679581782
transform 1 0 24576 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_267
timestamp 1679581782
transform 1 0 26784 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_274
timestamp 1679581782
transform 1 0 27456 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_281
timestamp 1679581782
transform 1 0 28128 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_288
timestamp 1677580104
transform 1 0 28800 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_290
timestamp 1677579658
transform 1 0 28992 0 -1 9072
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_295
timestamp 1677579658
transform 1 0 29472 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_300
timestamp 1679581782
transform 1 0 29952 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_307
timestamp 1679581782
transform 1 0 30624 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_314
timestamp 1679581782
transform 1 0 31296 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_321
timestamp 1677580104
transform 1 0 31968 0 -1 9072
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_351
timestamp 1677580104
transform 1 0 34848 0 -1 9072
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_361
timestamp 1679581782
transform 1 0 35808 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_368
timestamp 1679581782
transform 1 0 36480 0 -1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_375
timestamp 1679581782
transform 1 0 37152 0 -1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_382
timestamp 1677579658
transform 1 0 37824 0 -1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_24
timestamp 1679581782
transform 1 0 3456 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_31
timestamp 1679581782
transform 1 0 4128 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_38
timestamp 1679581782
transform 1 0 4800 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_45
timestamp 1679581782
transform 1 0 5472 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_52
timestamp 1679581782
transform 1 0 6144 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_59
timestamp 1679581782
transform 1 0 6816 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_66
timestamp 1679581782
transform 1 0 7488 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_73
timestamp 1679581782
transform 1 0 8160 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_80
timestamp 1679577901
transform 1 0 8832 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_84
timestamp 1677579658
transform 1 0 9216 0 1 9072
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_273
timestamp 1679581782
transform 1 0 27360 0 1 9072
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_280
timestamp 1677579658
transform 1 0 28032 0 1 9072
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_309
timestamp 1679577901
transform 1 0 30816 0 1 9072
box -48 -56 432 834
use sg13g2_decap_8  FILLER_10_369
timestamp 1679581782
transform 1 0 36576 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_376
timestamp 1679581782
transform 1 0 37248 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_383
timestamp 1679581782
transform 1 0 37920 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_390
timestamp 1679581782
transform 1 0 38592 0 1 9072
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_397
timestamp 1679581782
transform 1 0 39264 0 1 9072
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_404
timestamp 1679577901
transform 1 0 39936 0 1 9072
box -48 -56 432 834
use sg13g2_fill_1  FILLER_10_451
timestamp 1677579658
transform 1 0 44448 0 1 9072
box -48 -56 144 834
use sg13g2_buf_1  input1
timestamp 1676381911
transform 1 0 1440 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  input2
timestamp 1676381911
transform 1 0 1152 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input3
timestamp 1676381911
transform 1 0 1536 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  input4
timestamp 1676381911
transform 1 0 1152 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input5
timestamp 1676381911
transform 1 0 1536 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input6
timestamp 1676381911
transform 1 0 1920 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input7
timestamp 1676381911
transform 1 0 1152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input8
timestamp 1676381911
transform 1 0 2304 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input9
timestamp 1676381911
transform 1 0 3072 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input10
timestamp 1676381911
transform 1 0 1536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input11
timestamp 1676381911
transform 1 0 1920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input12
timestamp 1676381911
transform 1 0 2304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input13
timestamp 1676381911
transform 1 0 2688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input14
timestamp 1676381911
transform 1 0 20448 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input15
timestamp 1676381911
transform -1 0 21216 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input16
timestamp 1676381911
transform -1 0 21984 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input17
timestamp 1676381911
transform 1 0 21216 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input18
timestamp 1676381911
transform -1 0 23136 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input19
timestamp 1676381911
transform -1 0 23520 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input20
timestamp 1676381911
transform -1 0 23904 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input21
timestamp 1676381911
transform 1 0 23904 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input22
timestamp 1676381911
transform 1 0 24288 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input23
timestamp 1676381911
transform -1 0 25056 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input24
timestamp 1676381911
transform -1 0 25440 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input25
timestamp 1676381911
transform 1 0 25440 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input26
timestamp 1676381911
transform 1 0 21984 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input27
timestamp 1676381911
transform -1 0 21984 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input28
timestamp 1676381911
transform -1 0 22368 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input29
timestamp 1676381911
transform 1 0 22368 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input30
timestamp 1676381911
transform -1 0 26208 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input31
timestamp 1676381911
transform -1 0 25632 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input32
timestamp 1676381911
transform -1 0 26592 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input33
timestamp 1676381911
transform 1 0 25632 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input34
timestamp 1676381911
transform -1 0 26976 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input35
timestamp 1676381911
transform -1 0 26400 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input36
timestamp 1676381911
transform -1 0 27360 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input37
timestamp 1676381911
transform 1 0 26400 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input38
timestamp 1676381911
transform -1 0 28512 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input39
timestamp 1676381911
transform -1 0 28896 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input40
timestamp 1676381911
transform -1 0 29280 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input41
timestamp 1676381911
transform 1 0 29280 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input42
timestamp 1676381911
transform -1 0 30048 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input43
timestamp 1676381911
transform -1 0 29472 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  input44
timestamp 1676381911
transform -1 0 30432 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  input45
timestamp 1676381911
transform -1 0 30816 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output46
timestamp 1676381911
transform 1 0 44064 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output47
timestamp 1676381911
transform 1 0 44448 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output48
timestamp 1676381911
transform 1 0 44832 0 -1 4536
box -48 -56 432 834
use sg13g2_buf_1  output49
timestamp 1676381911
transform 1 0 44448 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output50
timestamp 1676381911
transform 1 0 44832 0 1 4536
box -48 -56 432 834
use sg13g2_buf_1  output51
timestamp 1676381911
transform 1 0 44448 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output52
timestamp 1676381911
transform 1 0 44832 0 -1 6048
box -48 -56 432 834
use sg13g2_buf_1  output53
timestamp 1676381911
transform 1 0 44448 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output54
timestamp 1676381911
transform 1 0 44832 0 1 6048
box -48 -56 432 834
use sg13g2_buf_1  output55
timestamp 1676381911
transform 1 0 44448 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output56
timestamp 1676381911
transform 1 0 44832 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output57
timestamp 1676381911
transform 1 0 43680 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output58
timestamp 1676381911
transform 1 0 44832 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output59
timestamp 1676381911
transform 1 0 44832 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output60
timestamp 1676381911
transform 1 0 44448 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output61
timestamp 1676381911
transform 1 0 44832 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output62
timestamp 1676381911
transform 1 0 44064 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output63
timestamp 1676381911
transform 1 0 41760 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output64
timestamp 1676381911
transform 1 0 44064 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output65
timestamp 1676381911
transform 1 0 43680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output66
timestamp 1676381911
transform 1 0 43296 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output67
timestamp 1676381911
transform 1 0 42912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output68
timestamp 1676381911
transform 1 0 43296 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output69
timestamp 1676381911
transform 1 0 42528 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output70
timestamp 1676381911
transform 1 0 42144 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output71
timestamp 1676381911
transform 1 0 44448 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output72
timestamp 1676381911
transform 1 0 44064 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output73
timestamp 1676381911
transform 1 0 44832 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output74
timestamp 1676381911
transform 1 0 44448 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output75
timestamp 1676381911
transform 1 0 44832 0 -1 3024
box -48 -56 432 834
use sg13g2_buf_1  output76
timestamp 1676381911
transform 1 0 44448 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output77
timestamp 1676381911
transform 1 0 44832 0 1 3024
box -48 -56 432 834
use sg13g2_buf_1  output78
timestamp 1676381911
transform -1 0 31968 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output79
timestamp 1676381911
transform -1 0 33696 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output80
timestamp 1676381911
transform -1 0 34656 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output81
timestamp 1676381911
transform -1 0 34080 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output82
timestamp 1676381911
transform -1 0 35040 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output83
timestamp 1676381911
transform -1 0 34464 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output84
timestamp 1676381911
transform -1 0 35424 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output85
timestamp 1676381911
transform -1 0 34848 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output86
timestamp 1676381911
transform -1 0 35808 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output87
timestamp 1676381911
transform -1 0 36192 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output88
timestamp 1676381911
transform -1 0 36576 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output89
timestamp 1676381911
transform -1 0 32352 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output90
timestamp 1676381911
transform -1 0 32736 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output91
timestamp 1676381911
transform -1 0 33120 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output92
timestamp 1676381911
transform -1 0 32544 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output93
timestamp 1676381911
transform -1 0 33504 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output94
timestamp 1676381911
transform -1 0 32928 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output95
timestamp 1676381911
transform -1 0 33888 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output96
timestamp 1676381911
transform -1 0 33312 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output97
timestamp 1676381911
transform -1 0 34272 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output98
timestamp 1676381911
transform -1 0 3552 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output99
timestamp 1676381911
transform -1 0 5280 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output100
timestamp 1676381911
transform -1 0 7008 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output101
timestamp 1676381911
transform -1 0 8736 0 1 1512
box -48 -56 432 834
use sg13g2_buf_1  output102
timestamp 1676381911
transform 1 0 9984 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output103
timestamp 1676381911
transform 1 0 9312 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output104
timestamp 1676381911
transform 1 0 10848 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output105
timestamp 1676381911
transform 1 0 10368 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output106
timestamp 1676381911
transform 1 0 9696 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output107
timestamp 1676381911
transform 1 0 10752 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output108
timestamp 1676381911
transform 1 0 10080 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output109
timestamp 1676381911
transform 1 0 11136 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output110
timestamp 1676381911
transform 1 0 10464 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output111
timestamp 1676381911
transform 1 0 11520 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output112
timestamp 1676381911
transform 1 0 10848 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output113
timestamp 1676381911
transform 1 0 11904 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output114
timestamp 1676381911
transform 1 0 11232 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output115
timestamp 1676381911
transform 1 0 12288 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output116
timestamp 1676381911
transform 1 0 11616 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output117
timestamp 1676381911
transform 1 0 12672 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output118
timestamp 1676381911
transform 1 0 12000 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output119
timestamp 1676381911
transform 1 0 13056 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output120
timestamp 1676381911
transform 1 0 13824 0 1 7560
box -48 -56 432 834
use sg13g2_buf_1  output121
timestamp 1676381911
transform 1 0 12384 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output122
timestamp 1676381911
transform 1 0 13440 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output123
timestamp 1676381911
transform 1 0 14688 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output124
timestamp 1676381911
transform 1 0 15552 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output125
timestamp 1676381911
transform 1 0 15072 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output126
timestamp 1676381911
transform 1 0 15456 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output127
timestamp 1676381911
transform 1 0 15840 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output128
timestamp 1676381911
transform 1 0 16224 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output129
timestamp 1676381911
transform 1 0 12768 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output130
timestamp 1676381911
transform 1 0 13824 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output131
timestamp 1676381911
transform -1 0 15840 0 -1 7560
box -48 -56 432 834
use sg13g2_buf_1  output132
timestamp 1676381911
transform 1 0 13152 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output133
timestamp 1676381911
transform 1 0 14208 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output134
timestamp 1676381911
transform 1 0 13536 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output135
timestamp 1676381911
transform 1 0 14592 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output136
timestamp 1676381911
transform 1 0 13920 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output137
timestamp 1676381911
transform 1 0 14304 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output138
timestamp 1676381911
transform 1 0 16608 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output139
timestamp 1676381911
transform 1 0 18912 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output140
timestamp 1676381911
transform -1 0 20352 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output141
timestamp 1676381911
transform 1 0 19296 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output142
timestamp 1676381911
transform -1 0 20736 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output143
timestamp 1676381911
transform 1 0 19680 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output144
timestamp 1676381911
transform -1 0 21120 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output145
timestamp 1676381911
transform 1 0 16992 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output146
timestamp 1676381911
transform 1 0 17376 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output147
timestamp 1676381911
transform -1 0 18816 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output148
timestamp 1676381911
transform 1 0 17760 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output149
timestamp 1676381911
transform -1 0 19200 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output150
timestamp 1676381911
transform 1 0 18144 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output151
timestamp 1676381911
transform -1 0 19584 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output152
timestamp 1676381911
transform 1 0 18528 0 1 9072
box -48 -56 432 834
use sg13g2_buf_1  output153
timestamp 1676381911
transform -1 0 19968 0 -1 9072
box -48 -56 432 834
use sg13g2_buf_1  output154
timestamp 1676381911
transform -1 0 31584 0 1 9072
box -48 -56 432 834
use sg13g2_tielo  S_CPU_IRQ_155
timestamp 1680000637
transform 1 0 20064 0 1 9072
box -48 -56 432 834
<< labels >>
flabel metal3 s 1400 0 1480 80 0 FreeSans 320 0 0 0 CONFIGURED_top
port 0 nsew signal input
flabel metal3 s 20984 11764 21064 11844 0 FreeSans 320 0 0 0 Co
port 1 nsew signal output
flabel metal2 s 0 548 90 628 0 FreeSans 320 0 0 0 FrameData[0]
port 2 nsew signal input
flabel metal2 s 0 3908 90 3988 0 FreeSans 320 0 0 0 FrameData[10]
port 3 nsew signal input
flabel metal2 s 0 4244 90 4324 0 FreeSans 320 0 0 0 FrameData[11]
port 4 nsew signal input
flabel metal2 s 0 4580 90 4660 0 FreeSans 320 0 0 0 FrameData[12]
port 5 nsew signal input
flabel metal2 s 0 4916 90 4996 0 FreeSans 320 0 0 0 FrameData[13]
port 6 nsew signal input
flabel metal2 s 0 5252 90 5332 0 FreeSans 320 0 0 0 FrameData[14]
port 7 nsew signal input
flabel metal2 s 0 5588 90 5668 0 FreeSans 320 0 0 0 FrameData[15]
port 8 nsew signal input
flabel metal2 s 0 5924 90 6004 0 FreeSans 320 0 0 0 FrameData[16]
port 9 nsew signal input
flabel metal2 s 0 6260 90 6340 0 FreeSans 320 0 0 0 FrameData[17]
port 10 nsew signal input
flabel metal2 s 0 6596 90 6676 0 FreeSans 320 0 0 0 FrameData[18]
port 11 nsew signal input
flabel metal2 s 0 6932 90 7012 0 FreeSans 320 0 0 0 FrameData[19]
port 12 nsew signal input
flabel metal2 s 0 884 90 964 0 FreeSans 320 0 0 0 FrameData[1]
port 13 nsew signal input
flabel metal2 s 0 7268 90 7348 0 FreeSans 320 0 0 0 FrameData[20]
port 14 nsew signal input
flabel metal2 s 0 7604 90 7684 0 FreeSans 320 0 0 0 FrameData[21]
port 15 nsew signal input
flabel metal2 s 0 7940 90 8020 0 FreeSans 320 0 0 0 FrameData[22]
port 16 nsew signal input
flabel metal2 s 0 8276 90 8356 0 FreeSans 320 0 0 0 FrameData[23]
port 17 nsew signal input
flabel metal2 s 0 8612 90 8692 0 FreeSans 320 0 0 0 FrameData[24]
port 18 nsew signal input
flabel metal2 s 0 8948 90 9028 0 FreeSans 320 0 0 0 FrameData[25]
port 19 nsew signal input
flabel metal2 s 0 9284 90 9364 0 FreeSans 320 0 0 0 FrameData[26]
port 20 nsew signal input
flabel metal2 s 0 9620 90 9700 0 FreeSans 320 0 0 0 FrameData[27]
port 21 nsew signal input
flabel metal2 s 0 9956 90 10036 0 FreeSans 320 0 0 0 FrameData[28]
port 22 nsew signal input
flabel metal2 s 0 10292 90 10372 0 FreeSans 320 0 0 0 FrameData[29]
port 23 nsew signal input
flabel metal2 s 0 1220 90 1300 0 FreeSans 320 0 0 0 FrameData[2]
port 24 nsew signal input
flabel metal2 s 0 10628 90 10708 0 FreeSans 320 0 0 0 FrameData[30]
port 25 nsew signal input
flabel metal2 s 0 10964 90 11044 0 FreeSans 320 0 0 0 FrameData[31]
port 26 nsew signal input
flabel metal2 s 0 1556 90 1636 0 FreeSans 320 0 0 0 FrameData[3]
port 27 nsew signal input
flabel metal2 s 0 1892 90 1972 0 FreeSans 320 0 0 0 FrameData[4]
port 28 nsew signal input
flabel metal2 s 0 2228 90 2308 0 FreeSans 320 0 0 0 FrameData[5]
port 29 nsew signal input
flabel metal2 s 0 2564 90 2644 0 FreeSans 320 0 0 0 FrameData[6]
port 30 nsew signal input
flabel metal2 s 0 2900 90 2980 0 FreeSans 320 0 0 0 FrameData[7]
port 31 nsew signal input
flabel metal2 s 0 3236 90 3316 0 FreeSans 320 0 0 0 FrameData[8]
port 32 nsew signal input
flabel metal2 s 0 3572 90 3652 0 FreeSans 320 0 0 0 FrameData[9]
port 33 nsew signal input
flabel metal2 s 46278 548 46368 628 0 FreeSans 320 0 0 0 FrameData_O[0]
port 34 nsew signal output
flabel metal2 s 46278 3908 46368 3988 0 FreeSans 320 0 0 0 FrameData_O[10]
port 35 nsew signal output
flabel metal2 s 46278 4244 46368 4324 0 FreeSans 320 0 0 0 FrameData_O[11]
port 36 nsew signal output
flabel metal2 s 46278 4580 46368 4660 0 FreeSans 320 0 0 0 FrameData_O[12]
port 37 nsew signal output
flabel metal2 s 46278 4916 46368 4996 0 FreeSans 320 0 0 0 FrameData_O[13]
port 38 nsew signal output
flabel metal2 s 46278 5252 46368 5332 0 FreeSans 320 0 0 0 FrameData_O[14]
port 39 nsew signal output
flabel metal2 s 46278 5588 46368 5668 0 FreeSans 320 0 0 0 FrameData_O[15]
port 40 nsew signal output
flabel metal2 s 46278 5924 46368 6004 0 FreeSans 320 0 0 0 FrameData_O[16]
port 41 nsew signal output
flabel metal2 s 46278 6260 46368 6340 0 FreeSans 320 0 0 0 FrameData_O[17]
port 42 nsew signal output
flabel metal2 s 46278 6596 46368 6676 0 FreeSans 320 0 0 0 FrameData_O[18]
port 43 nsew signal output
flabel metal2 s 46278 6932 46368 7012 0 FreeSans 320 0 0 0 FrameData_O[19]
port 44 nsew signal output
flabel metal2 s 46278 884 46368 964 0 FreeSans 320 0 0 0 FrameData_O[1]
port 45 nsew signal output
flabel metal2 s 46278 7268 46368 7348 0 FreeSans 320 0 0 0 FrameData_O[20]
port 46 nsew signal output
flabel metal2 s 46278 7604 46368 7684 0 FreeSans 320 0 0 0 FrameData_O[21]
port 47 nsew signal output
flabel metal2 s 46278 7940 46368 8020 0 FreeSans 320 0 0 0 FrameData_O[22]
port 48 nsew signal output
flabel metal2 s 46278 8276 46368 8356 0 FreeSans 320 0 0 0 FrameData_O[23]
port 49 nsew signal output
flabel metal2 s 46278 8612 46368 8692 0 FreeSans 320 0 0 0 FrameData_O[24]
port 50 nsew signal output
flabel metal2 s 46278 8948 46368 9028 0 FreeSans 320 0 0 0 FrameData_O[25]
port 51 nsew signal output
flabel metal2 s 46278 9284 46368 9364 0 FreeSans 320 0 0 0 FrameData_O[26]
port 52 nsew signal output
flabel metal2 s 46278 9620 46368 9700 0 FreeSans 320 0 0 0 FrameData_O[27]
port 53 nsew signal output
flabel metal2 s 46278 9956 46368 10036 0 FreeSans 320 0 0 0 FrameData_O[28]
port 54 nsew signal output
flabel metal2 s 46278 10292 46368 10372 0 FreeSans 320 0 0 0 FrameData_O[29]
port 55 nsew signal output
flabel metal2 s 46278 1220 46368 1300 0 FreeSans 320 0 0 0 FrameData_O[2]
port 56 nsew signal output
flabel metal2 s 46278 10628 46368 10708 0 FreeSans 320 0 0 0 FrameData_O[30]
port 57 nsew signal output
flabel metal2 s 46278 10964 46368 11044 0 FreeSans 320 0 0 0 FrameData_O[31]
port 58 nsew signal output
flabel metal2 s 46278 1556 46368 1636 0 FreeSans 320 0 0 0 FrameData_O[3]
port 59 nsew signal output
flabel metal2 s 46278 1892 46368 1972 0 FreeSans 320 0 0 0 FrameData_O[4]
port 60 nsew signal output
flabel metal2 s 46278 2228 46368 2308 0 FreeSans 320 0 0 0 FrameData_O[5]
port 61 nsew signal output
flabel metal2 s 46278 2564 46368 2644 0 FreeSans 320 0 0 0 FrameData_O[6]
port 62 nsew signal output
flabel metal2 s 46278 2900 46368 2980 0 FreeSans 320 0 0 0 FrameData_O[7]
port 63 nsew signal output
flabel metal2 s 46278 3236 46368 3316 0 FreeSans 320 0 0 0 FrameData_O[8]
port 64 nsew signal output
flabel metal2 s 46278 3572 46368 3652 0 FreeSans 320 0 0 0 FrameData_O[9]
port 65 nsew signal output
flabel metal3 s 11768 0 11848 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 66 nsew signal input
flabel metal3 s 29048 0 29128 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 67 nsew signal input
flabel metal3 s 30776 0 30856 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 68 nsew signal input
flabel metal3 s 32504 0 32584 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 69 nsew signal input
flabel metal3 s 34232 0 34312 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 70 nsew signal input
flabel metal3 s 35960 0 36040 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 71 nsew signal input
flabel metal3 s 37688 0 37768 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 72 nsew signal input
flabel metal3 s 39416 0 39496 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 73 nsew signal input
flabel metal3 s 41144 0 41224 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 74 nsew signal input
flabel metal3 s 42872 0 42952 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 75 nsew signal input
flabel metal3 s 44600 0 44680 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 76 nsew signal input
flabel metal3 s 13496 0 13576 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 77 nsew signal input
flabel metal3 s 15224 0 15304 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 78 nsew signal input
flabel metal3 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 79 nsew signal input
flabel metal3 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 80 nsew signal input
flabel metal3 s 20408 0 20488 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 81 nsew signal input
flabel metal3 s 22136 0 22216 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 82 nsew signal input
flabel metal3 s 23864 0 23944 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 83 nsew signal input
flabel metal3 s 25592 0 25672 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 84 nsew signal input
flabel metal3 s 27320 0 27400 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 85 nsew signal input
flabel metal3 s 31352 11764 31432 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 86 nsew signal output
flabel metal3 s 33272 11764 33352 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 87 nsew signal output
flabel metal3 s 33464 11764 33544 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 88 nsew signal output
flabel metal3 s 33656 11764 33736 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 89 nsew signal output
flabel metal3 s 33848 11764 33928 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 90 nsew signal output
flabel metal3 s 34040 11764 34120 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 91 nsew signal output
flabel metal3 s 34232 11764 34312 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 92 nsew signal output
flabel metal3 s 34424 11764 34504 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 93 nsew signal output
flabel metal3 s 34616 11764 34696 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 94 nsew signal output
flabel metal3 s 34808 11764 34888 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 95 nsew signal output
flabel metal3 s 35000 11764 35080 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 96 nsew signal output
flabel metal3 s 31544 11764 31624 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 97 nsew signal output
flabel metal3 s 31736 11764 31816 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 98 nsew signal output
flabel metal3 s 31928 11764 32008 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 99 nsew signal output
flabel metal3 s 32120 11764 32200 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 100 nsew signal output
flabel metal3 s 32312 11764 32392 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 101 nsew signal output
flabel metal3 s 32504 11764 32584 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 102 nsew signal output
flabel metal3 s 32696 11764 32776 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 103 nsew signal output
flabel metal3 s 32888 11764 32968 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 104 nsew signal output
flabel metal3 s 33080 11764 33160 11844 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 105 nsew signal output
flabel metal3 s 3128 0 3208 80 0 FreeSans 320 0 0 0 IRQ_top0
port 106 nsew signal output
flabel metal3 s 4856 0 4936 80 0 FreeSans 320 0 0 0 IRQ_top1
port 107 nsew signal output
flabel metal3 s 6584 0 6664 80 0 FreeSans 320 0 0 0 IRQ_top2
port 108 nsew signal output
flabel metal3 s 8312 0 8392 80 0 FreeSans 320 0 0 0 IRQ_top3
port 109 nsew signal output
flabel metal3 s 11000 11764 11080 11844 0 FreeSans 320 0 0 0 N1BEG[0]
port 110 nsew signal output
flabel metal3 s 11192 11764 11272 11844 0 FreeSans 320 0 0 0 N1BEG[1]
port 111 nsew signal output
flabel metal3 s 11384 11764 11464 11844 0 FreeSans 320 0 0 0 N1BEG[2]
port 112 nsew signal output
flabel metal3 s 11576 11764 11656 11844 0 FreeSans 320 0 0 0 N1BEG[3]
port 113 nsew signal output
flabel metal3 s 11768 11764 11848 11844 0 FreeSans 320 0 0 0 N2BEG[0]
port 114 nsew signal output
flabel metal3 s 11960 11764 12040 11844 0 FreeSans 320 0 0 0 N2BEG[1]
port 115 nsew signal output
flabel metal3 s 12152 11764 12232 11844 0 FreeSans 320 0 0 0 N2BEG[2]
port 116 nsew signal output
flabel metal3 s 12344 11764 12424 11844 0 FreeSans 320 0 0 0 N2BEG[3]
port 117 nsew signal output
flabel metal3 s 12536 11764 12616 11844 0 FreeSans 320 0 0 0 N2BEG[4]
port 118 nsew signal output
flabel metal3 s 12728 11764 12808 11844 0 FreeSans 320 0 0 0 N2BEG[5]
port 119 nsew signal output
flabel metal3 s 12920 11764 13000 11844 0 FreeSans 320 0 0 0 N2BEG[6]
port 120 nsew signal output
flabel metal3 s 13112 11764 13192 11844 0 FreeSans 320 0 0 0 N2BEG[7]
port 121 nsew signal output
flabel metal3 s 13304 11764 13384 11844 0 FreeSans 320 0 0 0 N2BEGb[0]
port 122 nsew signal output
flabel metal3 s 13496 11764 13576 11844 0 FreeSans 320 0 0 0 N2BEGb[1]
port 123 nsew signal output
flabel metal3 s 13688 11764 13768 11844 0 FreeSans 320 0 0 0 N2BEGb[2]
port 124 nsew signal output
flabel metal3 s 13880 11764 13960 11844 0 FreeSans 320 0 0 0 N2BEGb[3]
port 125 nsew signal output
flabel metal3 s 14072 11764 14152 11844 0 FreeSans 320 0 0 0 N2BEGb[4]
port 126 nsew signal output
flabel metal3 s 14264 11764 14344 11844 0 FreeSans 320 0 0 0 N2BEGb[5]
port 127 nsew signal output
flabel metal3 s 14456 11764 14536 11844 0 FreeSans 320 0 0 0 N2BEGb[6]
port 128 nsew signal output
flabel metal3 s 14648 11764 14728 11844 0 FreeSans 320 0 0 0 N2BEGb[7]
port 129 nsew signal output
flabel metal3 s 14840 11764 14920 11844 0 FreeSans 320 0 0 0 N4BEG[0]
port 130 nsew signal output
flabel metal3 s 16760 11764 16840 11844 0 FreeSans 320 0 0 0 N4BEG[10]
port 131 nsew signal output
flabel metal3 s 16952 11764 17032 11844 0 FreeSans 320 0 0 0 N4BEG[11]
port 132 nsew signal output
flabel metal3 s 17144 11764 17224 11844 0 FreeSans 320 0 0 0 N4BEG[12]
port 133 nsew signal output
flabel metal3 s 17336 11764 17416 11844 0 FreeSans 320 0 0 0 N4BEG[13]
port 134 nsew signal output
flabel metal3 s 17528 11764 17608 11844 0 FreeSans 320 0 0 0 N4BEG[14]
port 135 nsew signal output
flabel metal3 s 17720 11764 17800 11844 0 FreeSans 320 0 0 0 N4BEG[15]
port 136 nsew signal output
flabel metal3 s 15032 11764 15112 11844 0 FreeSans 320 0 0 0 N4BEG[1]
port 137 nsew signal output
flabel metal3 s 15224 11764 15304 11844 0 FreeSans 320 0 0 0 N4BEG[2]
port 138 nsew signal output
flabel metal3 s 15416 11764 15496 11844 0 FreeSans 320 0 0 0 N4BEG[3]
port 139 nsew signal output
flabel metal3 s 15608 11764 15688 11844 0 FreeSans 320 0 0 0 N4BEG[4]
port 140 nsew signal output
flabel metal3 s 15800 11764 15880 11844 0 FreeSans 320 0 0 0 N4BEG[5]
port 141 nsew signal output
flabel metal3 s 15992 11764 16072 11844 0 FreeSans 320 0 0 0 N4BEG[6]
port 142 nsew signal output
flabel metal3 s 16184 11764 16264 11844 0 FreeSans 320 0 0 0 N4BEG[7]
port 143 nsew signal output
flabel metal3 s 16376 11764 16456 11844 0 FreeSans 320 0 0 0 N4BEG[8]
port 144 nsew signal output
flabel metal3 s 16568 11764 16648 11844 0 FreeSans 320 0 0 0 N4BEG[9]
port 145 nsew signal output
flabel metal3 s 17912 11764 17992 11844 0 FreeSans 320 0 0 0 NN4BEG[0]
port 146 nsew signal output
flabel metal3 s 19832 11764 19912 11844 0 FreeSans 320 0 0 0 NN4BEG[10]
port 147 nsew signal output
flabel metal3 s 20024 11764 20104 11844 0 FreeSans 320 0 0 0 NN4BEG[11]
port 148 nsew signal output
flabel metal3 s 20216 11764 20296 11844 0 FreeSans 320 0 0 0 NN4BEG[12]
port 149 nsew signal output
flabel metal3 s 20408 11764 20488 11844 0 FreeSans 320 0 0 0 NN4BEG[13]
port 150 nsew signal output
flabel metal3 s 20600 11764 20680 11844 0 FreeSans 320 0 0 0 NN4BEG[14]
port 151 nsew signal output
flabel metal3 s 20792 11764 20872 11844 0 FreeSans 320 0 0 0 NN4BEG[15]
port 152 nsew signal output
flabel metal3 s 18104 11764 18184 11844 0 FreeSans 320 0 0 0 NN4BEG[1]
port 153 nsew signal output
flabel metal3 s 18296 11764 18376 11844 0 FreeSans 320 0 0 0 NN4BEG[2]
port 154 nsew signal output
flabel metal3 s 18488 11764 18568 11844 0 FreeSans 320 0 0 0 NN4BEG[3]
port 155 nsew signal output
flabel metal3 s 18680 11764 18760 11844 0 FreeSans 320 0 0 0 NN4BEG[4]
port 156 nsew signal output
flabel metal3 s 18872 11764 18952 11844 0 FreeSans 320 0 0 0 NN4BEG[5]
port 157 nsew signal output
flabel metal3 s 19064 11764 19144 11844 0 FreeSans 320 0 0 0 NN4BEG[6]
port 158 nsew signal output
flabel metal3 s 19256 11764 19336 11844 0 FreeSans 320 0 0 0 NN4BEG[7]
port 159 nsew signal output
flabel metal3 s 19448 11764 19528 11844 0 FreeSans 320 0 0 0 NN4BEG[8]
port 160 nsew signal output
flabel metal3 s 19640 11764 19720 11844 0 FreeSans 320 0 0 0 NN4BEG[9]
port 161 nsew signal output
flabel metal3 s 21176 11764 21256 11844 0 FreeSans 320 0 0 0 S1END[0]
port 162 nsew signal input
flabel metal3 s 21368 11764 21448 11844 0 FreeSans 320 0 0 0 S1END[1]
port 163 nsew signal input
flabel metal3 s 21560 11764 21640 11844 0 FreeSans 320 0 0 0 S1END[2]
port 164 nsew signal input
flabel metal3 s 21752 11764 21832 11844 0 FreeSans 320 0 0 0 S1END[3]
port 165 nsew signal input
flabel metal3 s 23480 11764 23560 11844 0 FreeSans 320 0 0 0 S2END[0]
port 166 nsew signal input
flabel metal3 s 23672 11764 23752 11844 0 FreeSans 320 0 0 0 S2END[1]
port 167 nsew signal input
flabel metal3 s 23864 11764 23944 11844 0 FreeSans 320 0 0 0 S2END[2]
port 168 nsew signal input
flabel metal3 s 24056 11764 24136 11844 0 FreeSans 320 0 0 0 S2END[3]
port 169 nsew signal input
flabel metal3 s 24248 11764 24328 11844 0 FreeSans 320 0 0 0 S2END[4]
port 170 nsew signal input
flabel metal3 s 24440 11764 24520 11844 0 FreeSans 320 0 0 0 S2END[5]
port 171 nsew signal input
flabel metal3 s 24632 11764 24712 11844 0 FreeSans 320 0 0 0 S2END[6]
port 172 nsew signal input
flabel metal3 s 24824 11764 24904 11844 0 FreeSans 320 0 0 0 S2END[7]
port 173 nsew signal input
flabel metal3 s 21944 11764 22024 11844 0 FreeSans 320 0 0 0 S2MID[0]
port 174 nsew signal input
flabel metal3 s 22136 11764 22216 11844 0 FreeSans 320 0 0 0 S2MID[1]
port 175 nsew signal input
flabel metal3 s 22328 11764 22408 11844 0 FreeSans 320 0 0 0 S2MID[2]
port 176 nsew signal input
flabel metal3 s 22520 11764 22600 11844 0 FreeSans 320 0 0 0 S2MID[3]
port 177 nsew signal input
flabel metal3 s 22712 11764 22792 11844 0 FreeSans 320 0 0 0 S2MID[4]
port 178 nsew signal input
flabel metal3 s 22904 11764 22984 11844 0 FreeSans 320 0 0 0 S2MID[5]
port 179 nsew signal input
flabel metal3 s 23096 11764 23176 11844 0 FreeSans 320 0 0 0 S2MID[6]
port 180 nsew signal input
flabel metal3 s 23288 11764 23368 11844 0 FreeSans 320 0 0 0 S2MID[7]
port 181 nsew signal input
flabel metal3 s 25016 11764 25096 11844 0 FreeSans 320 0 0 0 S4END[0]
port 182 nsew signal input
flabel metal3 s 26936 11764 27016 11844 0 FreeSans 320 0 0 0 S4END[10]
port 183 nsew signal input
flabel metal3 s 27128 11764 27208 11844 0 FreeSans 320 0 0 0 S4END[11]
port 184 nsew signal input
flabel metal3 s 27320 11764 27400 11844 0 FreeSans 320 0 0 0 S4END[12]
port 185 nsew signal input
flabel metal3 s 27512 11764 27592 11844 0 FreeSans 320 0 0 0 S4END[13]
port 186 nsew signal input
flabel metal3 s 27704 11764 27784 11844 0 FreeSans 320 0 0 0 S4END[14]
port 187 nsew signal input
flabel metal3 s 27896 11764 27976 11844 0 FreeSans 320 0 0 0 S4END[15]
port 188 nsew signal input
flabel metal3 s 25208 11764 25288 11844 0 FreeSans 320 0 0 0 S4END[1]
port 189 nsew signal input
flabel metal3 s 25400 11764 25480 11844 0 FreeSans 320 0 0 0 S4END[2]
port 190 nsew signal input
flabel metal3 s 25592 11764 25672 11844 0 FreeSans 320 0 0 0 S4END[3]
port 191 nsew signal input
flabel metal3 s 25784 11764 25864 11844 0 FreeSans 320 0 0 0 S4END[4]
port 192 nsew signal input
flabel metal3 s 25976 11764 26056 11844 0 FreeSans 320 0 0 0 S4END[5]
port 193 nsew signal input
flabel metal3 s 26168 11764 26248 11844 0 FreeSans 320 0 0 0 S4END[6]
port 194 nsew signal input
flabel metal3 s 26360 11764 26440 11844 0 FreeSans 320 0 0 0 S4END[7]
port 195 nsew signal input
flabel metal3 s 26552 11764 26632 11844 0 FreeSans 320 0 0 0 S4END[8]
port 196 nsew signal input
flabel metal3 s 26744 11764 26824 11844 0 FreeSans 320 0 0 0 S4END[9]
port 197 nsew signal input
flabel metal3 s 28088 11764 28168 11844 0 FreeSans 320 0 0 0 SS4END[0]
port 198 nsew signal input
flabel metal3 s 30008 11764 30088 11844 0 FreeSans 320 0 0 0 SS4END[10]
port 199 nsew signal input
flabel metal3 s 30200 11764 30280 11844 0 FreeSans 320 0 0 0 SS4END[11]
port 200 nsew signal input
flabel metal3 s 30392 11764 30472 11844 0 FreeSans 320 0 0 0 SS4END[12]
port 201 nsew signal input
flabel metal3 s 30584 11764 30664 11844 0 FreeSans 320 0 0 0 SS4END[13]
port 202 nsew signal input
flabel metal3 s 30776 11764 30856 11844 0 FreeSans 320 0 0 0 SS4END[14]
port 203 nsew signal input
flabel metal3 s 30968 11764 31048 11844 0 FreeSans 320 0 0 0 SS4END[15]
port 204 nsew signal input
flabel metal3 s 28280 11764 28360 11844 0 FreeSans 320 0 0 0 SS4END[1]
port 205 nsew signal input
flabel metal3 s 28472 11764 28552 11844 0 FreeSans 320 0 0 0 SS4END[2]
port 206 nsew signal input
flabel metal3 s 28664 11764 28744 11844 0 FreeSans 320 0 0 0 SS4END[3]
port 207 nsew signal input
flabel metal3 s 28856 11764 28936 11844 0 FreeSans 320 0 0 0 SS4END[4]
port 208 nsew signal input
flabel metal3 s 29048 11764 29128 11844 0 FreeSans 320 0 0 0 SS4END[5]
port 209 nsew signal input
flabel metal3 s 29240 11764 29320 11844 0 FreeSans 320 0 0 0 SS4END[6]
port 210 nsew signal input
flabel metal3 s 29432 11764 29512 11844 0 FreeSans 320 0 0 0 SS4END[7]
port 211 nsew signal input
flabel metal3 s 29624 11764 29704 11844 0 FreeSans 320 0 0 0 SS4END[8]
port 212 nsew signal input
flabel metal3 s 29816 11764 29896 11844 0 FreeSans 320 0 0 0 SS4END[9]
port 213 nsew signal input
flabel metal3 s 10040 0 10120 80 0 FreeSans 320 0 0 0 UserCLK
port 214 nsew signal input
flabel metal3 s 31160 11764 31240 11844 0 FreeSans 320 0 0 0 UserCLKo
port 215 nsew signal output
flabel metal5 s 4892 0 5332 11844 0 FreeSans 2560 90 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 4892 0 5332 40 0 FreeSans 320 0 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 4892 11804 5332 11844 0 FreeSans 320 0 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 20012 0 20452 11844 0 FreeSans 2560 90 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 20012 0 20452 40 0 FreeSans 320 0 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 20012 11804 20452 11844 0 FreeSans 320 0 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 35132 0 35572 11844 0 FreeSans 2560 90 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 35132 0 35572 40 0 FreeSans 320 0 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 35132 11804 35572 11844 0 FreeSans 320 0 0 0 VGND
port 216 nsew ground bidirectional
flabel metal5 s 3652 0 4092 11844 0 FreeSans 2560 90 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 3652 0 4092 40 0 FreeSans 320 0 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 3652 11804 4092 11844 0 FreeSans 320 0 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 18772 0 19212 11844 0 FreeSans 2560 90 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 18772 0 19212 40 0 FreeSans 320 0 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 18772 11804 19212 11844 0 FreeSans 320 0 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 33892 0 34332 11844 0 FreeSans 2560 90 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 33892 0 34332 40 0 FreeSans 320 0 0 0 VPWR
port 217 nsew power bidirectional
flabel metal5 s 33892 11804 34332 11844 0 FreeSans 320 0 0 0 VPWR
port 217 nsew power bidirectional
rlabel metal1 23184 9072 23184 9072 0 VGND
rlabel metal1 23184 9828 23184 9828 0 VPWR
rlabel metal3 1440 996 1440 996 0 CONFIGURED_top
rlabel metal3 42144 2016 42144 2016 0 FrameData[0]
rlabel metal2 752 3948 752 3948 0 FrameData[10]
rlabel metal2 752 4284 752 4284 0 FrameData[11]
rlabel metal3 38976 5418 38976 5418 0 FrameData[12]
rlabel metal2 21312 4914 21312 4914 0 FrameData[13]
rlabel metal2 752 5292 752 5292 0 FrameData[14]
rlabel metal2 704 5628 704 5628 0 FrameData[15]
rlabel metal4 34320 5880 34320 5880 0 FrameData[16]
rlabel metal2 35328 6300 35328 6300 0 FrameData[17]
rlabel metal2 464 6636 464 6636 0 FrameData[18]
rlabel metal2 416 6972 416 6972 0 FrameData[19]
rlabel metal3 42528 2184 42528 2184 0 FrameData[1]
rlabel metal2 656 7308 656 7308 0 FrameData[20]
rlabel metal2 464 7644 464 7644 0 FrameData[21]
rlabel metal2 368 7980 368 7980 0 FrameData[22]
rlabel metal2 848 8316 848 8316 0 FrameData[23]
rlabel metal2 320 8652 320 8652 0 FrameData[24]
rlabel metal2 656 8988 656 8988 0 FrameData[25]
rlabel metal2 128 9324 128 9324 0 FrameData[26]
rlabel metal2 512 9660 512 9660 0 FrameData[27]
rlabel metal2 272 9996 272 9996 0 FrameData[28]
rlabel metal2 560 10332 560 10332 0 FrameData[29]
rlabel metal2 42816 3444 42816 3444 0 FrameData[2]
rlabel metal2 608 10668 608 10668 0 FrameData[30]
rlabel metal2 752 11004 752 11004 0 FrameData[31]
rlabel metal3 41760 2520 41760 2520 0 FrameData[3]
rlabel metal2 128 1932 128 1932 0 FrameData[4]
rlabel metal3 42144 4074 42144 4074 0 FrameData[5]
rlabel metal2 35808 2982 35808 2982 0 FrameData[6]
rlabel metal2 752 2940 752 2940 0 FrameData[7]
rlabel metal2 128 3276 128 3276 0 FrameData[8]
rlabel metal2 656 3612 656 3612 0 FrameData[9]
rlabel metal2 45471 588 45471 588 0 FrameData_O[0]
rlabel metal2 45951 3948 45951 3948 0 FrameData_O[10]
rlabel metal2 45735 4284 45735 4284 0 FrameData_O[11]
rlabel metal2 45543 4620 45543 4620 0 FrameData_O[12]
rlabel metal2 45735 4956 45735 4956 0 FrameData_O[13]
rlabel via2 46287 5292 46287 5292 0 FrameData_O[14]
rlabel metal2 45735 5628 45735 5628 0 FrameData_O[15]
rlabel via2 46287 5964 46287 5964 0 FrameData_O[16]
rlabel metal2 45735 6300 45735 6300 0 FrameData_O[17]
rlabel via2 46287 6636 46287 6636 0 FrameData_O[18]
rlabel metal2 45735 6972 45735 6972 0 FrameData_O[19]
rlabel metal2 45951 924 45951 924 0 FrameData_O[1]
rlabel metal2 46095 7308 46095 7308 0 FrameData_O[20]
rlabel metal2 45999 7644 45999 7644 0 FrameData_O[21]
rlabel metal2 46047 7980 46047 7980 0 FrameData_O[22]
rlabel metal2 46095 8316 46095 8316 0 FrameData_O[23]
rlabel metal2 46239 8652 46239 8652 0 FrameData_O[24]
rlabel metal2 42624 9198 42624 9198 0 FrameData_O[25]
rlabel metal2 45351 9324 45351 9324 0 FrameData_O[26]
rlabel metal2 45159 9660 45159 9660 0 FrameData_O[27]
rlabel metal2 43752 9660 43752 9660 0 FrameData_O[28]
rlabel metal2 43272 9660 43272 9660 0 FrameData_O[29]
rlabel via2 46287 1260 46287 1260 0 FrameData_O[2]
rlabel metal2 42936 9660 42936 9660 0 FrameData_O[30]
rlabel metal3 44256 10164 44256 10164 0 FrameData_O[31]
rlabel metal2 45663 1596 45663 1596 0 FrameData_O[3]
rlabel metal2 45663 1932 45663 1932 0 FrameData_O[4]
rlabel metal2 45384 2100 45384 2100 0 FrameData_O[5]
rlabel metal2 46047 2604 46047 2604 0 FrameData_O[6]
rlabel metal2 45336 2856 45336 2856 0 FrameData_O[7]
rlabel metal2 45543 3276 45543 3276 0 FrameData_O[8]
rlabel metal2 45735 3612 45735 3612 0 FrameData_O[9]
rlabel metal2 20304 7140 20304 7140 0 FrameStrobe[0]
rlabel metal3 38016 3528 38016 3528 0 FrameStrobe[10]
rlabel metal4 36048 6300 36048 6300 0 FrameStrobe[11]
rlabel metal3 40416 7812 40416 7812 0 FrameStrobe[12]
rlabel metal3 34272 744 34272 744 0 FrameStrobe[13]
rlabel metal2 35616 7896 35616 7896 0 FrameStrobe[14]
rlabel metal2 36720 7140 36720 7140 0 FrameStrobe[15]
rlabel metal2 38832 7224 38832 7224 0 FrameStrobe[16]
rlabel metal2 38592 9156 38592 9156 0 FrameStrobe[17]
rlabel metal3 42912 1470 42912 1470 0 FrameStrobe[18]
rlabel metal3 44640 240 44640 240 0 FrameStrobe[19]
rlabel metal3 13536 114 13536 114 0 FrameStrobe[1]
rlabel metal3 15360 3108 15360 3108 0 FrameStrobe[2]
rlabel metal3 16992 2802 16992 2802 0 FrameStrobe[3]
rlabel metal3 18720 1500 18720 1500 0 FrameStrobe[4]
rlabel metal3 38496 3276 38496 3276 0 FrameStrobe[5]
rlabel metal3 22176 1122 22176 1122 0 FrameStrobe[6]
rlabel metal2 40896 4200 40896 4200 0 FrameStrobe[7]
rlabel metal3 25632 1080 25632 1080 0 FrameStrobe[8]
rlabel metal2 38592 4074 38592 4074 0 FrameStrobe[9]
rlabel metal2 31512 9576 31512 9576 0 FrameStrobe_O[0]
rlabel metal2 33336 8904 33336 8904 0 FrameStrobe_O[10]
rlabel metal2 34296 9240 34296 9240 0 FrameStrobe_O[11]
rlabel metal2 33720 8904 33720 8904 0 FrameStrobe_O[12]
rlabel metal2 34680 9492 34680 9492 0 FrameStrobe_O[13]
rlabel metal2 34248 8904 34248 8904 0 FrameStrobe_O[14]
rlabel metal2 34824 9324 34824 9324 0 FrameStrobe_O[15]
rlabel metal2 34488 8820 34488 8820 0 FrameStrobe_O[16]
rlabel metal2 35448 9660 35448 9660 0 FrameStrobe_O[17]
rlabel metal2 35352 9576 35352 9576 0 FrameStrobe_O[18]
rlabel metal2 36216 9660 36216 9660 0 FrameStrobe_O[19]
rlabel metal2 31800 9660 31800 9660 0 FrameStrobe_O[1]
rlabel metal2 32088 9576 32088 9576 0 FrameStrobe_O[2]
rlabel metal2 32568 9660 32568 9660 0 FrameStrobe_O[3]
rlabel metal2 32184 8904 32184 8904 0 FrameStrobe_O[4]
rlabel metal3 32352 10554 32352 10554 0 FrameStrobe_O[5]
rlabel metal2 32568 8904 32568 8904 0 FrameStrobe_O[6]
rlabel metal2 33528 9660 33528 9660 0 FrameStrobe_O[7]
rlabel metal2 32952 8904 32952 8904 0 FrameStrobe_O[8]
rlabel metal2 33576 9240 33576 9240 0 FrameStrobe_O[9]
rlabel metal3 3168 870 3168 870 0 IRQ_top0
rlabel metal3 4896 450 4896 450 0 IRQ_top1
rlabel metal3 6624 870 6624 870 0 IRQ_top2
rlabel metal3 8352 870 8352 870 0 IRQ_top3
rlabel metal2 20784 4200 20784 4200 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 25200 3360 25200 3360 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q
rlabel via2 23328 2688 23328 2688 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q
rlabel via2 13524 2688 13524 2688 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 13536 2772 13536 2772 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 14880 3444 14880 3444 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q
rlabel metal3 14688 7602 14688 7602 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 15840 7854 15840 7854 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q
rlabel metal3 18816 7560 18816 7560 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 29664 7350 29664 7350 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 30576 7224 30576 7224 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 29520 7896 29520 7896 0 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 10488 8904 10488 8904 0 N1BEG[0]
rlabel metal2 9960 9660 9960 9660 0 N1BEG[1]
rlabel metal2 11304 8148 11304 8148 0 N1BEG[2]
rlabel metal2 11016 8568 11016 8568 0 N1BEG[3]
rlabel metal2 10776 9576 10776 9576 0 N2BEG[0]
rlabel metal2 11544 8904 11544 8904 0 N2BEG[1]
rlabel metal2 10440 9492 10440 9492 0 N2BEG[2]
rlabel metal2 11784 8820 11784 8820 0 N2BEG[3]
rlabel metal2 11064 9240 11064 9240 0 N2BEG[4]
rlabel metal2 11880 8484 11880 8484 0 N2BEG[5]
rlabel metal3 13056 10752 13056 10752 0 N2BEG[6]
rlabel metal3 13152 10344 13152 10344 0 N2BEG[7]
rlabel metal3 13344 10722 13344 10722 0 N2BEGb[0]
rlabel metal2 12816 8904 12816 8904 0 N2BEGb[1]
rlabel metal3 13728 10554 13728 10554 0 N2BEGb[2]
rlabel metal2 13176 8820 13176 8820 0 N2BEGb[3]
rlabel metal3 14112 10470 14112 10470 0 N2BEGb[4]
rlabel metal2 13512 8568 13512 8568 0 N2BEGb[5]
rlabel metal2 14328 7812 14328 7812 0 N2BEGb[6]
rlabel metal3 14688 10764 14688 10764 0 N2BEGb[7]
rlabel metal2 13776 8694 13776 8694 0 N4BEG[0]
rlabel metal2 15048 9492 15048 9492 0 N4BEG[10]
rlabel metal2 16008 8904 16008 8904 0 N4BEG[11]
rlabel metal2 15528 9240 15528 9240 0 N4BEG[12]
rlabel metal2 16584 9240 16584 9240 0 N4BEG[13]
rlabel metal2 16248 9660 16248 9660 0 N4BEG[14]
rlabel metal2 17160 9324 17160 9324 0 N4BEG[15]
rlabel metal2 13320 9576 13320 9576 0 N4BEG[1]
rlabel metal2 14568 8904 14568 8904 0 N4BEG[2]
rlabel metal2 15480 7140 15480 7140 0 N4BEG[3]
rlabel metal2 13512 9492 13512 9492 0 N4BEG[4]
rlabel metal2 14568 8652 14568 8652 0 N4BEG[5]
rlabel metal2 13944 9660 13944 9660 0 N4BEG[6]
rlabel metal2 15432 8568 15432 8568 0 N4BEG[7]
rlabel metal2 14232 9324 14232 9324 0 N4BEG[8]
rlabel metal2 15528 9324 15528 9324 0 N4BEG[9]
rlabel metal2 16968 9492 16968 9492 0 NN4BEG[0]
rlabel metal2 19560 9576 19560 9576 0 NN4BEG[10]
rlabel metal2 19992 8904 19992 8904 0 NN4BEG[11]
rlabel metal2 19944 9660 19944 9660 0 NN4BEG[12]
rlabel metal2 20472 8904 20472 8904 0 NN4BEG[13]
rlabel metal2 20328 9324 20328 9324 0 NN4BEG[14]
rlabel metal2 20808 8904 20808 8904 0 NN4BEG[15]
rlabel metal2 17400 9660 17400 9660 0 NN4BEG[1]
rlabel metal2 18024 9660 18024 9660 0 NN4BEG[2]
rlabel metal2 18504 8904 18504 8904 0 NN4BEG[3]
rlabel metal2 18360 9576 18360 9576 0 NN4BEG[4]
rlabel metal2 18792 8904 18792 8904 0 NN4BEG[5]
rlabel metal2 18456 9660 18456 9660 0 NN4BEG[6]
rlabel metal2 19272 8904 19272 8904 0 NN4BEG[7]
rlabel metal2 19176 9660 19176 9660 0 NN4BEG[8]
rlabel metal2 19656 8904 19656 8904 0 NN4BEG[9]
rlabel metal3 21216 10722 21216 10722 0 S1END[0]
rlabel metal3 21408 10680 21408 10680 0 S1END[1]
rlabel metal3 21600 10218 21600 10218 0 S1END[2]
rlabel metal3 21792 10680 21792 10680 0 S1END[3]
rlabel metal2 23040 9534 23040 9534 0 S2END[0]
rlabel metal3 23712 10680 23712 10680 0 S2END[1]
rlabel metal3 23904 10680 23904 10680 0 S2END[2]
rlabel metal3 24096 10638 24096 10638 0 S2END[3]
rlabel metal3 24288 10638 24288 10638 0 S2END[4]
rlabel metal3 24480 10680 24480 10680 0 S2END[5]
rlabel metal3 24672 10680 24672 10680 0 S2END[6]
rlabel metal3 24864 10722 24864 10722 0 S2END[7]
rlabel metal3 21984 10260 21984 10260 0 S2MID[0]
rlabel metal3 22176 10680 22176 10680 0 S2MID[1]
rlabel metal3 22368 10680 22368 10680 0 S2MID[2]
rlabel metal3 22560 10638 22560 10638 0 S2MID[3]
rlabel metal3 22752 10722 22752 10722 0 S2MID[4]
rlabel metal3 22944 10890 22944 10890 0 S2MID[5]
rlabel metal3 17952 6636 17952 6636 0 S2MID[6]
rlabel metal3 8448 6720 8448 6720 0 S2MID[7]
rlabel metal3 25056 10596 25056 10596 0 S4END[0]
rlabel metal3 26976 10890 26976 10890 0 S4END[10]
rlabel metal2 41760 6552 41760 6552 0 S4END[11]
rlabel metal2 36672 8358 36672 8358 0 S4END[12]
rlabel metal3 35712 8358 35712 8358 0 S4END[13]
rlabel metal3 35040 6216 35040 6216 0 S4END[14]
rlabel metal3 42912 9366 42912 9366 0 S4END[15]
rlabel metal3 25248 10218 25248 10218 0 S4END[1]
rlabel metal3 25440 10764 25440 10764 0 S4END[2]
rlabel metal3 25632 10260 25632 10260 0 S4END[3]
rlabel metal3 25824 10764 25824 10764 0 S4END[4]
rlabel metal3 26016 10218 26016 10218 0 S4END[5]
rlabel metal3 26208 10596 26208 10596 0 S4END[6]
rlabel metal3 26400 10260 26400 10260 0 S4END[7]
rlabel metal2 23040 8694 23040 8694 0 S4END[8]
rlabel metal3 26784 10344 26784 10344 0 S4END[9]
rlabel metal3 28128 10638 28128 10638 0 SS4END[0]
rlabel metal3 35040 7770 35040 7770 0 SS4END[10]
rlabel metal3 38880 10248 38880 10248 0 SS4END[11]
rlabel metal3 37728 7938 37728 7938 0 SS4END[12]
rlabel metal3 38976 10080 38976 10080 0 SS4END[13]
rlabel metal2 36864 7854 36864 7854 0 SS4END[14]
rlabel metal3 42144 8106 42144 8106 0 SS4END[15]
rlabel metal3 28320 10680 28320 10680 0 SS4END[1]
rlabel metal3 28512 10722 28512 10722 0 SS4END[2]
rlabel metal3 28704 10596 28704 10596 0 SS4END[3]
rlabel metal3 28896 10764 28896 10764 0 SS4END[4]
rlabel metal3 29088 10218 29088 10218 0 SS4END[5]
rlabel metal3 29280 10680 29280 10680 0 SS4END[6]
rlabel metal3 29472 10806 29472 10806 0 SS4END[7]
rlabel metal3 43104 6930 43104 6930 0 SS4END[8]
rlabel metal2 35424 8526 35424 8526 0 SS4END[9]
rlabel metal3 40896 1764 40896 1764 0 UserCLK
rlabel metal2 31224 9660 31224 9660 0 UserCLKo
rlabel metal2 24096 3192 24096 3192 0 _000_
rlabel metal2 24768 4158 24768 4158 0 _001_
rlabel via1 24201 3360 24201 3360 0 _002_
rlabel metal3 24096 4032 24096 4032 0 _003_
rlabel metal2 24048 3612 24048 3612 0 _004_
rlabel metal3 22944 3528 22944 3528 0 _005_
rlabel metal2 23232 2562 23232 2562 0 _006_
rlabel metal3 23424 3444 23424 3444 0 _007_
rlabel metal2 24636 4200 24636 4200 0 _008_
rlabel metal2 14400 3192 14400 3192 0 _009_
rlabel metal2 15168 3360 15168 3360 0 _010_
rlabel metal2 13248 4242 13248 4242 0 _011_
rlabel via1 13151 4200 13151 4200 0 _012_
rlabel metal2 13728 4032 13728 4032 0 _013_
rlabel metal2 14517 3360 14517 3360 0 _014_
rlabel metal2 14304 2772 14304 2772 0 _015_
rlabel metal3 14976 3780 14976 3780 0 _016_
rlabel metal3 15456 3738 15456 3738 0 _017_
rlabel metal2 18528 7896 18528 7896 0 _018_
rlabel metal3 18624 8442 18624 8442 0 _019_
rlabel metal2 15264 7854 15264 7854 0 _020_
rlabel via1 15161 7896 15161 7896 0 _021_
rlabel metal2 16080 7938 16080 7938 0 _022_
rlabel metal2 16533 7224 16533 7224 0 _023_
rlabel metal2 16368 7140 16368 7140 0 _024_
rlabel metal2 16608 7392 16608 7392 0 _025_
rlabel metal3 16416 8274 16416 8274 0 _026_
rlabel metal2 30192 6384 30192 6384 0 _027_
rlabel metal2 30288 6636 30288 6636 0 _028_
rlabel metal2 29232 6972 29232 6972 0 _029_
rlabel metal2 28464 6972 28464 6972 0 _030_
rlabel metal2 29760 8064 29760 8064 0 _031_
rlabel metal3 29088 7602 29088 7602 0 _032_
rlabel metal3 29856 7560 29856 7560 0 _033_
rlabel metal2 29112 6468 29112 6468 0 _034_
rlabel metal2 28848 6216 28848 6216 0 _035_
rlabel metal3 15456 2616 15456 2616 0 net1
rlabel metal2 2760 8652 2760 8652 0 net10
rlabel metal2 8256 1974 8256 1974 0 net100
rlabel metal2 5184 2100 5184 2100 0 net101
rlabel metal2 17568 8484 17568 8484 0 net102
rlabel metal2 8640 1974 8640 1974 0 net103
rlabel metal3 29760 6174 29760 6174 0 net104
rlabel metal2 16968 8568 16968 8568 0 net105
rlabel metal2 12024 2772 12024 2772 0 net106
rlabel metal2 21240 3444 21240 3444 0 net107
rlabel metal2 4104 7140 4104 7140 0 net108
rlabel metal2 7272 6972 7272 6972 0 net109
rlabel metal3 11808 8568 11808 8568 0 net11
rlabel metal2 6696 8904 6696 8904 0 net110
rlabel metal3 11184 8652 11184 8652 0 net111
rlabel metal3 25872 8400 25872 8400 0 net112
rlabel metal2 11616 8610 11616 8610 0 net113
rlabel metal2 11256 3612 11256 3612 0 net114
rlabel metal2 20040 2436 20040 2436 0 net115
rlabel metal2 23040 7980 23040 7980 0 net116
rlabel metal2 17664 6930 17664 6930 0 net117
rlabel metal2 12840 2436 12840 2436 0 net118
rlabel metal3 20544 7518 20544 7518 0 net119
rlabel metal2 2376 9660 2376 9660 0 net12
rlabel metal3 28704 8190 28704 8190 0 net120
rlabel metal2 17448 7140 17448 7140 0 net121
rlabel metal2 13920 8022 13920 8022 0 net122
rlabel metal2 19656 3192 19656 3192 0 net123
rlabel metal2 42216 8652 42216 8652 0 net124
rlabel metal2 12984 4368 12984 4368 0 net125
rlabel metal2 19152 2688 19152 2688 0 net126
rlabel metal3 15168 9534 15168 9534 0 net127
rlabel metal2 15432 7056 15432 7056 0 net128
rlabel metal3 15936 9702 15936 9702 0 net129
rlabel metal2 3264 9282 3264 9282 0 net13
rlabel metal2 18528 9786 18528 9786 0 net130
rlabel metal2 34560 5754 34560 5754 0 net131
rlabel metal3 13920 8232 13920 8232 0 net132
rlabel metal3 15840 7350 15840 7350 0 net133
rlabel metal2 18240 6972 18240 6972 0 net134
rlabel metal3 14208 8862 14208 8862 0 net135
rlabel metal2 22944 8652 22944 8652 0 net136
rlabel metal2 14688 8694 14688 8694 0 net137
rlabel metal3 20928 8484 20928 8484 0 net138
rlabel metal2 14328 8148 14328 8148 0 net139
rlabel metal2 2712 9240 2712 9240 0 net14
rlabel metal3 16704 8778 16704 8778 0 net140
rlabel metal2 16440 2604 16440 2604 0 net141
rlabel metal2 21672 2772 21672 2772 0 net142
rlabel metal2 29400 6468 29400 6468 0 net143
rlabel metal2 20688 8652 20688 8652 0 net144
rlabel metal2 15240 3948 15240 3948 0 net145
rlabel metal2 21744 2520 21744 2520 0 net146
rlabel metal3 42240 7518 42240 7518 0 net147
rlabel metal3 17472 9450 17472 9450 0 net148
rlabel metal3 41760 7560 41760 7560 0 net149
rlabel metal2 16896 7560 16896 7560 0 net15
rlabel metal2 43416 8904 43416 8904 0 net150
rlabel metal3 43008 7686 43008 7686 0 net151
rlabel metal2 43272 8148 43272 8148 0 net152
rlabel metal3 19488 7602 19488 7602 0 net153
rlabel metal2 20832 8442 20832 8442 0 net154
rlabel metal2 19728 8652 19728 8652 0 net155
rlabel metal3 31872 6342 31872 6342 0 net156
rlabel metal3 21024 10512 21024 10512 0 net157
rlabel metal2 21120 9072 21120 9072 0 net16
rlabel metal4 15984 3780 15984 3780 0 net17
rlabel metal2 17280 8610 17280 8610 0 net18
rlabel metal2 21912 9660 21912 9660 0 net19
rlabel metal2 1728 7560 1728 7560 0 net2
rlabel metal3 22752 6300 22752 6300 0 net20
rlabel metal3 13824 2982 13824 2982 0 net21
rlabel metal2 17856 7140 17856 7140 0 net22
rlabel metal2 31824 7980 31824 7980 0 net23
rlabel metal2 25152 3486 25152 3486 0 net24
rlabel metal2 14160 2604 14160 2604 0 net25
rlabel metal3 17760 8526 17760 8526 0 net26
rlabel metal2 30960 7224 30960 7224 0 net27
rlabel metal2 22608 2604 22608 2604 0 net28
rlabel metal3 13536 3948 13536 3948 0 net29
rlabel metal2 17952 6636 17952 6636 0 net3
rlabel metal3 18240 8946 18240 8946 0 net30
rlabel metal3 31488 8988 31488 8988 0 net31
rlabel metal2 24432 4872 24432 4872 0 net32
rlabel metal3 24480 6972 24480 6972 0 net33
rlabel metal2 15456 8736 15456 8736 0 net34
rlabel metal3 29664 8736 29664 8736 0 net35
rlabel metal3 22992 9828 22992 9828 0 net36
rlabel metal3 13728 3780 13728 3780 0 net37
rlabel metal2 26760 9240 26760 9240 0 net38
rlabel metal2 27768 8652 27768 8652 0 net39
rlabel metal2 20832 4998 20832 4998 0 net4
rlabel metal2 27960 9240 27960 9240 0 net40
rlabel metal3 22752 3024 22752 3024 0 net41
rlabel metal2 28968 9576 28968 9576 0 net42
rlabel metal2 29832 9324 29832 9324 0 net43
rlabel metal2 28704 9324 28704 9324 0 net44
rlabel metal3 14496 2742 14496 2742 0 net45
rlabel metal3 16032 8694 16032 8694 0 net46
rlabel metal2 29712 9156 29712 9156 0 net47
rlabel metal2 43272 3528 43272 3528 0 net48
rlabel metal3 41088 6510 41088 6510 0 net49
rlabel metal2 16416 3402 16416 3402 0 net5
rlabel metal3 39072 7602 39072 7602 0 net50
rlabel metal3 41856 6090 41856 6090 0 net51
rlabel metal2 41664 7728 41664 7728 0 net52
rlabel metal3 41760 6258 41760 6258 0 net53
rlabel metal3 40224 6006 40224 6006 0 net54
rlabel metal2 37152 6174 37152 6174 0 net55
rlabel metal2 44640 6216 44640 6216 0 net56
rlabel metal2 36888 5628 36888 5628 0 net57
rlabel metal2 35976 4116 35976 4116 0 net58
rlabel metal2 43272 3276 43272 3276 0 net59
rlabel metal2 22440 6972 22440 6972 0 net6
rlabel metal2 17640 4284 17640 4284 0 net60
rlabel metal2 39456 3654 39456 3654 0 net61
rlabel metal2 22560 4746 22560 4746 0 net62
rlabel metal3 40704 6594 40704 6594 0 net63
rlabel metal2 42384 8736 42384 8736 0 net64
rlabel metal2 16200 3276 16200 3276 0 net65
rlabel metal2 11736 7728 11736 7728 0 net66
rlabel metal2 12504 7812 12504 7812 0 net67
rlabel metal2 25344 7518 25344 7518 0 net68
rlabel metal2 43008 9534 43008 9534 0 net69
rlabel metal2 1896 8820 1896 8820 0 net7
rlabel metal2 43272 3192 43272 3192 0 net70
rlabel metal2 36000 3864 36000 3864 0 net71
rlabel metal4 35424 6720 35424 6720 0 net72
rlabel metal2 44496 1932 44496 1932 0 net73
rlabel metal2 44160 2562 44160 2562 0 net74
rlabel metal2 43656 3948 43656 3948 0 net75
rlabel metal2 41856 3150 41856 3150 0 net76
rlabel metal2 44928 2688 44928 2688 0 net77
rlabel metal2 44544 3528 44544 3528 0 net78
rlabel metal2 44160 6426 44160 6426 0 net79
rlabel metal3 9408 6048 9408 6048 0 net8
rlabel metal2 23712 8736 23712 8736 0 net80
rlabel metal2 37128 3444 37128 3444 0 net81
rlabel metal2 40632 7140 40632 7140 0 net82
rlabel metal2 40152 7980 40152 7980 0 net83
rlabel metal2 34968 8148 34968 8148 0 net84
rlabel metal2 34776 8064 34776 8064 0 net85
rlabel metal2 35544 7056 35544 7056 0 net86
rlabel metal2 35352 8148 35352 8148 0 net87
rlabel metal2 35544 8820 35544 8820 0 net88
rlabel metal2 35784 8904 35784 8904 0 net89
rlabel metal2 1920 9156 1920 9156 0 net9
rlabel metal2 34920 6468 34920 6468 0 net90
rlabel metal2 40920 4032 40920 4032 0 net91
rlabel metal2 38712 3612 38712 3612 0 net92
rlabel metal2 42408 5628 42408 5628 0 net93
rlabel metal2 40152 4032 40152 4032 0 net94
rlabel metal2 35688 3192 35688 3192 0 net95
rlabel metal2 37080 2772 37080 2772 0 net96
rlabel metal2 40584 4032 40584 4032 0 net97
rlabel metal2 39048 2856 39048 2856 0 net98
rlabel metal2 37224 3948 37224 3948 0 net99
<< properties >>
string FIXED_BBOX 0 0 46368 11844
<< end >>
