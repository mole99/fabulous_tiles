magic
tech sky130A
magscale 1 2
timestamp 1740383537
<< viali >>
rect 5365 8585 5399 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 6837 8585 6871 8619
rect 7205 8585 7239 8619
rect 7481 8585 7515 8619
rect 7849 8585 7883 8619
rect 8309 8585 8343 8619
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11253 8585 11287 8619
rect 11989 8585 12023 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 13369 8585 13403 8619
rect 13737 8585 13771 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15209 8585 15243 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 16313 8585 16347 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 17785 8585 17819 8619
rect 18153 8585 18187 8619
rect 18521 8585 18555 8619
rect 18889 8585 18923 8619
rect 19717 8585 19751 8619
rect 34161 8585 34195 8619
rect 34897 8585 34931 8619
rect 35265 8585 35299 8619
rect 35633 8585 35667 8619
rect 36001 8585 36035 8619
rect 36369 8585 36403 8619
rect 37381 8585 37415 8619
rect 38577 8585 38611 8619
rect 40049 8585 40083 8619
rect 41797 8585 41831 8619
rect 42165 8585 42199 8619
rect 42717 8585 42751 8619
rect 5181 8449 5215 8483
rect 5549 8449 5583 8483
rect 5917 8449 5951 8483
rect 6653 8449 6687 8483
rect 7021 8449 7055 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8125 8449 8159 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11069 8449 11103 8483
rect 11805 8449 11839 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13553 8449 13587 8483
rect 13921 8449 13955 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 16129 8449 16163 8483
rect 16497 8449 16531 8483
rect 17233 8449 17267 8483
rect 17601 8449 17635 8483
rect 17969 8449 18003 8483
rect 18337 8449 18371 8483
rect 18705 8449 18739 8483
rect 19073 8449 19107 8483
rect 19533 8449 19567 8483
rect 19901 8449 19935 8483
rect 34345 8449 34379 8483
rect 34713 8449 34747 8483
rect 35081 8449 35115 8483
rect 35449 8449 35483 8483
rect 35817 8449 35851 8483
rect 36185 8449 36219 8483
rect 36553 8449 36587 8483
rect 37565 8449 37599 8483
rect 37657 8449 37691 8483
rect 38025 8449 38059 8483
rect 38393 8449 38427 8483
rect 38761 8449 38795 8483
rect 39129 8449 39163 8483
rect 39865 8449 39899 8483
rect 40233 8449 40267 8483
rect 41613 8449 41647 8483
rect 41981 8449 42015 8483
rect 42533 8449 42567 8483
rect 42901 8449 42935 8483
rect 43269 8449 43303 8483
rect 8585 8313 8619 8347
rect 20085 8313 20119 8347
rect 36737 8313 36771 8347
rect 37841 8313 37875 8347
rect 38209 8313 38243 8347
rect 38945 8313 38979 8347
rect 39313 8313 39347 8347
rect 40417 8313 40451 8347
rect 43085 8313 43119 8347
rect 43453 8313 43487 8347
rect 5917 8041 5951 8075
rect 6469 8041 6503 8075
rect 7021 8041 7055 8075
rect 8033 8041 8067 8075
rect 8585 8041 8619 8075
rect 9413 8041 9447 8075
rect 10241 8041 10275 8075
rect 11345 8041 11379 8075
rect 11989 8041 12023 8075
rect 12541 8041 12575 8075
rect 13185 8041 13219 8075
rect 13553 8041 13587 8075
rect 14197 8041 14231 8075
rect 14657 8041 14691 8075
rect 15393 8041 15427 8075
rect 15945 8041 15979 8075
rect 16589 8041 16623 8075
rect 17141 8041 17175 8075
rect 17417 8041 17451 8075
rect 17969 8041 18003 8075
rect 18429 8041 18463 8075
rect 20085 8041 20119 8075
rect 20729 8041 20763 8075
rect 22109 8041 22143 8075
rect 22477 8041 22511 8075
rect 23857 8041 23891 8075
rect 24225 8041 24259 8075
rect 26801 8041 26835 8075
rect 29009 8041 29043 8075
rect 36185 8041 36219 8075
rect 36553 8041 36587 8075
rect 36829 8041 36863 8075
rect 37657 8041 37691 8075
rect 38761 8041 38795 8075
rect 39129 8041 39163 8075
rect 39957 8041 39991 8075
rect 42349 8041 42383 8075
rect 42717 8041 42751 8075
rect 9873 7973 9907 8007
rect 15117 7973 15151 8007
rect 15761 7973 15795 8007
rect 26249 7973 26283 8007
rect 29101 7973 29135 8007
rect 28641 7905 28675 7939
rect 5733 7837 5767 7871
rect 6285 7837 6319 7871
rect 6837 7837 6871 7871
rect 8217 7837 8251 7871
rect 8769 7837 8803 7871
rect 9597 7837 9631 7871
rect 9689 7837 9723 7871
rect 10425 7837 10459 7871
rect 11529 7837 11563 7871
rect 11805 7837 11839 7871
rect 12357 7837 12391 7871
rect 12909 7837 12943 7871
rect 13369 7837 13403 7871
rect 13737 7837 13771 7871
rect 14381 7837 14415 7871
rect 14841 7837 14875 7871
rect 15025 7837 15059 7871
rect 15301 7837 15335 7871
rect 15577 7837 15611 7871
rect 15669 7837 15703 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 16773 7837 16807 7871
rect 17325 7837 17359 7871
rect 17601 7837 17635 7871
rect 18153 7837 18187 7871
rect 18245 7837 18279 7871
rect 20269 7837 20303 7871
rect 20821 7837 20855 7871
rect 20913 7837 20947 7871
rect 22109 7837 22143 7871
rect 22201 7837 22235 7871
rect 22661 7837 22695 7871
rect 23949 7837 23983 7871
rect 24041 7837 24075 7871
rect 24409 7837 24443 7871
rect 24685 7837 24719 7871
rect 26433 7837 26467 7871
rect 26985 7837 27019 7871
rect 27353 7837 27387 7871
rect 28825 7837 28859 7871
rect 29285 7837 29319 7871
rect 30205 7837 30239 7871
rect 36369 7837 36403 7871
rect 36737 7837 36771 7871
rect 37013 7837 37047 7871
rect 37473 7837 37507 7871
rect 38577 7837 38611 7871
rect 38945 7837 38979 7871
rect 39497 7837 39531 7871
rect 40141 7837 40175 7871
rect 42165 7837 42199 7871
rect 42533 7837 42567 7871
rect 42901 7837 42935 7871
rect 43269 7837 43303 7871
rect 13093 7701 13127 7735
rect 16221 7701 16255 7735
rect 21097 7701 21131 7735
rect 22385 7701 22419 7735
rect 24593 7701 24627 7735
rect 27169 7701 27203 7735
rect 30021 7701 30055 7735
rect 39313 7701 39347 7735
rect 43085 7701 43119 7735
rect 43453 7701 43487 7735
rect 4353 7497 4387 7531
rect 4629 7497 4663 7531
rect 5917 7497 5951 7531
rect 12633 7497 12667 7531
rect 15945 7497 15979 7531
rect 21833 7497 21867 7531
rect 38577 7497 38611 7531
rect 43085 7497 43119 7531
rect 4169 7361 4203 7395
rect 4445 7361 4479 7395
rect 5733 7361 5767 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 14933 7361 14967 7395
rect 15209 7361 15243 7395
rect 15853 7361 15887 7395
rect 16129 7361 16163 7395
rect 22017 7361 22051 7395
rect 24961 7361 24995 7395
rect 25053 7361 25087 7395
rect 30849 7361 30883 7395
rect 31401 7361 31435 7395
rect 32597 7361 32631 7395
rect 35357 7361 35391 7395
rect 38761 7361 38795 7395
rect 42901 7361 42935 7395
rect 43269 7361 43303 7395
rect 15025 7225 15059 7259
rect 24869 7225 24903 7259
rect 25237 7157 25271 7191
rect 30665 7157 30699 7191
rect 31217 7157 31251 7191
rect 32413 7157 32447 7191
rect 35173 7157 35207 7191
rect 43453 7157 43487 7191
rect 6285 6953 6319 6987
rect 7849 6953 7883 6987
rect 9597 6953 9631 6987
rect 13369 6953 13403 6987
rect 33057 6885 33091 6919
rect 26433 6817 26467 6851
rect 3893 6749 3927 6783
rect 4169 6749 4203 6783
rect 6101 6749 6135 6783
rect 6745 6749 6779 6783
rect 7205 6749 7239 6783
rect 8033 6749 8067 6783
rect 9781 6749 9815 6783
rect 13177 6749 13211 6783
rect 20085 6749 20119 6783
rect 22385 6749 22419 6783
rect 24409 6749 24443 6783
rect 24685 6749 24719 6783
rect 26525 6749 26559 6783
rect 26617 6749 26651 6783
rect 33241 6749 33275 6783
rect 34897 6749 34931 6783
rect 40877 6749 40911 6783
rect 42901 6749 42935 6783
rect 43269 6749 43303 6783
rect 4261 6681 4295 6715
rect 4077 6613 4111 6647
rect 6561 6613 6595 6647
rect 7021 6613 7055 6647
rect 19901 6613 19935 6647
rect 22201 6613 22235 6647
rect 24593 6613 24627 6647
rect 26801 6613 26835 6647
rect 34713 6613 34747 6647
rect 40693 6613 40727 6647
rect 43085 6613 43119 6647
rect 43453 6613 43487 6647
rect 7941 6409 7975 6443
rect 8953 6409 8987 6443
rect 9505 6409 9539 6443
rect 10701 6409 10735 6443
rect 11621 6409 11655 6443
rect 11989 6409 12023 6443
rect 15853 6409 15887 6443
rect 19257 6409 19291 6443
rect 36737 6409 36771 6443
rect 43453 6409 43487 6443
rect 7757 6273 7791 6307
rect 9137 6273 9171 6307
rect 9689 6273 9723 6307
rect 10149 6273 10183 6307
rect 10517 6273 10551 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 12817 6273 12851 6307
rect 16037 6273 16071 6307
rect 19441 6273 19475 6307
rect 36553 6273 36587 6307
rect 42901 6273 42935 6307
rect 43269 6273 43303 6307
rect 9965 6137 9999 6171
rect 12633 6069 12667 6103
rect 43085 6069 43119 6103
rect 4997 5865 5031 5899
rect 11161 5865 11195 5899
rect 18613 5865 18647 5899
rect 22201 5797 22235 5831
rect 39405 5797 39439 5831
rect 43453 5797 43487 5831
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 11345 5661 11379 5695
rect 18705 5661 18739 5695
rect 18797 5661 18831 5695
rect 21925 5661 21959 5695
rect 22017 5661 22051 5695
rect 26433 5661 26467 5695
rect 39589 5661 39623 5695
rect 42901 5661 42935 5695
rect 43269 5661 43303 5695
rect 18981 5525 19015 5559
rect 21833 5525 21867 5559
rect 26617 5525 26651 5559
rect 43085 5525 43119 5559
rect 10241 5321 10275 5355
rect 12909 5321 12943 5355
rect 29653 5321 29687 5355
rect 43453 5321 43487 5355
rect 10057 5185 10091 5219
rect 13093 5185 13127 5219
rect 20269 5185 20303 5219
rect 20453 5185 20487 5219
rect 24501 5185 24535 5219
rect 27077 5185 27111 5219
rect 29469 5185 29503 5219
rect 42901 5185 42935 5219
rect 43269 5185 43303 5219
rect 24685 5049 24719 5083
rect 27261 5049 27295 5083
rect 20637 4981 20671 5015
rect 43085 4981 43119 5015
rect 9137 4777 9171 4811
rect 32413 4777 32447 4811
rect 33701 4777 33735 4811
rect 36645 4777 36679 4811
rect 38761 4777 38795 4811
rect 31493 4709 31527 4743
rect 43453 4709 43487 4743
rect 8953 4573 8987 4607
rect 22569 4573 22603 4607
rect 22661 4573 22695 4607
rect 31309 4573 31343 4607
rect 32229 4573 32263 4607
rect 33517 4573 33551 4607
rect 36461 4573 36495 4607
rect 38577 4573 38611 4607
rect 42901 4573 42935 4607
rect 43269 4573 43303 4607
rect 22477 4505 22511 4539
rect 22845 4437 22879 4471
rect 43085 4437 43119 4471
rect 15577 4233 15611 4267
rect 15669 4165 15703 4199
rect 15853 4165 15887 4199
rect 21833 4097 21867 4131
rect 22109 4097 22143 4131
rect 22845 4097 22879 4131
rect 25697 4097 25731 4131
rect 35081 4097 35115 4131
rect 40877 4097 40911 4131
rect 42901 4097 42935 4131
rect 43269 4097 43303 4131
rect 16037 4029 16071 4063
rect 22017 3961 22051 3995
rect 23029 3961 23063 3995
rect 25881 3961 25915 3995
rect 35265 3961 35299 3995
rect 40693 3961 40727 3995
rect 43453 3961 43487 3995
rect 43085 3893 43119 3927
rect 17233 3689 17267 3723
rect 18521 3689 18555 3723
rect 34897 3689 34931 3723
rect 22937 3621 22971 3655
rect 43453 3621 43487 3655
rect 24869 3553 24903 3587
rect 17325 3485 17359 3519
rect 17417 3485 17451 3519
rect 18153 3485 18187 3519
rect 18337 3485 18371 3519
rect 23121 3485 23155 3519
rect 24961 3485 24995 3519
rect 25053 3485 25087 3519
rect 34713 3485 34747 3519
rect 42901 3485 42935 3519
rect 43269 3485 43303 3519
rect 17601 3349 17635 3383
rect 25237 3349 25271 3383
rect 43085 3349 43119 3383
rect 12449 3145 12483 3179
rect 23765 3145 23799 3179
rect 24133 3145 24167 3179
rect 31125 3145 31159 3179
rect 43453 3145 43487 3179
rect 12357 3077 12391 3111
rect 14013 3077 14047 3111
rect 16773 3077 16807 3111
rect 16957 3077 16991 3111
rect 9689 3009 9723 3043
rect 9873 3009 9907 3043
rect 11805 3009 11839 3043
rect 11989 3009 12023 3043
rect 14381 3009 14415 3043
rect 17049 3009 17083 3043
rect 17877 3009 17911 3043
rect 17969 3009 18003 3043
rect 19993 3009 20027 3043
rect 20361 3009 20395 3043
rect 20453 3009 20487 3043
rect 20729 3009 20763 3043
rect 21005 3009 21039 3043
rect 23857 3009 23891 3043
rect 23949 3009 23983 3043
rect 25145 3009 25179 3043
rect 25237 3009 25271 3043
rect 25329 3009 25363 3043
rect 27353 3009 27387 3043
rect 27445 3009 27479 3043
rect 27721 3009 27755 3043
rect 27905 3009 27939 3043
rect 28541 3009 28575 3043
rect 30941 3009 30975 3043
rect 42533 3009 42567 3043
rect 42901 3009 42935 3043
rect 43269 3009 43303 3043
rect 14565 2941 14599 2975
rect 11713 2873 11747 2907
rect 12173 2873 12207 2907
rect 14197 2873 14231 2907
rect 17785 2873 17819 2907
rect 20177 2873 20211 2907
rect 20913 2873 20947 2907
rect 18153 2805 18187 2839
rect 20637 2805 20671 2839
rect 25513 2805 25547 2839
rect 27261 2805 27295 2839
rect 27629 2805 27663 2839
rect 28089 2805 28123 2839
rect 28733 2805 28767 2839
rect 42717 2805 42751 2839
rect 43085 2805 43119 2839
rect 42165 2533 42199 2567
rect 43453 2533 43487 2567
rect 41969 2397 42003 2431
rect 42533 2397 42567 2431
rect 42901 2397 42935 2431
rect 43269 2397 43303 2431
rect 42717 2261 42751 2295
rect 43085 2261 43119 2295
<< metal1 >>
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 24946 11200 24952 11212
rect 7708 11172 24952 11200
rect 7708 11160 7714 11172
rect 24946 11160 24952 11172
rect 25004 11160 25010 11212
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 27982 11132 27988 11144
rect 11572 11104 27988 11132
rect 11572 11092 11578 11104
rect 27982 11092 27988 11104
rect 28040 11092 28046 11144
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 29638 11064 29644 11076
rect 14884 11036 29644 11064
rect 14884 11024 14890 11036
rect 29638 11024 29644 11036
rect 29696 11024 29702 11076
rect 19058 10956 19064 11008
rect 19116 10996 19122 11008
rect 29914 10996 29920 11008
rect 19116 10968 29920 10996
rect 19116 10956 19122 10968
rect 29914 10956 29920 10968
rect 29972 10956 29978 11008
rect 18782 10684 18788 10736
rect 18840 10724 18846 10736
rect 23842 10724 23848 10736
rect 18840 10696 23848 10724
rect 18840 10684 18846 10696
rect 23842 10684 23848 10696
rect 23900 10684 23906 10736
rect 17310 9664 17316 9716
rect 17368 9704 17374 9716
rect 24394 9704 24400 9716
rect 17368 9676 24400 9704
rect 17368 9664 17374 9676
rect 24394 9664 24400 9676
rect 24452 9664 24458 9716
rect 18414 9636 18420 9648
rect 12406 9608 18420 9636
rect 10962 9392 10968 9444
rect 11020 9432 11026 9444
rect 12406 9432 12434 9608
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 17126 9528 17132 9580
rect 17184 9568 17190 9580
rect 22738 9568 22744 9580
rect 17184 9540 22744 9568
rect 17184 9528 17190 9540
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 14642 9460 14648 9512
rect 14700 9500 14706 9512
rect 19794 9500 19800 9512
rect 14700 9472 19800 9500
rect 14700 9460 14706 9472
rect 19794 9460 19800 9472
rect 19852 9460 19858 9512
rect 19702 9432 19708 9444
rect 11020 9404 12434 9432
rect 16132 9404 19708 9432
rect 11020 9392 11026 9404
rect 16132 9364 16160 9404
rect 19702 9392 19708 9404
rect 19760 9392 19766 9444
rect 24210 9392 24216 9444
rect 24268 9432 24274 9444
rect 41690 9432 41696 9444
rect 24268 9404 41696 9432
rect 24268 9392 24274 9404
rect 41690 9392 41696 9404
rect 41748 9392 41754 9444
rect 12406 9336 16160 9364
rect 10778 9188 10784 9240
rect 10836 9228 10842 9240
rect 12406 9228 12434 9336
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 34422 9364 34428 9376
rect 16816 9336 34428 9364
rect 16816 9324 16822 9336
rect 34422 9324 34428 9336
rect 34480 9324 34486 9376
rect 19702 9256 19708 9308
rect 19760 9296 19766 9308
rect 20254 9296 20260 9308
rect 19760 9268 20260 9296
rect 19760 9256 19766 9268
rect 20254 9256 20260 9268
rect 20312 9256 20318 9308
rect 28718 9256 28724 9308
rect 28776 9296 28782 9308
rect 36170 9296 36176 9308
rect 28776 9268 36176 9296
rect 28776 9256 28782 9268
rect 36170 9256 36176 9268
rect 36228 9256 36234 9308
rect 10836 9200 12434 9228
rect 10836 9188 10842 9200
rect 17034 9188 17040 9240
rect 17092 9228 17098 9240
rect 32306 9228 32312 9240
rect 17092 9200 32312 9228
rect 17092 9188 17098 9200
rect 32306 9188 32312 9200
rect 32364 9188 32370 9240
rect 32582 9188 32588 9240
rect 32640 9228 32646 9240
rect 38010 9228 38016 9240
rect 32640 9200 38016 9228
rect 32640 9188 32646 9200
rect 38010 9188 38016 9200
rect 38068 9188 38074 9240
rect 24486 9120 24492 9172
rect 24544 9160 24550 9172
rect 30190 9160 30196 9172
rect 24544 9132 30196 9160
rect 24544 9120 24550 9132
rect 30190 9120 30196 9132
rect 30248 9120 30254 9172
rect 32766 9120 32772 9172
rect 32824 9160 32830 9172
rect 38378 9160 38384 9172
rect 32824 9132 38384 9160
rect 32824 9120 32830 9132
rect 38378 9120 38384 9132
rect 38436 9120 38442 9172
rect 18506 9052 18512 9104
rect 18564 9092 18570 9104
rect 24670 9092 24676 9104
rect 18564 9064 24676 9092
rect 18564 9052 18570 9064
rect 24670 9052 24676 9064
rect 24728 9052 24734 9104
rect 27706 9092 27712 9104
rect 25240 9064 27712 9092
rect 16574 9024 16580 9036
rect 12406 8996 16580 9024
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 12406 8820 12434 8996
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 18138 8984 18144 9036
rect 18196 9024 18202 9036
rect 25240 9024 25268 9064
rect 27706 9052 27712 9064
rect 27764 9052 27770 9104
rect 34606 9052 34612 9104
rect 34664 9092 34670 9104
rect 35250 9092 35256 9104
rect 34664 9064 35256 9092
rect 34664 9052 34670 9064
rect 35250 9052 35256 9064
rect 35308 9052 35314 9104
rect 35710 9052 35716 9104
rect 35768 9092 35774 9104
rect 36722 9092 36728 9104
rect 35768 9064 36728 9092
rect 35768 9052 35774 9064
rect 36722 9052 36728 9064
rect 36780 9052 36786 9104
rect 37918 9052 37924 9104
rect 37976 9092 37982 9104
rect 38562 9092 38568 9104
rect 37976 9064 38568 9092
rect 37976 9052 37982 9064
rect 38562 9052 38568 9064
rect 38620 9052 38626 9104
rect 18196 8996 25268 9024
rect 18196 8984 18202 8996
rect 25314 8984 25320 9036
rect 25372 9024 25378 9036
rect 41874 9024 41880 9036
rect 25372 8996 41880 9024
rect 25372 8984 25378 8996
rect 41874 8984 41880 8996
rect 41932 8984 41938 9036
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 22462 8956 22468 8968
rect 18288 8928 22468 8956
rect 18288 8916 18294 8928
rect 22462 8916 22468 8928
rect 22520 8916 22526 8968
rect 26602 8916 26608 8968
rect 26660 8956 26666 8968
rect 34698 8956 34704 8968
rect 26660 8928 34704 8956
rect 26660 8916 26666 8928
rect 34698 8916 34704 8928
rect 34756 8916 34762 8968
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 38838 8956 38844 8968
rect 34848 8928 38844 8956
rect 34848 8916 34854 8928
rect 38838 8916 38844 8928
rect 38896 8916 38902 8968
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 41598 8888 41604 8900
rect 29052 8860 41604 8888
rect 29052 8848 29058 8860
rect 41598 8848 41604 8860
rect 41656 8848 41662 8900
rect 10560 8792 12434 8820
rect 10560 8780 10566 8792
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 16666 8820 16672 8832
rect 16356 8792 16672 8820
rect 16356 8780 16362 8792
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 29270 8820 29276 8832
rect 17644 8792 29276 8820
rect 17644 8780 17650 8792
rect 29270 8780 29276 8792
rect 29328 8780 29334 8832
rect 35158 8780 35164 8832
rect 35216 8820 35222 8832
rect 35802 8820 35808 8832
rect 35216 8792 35808 8820
rect 35216 8780 35222 8792
rect 35802 8780 35808 8792
rect 35860 8780 35866 8832
rect 37826 8780 37832 8832
rect 37884 8820 37890 8832
rect 41966 8820 41972 8832
rect 37884 8792 41972 8820
rect 37884 8780 37890 8792
rect 41966 8780 41972 8792
rect 42024 8780 42030 8832
rect 1104 8730 43884 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 43884 8730
rect 1104 8656 43884 8678
rect 5350 8576 5356 8628
rect 5408 8576 5414 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5902 8616 5908 8628
rect 5767 8588 5908 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6454 8616 6460 8628
rect 6135 8588 6460 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 6825 8619 6883 8625
rect 6825 8585 6837 8619
rect 6871 8616 6883 8619
rect 7006 8616 7012 8628
rect 6871 8588 7012 8616
rect 6871 8585 6883 8588
rect 6825 8579 6883 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7282 8616 7288 8628
rect 7239 8588 7288 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7558 8616 7564 8628
rect 7515 8588 7564 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8110 8616 8116 8628
rect 7883 8588 8116 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8662 8616 8668 8628
rect 8343 8588 8668 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9490 8616 9496 8628
rect 9355 8588 9496 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9766 8616 9772 8628
rect 9723 8588 9772 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10318 8616 10324 8628
rect 10091 8588 10324 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10594 8616 10600 8628
rect 10459 8588 10600 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10870 8616 10876 8628
rect 10827 8588 10876 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11422 8616 11428 8628
rect 11287 8588 11428 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12526 8616 12532 8628
rect 12299 8588 12532 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 12802 8616 12808 8628
rect 12667 8588 12808 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13078 8616 13084 8628
rect 13035 8588 13084 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13630 8616 13636 8628
rect 13403 8588 13636 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 14182 8616 14188 8628
rect 13771 8588 14188 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14734 8616 14740 8628
rect 14507 8588 14740 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15838 8616 15844 8628
rect 15611 8588 15844 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16114 8616 16120 8628
rect 15979 8588 16120 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17218 8616 17224 8628
rect 17083 8588 17224 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 17405 8619 17463 8625
rect 17405 8585 17417 8619
rect 17451 8616 17463 8619
rect 17494 8616 17500 8628
rect 17451 8588 17500 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8616 17831 8619
rect 18046 8616 18052 8628
rect 17819 8588 18052 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18322 8616 18328 8628
rect 18187 8588 18328 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18509 8619 18567 8625
rect 18509 8585 18521 8619
rect 18555 8616 18567 8619
rect 18598 8616 18604 8628
rect 18555 8588 18604 8616
rect 18555 8585 18567 8588
rect 18509 8579 18567 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18874 8576 18880 8628
rect 18932 8576 18938 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 19484 8588 19717 8616
rect 19484 8576 19490 8588
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 19705 8579 19763 8585
rect 34054 8576 34060 8628
rect 34112 8616 34118 8628
rect 34149 8619 34207 8625
rect 34149 8616 34161 8619
rect 34112 8588 34161 8616
rect 34112 8576 34118 8588
rect 34149 8585 34161 8588
rect 34195 8585 34207 8619
rect 34149 8579 34207 8585
rect 34330 8576 34336 8628
rect 34388 8616 34394 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 34388 8588 34897 8616
rect 34388 8576 34394 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 34974 8576 34980 8628
rect 35032 8616 35038 8628
rect 35032 8588 35204 8616
rect 35032 8576 35038 8588
rect 13446 8548 13452 8560
rect 10244 8520 13452 8548
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 5552 8412 5580 8443
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 6546 8440 6552 8492
rect 6604 8480 6610 8492
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6604 8452 6653 8480
rect 6604 8440 6610 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7834 8480 7840 8492
rect 7699 8452 7840 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 4120 8384 5580 8412
rect 4120 8372 4126 8384
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 8036 8412 8064 8443
rect 7524 8384 8064 8412
rect 7524 8372 7530 8384
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 8128 8344 8156 8443
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10244 8489 10272 8520
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 16758 8548 16764 8560
rect 13924 8520 14964 8548
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 10597 8483 10655 8489
rect 10597 8480 10609 8483
rect 10560 8452 10609 8480
rect 10560 8440 10566 8452
rect 10597 8449 10609 8452
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 11072 8412 11100 8443
rect 10744 8384 11100 8412
rect 10744 8372 10750 8384
rect 7432 8316 8156 8344
rect 8573 8347 8631 8353
rect 7432 8304 7438 8316
rect 8573 8313 8585 8347
rect 8619 8344 8631 8347
rect 8846 8344 8852 8356
rect 8619 8316 8852 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 8846 8304 8852 8316
rect 8904 8304 8910 8356
rect 10318 8304 10324 8356
rect 10376 8344 10382 8356
rect 11808 8344 11836 8443
rect 12434 8440 12440 8492
rect 12492 8440 12498 8492
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13924 8489 13952 8520
rect 14936 8492 14964 8520
rect 15028 8520 15700 8548
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 10376 8316 11836 8344
rect 13188 8344 13216 8443
rect 13556 8412 13584 8443
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 14918 8440 14924 8492
rect 14976 8440 14982 8492
rect 15028 8489 15056 8520
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 15286 8412 15292 8424
rect 13556 8384 15292 8412
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 15672 8412 15700 8520
rect 15764 8520 16764 8548
rect 15764 8489 15792 8520
rect 16758 8508 16764 8520
rect 16816 8508 16822 8560
rect 18230 8548 18236 8560
rect 17144 8520 18236 8548
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 17034 8480 17040 8492
rect 16531 8452 17040 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17144 8412 17172 8520
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 18340 8520 24624 8548
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 15672 8384 17172 8412
rect 17236 8412 17264 8443
rect 17586 8440 17592 8492
rect 17644 8440 17650 8492
rect 18340 8489 18368 8520
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 17862 8412 17868 8424
rect 17236 8384 17868 8412
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 14918 8344 14924 8356
rect 13188 8316 14924 8344
rect 10376 8304 10382 8316
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 17402 8344 17408 8356
rect 15068 8316 17408 8344
rect 15068 8304 15074 8316
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 17678 8276 17684 8288
rect 13688 8248 17684 8276
rect 13688 8236 13694 8248
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 17972 8276 18000 8443
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 19076 8412 19104 8443
rect 19518 8440 19524 8492
rect 19576 8440 19582 8492
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19668 8452 19901 8480
rect 19668 8440 19674 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 24596 8480 24624 8520
rect 24670 8508 24676 8560
rect 24728 8548 24734 8560
rect 35176 8548 35204 8588
rect 35250 8576 35256 8628
rect 35308 8576 35314 8628
rect 35621 8619 35679 8625
rect 35621 8585 35633 8619
rect 35667 8585 35679 8619
rect 35621 8579 35679 8585
rect 35636 8548 35664 8579
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 35989 8619 36047 8625
rect 35989 8616 36001 8619
rect 35860 8588 36001 8616
rect 35860 8576 35866 8588
rect 35989 8585 36001 8588
rect 36035 8585 36047 8619
rect 35989 8579 36047 8585
rect 36357 8619 36415 8625
rect 36357 8585 36369 8619
rect 36403 8585 36415 8619
rect 36357 8579 36415 8585
rect 36372 8548 36400 8579
rect 36538 8576 36544 8628
rect 36596 8616 36602 8628
rect 37369 8619 37427 8625
rect 37369 8616 37381 8619
rect 36596 8588 37381 8616
rect 36596 8576 36602 8588
rect 37369 8585 37381 8588
rect 37415 8585 37427 8619
rect 37369 8579 37427 8585
rect 37642 8576 37648 8628
rect 37700 8616 37706 8628
rect 38565 8619 38623 8625
rect 38565 8616 38577 8619
rect 37700 8588 38577 8616
rect 37700 8576 37706 8588
rect 38565 8585 38577 8588
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 38930 8576 38936 8628
rect 38988 8616 38994 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 38988 8588 40049 8616
rect 38988 8576 38994 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 41782 8576 41788 8628
rect 41840 8576 41846 8628
rect 42150 8576 42156 8628
rect 42208 8576 42214 8628
rect 42702 8576 42708 8628
rect 42760 8576 42766 8628
rect 24728 8520 35112 8548
rect 35176 8520 35664 8548
rect 35728 8520 36400 8548
rect 24728 8508 24734 8520
rect 25866 8480 25872 8492
rect 20404 8452 22094 8480
rect 24596 8452 25872 8480
rect 20404 8440 20410 8452
rect 21818 8412 21824 8424
rect 19076 8384 21824 8412
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 19150 8304 19156 8356
rect 19208 8344 19214 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19208 8316 20085 8344
rect 19208 8304 19214 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 22066 8344 22094 8452
rect 25866 8440 25872 8452
rect 25924 8440 25930 8492
rect 32398 8440 32404 8492
rect 32456 8480 32462 8492
rect 34333 8483 34391 8489
rect 34333 8480 34345 8483
rect 32456 8452 34345 8480
rect 32456 8440 32462 8452
rect 34333 8449 34345 8452
rect 34379 8449 34391 8483
rect 34333 8443 34391 8449
rect 34698 8440 34704 8492
rect 34756 8440 34762 8492
rect 35084 8489 35112 8520
rect 35069 8483 35127 8489
rect 35069 8449 35081 8483
rect 35115 8449 35127 8483
rect 35069 8443 35127 8449
rect 35437 8483 35495 8489
rect 35437 8449 35449 8483
rect 35483 8449 35495 8483
rect 35437 8443 35495 8449
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 28626 8412 28632 8424
rect 23440 8384 28632 8412
rect 23440 8372 23446 8384
rect 28626 8372 28632 8384
rect 28684 8372 28690 8424
rect 33594 8372 33600 8424
rect 33652 8412 33658 8424
rect 35452 8412 35480 8443
rect 35526 8440 35532 8492
rect 35584 8480 35590 8492
rect 35728 8480 35756 8520
rect 36630 8508 36636 8560
rect 36688 8548 36694 8560
rect 36688 8520 39896 8548
rect 36688 8508 36694 8520
rect 35584 8452 35756 8480
rect 35805 8483 35863 8489
rect 35584 8440 35590 8452
rect 35805 8449 35817 8483
rect 35851 8449 35863 8483
rect 35805 8443 35863 8449
rect 33652 8384 35480 8412
rect 33652 8372 33658 8384
rect 26878 8344 26884 8356
rect 22066 8316 26884 8344
rect 20073 8307 20131 8313
rect 26878 8304 26884 8316
rect 26936 8304 26942 8356
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 35820 8344 35848 8443
rect 36170 8440 36176 8492
rect 36228 8440 36234 8492
rect 36541 8483 36599 8489
rect 36541 8449 36553 8483
rect 36587 8449 36599 8483
rect 36541 8443 36599 8449
rect 36556 8412 36584 8443
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37642 8440 37648 8492
rect 37700 8440 37706 8492
rect 38010 8440 38016 8492
rect 38068 8440 38074 8492
rect 38194 8440 38200 8492
rect 38252 8480 38258 8492
rect 38252 8452 38332 8480
rect 38252 8440 38258 8452
rect 27672 8316 35848 8344
rect 36280 8384 36584 8412
rect 27672 8304 27678 8316
rect 19242 8276 19248 8288
rect 17972 8248 19248 8276
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 22278 8236 22284 8288
rect 22336 8276 22342 8288
rect 25498 8276 25504 8288
rect 22336 8248 25504 8276
rect 22336 8236 22342 8248
rect 25498 8236 25504 8248
rect 25556 8236 25562 8288
rect 26418 8236 26424 8288
rect 26476 8276 26482 8288
rect 30466 8276 30472 8288
rect 26476 8248 30472 8276
rect 26476 8236 26482 8248
rect 30466 8236 30472 8248
rect 30524 8236 30530 8288
rect 31754 8236 31760 8288
rect 31812 8276 31818 8288
rect 32122 8276 32128 8288
rect 31812 8248 32128 8276
rect 31812 8236 31818 8248
rect 32122 8236 32128 8248
rect 32180 8236 32186 8288
rect 35802 8236 35808 8288
rect 35860 8276 35866 8288
rect 36280 8276 36308 8384
rect 37090 8372 37096 8424
rect 37148 8412 37154 8424
rect 38304 8412 38332 8452
rect 38378 8440 38384 8492
rect 38436 8440 38442 8492
rect 38654 8440 38660 8492
rect 38712 8480 38718 8492
rect 38749 8483 38807 8489
rect 38749 8480 38761 8483
rect 38712 8452 38761 8480
rect 38712 8440 38718 8452
rect 38749 8449 38761 8452
rect 38795 8449 38807 8483
rect 38749 8443 38807 8449
rect 38838 8440 38844 8492
rect 38896 8480 38902 8492
rect 39868 8489 39896 8520
rect 42058 8508 42064 8560
rect 42116 8548 42122 8560
rect 42116 8520 42932 8548
rect 42116 8508 42122 8520
rect 39117 8483 39175 8489
rect 39117 8480 39129 8483
rect 38896 8452 39129 8480
rect 38896 8440 38902 8452
rect 39117 8449 39129 8452
rect 39163 8449 39175 8483
rect 39117 8443 39175 8449
rect 39853 8483 39911 8489
rect 39853 8449 39865 8483
rect 39899 8449 39911 8483
rect 39853 8443 39911 8449
rect 39942 8440 39948 8492
rect 40000 8480 40006 8492
rect 40221 8483 40279 8489
rect 40221 8480 40233 8483
rect 40000 8452 40233 8480
rect 40000 8440 40006 8452
rect 40221 8449 40233 8452
rect 40267 8449 40279 8483
rect 40221 8443 40279 8449
rect 41598 8440 41604 8492
rect 41656 8440 41662 8492
rect 41690 8440 41696 8492
rect 41748 8480 41754 8492
rect 41969 8483 42027 8489
rect 41969 8480 41981 8483
rect 41748 8452 41981 8480
rect 41748 8440 41754 8452
rect 41969 8449 41981 8452
rect 42015 8449 42027 8483
rect 41969 8443 42027 8449
rect 42150 8440 42156 8492
rect 42208 8480 42214 8492
rect 42904 8489 42932 8520
rect 42521 8483 42579 8489
rect 42521 8480 42533 8483
rect 42208 8452 42533 8480
rect 42208 8440 42214 8452
rect 42521 8449 42533 8452
rect 42567 8449 42579 8483
rect 42521 8443 42579 8449
rect 42889 8483 42947 8489
rect 42889 8449 42901 8483
rect 42935 8449 42947 8483
rect 42889 8443 42947 8449
rect 43257 8483 43315 8489
rect 43257 8449 43269 8483
rect 43303 8449 43315 8483
rect 43257 8443 43315 8449
rect 37148 8384 38240 8412
rect 38304 8384 39344 8412
rect 37148 8372 37154 8384
rect 36722 8304 36728 8356
rect 36780 8304 36786 8356
rect 36814 8304 36820 8356
rect 36872 8344 36878 8356
rect 38212 8353 38240 8384
rect 37829 8347 37887 8353
rect 37829 8344 37841 8347
rect 36872 8316 37841 8344
rect 36872 8304 36878 8316
rect 37829 8313 37841 8316
rect 37875 8313 37887 8347
rect 37829 8307 37887 8313
rect 38197 8347 38255 8353
rect 38197 8313 38209 8347
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 38562 8304 38568 8356
rect 38620 8344 38626 8356
rect 39316 8353 39344 8384
rect 40310 8372 40316 8424
rect 40368 8412 40374 8424
rect 43272 8412 43300 8443
rect 40368 8384 43300 8412
rect 40368 8372 40374 8384
rect 38933 8347 38991 8353
rect 38933 8344 38945 8347
rect 38620 8316 38945 8344
rect 38620 8304 38626 8316
rect 38933 8313 38945 8316
rect 38979 8313 38991 8347
rect 38933 8307 38991 8313
rect 39301 8347 39359 8353
rect 39301 8313 39313 8347
rect 39347 8313 39359 8347
rect 39301 8307 39359 8313
rect 39390 8304 39396 8356
rect 39448 8344 39454 8356
rect 40405 8347 40463 8353
rect 40405 8344 40417 8347
rect 39448 8316 40417 8344
rect 39448 8304 39454 8316
rect 40405 8313 40417 8316
rect 40451 8313 40463 8347
rect 40405 8307 40463 8313
rect 43070 8304 43076 8356
rect 43128 8304 43134 8356
rect 43438 8304 43444 8356
rect 43496 8304 43502 8356
rect 35860 8248 36308 8276
rect 35860 8236 35866 8248
rect 1104 8186 43884 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 43884 8186
rect 1104 8112 43884 8134
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5684 8044 5917 8072
rect 5684 8032 5690 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 5905 8035 5963 8041
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 6236 8044 6469 8072
rect 6236 8032 6242 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7009 8075 7067 8081
rect 7009 8072 7021 8075
rect 6788 8044 7021 8072
rect 6788 8032 6794 8044
rect 7009 8041 7021 8044
rect 7055 8041 7067 8075
rect 7009 8035 7067 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7800 8044 8033 8072
rect 7800 8032 7806 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8444 8044 8585 8072
rect 8444 8032 8450 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 9398 8032 9404 8084
rect 9456 8032 9462 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10229 8075 10287 8081
rect 10229 8072 10241 8075
rect 10100 8044 10241 8072
rect 10100 8032 10106 8044
rect 10229 8041 10241 8044
rect 10275 8041 10287 8075
rect 10229 8035 10287 8041
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 11204 8044 11345 8072
rect 11204 8032 11210 8044
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11756 8044 11989 8072
rect 11756 8032 11762 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12308 8044 12541 8072
rect 12308 8032 12314 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 12529 8035 12587 8041
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 12860 8044 13185 8072
rect 12860 8032 12866 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 13173 8035 13231 8041
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13412 8044 13553 8072
rect 13412 8032 13418 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13872 8044 14197 8072
rect 13872 8032 13878 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14516 8044 14657 8072
rect 14516 8032 14522 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 15381 8075 15439 8081
rect 15381 8072 15393 8075
rect 15344 8044 15393 8072
rect 15344 8032 15350 8044
rect 15381 8041 15393 8044
rect 15427 8041 15439 8075
rect 15381 8035 15439 8041
rect 15562 8032 15568 8084
rect 15620 8072 15626 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15620 8044 15945 8072
rect 15620 8032 15626 8044
rect 15933 8041 15945 8044
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 16577 8075 16635 8081
rect 16577 8072 16589 8075
rect 16448 8044 16589 8072
rect 16448 8032 16454 8044
rect 16577 8041 16589 8044
rect 16623 8041 16635 8075
rect 16577 8035 16635 8041
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 17000 8044 17141 8072
rect 17000 8032 17006 8044
rect 17129 8041 17141 8044
rect 17175 8041 17187 8075
rect 17129 8035 17187 8041
rect 17402 8032 17408 8084
rect 17460 8032 17466 8084
rect 17770 8032 17776 8084
rect 17828 8072 17834 8084
rect 17957 8075 18015 8081
rect 17957 8072 17969 8075
rect 17828 8044 17969 8072
rect 17828 8032 17834 8044
rect 17957 8041 17969 8044
rect 18003 8041 18015 8075
rect 17957 8035 18015 8041
rect 18417 8075 18475 8081
rect 18417 8041 18429 8075
rect 18463 8072 18475 8075
rect 19610 8072 19616 8084
rect 18463 8044 19616 8072
rect 18463 8041 18475 8044
rect 18417 8035 18475 8041
rect 19610 8032 19616 8044
rect 19668 8032 19674 8084
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 20073 8075 20131 8081
rect 20073 8072 20085 8075
rect 19852 8044 20085 8072
rect 19852 8032 19858 8044
rect 20073 8041 20085 8044
rect 20119 8041 20131 8075
rect 20073 8035 20131 8041
rect 20714 8032 20720 8084
rect 20772 8032 20778 8084
rect 22094 8032 22100 8084
rect 22152 8032 22158 8084
rect 22462 8032 22468 8084
rect 22520 8032 22526 8084
rect 23842 8032 23848 8084
rect 23900 8032 23906 8084
rect 24210 8032 24216 8084
rect 24268 8032 24274 8084
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 26789 8075 26847 8081
rect 26789 8072 26801 8075
rect 25924 8044 26801 8072
rect 25924 8032 25930 8044
rect 26789 8041 26801 8044
rect 26835 8041 26847 8075
rect 26789 8035 26847 8041
rect 28994 8032 29000 8084
rect 29052 8032 29058 8084
rect 29178 8032 29184 8084
rect 29236 8072 29242 8084
rect 30742 8072 30748 8084
rect 29236 8044 30748 8072
rect 29236 8032 29242 8044
rect 30742 8032 30748 8044
rect 30800 8032 30806 8084
rect 35986 8032 35992 8084
rect 36044 8072 36050 8084
rect 36173 8075 36231 8081
rect 36173 8072 36185 8075
rect 36044 8044 36185 8072
rect 36044 8032 36050 8044
rect 36173 8041 36185 8044
rect 36219 8041 36231 8075
rect 36173 8035 36231 8041
rect 36262 8032 36268 8084
rect 36320 8072 36326 8084
rect 36541 8075 36599 8081
rect 36541 8072 36553 8075
rect 36320 8044 36553 8072
rect 36320 8032 36326 8044
rect 36541 8041 36553 8044
rect 36587 8041 36599 8075
rect 36541 8035 36599 8041
rect 36814 8032 36820 8084
rect 36872 8032 36878 8084
rect 37366 8032 37372 8084
rect 37424 8072 37430 8084
rect 37645 8075 37703 8081
rect 37645 8072 37657 8075
rect 37424 8044 37657 8072
rect 37424 8032 37430 8044
rect 37645 8041 37657 8044
rect 37691 8041 37703 8075
rect 37645 8035 37703 8041
rect 38470 8032 38476 8084
rect 38528 8072 38534 8084
rect 38749 8075 38807 8081
rect 38749 8072 38761 8075
rect 38528 8044 38761 8072
rect 38528 8032 38534 8044
rect 38749 8041 38761 8044
rect 38795 8041 38807 8075
rect 38749 8035 38807 8041
rect 38838 8032 38844 8084
rect 38896 8072 38902 8084
rect 39117 8075 39175 8081
rect 39117 8072 39129 8075
rect 38896 8044 39129 8072
rect 38896 8032 38902 8044
rect 39117 8041 39129 8044
rect 39163 8041 39175 8075
rect 39117 8035 39175 8041
rect 39574 8032 39580 8084
rect 39632 8072 39638 8084
rect 39945 8075 40003 8081
rect 39945 8072 39957 8075
rect 39632 8044 39957 8072
rect 39632 8032 39638 8044
rect 39945 8041 39957 8044
rect 39991 8041 40003 8075
rect 39945 8035 40003 8041
rect 42334 8032 42340 8084
rect 42392 8032 42398 8084
rect 42610 8032 42616 8084
rect 42668 8072 42674 8084
rect 42705 8075 42763 8081
rect 42705 8072 42717 8075
rect 42668 8044 42717 8072
rect 42668 8032 42674 8044
rect 42705 8041 42717 8044
rect 42751 8041 42763 8075
rect 42705 8035 42763 8041
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 9950 8004 9956 8016
rect 9907 7976 9956 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 9950 7964 9956 7976
rect 10008 7964 10014 8016
rect 14826 8004 14832 8016
rect 12912 7976 14832 8004
rect 9398 7896 9404 7948
rect 9456 7936 9462 7948
rect 9456 7908 11836 7936
rect 9456 7896 9462 7908
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 4396 7840 5733 7868
rect 4396 7828 4402 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7868 8263 7871
rect 8662 7868 8668 7880
rect 8251 7840 8668 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8846 7868 8852 7880
rect 8803 7840 8852 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9766 7868 9772 7880
rect 9723 7840 9772 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 11808 7877 11836 7908
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 10428 7732 10456 7831
rect 11532 7800 11560 7831
rect 12342 7828 12348 7880
rect 12400 7828 12406 7880
rect 12912 7877 12940 7976
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 15105 8007 15163 8013
rect 15105 7973 15117 8007
rect 15151 7973 15163 8007
rect 15105 7967 15163 7973
rect 15120 7936 15148 7967
rect 15746 7964 15752 8016
rect 15804 7964 15810 8016
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 26237 8007 26295 8013
rect 26237 8004 26249 8007
rect 18748 7976 26249 8004
rect 18748 7964 18754 7976
rect 26237 7973 26249 7976
rect 26283 7973 26295 8007
rect 26237 7967 26295 7973
rect 29089 8007 29147 8013
rect 29089 7973 29101 8007
rect 29135 7973 29147 8007
rect 29089 7967 29147 7973
rect 22554 7936 22560 7948
rect 13740 7908 15148 7936
rect 15304 7908 16620 7936
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13630 7868 13636 7880
rect 13403 7840 13636 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 13740 7877 13768 7908
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 14366 7828 14372 7880
rect 14424 7828 14430 7880
rect 15304 7877 15332 7908
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15059 7840 15301 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7868 15623 7871
rect 15657 7871 15715 7877
rect 15657 7868 15669 7871
rect 15611 7840 15669 7868
rect 15611 7837 15623 7840
rect 15565 7831 15623 7837
rect 15657 7837 15669 7840
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16298 7868 16304 7880
rect 16163 7840 16304 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 13538 7800 13544 7812
rect 11532 7772 13544 7800
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 14844 7800 14872 7831
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7868 16451 7871
rect 16482 7868 16488 7880
rect 16439 7840 16488 7868
rect 16439 7837 16451 7840
rect 16393 7831 16451 7837
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 14844 7772 16252 7800
rect 12894 7732 12900 7744
rect 10428 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13078 7692 13084 7744
rect 13136 7692 13142 7744
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15378 7732 15384 7744
rect 15252 7704 15384 7732
rect 15252 7692 15258 7704
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 16224 7741 16252 7772
rect 16209 7735 16267 7741
rect 16209 7701 16221 7735
rect 16255 7701 16267 7735
rect 16592 7732 16620 7908
rect 18156 7908 22560 7936
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7837 17371 7871
rect 17313 7831 17371 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 18046 7868 18052 7880
rect 17635 7840 18052 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17328 7800 17356 7831
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18156 7877 18184 7908
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 25222 7936 25228 7948
rect 22664 7908 25228 7936
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 19058 7868 19064 7880
rect 18279 7840 19064 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 20254 7828 20260 7880
rect 20312 7828 20318 7880
rect 22664 7877 22692 7908
rect 25222 7896 25228 7908
rect 25280 7896 25286 7948
rect 28626 7896 28632 7948
rect 28684 7936 28690 7948
rect 28684 7908 28856 7936
rect 28684 7896 28690 7908
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20855 7840 20913 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22189 7871 22247 7877
rect 22189 7868 22201 7871
rect 22143 7840 22201 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 22189 7837 22201 7840
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22649 7871 22707 7877
rect 22649 7837 22661 7871
rect 22695 7837 22707 7871
rect 22649 7831 22707 7837
rect 23937 7871 23995 7877
rect 23937 7837 23949 7871
rect 23983 7868 23995 7871
rect 24029 7871 24087 7877
rect 24029 7868 24041 7871
rect 23983 7840 24041 7868
rect 23983 7837 23995 7840
rect 23937 7831 23995 7837
rect 24029 7837 24041 7840
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24394 7828 24400 7880
rect 24452 7868 24458 7880
rect 24673 7871 24731 7877
rect 24673 7868 24685 7871
rect 24452 7840 24685 7868
rect 24452 7828 24458 7840
rect 24673 7837 24685 7840
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 26418 7828 26424 7880
rect 26476 7828 26482 7880
rect 26970 7828 26976 7880
rect 27028 7828 27034 7880
rect 27341 7871 27399 7877
rect 27341 7837 27353 7871
rect 27387 7868 27399 7871
rect 28442 7868 28448 7880
rect 27387 7840 28448 7868
rect 27387 7837 27399 7840
rect 27341 7831 27399 7837
rect 28442 7828 28448 7840
rect 28500 7828 28506 7880
rect 28828 7877 28856 7908
rect 28813 7871 28871 7877
rect 28813 7837 28825 7871
rect 28859 7837 28871 7871
rect 28813 7831 28871 7837
rect 19702 7800 19708 7812
rect 17328 7772 19708 7800
rect 19702 7760 19708 7772
rect 19760 7760 19766 7812
rect 28626 7800 28632 7812
rect 22388 7772 28632 7800
rect 20346 7732 20352 7744
rect 16592 7704 20352 7732
rect 16209 7695 16267 7701
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 21085 7735 21143 7741
rect 21085 7701 21097 7735
rect 21131 7732 21143 7735
rect 21910 7732 21916 7744
rect 21131 7704 21916 7732
rect 21131 7701 21143 7704
rect 21085 7695 21143 7701
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22388 7741 22416 7772
rect 28626 7760 28632 7772
rect 28684 7760 28690 7812
rect 29104 7800 29132 7967
rect 29454 7964 29460 8016
rect 29512 8004 29518 8016
rect 31018 8004 31024 8016
rect 29512 7976 31024 8004
rect 29512 7964 29518 7976
rect 31018 7964 31024 7976
rect 31076 7964 31082 8016
rect 38562 8004 38568 8016
rect 36372 7976 38568 8004
rect 31294 7936 31300 7948
rect 29288 7908 31300 7936
rect 29288 7877 29316 7908
rect 31294 7896 31300 7908
rect 31352 7896 31358 7948
rect 29273 7871 29331 7877
rect 29273 7837 29285 7871
rect 29319 7837 29331 7871
rect 29273 7831 29331 7837
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7868 30251 7871
rect 31570 7868 31576 7880
rect 30239 7840 31576 7868
rect 30239 7837 30251 7840
rect 30193 7831 30251 7837
rect 31570 7828 31576 7840
rect 31628 7828 31634 7880
rect 36372 7877 36400 7976
rect 38562 7964 38568 7976
rect 38620 7964 38626 8016
rect 38470 7936 38476 7948
rect 36740 7908 38476 7936
rect 36740 7877 36768 7908
rect 38470 7896 38476 7908
rect 38528 7896 38534 7948
rect 38672 7908 42932 7936
rect 36357 7871 36415 7877
rect 36357 7837 36369 7871
rect 36403 7837 36415 7871
rect 36357 7831 36415 7837
rect 36725 7871 36783 7877
rect 36725 7837 36737 7871
rect 36771 7837 36783 7871
rect 37001 7871 37059 7877
rect 37001 7868 37013 7871
rect 36725 7831 36783 7837
rect 36924 7840 37013 7868
rect 28920 7772 29132 7800
rect 28920 7744 28948 7772
rect 29178 7760 29184 7812
rect 29236 7800 29242 7812
rect 36446 7800 36452 7812
rect 29236 7772 36452 7800
rect 29236 7760 29242 7772
rect 36446 7760 36452 7772
rect 36504 7760 36510 7812
rect 22373 7735 22431 7741
rect 22373 7701 22385 7735
rect 22419 7701 22431 7735
rect 22373 7695 22431 7701
rect 24578 7692 24584 7744
rect 24636 7692 24642 7744
rect 26878 7692 26884 7744
rect 26936 7732 26942 7744
rect 27157 7735 27215 7741
rect 27157 7732 27169 7735
rect 26936 7704 27169 7732
rect 26936 7692 26942 7704
rect 27157 7701 27169 7704
rect 27203 7701 27215 7735
rect 27157 7695 27215 7701
rect 28902 7692 28908 7744
rect 28960 7692 28966 7744
rect 29270 7692 29276 7744
rect 29328 7732 29334 7744
rect 30009 7735 30067 7741
rect 30009 7732 30021 7735
rect 29328 7704 30021 7732
rect 29328 7692 29334 7704
rect 30009 7701 30021 7704
rect 30055 7701 30067 7735
rect 30009 7695 30067 7701
rect 33502 7692 33508 7744
rect 33560 7732 33566 7744
rect 36924 7732 36952 7840
rect 37001 7837 37013 7840
rect 37047 7837 37059 7871
rect 37001 7831 37059 7837
rect 37458 7828 37464 7880
rect 37516 7828 37522 7880
rect 37734 7828 37740 7880
rect 37792 7868 37798 7880
rect 38565 7871 38623 7877
rect 38565 7868 38577 7871
rect 37792 7840 38577 7868
rect 37792 7828 37798 7840
rect 38565 7837 38577 7840
rect 38611 7837 38623 7871
rect 38565 7831 38623 7837
rect 33560 7704 36952 7732
rect 33560 7692 33566 7704
rect 37274 7692 37280 7744
rect 37332 7732 37338 7744
rect 38672 7732 38700 7908
rect 38930 7828 38936 7880
rect 38988 7828 38994 7880
rect 39482 7828 39488 7880
rect 39540 7828 39546 7880
rect 40129 7871 40187 7877
rect 40129 7837 40141 7871
rect 40175 7868 40187 7871
rect 40678 7868 40684 7880
rect 40175 7840 40684 7868
rect 40175 7837 40187 7840
rect 40129 7831 40187 7837
rect 40678 7828 40684 7840
rect 40736 7828 40742 7880
rect 42153 7871 42211 7877
rect 42153 7868 42165 7871
rect 41386 7840 42165 7868
rect 38838 7760 38844 7812
rect 38896 7800 38902 7812
rect 41386 7800 41414 7840
rect 42153 7837 42165 7840
rect 42199 7837 42211 7871
rect 42153 7831 42211 7837
rect 42518 7828 42524 7880
rect 42576 7828 42582 7880
rect 42904 7877 42932 7908
rect 42889 7871 42947 7877
rect 42889 7837 42901 7871
rect 42935 7837 42947 7871
rect 42889 7831 42947 7837
rect 43254 7828 43260 7880
rect 43312 7828 43318 7880
rect 38896 7772 41414 7800
rect 38896 7760 38902 7772
rect 37332 7704 38700 7732
rect 37332 7692 37338 7704
rect 39298 7692 39304 7744
rect 39356 7692 39362 7744
rect 43070 7692 43076 7744
rect 43128 7692 43134 7744
rect 43438 7692 43444 7744
rect 43496 7692 43502 7744
rect 1104 7642 43884 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 43884 7642
rect 1104 7568 43884 7590
rect 4338 7488 4344 7540
rect 4396 7488 4402 7540
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 5166 7528 5172 7540
rect 4663 7500 5172 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5902 7488 5908 7540
rect 5960 7488 5966 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12621 7531 12679 7537
rect 12621 7528 12633 7531
rect 12492 7500 12633 7528
rect 12492 7488 12498 7500
rect 12621 7497 12633 7500
rect 12667 7497 12679 7531
rect 12621 7491 12679 7497
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 14424 7500 15945 7528
rect 14424 7488 14430 7500
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 15933 7491 15991 7497
rect 21818 7488 21824 7540
rect 21876 7488 21882 7540
rect 24486 7528 24492 7540
rect 22388 7500 24492 7528
rect 11606 7460 11612 7472
rect 4172 7432 11612 7460
rect 4172 7401 4200 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 12452 7432 12940 7460
rect 12452 7404 12480 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 11698 7392 11704 7404
rect 5767 7364 11704 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 4448 7324 4476 7355
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12434 7352 12440 7404
rect 12492 7352 12498 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12805 7395 12863 7401
rect 12805 7392 12817 7395
rect 12575 7364 12817 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12805 7361 12817 7364
rect 12851 7361 12863 7395
rect 12912 7392 12940 7432
rect 13078 7420 13084 7472
rect 13136 7460 13142 7472
rect 19518 7460 19524 7472
rect 13136 7432 19524 7460
rect 13136 7420 13142 7432
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 20254 7420 20260 7472
rect 20312 7460 20318 7472
rect 22278 7460 22284 7472
rect 20312 7432 22284 7460
rect 20312 7420 20318 7432
rect 22278 7420 22284 7432
rect 22336 7420 22342 7472
rect 14826 7392 14832 7404
rect 12912 7364 14832 7392
rect 12805 7355 12863 7361
rect 12820 7324 12848 7355
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 15194 7392 15200 7404
rect 14967 7364 15200 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16022 7392 16028 7404
rect 15887 7364 16028 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16022 7352 16028 7364
rect 16080 7392 16086 7404
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 16080 7364 16129 7392
rect 16080 7352 16086 7364
rect 16117 7361 16129 7364
rect 16163 7361 16175 7395
rect 18138 7392 18144 7404
rect 16117 7355 16175 7361
rect 16224 7364 18144 7392
rect 16224 7324 16252 7364
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7392 22063 7395
rect 22388 7392 22416 7500
rect 24486 7488 24492 7500
rect 24544 7488 24550 7540
rect 24578 7488 24584 7540
rect 24636 7528 24642 7540
rect 36538 7528 36544 7540
rect 24636 7500 36544 7528
rect 24636 7488 24642 7500
rect 36538 7488 36544 7500
rect 36596 7488 36602 7540
rect 37550 7488 37556 7540
rect 37608 7528 37614 7540
rect 38565 7531 38623 7537
rect 38565 7528 38577 7531
rect 37608 7500 38577 7528
rect 37608 7488 37614 7500
rect 38565 7497 38577 7500
rect 38611 7497 38623 7531
rect 38565 7491 38623 7497
rect 43073 7531 43131 7537
rect 43073 7497 43085 7531
rect 43119 7528 43131 7531
rect 43162 7528 43168 7540
rect 43119 7500 43168 7528
rect 43119 7497 43131 7500
rect 43073 7491 43131 7497
rect 43162 7488 43168 7500
rect 43220 7488 43226 7540
rect 22554 7420 22560 7472
rect 22612 7460 22618 7472
rect 28902 7460 28908 7472
rect 22612 7432 28908 7460
rect 22612 7420 22618 7432
rect 28902 7420 28908 7432
rect 28960 7420 28966 7472
rect 31846 7460 31852 7472
rect 30852 7432 31852 7460
rect 30852 7401 30880 7432
rect 31846 7420 31852 7432
rect 31904 7420 31910 7472
rect 33686 7420 33692 7472
rect 33744 7460 33750 7472
rect 37734 7460 37740 7472
rect 33744 7432 37740 7460
rect 33744 7420 33750 7432
rect 37734 7420 37740 7432
rect 37792 7420 37798 7472
rect 38838 7460 38844 7472
rect 37844 7432 38844 7460
rect 22051 7364 22416 7392
rect 24949 7395 25007 7401
rect 22051 7361 22063 7364
rect 22005 7355 22063 7361
rect 24949 7361 24961 7395
rect 24995 7392 25007 7395
rect 25041 7395 25099 7401
rect 25041 7392 25053 7395
rect 24995 7364 25053 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 25041 7361 25053 7364
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 30837 7395 30895 7401
rect 30837 7361 30849 7395
rect 30883 7361 30895 7395
rect 30837 7355 30895 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7392 31447 7395
rect 31754 7392 31760 7404
rect 31435 7364 31760 7392
rect 31435 7361 31447 7364
rect 31389 7355 31447 7361
rect 31754 7352 31760 7364
rect 31812 7352 31818 7404
rect 32490 7352 32496 7404
rect 32548 7392 32554 7404
rect 32585 7395 32643 7401
rect 32585 7392 32597 7395
rect 32548 7364 32597 7392
rect 32548 7352 32554 7364
rect 32585 7361 32597 7364
rect 32631 7361 32643 7395
rect 32585 7355 32643 7361
rect 33410 7352 33416 7404
rect 33468 7392 33474 7404
rect 35345 7395 35403 7401
rect 35345 7392 35357 7395
rect 33468 7364 35357 7392
rect 33468 7352 33474 7364
rect 35345 7361 35357 7364
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 36446 7352 36452 7404
rect 36504 7392 36510 7404
rect 37844 7392 37872 7432
rect 38838 7420 38844 7432
rect 38896 7420 38902 7472
rect 36504 7364 37872 7392
rect 36504 7352 36510 7364
rect 38654 7352 38660 7404
rect 38712 7392 38718 7404
rect 38749 7395 38807 7401
rect 38749 7392 38761 7395
rect 38712 7364 38761 7392
rect 38712 7352 38718 7364
rect 38749 7361 38761 7364
rect 38795 7361 38807 7395
rect 42889 7395 42947 7401
rect 42889 7392 42901 7395
rect 38749 7355 38807 7361
rect 41386 7364 42901 7392
rect 4448 7296 12756 7324
rect 12820 7296 16252 7324
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 12728 7256 12756 7296
rect 16298 7284 16304 7336
rect 16356 7324 16362 7336
rect 36814 7324 36820 7336
rect 16356 7296 36820 7324
rect 16356 7284 16362 7296
rect 36814 7284 36820 7296
rect 36872 7284 36878 7336
rect 14642 7256 14648 7268
rect 11664 7228 12664 7256
rect 12728 7228 14648 7256
rect 11664 7216 11670 7228
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 12434 7188 12440 7200
rect 11756 7160 12440 7188
rect 11756 7148 11762 7160
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 12636 7188 12664 7228
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 14918 7216 14924 7268
rect 14976 7256 14982 7268
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14976 7228 15025 7256
rect 14976 7216 14982 7228
rect 15013 7225 15025 7228
rect 15059 7225 15071 7259
rect 15013 7219 15071 7225
rect 24854 7216 24860 7268
rect 24912 7216 24918 7268
rect 41386 7256 41414 7364
rect 42889 7361 42901 7364
rect 42935 7361 42947 7395
rect 42889 7355 42947 7361
rect 43257 7395 43315 7401
rect 43257 7361 43269 7395
rect 43303 7361 43315 7395
rect 43257 7355 43315 7361
rect 41782 7284 41788 7336
rect 41840 7324 41846 7336
rect 43272 7324 43300 7355
rect 41840 7296 43300 7324
rect 41840 7284 41846 7296
rect 25148 7228 41414 7256
rect 14734 7188 14740 7200
rect 12636 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 14826 7148 14832 7200
rect 14884 7188 14890 7200
rect 17126 7188 17132 7200
rect 14884 7160 17132 7188
rect 14884 7148 14890 7160
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 21910 7148 21916 7200
rect 21968 7188 21974 7200
rect 25148 7188 25176 7228
rect 21968 7160 25176 7188
rect 25225 7191 25283 7197
rect 21968 7148 21974 7160
rect 25225 7157 25237 7191
rect 25271 7188 25283 7191
rect 25314 7188 25320 7200
rect 25271 7160 25320 7188
rect 25271 7157 25283 7160
rect 25225 7151 25283 7157
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 30650 7148 30656 7200
rect 30708 7148 30714 7200
rect 31202 7148 31208 7200
rect 31260 7148 31266 7200
rect 32306 7148 32312 7200
rect 32364 7188 32370 7200
rect 32401 7191 32459 7197
rect 32401 7188 32413 7191
rect 32364 7160 32413 7188
rect 32364 7148 32370 7160
rect 32401 7157 32413 7160
rect 32447 7157 32459 7191
rect 32401 7151 32459 7157
rect 34422 7148 34428 7200
rect 34480 7188 34486 7200
rect 35161 7191 35219 7197
rect 35161 7188 35173 7191
rect 34480 7160 35173 7188
rect 34480 7148 34486 7160
rect 35161 7157 35173 7160
rect 35207 7157 35219 7191
rect 35161 7151 35219 7157
rect 36538 7148 36544 7200
rect 36596 7188 36602 7200
rect 42518 7188 42524 7200
rect 36596 7160 42524 7188
rect 36596 7148 36602 7160
rect 42518 7148 42524 7160
rect 42576 7148 42582 7200
rect 43438 7148 43444 7200
rect 43496 7148 43502 7200
rect 1104 7098 43884 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 43884 7098
rect 1104 7024 43884 7046
rect 6273 6987 6331 6993
rect 6273 6953 6285 6987
rect 6319 6984 6331 6987
rect 6822 6984 6828 6996
rect 6319 6956 6828 6984
rect 6319 6953 6331 6956
rect 6273 6947 6331 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7834 6944 7840 6996
rect 7892 6944 7898 6996
rect 8662 6944 8668 6996
rect 8720 6984 8726 6996
rect 9585 6987 9643 6993
rect 9585 6984 9597 6987
rect 8720 6956 9597 6984
rect 8720 6944 8726 6956
rect 9585 6953 9597 6956
rect 9631 6953 9643 6987
rect 9585 6947 9643 6953
rect 13354 6944 13360 6996
rect 13412 6944 13418 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 23382 6984 23388 6996
rect 15252 6956 23388 6984
rect 15252 6944 15258 6956
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 33778 6944 33784 6996
rect 33836 6984 33842 6996
rect 39482 6984 39488 6996
rect 33836 6956 39488 6984
rect 33836 6944 33842 6956
rect 39482 6944 39488 6956
rect 39540 6944 39546 6996
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 7650 6916 7656 6928
rect 7432 6888 7656 6916
rect 7432 6876 7438 6888
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 19242 6916 19248 6928
rect 8904 6888 19248 6916
rect 8904 6876 8910 6888
rect 19242 6876 19248 6888
rect 19300 6876 19306 6928
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 26878 6916 26884 6928
rect 19392 6888 26884 6916
rect 19392 6876 19398 6888
rect 26878 6876 26884 6888
rect 26936 6876 26942 6928
rect 33045 6919 33103 6925
rect 33045 6916 33057 6919
rect 32784 6888 33057 6916
rect 22186 6848 22192 6860
rect 6886 6820 13308 6848
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3927 6752 4169 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6454 6780 6460 6792
rect 6135 6752 6460 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 6886 6780 6914 6820
rect 6779 6752 6914 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 9674 6780 9680 6792
rect 8067 6752 9680 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 4249 6715 4307 6721
rect 4249 6681 4261 6715
rect 4295 6712 4307 6715
rect 9784 6712 9812 6743
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 13165 6783 13223 6789
rect 13165 6780 13177 6783
rect 10100 6752 13177 6780
rect 10100 6740 10106 6752
rect 13165 6749 13177 6752
rect 13211 6749 13223 6783
rect 13165 6743 13223 6749
rect 13280 6776 13308 6820
rect 13464 6820 22192 6848
rect 13464 6776 13492 6820
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 23014 6848 23020 6860
rect 22296 6820 23020 6848
rect 19978 6780 19984 6792
rect 13280 6748 13492 6776
rect 18340 6752 19984 6780
rect 18340 6712 18368 6752
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6780 20131 6783
rect 22296 6780 22324 6820
rect 23014 6808 23020 6820
rect 23072 6808 23078 6860
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 26421 6851 26479 6857
rect 26421 6848 26433 6851
rect 26384 6820 26433 6848
rect 26384 6808 26390 6820
rect 26421 6817 26433 6820
rect 26467 6817 26479 6851
rect 26421 6811 26479 6817
rect 26786 6808 26792 6860
rect 26844 6848 26850 6860
rect 32784 6848 32812 6888
rect 33045 6885 33057 6888
rect 33091 6885 33103 6919
rect 33045 6879 33103 6885
rect 26844 6820 32812 6848
rect 26844 6808 26850 6820
rect 32858 6808 32864 6860
rect 32916 6848 32922 6860
rect 32916 6820 34928 6848
rect 32916 6808 32922 6820
rect 20119 6752 22324 6780
rect 22373 6783 22431 6789
rect 20119 6749 20131 6752
rect 20073 6743 20131 6749
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 4295 6684 9720 6712
rect 9784 6684 18368 6712
rect 4295 6681 4307 6684
rect 4249 6675 4307 6681
rect 4062 6604 4068 6656
rect 4120 6604 4126 6656
rect 6546 6604 6552 6656
rect 6604 6604 6610 6656
rect 7006 6604 7012 6656
rect 7064 6604 7070 6656
rect 9692 6644 9720 6684
rect 18414 6672 18420 6724
rect 18472 6712 18478 6724
rect 22388 6712 22416 6743
rect 24394 6740 24400 6792
rect 24452 6780 24458 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 24452 6752 24685 6780
rect 24452 6740 24458 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6780 26571 6783
rect 26605 6783 26663 6789
rect 26605 6780 26617 6783
rect 26559 6752 26617 6780
rect 26559 6749 26571 6752
rect 26513 6743 26571 6749
rect 26605 6749 26617 6752
rect 26651 6749 26663 6783
rect 26605 6743 26663 6749
rect 32674 6740 32680 6792
rect 32732 6780 32738 6792
rect 34900 6789 34928 6820
rect 36446 6808 36452 6860
rect 36504 6848 36510 6860
rect 36504 6820 41414 6848
rect 36504 6808 36510 6820
rect 33229 6783 33287 6789
rect 33229 6780 33241 6783
rect 32732 6752 33241 6780
rect 32732 6740 32738 6752
rect 33229 6749 33241 6752
rect 33275 6749 33287 6783
rect 33229 6743 33287 6749
rect 34885 6783 34943 6789
rect 34885 6749 34897 6783
rect 34931 6749 34943 6783
rect 34885 6743 34943 6749
rect 40862 6740 40868 6792
rect 40920 6740 40926 6792
rect 41386 6780 41414 6820
rect 42889 6783 42947 6789
rect 42889 6780 42901 6783
rect 41386 6752 42901 6780
rect 42889 6749 42901 6752
rect 42935 6749 42947 6783
rect 42889 6743 42947 6749
rect 42978 6740 42984 6792
rect 43036 6780 43042 6792
rect 43257 6783 43315 6789
rect 43257 6780 43269 6783
rect 43036 6752 43269 6780
rect 43036 6740 43042 6752
rect 43257 6749 43269 6752
rect 43303 6749 43315 6783
rect 43257 6743 43315 6749
rect 29362 6712 29368 6724
rect 18472 6684 22094 6712
rect 22388 6684 29368 6712
rect 18472 6672 18478 6684
rect 15930 6644 15936 6656
rect 9692 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 16632 6616 19901 6644
rect 16632 6604 16638 6616
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 22066 6644 22094 6684
rect 29362 6672 29368 6684
rect 29420 6672 29426 6724
rect 37826 6712 37832 6724
rect 33152 6684 37832 6712
rect 22189 6647 22247 6653
rect 22189 6644 22201 6647
rect 22066 6616 22201 6644
rect 19889 6607 19947 6613
rect 22189 6613 22201 6616
rect 22235 6613 22247 6647
rect 22189 6607 22247 6613
rect 24578 6604 24584 6656
rect 24636 6604 24642 6656
rect 26789 6647 26847 6653
rect 26789 6613 26801 6647
rect 26835 6644 26847 6647
rect 33152 6644 33180 6684
rect 37826 6672 37832 6684
rect 37884 6672 37890 6724
rect 26835 6616 33180 6644
rect 26835 6613 26847 6616
rect 26789 6607 26847 6613
rect 33226 6604 33232 6656
rect 33284 6644 33290 6656
rect 34701 6647 34759 6653
rect 34701 6644 34713 6647
rect 33284 6616 34713 6644
rect 33284 6604 33290 6616
rect 34701 6613 34713 6616
rect 34747 6613 34759 6647
rect 34701 6607 34759 6613
rect 38470 6604 38476 6656
rect 38528 6644 38534 6656
rect 40681 6647 40739 6653
rect 40681 6644 40693 6647
rect 38528 6616 40693 6644
rect 38528 6604 38534 6616
rect 40681 6613 40693 6616
rect 40727 6613 40739 6647
rect 40681 6607 40739 6613
rect 43070 6604 43076 6656
rect 43128 6604 43134 6656
rect 43438 6604 43444 6656
rect 43496 6604 43502 6656
rect 1104 6554 43884 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 43884 6554
rect 1104 6480 43884 6502
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7708 6412 7941 6440
rect 7708 6400 7714 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8812 6412 8953 6440
rect 8812 6400 8818 6412
rect 8941 6409 8953 6412
rect 8987 6409 8999 6443
rect 8941 6403 8999 6409
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 9582 6440 9588 6452
rect 9539 6412 9588 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 10686 6400 10692 6452
rect 10744 6400 10750 6452
rect 11606 6400 11612 6452
rect 11664 6400 11670 6452
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12342 6440 12348 6452
rect 12023 6412 12348 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 13504 6412 15853 6440
rect 13504 6400 13510 6412
rect 15841 6409 15853 6412
rect 15887 6409 15899 6443
rect 15841 6403 15899 6409
rect 19242 6400 19248 6452
rect 19300 6400 19306 6452
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 24394 6440 24400 6452
rect 20956 6412 24400 6440
rect 20956 6400 20962 6412
rect 24394 6400 24400 6412
rect 24452 6400 24458 6452
rect 24578 6400 24584 6452
rect 24636 6440 24642 6452
rect 36725 6443 36783 6449
rect 24636 6412 36676 6440
rect 24636 6400 24642 6412
rect 1210 6332 1216 6384
rect 1268 6372 1274 6384
rect 8846 6372 8852 6384
rect 1268 6344 8852 6372
rect 1268 6332 1274 6344
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 10042 6372 10048 6384
rect 9600 6344 10048 6372
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 9600 6236 9628 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 21358 6372 21364 6384
rect 12820 6344 21364 6372
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 5684 6208 9628 6236
rect 9692 6236 9720 6267
rect 10134 6264 10140 6316
rect 10192 6264 10198 6316
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 12820 6313 12848 6344
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 30374 6332 30380 6384
rect 30432 6372 30438 6384
rect 36446 6372 36452 6384
rect 30432 6344 36452 6372
rect 30432 6332 30438 6344
rect 36446 6332 36452 6344
rect 36504 6332 36510 6384
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 11793 6307 11851 6313
rect 11793 6304 11805 6307
rect 11747 6276 11805 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 11793 6273 11805 6276
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6304 16083 6307
rect 19058 6304 19064 6316
rect 16071 6276 19064 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 19058 6264 19064 6276
rect 19116 6264 19122 6316
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6304 19487 6307
rect 20806 6304 20812 6316
rect 19475 6276 20812 6304
rect 19475 6273 19487 6276
rect 19429 6267 19487 6273
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 22462 6264 22468 6316
rect 22520 6304 22526 6316
rect 36541 6307 36599 6313
rect 36541 6304 36553 6307
rect 22520 6276 36553 6304
rect 22520 6264 22526 6276
rect 36541 6273 36553 6276
rect 36587 6273 36599 6307
rect 36541 6267 36599 6273
rect 17310 6236 17316 6248
rect 9692 6208 17316 6236
rect 5684 6196 5690 6208
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 36648 6236 36676 6412
rect 36725 6409 36737 6443
rect 36771 6440 36783 6443
rect 37642 6440 37648 6452
rect 36771 6412 37648 6440
rect 36771 6409 36783 6412
rect 36725 6403 36783 6409
rect 37642 6400 37648 6412
rect 37700 6400 37706 6452
rect 43438 6400 43444 6452
rect 43496 6400 43502 6452
rect 40126 6264 40132 6316
rect 40184 6304 40190 6316
rect 42889 6307 42947 6313
rect 42889 6304 42901 6307
rect 40184 6276 42901 6304
rect 40184 6264 40190 6276
rect 42889 6273 42901 6276
rect 42935 6273 42947 6307
rect 42889 6267 42947 6273
rect 43257 6307 43315 6313
rect 43257 6273 43269 6307
rect 43303 6304 43315 6307
rect 43303 6276 43944 6304
rect 43303 6273 43315 6276
rect 43257 6267 43315 6273
rect 43162 6236 43168 6248
rect 36648 6208 43168 6236
rect 43162 6196 43168 6208
rect 43220 6196 43226 6248
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 9953 6171 10011 6177
rect 9953 6168 9965 6171
rect 9548 6140 9965 6168
rect 9548 6128 9554 6140
rect 9953 6137 9965 6140
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 30650 6168 30656 6180
rect 18012 6140 30656 6168
rect 18012 6128 18018 6140
rect 30650 6128 30656 6140
rect 30708 6128 30714 6180
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 12621 6103 12679 6109
rect 12621 6100 12633 6103
rect 7524 6072 12633 6100
rect 7524 6060 7530 6072
rect 12621 6069 12633 6072
rect 12667 6069 12679 6103
rect 12621 6063 12679 6069
rect 16758 6060 16764 6112
rect 16816 6100 16822 6112
rect 26786 6100 26792 6112
rect 16816 6072 26792 6100
rect 16816 6060 16822 6072
rect 26786 6060 26792 6072
rect 26844 6060 26850 6112
rect 43070 6060 43076 6112
rect 43128 6060 43134 6112
rect 1104 6010 43884 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 43884 6010
rect 1104 5936 43884 5958
rect 4985 5899 5043 5905
rect 4985 5865 4997 5899
rect 5031 5896 5043 5899
rect 6270 5896 6276 5908
rect 5031 5868 6276 5896
rect 5031 5865 5043 5868
rect 4985 5859 5043 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 6512 5868 6914 5896
rect 6512 5856 6518 5868
rect 6886 5828 6914 5868
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 11149 5899 11207 5905
rect 11149 5896 11161 5899
rect 9916 5868 11161 5896
rect 9916 5856 9922 5868
rect 11149 5865 11161 5868
rect 11195 5865 11207 5899
rect 11149 5859 11207 5865
rect 18598 5856 18604 5908
rect 18656 5856 18662 5908
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 43916 5896 43944 6276
rect 20772 5868 43944 5896
rect 20772 5856 20778 5868
rect 22189 5831 22247 5837
rect 6886 5800 22094 5828
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 21726 5760 21732 5772
rect 7248 5732 21732 5760
rect 7248 5720 7254 5732
rect 21726 5720 21732 5732
rect 21784 5720 21790 5772
rect 22066 5760 22094 5800
rect 22189 5797 22201 5831
rect 22235 5828 22247 5831
rect 33594 5828 33600 5840
rect 22235 5800 33600 5828
rect 22235 5797 22247 5800
rect 22189 5791 22247 5797
rect 33594 5788 33600 5800
rect 33652 5788 33658 5840
rect 38562 5788 38568 5840
rect 38620 5828 38626 5840
rect 39393 5831 39451 5837
rect 39393 5828 39405 5831
rect 38620 5800 39405 5828
rect 38620 5788 38626 5800
rect 39393 5797 39405 5800
rect 39439 5797 39451 5831
rect 39393 5791 39451 5797
rect 43438 5788 43444 5840
rect 43496 5788 43502 5840
rect 22370 5760 22376 5772
rect 22066 5732 22376 5760
rect 22370 5720 22376 5732
rect 22428 5720 22434 5772
rect 23290 5720 23296 5772
rect 23348 5760 23354 5772
rect 23348 5732 30374 5760
rect 23348 5720 23354 5732
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 4801 5695 4859 5701
rect 4801 5692 4813 5695
rect 4755 5664 4813 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 4801 5661 4813 5664
rect 4847 5692 4859 5695
rect 10870 5692 10876 5704
rect 4847 5664 10876 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 18598 5692 18604 5704
rect 11379 5664 18604 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5692 18751 5695
rect 18785 5695 18843 5701
rect 18785 5692 18797 5695
rect 18739 5664 18797 5692
rect 18739 5661 18751 5664
rect 18693 5655 18751 5661
rect 18785 5661 18797 5664
rect 18831 5661 18843 5695
rect 21634 5692 21640 5704
rect 18785 5655 18843 5661
rect 18892 5664 21640 5692
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 18892 5624 18920 5664
rect 21634 5652 21640 5664
rect 21692 5652 21698 5704
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5692 21971 5695
rect 22005 5695 22063 5701
rect 22005 5692 22017 5695
rect 21959 5664 22017 5692
rect 21959 5661 21971 5664
rect 21913 5655 21971 5661
rect 22005 5661 22017 5664
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 26418 5652 26424 5704
rect 26476 5652 26482 5704
rect 30346 5692 30374 5732
rect 32508 5732 41414 5760
rect 32508 5692 32536 5732
rect 30346 5664 32536 5692
rect 39574 5652 39580 5704
rect 39632 5652 39638 5704
rect 41386 5692 41414 5732
rect 42889 5695 42947 5701
rect 42889 5692 42901 5695
rect 41386 5664 42901 5692
rect 42889 5661 42901 5664
rect 42935 5661 42947 5695
rect 42889 5655 42947 5661
rect 43257 5695 43315 5701
rect 43257 5661 43269 5695
rect 43303 5692 43315 5695
rect 43346 5692 43352 5704
rect 43303 5664 43352 5692
rect 43303 5661 43315 5664
rect 43257 5655 43315 5661
rect 43346 5652 43352 5664
rect 43404 5652 43410 5704
rect 42978 5624 42984 5636
rect 9732 5596 18920 5624
rect 18984 5596 42984 5624
rect 9732 5584 9738 5596
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 18506 5556 18512 5568
rect 9180 5528 18512 5556
rect 9180 5516 9186 5528
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 18984 5565 19012 5596
rect 42978 5584 42984 5596
rect 43036 5584 43042 5636
rect 18969 5559 19027 5565
rect 18969 5525 18981 5559
rect 19015 5525 19027 5559
rect 18969 5519 19027 5525
rect 21818 5516 21824 5568
rect 21876 5516 21882 5568
rect 26602 5516 26608 5568
rect 26660 5516 26666 5568
rect 43070 5516 43076 5568
rect 43128 5516 43134 5568
rect 1104 5466 43884 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 43884 5466
rect 1104 5392 43884 5414
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5352 10287 5355
rect 10318 5352 10324 5364
rect 10275 5324 10324 5352
rect 10275 5321 10287 5324
rect 10229 5315 10287 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 12894 5312 12900 5364
rect 12952 5312 12958 5364
rect 17034 5312 17040 5364
rect 17092 5352 17098 5364
rect 28258 5352 28264 5364
rect 17092 5324 28264 5352
rect 17092 5312 17098 5324
rect 28258 5312 28264 5324
rect 28316 5312 28322 5364
rect 29641 5355 29699 5361
rect 29641 5321 29653 5355
rect 29687 5352 29699 5355
rect 38746 5352 38752 5364
rect 29687 5324 38752 5352
rect 29687 5321 29699 5324
rect 29641 5315 29699 5321
rect 38746 5312 38752 5324
rect 38804 5312 38810 5364
rect 43438 5312 43444 5364
rect 43496 5312 43502 5364
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 8904 5256 10180 5284
rect 8904 5244 8910 5256
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 10060 5080 10088 5179
rect 10152 5148 10180 5256
rect 12406 5256 27108 5284
rect 12406 5148 12434 5256
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 10152 5120 12434 5148
rect 13096 5148 13124 5179
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 27080 5225 27108 5256
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 13780 5188 20269 5216
rect 13780 5176 13786 5188
rect 20257 5185 20269 5188
rect 20303 5216 20315 5219
rect 20441 5219 20499 5225
rect 20441 5216 20453 5219
rect 20303 5188 20453 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 20441 5185 20453 5188
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5185 24547 5219
rect 24489 5179 24547 5185
rect 27065 5219 27123 5225
rect 27065 5185 27077 5219
rect 27111 5185 27123 5219
rect 27065 5179 27123 5185
rect 29457 5219 29515 5225
rect 29457 5185 29469 5219
rect 29503 5216 29515 5219
rect 30926 5216 30932 5228
rect 29503 5188 30932 5216
rect 29503 5185 29515 5188
rect 29457 5179 29515 5185
rect 23566 5148 23572 5160
rect 13096 5120 23572 5148
rect 23566 5108 23572 5120
rect 23624 5108 23630 5160
rect 17034 5080 17040 5092
rect 10060 5052 17040 5080
rect 17034 5040 17040 5052
rect 17092 5040 17098 5092
rect 20622 4972 20628 5024
rect 20680 4972 20686 5024
rect 24504 5012 24532 5179
rect 30926 5176 30932 5188
rect 30984 5176 30990 5228
rect 40034 5176 40040 5228
rect 40092 5216 40098 5228
rect 42889 5219 42947 5225
rect 42889 5216 42901 5219
rect 40092 5188 42901 5216
rect 40092 5176 40098 5188
rect 42889 5185 42901 5188
rect 42935 5185 42947 5219
rect 42889 5179 42947 5185
rect 43257 5219 43315 5225
rect 43257 5185 43269 5219
rect 43303 5185 43315 5219
rect 43257 5179 43315 5185
rect 32766 5148 32772 5160
rect 24688 5120 32772 5148
rect 24688 5089 24716 5120
rect 32766 5108 32772 5120
rect 32824 5108 32830 5160
rect 42334 5108 42340 5160
rect 42392 5148 42398 5160
rect 43272 5148 43300 5179
rect 42392 5120 43300 5148
rect 42392 5108 42398 5120
rect 24673 5083 24731 5089
rect 24673 5049 24685 5083
rect 24719 5049 24731 5083
rect 24673 5043 24731 5049
rect 27249 5083 27307 5089
rect 27249 5049 27261 5083
rect 27295 5080 27307 5083
rect 40310 5080 40316 5092
rect 27295 5052 40316 5080
rect 27295 5049 27307 5052
rect 27249 5043 27307 5049
rect 40310 5040 40316 5052
rect 40368 5040 40374 5092
rect 28810 5012 28816 5024
rect 24504 4984 28816 5012
rect 28810 4972 28816 4984
rect 28868 4972 28874 5024
rect 43070 4972 43076 5024
rect 43128 4972 43134 5024
rect 1104 4922 43884 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 43884 4922
rect 1104 4848 43884 4870
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9398 4808 9404 4820
rect 9171 4780 9404 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 25130 4808 25136 4820
rect 11020 4780 25136 4808
rect 11020 4768 11026 4780
rect 25130 4768 25136 4780
rect 25188 4768 25194 4820
rect 32398 4768 32404 4820
rect 32456 4768 32462 4820
rect 33686 4768 33692 4820
rect 33744 4768 33750 4820
rect 36630 4768 36636 4820
rect 36688 4768 36694 4820
rect 38749 4811 38807 4817
rect 38749 4777 38761 4811
rect 38795 4808 38807 4811
rect 39942 4808 39948 4820
rect 38795 4780 39948 4808
rect 38795 4777 38807 4780
rect 38749 4771 38807 4777
rect 39942 4768 39948 4780
rect 40000 4768 40006 4820
rect 20622 4700 20628 4752
rect 20680 4740 20686 4752
rect 30374 4740 30380 4752
rect 20680 4712 30380 4740
rect 20680 4700 20686 4712
rect 30374 4700 30380 4712
rect 30432 4700 30438 4752
rect 31481 4743 31539 4749
rect 31481 4709 31493 4743
rect 31527 4740 31539 4743
rect 34790 4740 34796 4752
rect 31527 4712 34796 4740
rect 31527 4709 31539 4712
rect 31481 4703 31539 4709
rect 34790 4700 34796 4712
rect 34848 4700 34854 4752
rect 37274 4740 37280 4752
rect 36372 4712 37280 4740
rect 12406 4644 28028 4672
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4604 8999 4607
rect 12406 4604 12434 4644
rect 8987 4576 12434 4604
rect 22557 4607 22615 4613
rect 8987 4573 8999 4576
rect 8941 4567 8999 4573
rect 22557 4573 22569 4607
rect 22603 4604 22615 4607
rect 22649 4607 22707 4613
rect 22649 4604 22661 4607
rect 22603 4576 22661 4604
rect 22603 4573 22615 4576
rect 22557 4567 22615 4573
rect 22649 4573 22661 4576
rect 22695 4573 22707 4607
rect 28000 4604 28028 4644
rect 28074 4632 28080 4684
rect 28132 4672 28138 4684
rect 36372 4672 36400 4712
rect 37274 4700 37280 4712
rect 37332 4700 37338 4752
rect 43438 4700 43444 4752
rect 43496 4700 43502 4752
rect 39390 4672 39396 4684
rect 28132 4644 36400 4672
rect 36464 4644 39396 4672
rect 28132 4632 28138 4644
rect 28534 4604 28540 4616
rect 28000 4576 28540 4604
rect 22649 4567 22707 4573
rect 28534 4564 28540 4576
rect 28592 4564 28598 4616
rect 31297 4607 31355 4613
rect 31297 4573 31309 4607
rect 31343 4573 31355 4607
rect 31297 4567 31355 4573
rect 19334 4496 19340 4548
rect 19392 4536 19398 4548
rect 22465 4539 22523 4545
rect 22465 4536 22477 4539
rect 19392 4508 22477 4536
rect 19392 4496 19398 4508
rect 22465 4505 22477 4508
rect 22511 4505 22523 4539
rect 31312 4536 31340 4567
rect 31754 4564 31760 4616
rect 31812 4604 31818 4616
rect 32217 4607 32275 4613
rect 32217 4604 32229 4607
rect 31812 4576 32229 4604
rect 31812 4564 31818 4576
rect 32217 4573 32229 4576
rect 32263 4573 32275 4607
rect 32217 4567 32275 4573
rect 33505 4607 33563 4613
rect 33505 4573 33517 4607
rect 33551 4604 33563 4607
rect 35158 4604 35164 4616
rect 33551 4576 35164 4604
rect 33551 4573 33563 4576
rect 33505 4567 33563 4573
rect 35158 4564 35164 4576
rect 35216 4564 35222 4616
rect 36464 4613 36492 4644
rect 39390 4632 39396 4644
rect 39448 4632 39454 4684
rect 36449 4607 36507 4613
rect 36449 4573 36461 4607
rect 36495 4573 36507 4607
rect 36449 4567 36507 4573
rect 38565 4607 38623 4613
rect 38565 4573 38577 4607
rect 38611 4604 38623 4607
rect 41506 4604 41512 4616
rect 38611 4576 41512 4604
rect 38611 4573 38623 4576
rect 38565 4567 38623 4573
rect 41506 4564 41512 4576
rect 41564 4564 41570 4616
rect 42886 4564 42892 4616
rect 42944 4564 42950 4616
rect 43257 4607 43315 4613
rect 43257 4573 43269 4607
rect 43303 4573 43315 4607
rect 43257 4567 43315 4573
rect 32766 4536 32772 4548
rect 31312 4508 32772 4536
rect 22465 4499 22523 4505
rect 32766 4496 32772 4508
rect 32824 4496 32830 4548
rect 43272 4536 43300 4567
rect 33612 4508 43300 4536
rect 22830 4428 22836 4480
rect 22888 4428 22894 4480
rect 30374 4428 30380 4480
rect 30432 4468 30438 4480
rect 33612 4468 33640 4508
rect 30432 4440 33640 4468
rect 30432 4428 30438 4440
rect 43070 4428 43076 4480
rect 43128 4428 43134 4480
rect 1104 4378 43884 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 43884 4378
rect 1104 4304 43884 4326
rect 15562 4224 15568 4276
rect 15620 4224 15626 4276
rect 22830 4224 22836 4276
rect 22888 4264 22894 4276
rect 42886 4264 42892 4276
rect 22888 4236 42892 4264
rect 22888 4224 22894 4236
rect 42886 4224 42892 4236
rect 42944 4224 42950 4276
rect 15657 4199 15715 4205
rect 15657 4165 15669 4199
rect 15703 4196 15715 4199
rect 15841 4199 15899 4205
rect 15841 4196 15853 4199
rect 15703 4168 15853 4196
rect 15703 4165 15715 4168
rect 15657 4159 15715 4165
rect 15841 4165 15853 4168
rect 15887 4165 15899 4199
rect 15841 4159 15899 4165
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 19484 4100 21833 4128
rect 19484 4088 19490 4100
rect 21821 4097 21833 4100
rect 21867 4128 21879 4131
rect 22097 4131 22155 4137
rect 22097 4128 22109 4131
rect 21867 4100 22109 4128
rect 21867 4097 21879 4100
rect 21821 4091 21879 4097
rect 22097 4097 22109 4100
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 22830 4088 22836 4140
rect 22888 4088 22894 4140
rect 24578 4088 24584 4140
rect 24636 4128 24642 4140
rect 25685 4131 25743 4137
rect 25685 4128 25697 4131
rect 24636 4100 25697 4128
rect 24636 4088 24642 4100
rect 25685 4097 25697 4100
rect 25731 4097 25743 4131
rect 25685 4091 25743 4097
rect 35069 4131 35127 4137
rect 35069 4097 35081 4131
rect 35115 4128 35127 4131
rect 37274 4128 37280 4140
rect 35115 4100 37280 4128
rect 35115 4097 35127 4100
rect 35069 4091 35127 4097
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 40865 4131 40923 4137
rect 40865 4097 40877 4131
rect 40911 4097 40923 4131
rect 40865 4091 40923 4097
rect 16025 4063 16083 4069
rect 16025 4029 16037 4063
rect 16071 4060 16083 4063
rect 20714 4060 20720 4072
rect 16071 4032 20720 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 30374 4060 30380 4072
rect 22020 4032 30380 4060
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 21818 3992 21824 4004
rect 18288 3964 21824 3992
rect 18288 3952 18294 3964
rect 21818 3952 21824 3964
rect 21876 3952 21882 4004
rect 22020 4001 22048 4032
rect 30374 4020 30380 4032
rect 30432 4020 30438 4072
rect 40880 4060 40908 4091
rect 40954 4088 40960 4140
rect 41012 4128 41018 4140
rect 42889 4131 42947 4137
rect 42889 4128 42901 4131
rect 41012 4100 42901 4128
rect 41012 4088 41018 4100
rect 42889 4097 42901 4100
rect 42935 4097 42947 4131
rect 42889 4091 42947 4097
rect 43162 4088 43168 4140
rect 43220 4128 43226 4140
rect 43257 4131 43315 4137
rect 43257 4128 43269 4131
rect 43220 4100 43269 4128
rect 43220 4088 43226 4100
rect 43257 4097 43269 4100
rect 43303 4097 43315 4131
rect 43257 4091 43315 4097
rect 43622 4060 43628 4072
rect 40880 4032 43628 4060
rect 43622 4020 43628 4032
rect 43680 4020 43686 4072
rect 22005 3995 22063 4001
rect 22005 3961 22017 3995
rect 22051 3961 22063 3995
rect 22005 3955 22063 3961
rect 23014 3952 23020 4004
rect 23072 3952 23078 4004
rect 25866 3952 25872 4004
rect 25924 3952 25930 4004
rect 35253 3995 35311 4001
rect 35253 3961 35265 3995
rect 35299 3992 35311 3995
rect 38930 3992 38936 4004
rect 35299 3964 38936 3992
rect 35299 3961 35311 3964
rect 35253 3955 35311 3961
rect 38930 3952 38936 3964
rect 38988 3952 38994 4004
rect 40678 3952 40684 4004
rect 40736 3952 40742 4004
rect 43438 3952 43444 4004
rect 43496 3952 43502 4004
rect 13538 3884 13544 3936
rect 13596 3924 13602 3936
rect 21910 3924 21916 3936
rect 13596 3896 21916 3924
rect 13596 3884 13602 3896
rect 21910 3884 21916 3896
rect 21968 3884 21974 3936
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 26694 3924 26700 3936
rect 22796 3896 26700 3924
rect 22796 3884 22802 3896
rect 26694 3884 26700 3896
rect 26752 3884 26758 3936
rect 43070 3884 43076 3936
rect 43128 3884 43134 3936
rect 1104 3834 43884 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 43884 3834
rect 1104 3760 43884 3782
rect 17218 3680 17224 3732
rect 17276 3680 17282 3732
rect 18506 3680 18512 3732
rect 18564 3680 18570 3732
rect 19978 3680 19984 3732
rect 20036 3720 20042 3732
rect 22738 3720 22744 3732
rect 20036 3692 22744 3720
rect 20036 3680 20042 3692
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 34885 3723 34943 3729
rect 23032 3692 31754 3720
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 22925 3655 22983 3661
rect 22925 3652 22937 3655
rect 9916 3624 18460 3652
rect 9916 3612 9922 3624
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 18230 3584 18236 3596
rect 7708 3556 18236 3584
rect 7708 3544 7714 3556
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 17313 3519 17371 3525
rect 17313 3485 17325 3519
rect 17359 3516 17371 3519
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 17359 3488 17417 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 17405 3485 17417 3488
rect 17451 3485 17463 3519
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17405 3479 17463 3485
rect 17512 3488 18153 3516
rect 15378 3408 15384 3460
rect 15436 3448 15442 3460
rect 17512 3448 17540 3488
rect 18141 3485 18153 3488
rect 18187 3516 18199 3519
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 18187 3488 18337 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18432 3516 18460 3624
rect 22066 3624 22937 3652
rect 21910 3544 21916 3596
rect 21968 3584 21974 3596
rect 22066 3584 22094 3624
rect 22925 3621 22937 3624
rect 22971 3621 22983 3655
rect 22925 3615 22983 3621
rect 21968 3556 22094 3584
rect 21968 3544 21974 3556
rect 23032 3516 23060 3692
rect 31726 3652 31754 3692
rect 34885 3689 34897 3723
rect 34931 3720 34943 3723
rect 35802 3720 35808 3732
rect 34931 3692 35808 3720
rect 34931 3689 34943 3692
rect 34885 3683 34943 3689
rect 35802 3680 35808 3692
rect 35860 3680 35866 3732
rect 36538 3680 36544 3732
rect 36596 3720 36602 3732
rect 36596 3692 42932 3720
rect 36596 3680 36602 3692
rect 42334 3652 42340 3664
rect 31726 3624 42340 3652
rect 42334 3612 42340 3624
rect 42392 3612 42398 3664
rect 24854 3544 24860 3596
rect 24912 3544 24918 3596
rect 25406 3584 25412 3596
rect 25148 3556 25412 3584
rect 18432 3488 23060 3516
rect 18325 3479 18383 3485
rect 23106 3476 23112 3528
rect 23164 3476 23170 3528
rect 24949 3519 25007 3525
rect 24949 3485 24961 3519
rect 24995 3516 25007 3519
rect 25041 3519 25099 3525
rect 25041 3516 25053 3519
rect 24995 3488 25053 3516
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 25041 3485 25053 3488
rect 25087 3485 25099 3519
rect 25041 3479 25099 3485
rect 25148 3448 25176 3556
rect 25406 3544 25412 3556
rect 25464 3544 25470 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 40126 3584 40132 3596
rect 25556 3556 40132 3584
rect 25556 3544 25562 3556
rect 40126 3544 40132 3556
rect 40184 3544 40190 3596
rect 15436 3420 17540 3448
rect 17604 3420 25176 3448
rect 25240 3488 34652 3516
rect 15436 3408 15442 3420
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 13998 3380 14004 3392
rect 9640 3352 14004 3380
rect 9640 3340 9646 3352
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 17604 3389 17632 3420
rect 25240 3389 25268 3488
rect 34624 3448 34652 3488
rect 34698 3476 34704 3528
rect 34756 3476 34762 3528
rect 42904 3525 42932 3692
rect 43438 3612 43444 3664
rect 43496 3612 43502 3664
rect 42889 3519 42947 3525
rect 42889 3485 42901 3519
rect 42935 3485 42947 3519
rect 42889 3479 42947 3485
rect 43257 3519 43315 3525
rect 43257 3485 43269 3519
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 43272 3448 43300 3479
rect 34624 3420 43300 3448
rect 17589 3383 17647 3389
rect 17589 3349 17601 3383
rect 17635 3349 17647 3383
rect 17589 3343 17647 3349
rect 25225 3383 25283 3389
rect 25225 3349 25237 3383
rect 25271 3349 25283 3383
rect 25225 3343 25283 3349
rect 25406 3340 25412 3392
rect 25464 3380 25470 3392
rect 40034 3380 40040 3392
rect 25464 3352 40040 3380
rect 25464 3340 25470 3352
rect 40034 3340 40040 3352
rect 40092 3340 40098 3392
rect 43070 3340 43076 3392
rect 43128 3340 43134 3392
rect 1104 3290 43884 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 43884 3290
rect 1104 3216 43884 3238
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 12437 3179 12495 3185
rect 7892 3148 12388 3176
rect 7892 3136 7898 3148
rect 12360 3117 12388 3148
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 23290 3176 23296 3188
rect 12483 3148 23296 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 23382 3136 23388 3188
rect 23440 3176 23446 3188
rect 23753 3179 23811 3185
rect 23753 3176 23765 3179
rect 23440 3148 23765 3176
rect 23440 3136 23446 3148
rect 23753 3145 23765 3148
rect 23799 3145 23811 3179
rect 23753 3139 23811 3145
rect 24121 3179 24179 3185
rect 24121 3145 24133 3179
rect 24167 3176 24179 3179
rect 28902 3176 28908 3188
rect 24167 3148 26832 3176
rect 24167 3145 24179 3148
rect 24121 3139 24179 3145
rect 12345 3111 12403 3117
rect 12345 3077 12357 3111
rect 12391 3077 12403 3111
rect 12345 3071 12403 3077
rect 13998 3068 14004 3120
rect 14056 3068 14062 3120
rect 16482 3068 16488 3120
rect 16540 3108 16546 3120
rect 16761 3111 16819 3117
rect 16761 3108 16773 3111
rect 16540 3080 16773 3108
rect 16540 3068 16546 3080
rect 16761 3077 16773 3080
rect 16807 3077 16819 3111
rect 16761 3071 16819 3077
rect 16945 3111 17003 3117
rect 16945 3077 16957 3111
rect 16991 3108 17003 3111
rect 16991 3080 22094 3108
rect 16991 3077 17003 3080
rect 16945 3071 17003 3077
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 7064 3012 9689 3040
rect 7064 3000 7070 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 9858 3000 9864 3052
rect 9916 3000 9922 3052
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11839 3012 11989 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 11977 3003 12035 3009
rect 12406 3012 14381 3040
rect 9490 2932 9496 2984
rect 9548 2972 9554 2984
rect 12406 2972 12434 3012
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 16776 3040 16804 3071
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16776 3012 17049 3040
rect 14369 3003 14427 3009
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 17957 3043 18015 3049
rect 17957 3040 17969 3043
rect 17911 3012 17969 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 17957 3009 17969 3012
rect 18003 3009 18015 3043
rect 17957 3003 18015 3009
rect 19978 3000 19984 3052
rect 20036 3000 20042 3052
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20404 3012 20453 3040
rect 20404 3000 20410 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 20772 3012 21005 3040
rect 20772 3000 20778 3012
rect 20993 3009 21005 3012
rect 21039 3009 21051 3043
rect 20993 3003 21051 3009
rect 9548 2944 12434 2972
rect 14553 2975 14611 2981
rect 9548 2932 9554 2944
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 22066 2972 22094 3080
rect 23845 3043 23903 3049
rect 23845 3009 23857 3043
rect 23891 3040 23903 3043
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23891 3012 23949 3040
rect 23891 3009 23903 3012
rect 23845 3003 23903 3009
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 25130 3000 25136 3052
rect 25188 3000 25194 3052
rect 25225 3043 25283 3049
rect 25225 3009 25237 3043
rect 25271 3040 25283 3043
rect 25317 3043 25375 3049
rect 25317 3040 25329 3043
rect 25271 3012 25329 3040
rect 25271 3009 25283 3012
rect 25225 3003 25283 3009
rect 25317 3009 25329 3012
rect 25363 3009 25375 3043
rect 26804 3040 26832 3148
rect 27264 3148 28908 3176
rect 27264 3040 27292 3148
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 31113 3179 31171 3185
rect 31113 3145 31125 3179
rect 31159 3176 31171 3179
rect 35802 3176 35808 3188
rect 31159 3148 35808 3176
rect 31159 3145 31171 3148
rect 31113 3139 31171 3145
rect 35802 3136 35808 3148
rect 35860 3136 35866 3188
rect 43438 3136 43444 3188
rect 43496 3136 43502 3188
rect 27614 3068 27620 3120
rect 27672 3108 27678 3120
rect 27672 3080 43300 3108
rect 27672 3068 27678 3080
rect 26804 3012 27292 3040
rect 27341 3043 27399 3049
rect 25317 3003 25375 3009
rect 27341 3009 27353 3043
rect 27387 3040 27399 3043
rect 27433 3043 27491 3049
rect 27433 3040 27445 3043
rect 27387 3012 27445 3040
rect 27387 3009 27399 3012
rect 27341 3003 27399 3009
rect 27433 3009 27445 3012
rect 27479 3009 27491 3043
rect 27433 3003 27491 3009
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 28534 3049 28540 3052
rect 27893 3043 27951 3049
rect 27893 3040 27905 3043
rect 27764 3012 27905 3040
rect 27764 3000 27770 3012
rect 27893 3009 27905 3012
rect 27939 3009 27951 3043
rect 27893 3003 27951 3009
rect 28529 3003 28540 3049
rect 28534 3000 28540 3003
rect 28592 3000 28598 3052
rect 30374 3000 30380 3052
rect 30432 3040 30438 3052
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30432 3012 30941 3040
rect 30432 3000 30438 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 42521 3043 42579 3049
rect 42521 3040 42533 3043
rect 37424 3012 42533 3040
rect 37424 3000 37430 3012
rect 42521 3009 42533 3012
rect 42567 3009 42579 3043
rect 42521 3003 42579 3009
rect 42886 3000 42892 3052
rect 42944 3000 42950 3052
rect 43272 3049 43300 3080
rect 43257 3043 43315 3049
rect 43257 3009 43269 3043
rect 43303 3009 43315 3043
rect 43257 3003 43315 3009
rect 43346 2972 43352 2984
rect 14599 2944 21864 2972
rect 22066 2944 43352 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 9456 2876 11713 2904
rect 9456 2864 9462 2876
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 11701 2867 11759 2873
rect 12158 2864 12164 2916
rect 12216 2864 12222 2916
rect 14185 2907 14243 2913
rect 12406 2876 14136 2904
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 12406 2836 12434 2876
rect 9548 2808 12434 2836
rect 14108 2836 14136 2876
rect 14185 2873 14197 2907
rect 14231 2904 14243 2907
rect 14366 2904 14372 2916
rect 14231 2876 14372 2904
rect 14231 2873 14243 2876
rect 14185 2867 14243 2873
rect 14366 2864 14372 2876
rect 14424 2864 14430 2916
rect 17773 2907 17831 2913
rect 17773 2904 17785 2907
rect 16040 2876 17785 2904
rect 16040 2836 16068 2876
rect 17773 2873 17785 2876
rect 17819 2873 17831 2907
rect 17773 2867 17831 2873
rect 20162 2864 20168 2916
rect 20220 2864 20226 2916
rect 20901 2907 20959 2913
rect 20901 2873 20913 2907
rect 20947 2904 20959 2907
rect 21836 2904 21864 2944
rect 43346 2932 43352 2944
rect 43404 2932 43410 2984
rect 40954 2904 40960 2916
rect 20947 2876 21772 2904
rect 21836 2876 27752 2904
rect 20947 2873 20959 2876
rect 20901 2867 20959 2873
rect 14108 2808 16068 2836
rect 9548 2796 9554 2808
rect 18138 2796 18144 2848
rect 18196 2796 18202 2848
rect 20622 2796 20628 2848
rect 20680 2796 20686 2848
rect 21744 2836 21772 2876
rect 24762 2836 24768 2848
rect 21744 2808 24768 2836
rect 24762 2796 24768 2808
rect 24820 2796 24826 2848
rect 25498 2796 25504 2848
rect 25556 2796 25562 2848
rect 27062 2796 27068 2848
rect 27120 2836 27126 2848
rect 27249 2839 27307 2845
rect 27249 2836 27261 2839
rect 27120 2808 27261 2836
rect 27120 2796 27126 2808
rect 27249 2805 27261 2808
rect 27295 2805 27307 2839
rect 27249 2799 27307 2805
rect 27614 2796 27620 2848
rect 27672 2796 27678 2848
rect 27724 2836 27752 2876
rect 28000 2876 40960 2904
rect 28000 2836 28028 2876
rect 40954 2864 40960 2876
rect 41012 2864 41018 2916
rect 27724 2808 28028 2836
rect 28074 2796 28080 2848
rect 28132 2796 28138 2848
rect 28718 2796 28724 2848
rect 28776 2796 28782 2848
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 36538 2836 36544 2848
rect 28960 2808 36544 2836
rect 28960 2796 28966 2808
rect 36538 2796 36544 2808
rect 36596 2796 36602 2848
rect 42705 2839 42763 2845
rect 42705 2805 42717 2839
rect 42751 2836 42763 2839
rect 42978 2836 42984 2848
rect 42751 2808 42984 2836
rect 42751 2805 42763 2808
rect 42705 2799 42763 2805
rect 42978 2796 42984 2808
rect 43036 2796 43042 2848
rect 43070 2796 43076 2848
rect 43128 2796 43134 2848
rect 1104 2746 43884 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 43884 2746
rect 1104 2672 43884 2694
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 20680 2604 42748 2632
rect 20680 2592 20686 2604
rect 18138 2524 18144 2576
rect 18196 2564 18202 2576
rect 18196 2536 41920 2564
rect 18196 2524 18202 2536
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 26142 2496 26148 2508
rect 14424 2468 26148 2496
rect 14424 2456 14430 2468
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 27080 2468 31754 2496
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 27080 2428 27108 2468
rect 12216 2400 27108 2428
rect 31726 2428 31754 2468
rect 41892 2428 41920 2536
rect 42150 2524 42156 2576
rect 42208 2524 42214 2576
rect 41957 2431 42015 2437
rect 41957 2428 41969 2431
rect 31726 2400 41414 2428
rect 41892 2400 41969 2428
rect 12216 2388 12222 2400
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 27062 2360 27068 2372
rect 11020 2332 27068 2360
rect 11020 2320 11026 2332
rect 27062 2320 27068 2332
rect 27120 2320 27126 2372
rect 27154 2320 27160 2372
rect 27212 2360 27218 2372
rect 41386 2360 41414 2400
rect 41957 2397 41969 2400
rect 42003 2397 42015 2431
rect 41957 2391 42015 2397
rect 42521 2431 42579 2437
rect 42521 2397 42533 2431
rect 42567 2397 42579 2431
rect 42720 2428 42748 2604
rect 43438 2524 43444 2576
rect 43496 2524 43502 2576
rect 42889 2431 42947 2437
rect 42889 2428 42901 2431
rect 42720 2400 42901 2428
rect 42521 2391 42579 2397
rect 42889 2397 42901 2400
rect 42935 2397 42947 2431
rect 42889 2391 42947 2397
rect 43257 2431 43315 2437
rect 43257 2397 43269 2431
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 42536 2360 42564 2391
rect 43272 2360 43300 2391
rect 27212 2332 31754 2360
rect 41386 2332 42564 2360
rect 42628 2332 43300 2360
rect 27212 2320 27218 2332
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 30374 2292 30380 2304
rect 5592 2264 30380 2292
rect 5592 2252 5598 2264
rect 30374 2252 30380 2264
rect 30432 2252 30438 2304
rect 31726 2292 31754 2332
rect 42628 2292 42656 2332
rect 31726 2264 42656 2292
rect 42702 2252 42708 2304
rect 42760 2252 42766 2304
rect 43070 2252 43076 2304
rect 43128 2252 43134 2304
rect 1104 2202 43884 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 43884 2202
rect 1104 2128 43884 2150
rect 1118 2048 1124 2100
rect 1176 2088 1182 2100
rect 22830 2088 22836 2100
rect 1176 2060 22836 2088
rect 1176 2048 1182 2060
rect 22830 2048 22836 2060
rect 22888 2048 22894 2100
rect 20346 348 20352 400
rect 20404 388 20410 400
rect 38654 388 38660 400
rect 20404 360 38660 388
rect 20404 348 20410 360
rect 38654 348 38660 360
rect 38712 348 38718 400
rect 13998 280 14004 332
rect 14056 320 14062 332
rect 34698 320 34704 332
rect 14056 292 34704 320
rect 14056 280 14062 292
rect 34698 280 34704 292
rect 34756 280 34762 332
rect 18230 212 18236 264
rect 18288 252 18294 264
rect 40862 252 40868 264
rect 18288 224 40868 252
rect 18288 212 18294 224
rect 40862 212 40868 224
rect 40920 212 40926 264
rect 1302 144 1308 196
rect 1360 144 1366 196
rect 3418 144 3424 196
rect 3476 184 3482 196
rect 26418 184 26424 196
rect 3476 156 26424 184
rect 3476 144 3482 156
rect 26418 144 26424 156
rect 26476 144 26482 196
rect 1320 116 1348 144
rect 1320 88 6914 116
rect 6886 48 6914 88
rect 16206 76 16212 128
rect 16264 116 16270 128
rect 39574 116 39580 128
rect 16264 88 39580 116
rect 16264 76 16270 88
rect 39574 76 39580 88
rect 39632 76 39638 128
rect 31754 48 31760 60
rect 6886 20 31760 48
rect 31754 8 31760 20
rect 31812 8 31818 60
<< via1 >>
rect 7656 11160 7708 11212
rect 24952 11160 25004 11212
rect 11520 11092 11572 11144
rect 27988 11092 28040 11144
rect 14832 11024 14884 11076
rect 29644 11024 29696 11076
rect 19064 10956 19116 11008
rect 29920 10956 29972 11008
rect 18788 10684 18840 10736
rect 23848 10684 23900 10736
rect 17316 9664 17368 9716
rect 24400 9664 24452 9716
rect 10968 9392 11020 9444
rect 18420 9596 18472 9648
rect 17132 9528 17184 9580
rect 22744 9528 22796 9580
rect 14648 9460 14700 9512
rect 19800 9460 19852 9512
rect 19708 9392 19760 9444
rect 24216 9392 24268 9444
rect 41696 9392 41748 9444
rect 10784 9188 10836 9240
rect 16764 9324 16816 9376
rect 34428 9324 34480 9376
rect 19708 9256 19760 9308
rect 20260 9256 20312 9308
rect 28724 9256 28776 9308
rect 36176 9256 36228 9308
rect 17040 9188 17092 9240
rect 32312 9188 32364 9240
rect 32588 9188 32640 9240
rect 38016 9188 38068 9240
rect 24492 9120 24544 9172
rect 30196 9120 30248 9172
rect 32772 9120 32824 9172
rect 38384 9120 38436 9172
rect 18512 9052 18564 9104
rect 24676 9052 24728 9104
rect 10508 8780 10560 8832
rect 16580 8984 16632 9036
rect 18144 8984 18196 9036
rect 27712 9052 27764 9104
rect 34612 9052 34664 9104
rect 35256 9052 35308 9104
rect 35716 9052 35768 9104
rect 36728 9052 36780 9104
rect 37924 9052 37976 9104
rect 38568 9052 38620 9104
rect 25320 8984 25372 9036
rect 41880 8984 41932 9036
rect 18236 8916 18288 8968
rect 22468 8916 22520 8968
rect 26608 8916 26660 8968
rect 34704 8916 34756 8968
rect 34796 8916 34848 8968
rect 38844 8916 38896 8968
rect 29000 8848 29052 8900
rect 41604 8848 41656 8900
rect 16304 8780 16356 8832
rect 16672 8780 16724 8832
rect 17592 8780 17644 8832
rect 29276 8780 29328 8832
rect 35164 8780 35216 8832
rect 35808 8780 35860 8832
rect 37832 8780 37884 8832
rect 41972 8780 42024 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 5908 8576 5960 8628
rect 6460 8576 6512 8628
rect 7012 8576 7064 8628
rect 7288 8576 7340 8628
rect 7564 8576 7616 8628
rect 8116 8576 8168 8628
rect 8668 8576 8720 8628
rect 9496 8576 9548 8628
rect 9772 8576 9824 8628
rect 10324 8576 10376 8628
rect 10600 8576 10652 8628
rect 10876 8576 10928 8628
rect 11428 8576 11480 8628
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 12532 8576 12584 8628
rect 12808 8576 12860 8628
rect 13084 8576 13136 8628
rect 13636 8576 13688 8628
rect 14188 8576 14240 8628
rect 14740 8576 14792 8628
rect 14924 8576 14976 8628
rect 15384 8576 15436 8628
rect 15844 8576 15896 8628
rect 16120 8576 16172 8628
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 17224 8576 17276 8628
rect 17500 8576 17552 8628
rect 18052 8576 18104 8628
rect 18328 8576 18380 8628
rect 18604 8576 18656 8628
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 19432 8576 19484 8628
rect 34060 8576 34112 8628
rect 34336 8576 34388 8628
rect 34980 8576 35032 8628
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 4068 8372 4120 8424
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6552 8440 6604 8492
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7840 8440 7892 8492
rect 7472 8372 7524 8424
rect 7380 8304 7432 8356
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 13452 8508 13504 8560
rect 10508 8440 10560 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 10692 8372 10744 8424
rect 8852 8304 8904 8356
rect 10324 8304 10376 8356
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14924 8440 14976 8492
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 15292 8372 15344 8424
rect 16764 8508 16816 8560
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 17040 8440 17092 8492
rect 18236 8508 18288 8560
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 17868 8372 17920 8424
rect 14924 8304 14976 8356
rect 15016 8304 15068 8356
rect 17408 8304 17460 8356
rect 13636 8236 13688 8288
rect 17684 8236 17736 8288
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 19616 8440 19668 8492
rect 20352 8440 20404 8492
rect 24676 8508 24728 8560
rect 35256 8619 35308 8628
rect 35256 8585 35265 8619
rect 35265 8585 35299 8619
rect 35299 8585 35308 8619
rect 35256 8576 35308 8585
rect 35808 8576 35860 8628
rect 36544 8576 36596 8628
rect 37648 8576 37700 8628
rect 38936 8576 38988 8628
rect 41788 8619 41840 8628
rect 41788 8585 41797 8619
rect 41797 8585 41831 8619
rect 41831 8585 41840 8619
rect 41788 8576 41840 8585
rect 42156 8619 42208 8628
rect 42156 8585 42165 8619
rect 42165 8585 42199 8619
rect 42199 8585 42208 8619
rect 42156 8576 42208 8585
rect 42708 8619 42760 8628
rect 42708 8585 42717 8619
rect 42717 8585 42751 8619
rect 42751 8585 42760 8619
rect 42708 8576 42760 8585
rect 21824 8372 21876 8424
rect 19156 8304 19208 8356
rect 25872 8440 25924 8492
rect 32404 8440 32456 8492
rect 34704 8483 34756 8492
rect 34704 8449 34713 8483
rect 34713 8449 34747 8483
rect 34747 8449 34756 8483
rect 34704 8440 34756 8449
rect 23388 8372 23440 8424
rect 28632 8372 28684 8424
rect 33600 8372 33652 8424
rect 35532 8440 35584 8492
rect 36636 8508 36688 8560
rect 26884 8304 26936 8356
rect 27620 8304 27672 8356
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37648 8483 37700 8492
rect 37648 8449 37657 8483
rect 37657 8449 37691 8483
rect 37691 8449 37700 8483
rect 37648 8440 37700 8449
rect 38016 8483 38068 8492
rect 38016 8449 38025 8483
rect 38025 8449 38059 8483
rect 38059 8449 38068 8483
rect 38016 8440 38068 8449
rect 38200 8440 38252 8492
rect 19248 8236 19300 8288
rect 22284 8236 22336 8288
rect 25504 8236 25556 8288
rect 26424 8236 26476 8288
rect 30472 8236 30524 8288
rect 31760 8236 31812 8288
rect 32128 8236 32180 8288
rect 35808 8236 35860 8288
rect 37096 8372 37148 8424
rect 38384 8483 38436 8492
rect 38384 8449 38393 8483
rect 38393 8449 38427 8483
rect 38427 8449 38436 8483
rect 38384 8440 38436 8449
rect 38660 8440 38712 8492
rect 38844 8440 38896 8492
rect 42064 8508 42116 8560
rect 39948 8440 40000 8492
rect 41604 8483 41656 8492
rect 41604 8449 41613 8483
rect 41613 8449 41647 8483
rect 41647 8449 41656 8483
rect 41604 8440 41656 8449
rect 41696 8440 41748 8492
rect 42156 8440 42208 8492
rect 36728 8347 36780 8356
rect 36728 8313 36737 8347
rect 36737 8313 36771 8347
rect 36771 8313 36780 8347
rect 36728 8304 36780 8313
rect 36820 8304 36872 8356
rect 38568 8304 38620 8356
rect 40316 8372 40368 8424
rect 39396 8304 39448 8356
rect 43076 8347 43128 8356
rect 43076 8313 43085 8347
rect 43085 8313 43119 8347
rect 43119 8313 43128 8347
rect 43076 8304 43128 8313
rect 43444 8347 43496 8356
rect 43444 8313 43453 8347
rect 43453 8313 43487 8347
rect 43487 8313 43496 8347
rect 43444 8304 43496 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 5632 8032 5684 8084
rect 6184 8032 6236 8084
rect 6736 8032 6788 8084
rect 7748 8032 7800 8084
rect 8392 8032 8444 8084
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 10048 8032 10100 8084
rect 11152 8032 11204 8084
rect 11704 8032 11756 8084
rect 12256 8032 12308 8084
rect 12808 8032 12860 8084
rect 13360 8032 13412 8084
rect 13820 8032 13872 8084
rect 14464 8032 14516 8084
rect 15292 8032 15344 8084
rect 15568 8032 15620 8084
rect 16396 8032 16448 8084
rect 16948 8032 17000 8084
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 17776 8032 17828 8084
rect 19616 8032 19668 8084
rect 19800 8032 19852 8084
rect 20720 8075 20772 8084
rect 20720 8041 20729 8075
rect 20729 8041 20763 8075
rect 20763 8041 20772 8075
rect 20720 8032 20772 8041
rect 22100 8075 22152 8084
rect 22100 8041 22109 8075
rect 22109 8041 22143 8075
rect 22143 8041 22152 8075
rect 22100 8032 22152 8041
rect 22468 8075 22520 8084
rect 22468 8041 22477 8075
rect 22477 8041 22511 8075
rect 22511 8041 22520 8075
rect 22468 8032 22520 8041
rect 23848 8075 23900 8084
rect 23848 8041 23857 8075
rect 23857 8041 23891 8075
rect 23891 8041 23900 8075
rect 23848 8032 23900 8041
rect 24216 8075 24268 8084
rect 24216 8041 24225 8075
rect 24225 8041 24259 8075
rect 24259 8041 24268 8075
rect 24216 8032 24268 8041
rect 25872 8032 25924 8084
rect 29000 8075 29052 8084
rect 29000 8041 29009 8075
rect 29009 8041 29043 8075
rect 29043 8041 29052 8075
rect 29000 8032 29052 8041
rect 29184 8032 29236 8084
rect 30748 8032 30800 8084
rect 35992 8032 36044 8084
rect 36268 8032 36320 8084
rect 36820 8075 36872 8084
rect 36820 8041 36829 8075
rect 36829 8041 36863 8075
rect 36863 8041 36872 8075
rect 36820 8032 36872 8041
rect 37372 8032 37424 8084
rect 38476 8032 38528 8084
rect 38844 8032 38896 8084
rect 39580 8032 39632 8084
rect 42340 8075 42392 8084
rect 42340 8041 42349 8075
rect 42349 8041 42383 8075
rect 42383 8041 42392 8075
rect 42340 8032 42392 8041
rect 42616 8032 42668 8084
rect 9956 7964 10008 8016
rect 9404 7896 9456 7948
rect 4344 7828 4396 7880
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 8668 7828 8720 7880
rect 8852 7828 8904 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 9772 7828 9824 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 14832 7964 14884 8016
rect 15752 8007 15804 8016
rect 15752 7973 15761 8007
rect 15761 7973 15795 8007
rect 15795 7973 15804 8007
rect 15752 7964 15804 7973
rect 18696 7964 18748 8016
rect 13636 7828 13688 7880
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 13544 7760 13596 7812
rect 16304 7828 16356 7880
rect 16488 7828 16540 7880
rect 12900 7692 12952 7744
rect 13084 7735 13136 7744
rect 13084 7701 13093 7735
rect 13093 7701 13127 7735
rect 13127 7701 13136 7735
rect 13084 7692 13136 7701
rect 15200 7692 15252 7744
rect 15384 7692 15436 7744
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 18052 7828 18104 7880
rect 22560 7896 22612 7948
rect 19064 7828 19116 7880
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 25228 7896 25280 7948
rect 28632 7939 28684 7948
rect 28632 7905 28641 7939
rect 28641 7905 28675 7939
rect 28675 7905 28684 7939
rect 28632 7896 28684 7905
rect 24400 7871 24452 7880
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 26424 7871 26476 7880
rect 26424 7837 26433 7871
rect 26433 7837 26467 7871
rect 26467 7837 26476 7871
rect 26424 7828 26476 7837
rect 26976 7871 27028 7880
rect 26976 7837 26985 7871
rect 26985 7837 27019 7871
rect 27019 7837 27028 7871
rect 26976 7828 27028 7837
rect 28448 7828 28500 7880
rect 19708 7760 19760 7812
rect 20352 7692 20404 7744
rect 21916 7692 21968 7744
rect 28632 7760 28684 7812
rect 29460 7964 29512 8016
rect 31024 7964 31076 8016
rect 31300 7896 31352 7948
rect 31576 7828 31628 7880
rect 38568 7964 38620 8016
rect 38476 7896 38528 7948
rect 29184 7760 29236 7812
rect 36452 7760 36504 7812
rect 24584 7735 24636 7744
rect 24584 7701 24593 7735
rect 24593 7701 24627 7735
rect 24627 7701 24636 7735
rect 24584 7692 24636 7701
rect 26884 7692 26936 7744
rect 28908 7692 28960 7744
rect 29276 7692 29328 7744
rect 33508 7692 33560 7744
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 37740 7828 37792 7880
rect 37280 7692 37332 7744
rect 38936 7871 38988 7880
rect 38936 7837 38945 7871
rect 38945 7837 38979 7871
rect 38979 7837 38988 7871
rect 38936 7828 38988 7837
rect 39488 7871 39540 7880
rect 39488 7837 39497 7871
rect 39497 7837 39531 7871
rect 39531 7837 39540 7871
rect 39488 7828 39540 7837
rect 40684 7828 40736 7880
rect 38844 7760 38896 7812
rect 42524 7871 42576 7880
rect 42524 7837 42533 7871
rect 42533 7837 42567 7871
rect 42567 7837 42576 7871
rect 42524 7828 42576 7837
rect 43260 7871 43312 7880
rect 43260 7837 43269 7871
rect 43269 7837 43303 7871
rect 43303 7837 43312 7871
rect 43260 7828 43312 7837
rect 39304 7735 39356 7744
rect 39304 7701 39313 7735
rect 39313 7701 39347 7735
rect 39347 7701 39356 7735
rect 39304 7692 39356 7701
rect 43076 7735 43128 7744
rect 43076 7701 43085 7735
rect 43085 7701 43119 7735
rect 43119 7701 43128 7735
rect 43076 7692 43128 7701
rect 43444 7735 43496 7744
rect 43444 7701 43453 7735
rect 43453 7701 43487 7735
rect 43487 7701 43496 7735
rect 43444 7692 43496 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 5172 7488 5224 7540
rect 5908 7531 5960 7540
rect 5908 7497 5917 7531
rect 5917 7497 5951 7531
rect 5951 7497 5960 7531
rect 5908 7488 5960 7497
rect 12440 7488 12492 7540
rect 14372 7488 14424 7540
rect 21824 7531 21876 7540
rect 21824 7497 21833 7531
rect 21833 7497 21867 7531
rect 21867 7497 21876 7531
rect 21824 7488 21876 7497
rect 11612 7420 11664 7472
rect 11704 7352 11756 7404
rect 12440 7352 12492 7404
rect 13084 7420 13136 7472
rect 19524 7420 19576 7472
rect 20260 7420 20312 7472
rect 22284 7420 22336 7472
rect 14832 7352 14884 7404
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 16028 7352 16080 7404
rect 18144 7352 18196 7404
rect 24492 7488 24544 7540
rect 24584 7488 24636 7540
rect 36544 7488 36596 7540
rect 37556 7488 37608 7540
rect 43168 7488 43220 7540
rect 22560 7420 22612 7472
rect 28908 7420 28960 7472
rect 31852 7420 31904 7472
rect 33692 7420 33744 7472
rect 37740 7420 37792 7472
rect 31760 7352 31812 7404
rect 32496 7352 32548 7404
rect 33416 7352 33468 7404
rect 36452 7352 36504 7404
rect 38844 7420 38896 7472
rect 38660 7352 38712 7404
rect 11612 7216 11664 7268
rect 16304 7284 16356 7336
rect 36820 7284 36872 7336
rect 11704 7148 11756 7200
rect 12440 7148 12492 7200
rect 14648 7216 14700 7268
rect 14924 7216 14976 7268
rect 24860 7259 24912 7268
rect 24860 7225 24869 7259
rect 24869 7225 24903 7259
rect 24903 7225 24912 7259
rect 24860 7216 24912 7225
rect 41788 7284 41840 7336
rect 14740 7148 14792 7200
rect 14832 7148 14884 7200
rect 17132 7148 17184 7200
rect 21916 7148 21968 7200
rect 25320 7148 25372 7200
rect 30656 7191 30708 7200
rect 30656 7157 30665 7191
rect 30665 7157 30699 7191
rect 30699 7157 30708 7191
rect 30656 7148 30708 7157
rect 31208 7191 31260 7200
rect 31208 7157 31217 7191
rect 31217 7157 31251 7191
rect 31251 7157 31260 7191
rect 31208 7148 31260 7157
rect 32312 7148 32364 7200
rect 34428 7148 34480 7200
rect 36544 7148 36596 7200
rect 42524 7148 42576 7200
rect 43444 7191 43496 7200
rect 43444 7157 43453 7191
rect 43453 7157 43487 7191
rect 43487 7157 43496 7191
rect 43444 7148 43496 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 6828 6944 6880 6996
rect 7840 6987 7892 6996
rect 7840 6953 7849 6987
rect 7849 6953 7883 6987
rect 7883 6953 7892 6987
rect 7840 6944 7892 6953
rect 8668 6944 8720 6996
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 15200 6944 15252 6996
rect 23388 6944 23440 6996
rect 33784 6944 33836 6996
rect 39488 6944 39540 6996
rect 7380 6876 7432 6928
rect 7656 6876 7708 6928
rect 8852 6876 8904 6928
rect 19248 6876 19300 6928
rect 19340 6876 19392 6928
rect 26884 6876 26936 6928
rect 6460 6740 6512 6792
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 9680 6740 9732 6792
rect 10048 6740 10100 6792
rect 22192 6808 22244 6860
rect 19984 6740 20036 6792
rect 23020 6808 23072 6860
rect 26332 6808 26384 6860
rect 26792 6808 26844 6860
rect 32864 6808 32916 6860
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 18420 6672 18472 6724
rect 24400 6783 24452 6792
rect 24400 6749 24409 6783
rect 24409 6749 24443 6783
rect 24443 6749 24452 6783
rect 24400 6740 24452 6749
rect 32680 6740 32732 6792
rect 36452 6808 36504 6860
rect 40868 6783 40920 6792
rect 40868 6749 40877 6783
rect 40877 6749 40911 6783
rect 40911 6749 40920 6783
rect 40868 6740 40920 6749
rect 42984 6740 43036 6792
rect 15936 6604 15988 6656
rect 16580 6604 16632 6656
rect 29368 6672 29420 6724
rect 24584 6647 24636 6656
rect 24584 6613 24593 6647
rect 24593 6613 24627 6647
rect 24627 6613 24636 6647
rect 24584 6604 24636 6613
rect 37832 6672 37884 6724
rect 33232 6604 33284 6656
rect 38476 6604 38528 6656
rect 43076 6647 43128 6656
rect 43076 6613 43085 6647
rect 43085 6613 43119 6647
rect 43119 6613 43128 6647
rect 43076 6604 43128 6613
rect 43444 6647 43496 6656
rect 43444 6613 43453 6647
rect 43453 6613 43487 6647
rect 43487 6613 43496 6647
rect 43444 6604 43496 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 7656 6400 7708 6452
rect 8760 6400 8812 6452
rect 9588 6400 9640 6452
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 11612 6443 11664 6452
rect 11612 6409 11621 6443
rect 11621 6409 11655 6443
rect 11655 6409 11664 6443
rect 11612 6400 11664 6409
rect 12348 6400 12400 6452
rect 13452 6400 13504 6452
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 20904 6400 20956 6452
rect 24400 6400 24452 6452
rect 24584 6400 24636 6452
rect 1216 6332 1268 6384
rect 8852 6332 8904 6384
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 5632 6196 5684 6248
rect 10048 6332 10100 6384
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 21364 6332 21416 6384
rect 30380 6332 30432 6384
rect 36452 6332 36504 6384
rect 19064 6264 19116 6316
rect 20812 6264 20864 6316
rect 22468 6264 22520 6316
rect 17316 6196 17368 6248
rect 37648 6400 37700 6452
rect 43444 6443 43496 6452
rect 43444 6409 43453 6443
rect 43453 6409 43487 6443
rect 43487 6409 43496 6443
rect 43444 6400 43496 6409
rect 40132 6264 40184 6316
rect 43168 6196 43220 6248
rect 9496 6128 9548 6180
rect 17960 6128 18012 6180
rect 30656 6128 30708 6180
rect 7472 6060 7524 6112
rect 16764 6060 16816 6112
rect 26792 6060 26844 6112
rect 43076 6103 43128 6112
rect 43076 6069 43085 6103
rect 43085 6069 43119 6103
rect 43119 6069 43128 6103
rect 43076 6060 43128 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 6276 5856 6328 5908
rect 6460 5856 6512 5908
rect 9864 5856 9916 5908
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 20720 5856 20772 5908
rect 7196 5720 7248 5772
rect 21732 5720 21784 5772
rect 33600 5788 33652 5840
rect 38568 5788 38620 5840
rect 43444 5831 43496 5840
rect 43444 5797 43453 5831
rect 43453 5797 43487 5831
rect 43487 5797 43496 5831
rect 43444 5788 43496 5797
rect 22376 5720 22428 5772
rect 23296 5720 23348 5772
rect 10876 5652 10928 5704
rect 18604 5652 18656 5704
rect 9680 5584 9732 5636
rect 21640 5652 21692 5704
rect 26424 5695 26476 5704
rect 26424 5661 26433 5695
rect 26433 5661 26467 5695
rect 26467 5661 26476 5695
rect 26424 5652 26476 5661
rect 39580 5695 39632 5704
rect 39580 5661 39589 5695
rect 39589 5661 39623 5695
rect 39623 5661 39632 5695
rect 39580 5652 39632 5661
rect 43352 5652 43404 5704
rect 9128 5516 9180 5568
rect 18512 5516 18564 5568
rect 42984 5584 43036 5636
rect 21824 5559 21876 5568
rect 21824 5525 21833 5559
rect 21833 5525 21867 5559
rect 21867 5525 21876 5559
rect 21824 5516 21876 5525
rect 26608 5559 26660 5568
rect 26608 5525 26617 5559
rect 26617 5525 26651 5559
rect 26651 5525 26660 5559
rect 26608 5516 26660 5525
rect 43076 5559 43128 5568
rect 43076 5525 43085 5559
rect 43085 5525 43119 5559
rect 43119 5525 43128 5559
rect 43076 5516 43128 5525
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 10324 5312 10376 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 17040 5312 17092 5364
rect 28264 5312 28316 5364
rect 38752 5312 38804 5364
rect 43444 5355 43496 5364
rect 43444 5321 43453 5355
rect 43453 5321 43487 5355
rect 43487 5321 43496 5355
rect 43444 5312 43496 5321
rect 8852 5244 8904 5296
rect 13728 5176 13780 5228
rect 23572 5108 23624 5160
rect 17040 5040 17092 5092
rect 20628 5015 20680 5024
rect 20628 4981 20637 5015
rect 20637 4981 20671 5015
rect 20671 4981 20680 5015
rect 20628 4972 20680 4981
rect 30932 5176 30984 5228
rect 40040 5176 40092 5228
rect 32772 5108 32824 5160
rect 42340 5108 42392 5160
rect 40316 5040 40368 5092
rect 28816 4972 28868 5024
rect 43076 5015 43128 5024
rect 43076 4981 43085 5015
rect 43085 4981 43119 5015
rect 43119 4981 43128 5015
rect 43076 4972 43128 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 9404 4768 9456 4820
rect 10968 4768 11020 4820
rect 25136 4768 25188 4820
rect 32404 4811 32456 4820
rect 32404 4777 32413 4811
rect 32413 4777 32447 4811
rect 32447 4777 32456 4811
rect 32404 4768 32456 4777
rect 33692 4811 33744 4820
rect 33692 4777 33701 4811
rect 33701 4777 33735 4811
rect 33735 4777 33744 4811
rect 33692 4768 33744 4777
rect 36636 4811 36688 4820
rect 36636 4777 36645 4811
rect 36645 4777 36679 4811
rect 36679 4777 36688 4811
rect 36636 4768 36688 4777
rect 39948 4768 40000 4820
rect 20628 4700 20680 4752
rect 30380 4700 30432 4752
rect 34796 4700 34848 4752
rect 28080 4632 28132 4684
rect 37280 4700 37332 4752
rect 43444 4743 43496 4752
rect 43444 4709 43453 4743
rect 43453 4709 43487 4743
rect 43487 4709 43496 4743
rect 43444 4700 43496 4709
rect 28540 4564 28592 4616
rect 19340 4496 19392 4548
rect 31760 4564 31812 4616
rect 35164 4564 35216 4616
rect 39396 4632 39448 4684
rect 41512 4564 41564 4616
rect 42892 4607 42944 4616
rect 42892 4573 42901 4607
rect 42901 4573 42935 4607
rect 42935 4573 42944 4607
rect 42892 4564 42944 4573
rect 32772 4496 32824 4548
rect 22836 4471 22888 4480
rect 22836 4437 22845 4471
rect 22845 4437 22879 4471
rect 22879 4437 22888 4471
rect 22836 4428 22888 4437
rect 30380 4428 30432 4480
rect 43076 4471 43128 4480
rect 43076 4437 43085 4471
rect 43085 4437 43119 4471
rect 43119 4437 43128 4471
rect 43076 4428 43128 4437
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 15568 4267 15620 4276
rect 15568 4233 15577 4267
rect 15577 4233 15611 4267
rect 15611 4233 15620 4267
rect 15568 4224 15620 4233
rect 22836 4224 22888 4276
rect 42892 4224 42944 4276
rect 19432 4088 19484 4140
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 24584 4088 24636 4140
rect 37280 4088 37332 4140
rect 20720 4020 20772 4072
rect 18236 3952 18288 4004
rect 21824 3952 21876 4004
rect 30380 4020 30432 4072
rect 40960 4088 41012 4140
rect 43168 4088 43220 4140
rect 43628 4020 43680 4072
rect 23020 3995 23072 4004
rect 23020 3961 23029 3995
rect 23029 3961 23063 3995
rect 23063 3961 23072 3995
rect 23020 3952 23072 3961
rect 25872 3995 25924 4004
rect 25872 3961 25881 3995
rect 25881 3961 25915 3995
rect 25915 3961 25924 3995
rect 25872 3952 25924 3961
rect 38936 3952 38988 4004
rect 40684 3995 40736 4004
rect 40684 3961 40693 3995
rect 40693 3961 40727 3995
rect 40727 3961 40736 3995
rect 40684 3952 40736 3961
rect 43444 3995 43496 4004
rect 43444 3961 43453 3995
rect 43453 3961 43487 3995
rect 43487 3961 43496 3995
rect 43444 3952 43496 3961
rect 13544 3884 13596 3936
rect 21916 3884 21968 3936
rect 22744 3884 22796 3936
rect 26700 3884 26752 3936
rect 43076 3927 43128 3936
rect 43076 3893 43085 3927
rect 43085 3893 43119 3927
rect 43119 3893 43128 3927
rect 43076 3884 43128 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 18512 3723 18564 3732
rect 18512 3689 18521 3723
rect 18521 3689 18555 3723
rect 18555 3689 18564 3723
rect 18512 3680 18564 3689
rect 19984 3680 20036 3732
rect 22744 3680 22796 3732
rect 9864 3612 9916 3664
rect 7656 3544 7708 3596
rect 18236 3544 18288 3596
rect 15384 3408 15436 3460
rect 21916 3544 21968 3596
rect 35808 3680 35860 3732
rect 36544 3680 36596 3732
rect 42340 3612 42392 3664
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 25412 3544 25464 3596
rect 25504 3544 25556 3596
rect 40132 3544 40184 3596
rect 9588 3340 9640 3392
rect 14004 3340 14056 3392
rect 34704 3519 34756 3528
rect 34704 3485 34713 3519
rect 34713 3485 34747 3519
rect 34747 3485 34756 3519
rect 34704 3476 34756 3485
rect 43444 3655 43496 3664
rect 43444 3621 43453 3655
rect 43453 3621 43487 3655
rect 43487 3621 43496 3655
rect 43444 3612 43496 3621
rect 25412 3340 25464 3392
rect 40040 3340 40092 3392
rect 43076 3383 43128 3392
rect 43076 3349 43085 3383
rect 43085 3349 43119 3383
rect 43119 3349 43128 3383
rect 43076 3340 43128 3349
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 7840 3136 7892 3188
rect 23296 3136 23348 3188
rect 23388 3136 23440 3188
rect 14004 3111 14056 3120
rect 14004 3077 14013 3111
rect 14013 3077 14047 3111
rect 14047 3077 14056 3111
rect 14004 3068 14056 3077
rect 16488 3068 16540 3120
rect 7012 3000 7064 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 9496 2932 9548 2984
rect 19984 3043 20036 3052
rect 19984 3009 19993 3043
rect 19993 3009 20027 3043
rect 20027 3009 20036 3043
rect 19984 3000 20036 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 25136 3043 25188 3052
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 28908 3136 28960 3188
rect 35808 3136 35860 3188
rect 43444 3179 43496 3188
rect 43444 3145 43453 3179
rect 43453 3145 43487 3179
rect 43487 3145 43496 3179
rect 43444 3136 43496 3145
rect 27620 3068 27672 3120
rect 27712 3043 27764 3052
rect 27712 3009 27721 3043
rect 27721 3009 27755 3043
rect 27755 3009 27764 3043
rect 27712 3000 27764 3009
rect 28540 3043 28592 3052
rect 28540 3009 28541 3043
rect 28541 3009 28575 3043
rect 28575 3009 28592 3043
rect 28540 3000 28592 3009
rect 30380 3000 30432 3052
rect 37372 3000 37424 3052
rect 42892 3043 42944 3052
rect 42892 3009 42901 3043
rect 42901 3009 42935 3043
rect 42935 3009 42944 3043
rect 42892 3000 42944 3009
rect 9404 2864 9456 2916
rect 12164 2907 12216 2916
rect 12164 2873 12173 2907
rect 12173 2873 12207 2907
rect 12207 2873 12216 2907
rect 12164 2864 12216 2873
rect 9496 2796 9548 2848
rect 14372 2864 14424 2916
rect 20168 2907 20220 2916
rect 20168 2873 20177 2907
rect 20177 2873 20211 2907
rect 20211 2873 20220 2907
rect 20168 2864 20220 2873
rect 43352 2932 43404 2984
rect 18144 2839 18196 2848
rect 18144 2805 18153 2839
rect 18153 2805 18187 2839
rect 18187 2805 18196 2839
rect 18144 2796 18196 2805
rect 20628 2839 20680 2848
rect 20628 2805 20637 2839
rect 20637 2805 20671 2839
rect 20671 2805 20680 2839
rect 20628 2796 20680 2805
rect 24768 2796 24820 2848
rect 25504 2839 25556 2848
rect 25504 2805 25513 2839
rect 25513 2805 25547 2839
rect 25547 2805 25556 2839
rect 25504 2796 25556 2805
rect 27068 2796 27120 2848
rect 27620 2839 27672 2848
rect 27620 2805 27629 2839
rect 27629 2805 27663 2839
rect 27663 2805 27672 2839
rect 27620 2796 27672 2805
rect 40960 2864 41012 2916
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 28724 2839 28776 2848
rect 28724 2805 28733 2839
rect 28733 2805 28767 2839
rect 28767 2805 28776 2839
rect 28724 2796 28776 2805
rect 28908 2796 28960 2848
rect 36544 2796 36596 2848
rect 42984 2796 43036 2848
rect 43076 2839 43128 2848
rect 43076 2805 43085 2839
rect 43085 2805 43119 2839
rect 43119 2805 43128 2839
rect 43076 2796 43128 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 20628 2592 20680 2644
rect 18144 2524 18196 2576
rect 14372 2456 14424 2508
rect 26148 2456 26200 2508
rect 12164 2388 12216 2440
rect 42156 2567 42208 2576
rect 42156 2533 42165 2567
rect 42165 2533 42199 2567
rect 42199 2533 42208 2567
rect 42156 2524 42208 2533
rect 10968 2320 11020 2372
rect 27068 2320 27120 2372
rect 27160 2320 27212 2372
rect 43444 2567 43496 2576
rect 43444 2533 43453 2567
rect 43453 2533 43487 2567
rect 43487 2533 43496 2567
rect 43444 2524 43496 2533
rect 5540 2252 5592 2304
rect 30380 2252 30432 2304
rect 42708 2295 42760 2304
rect 42708 2261 42717 2295
rect 42717 2261 42751 2295
rect 42751 2261 42760 2295
rect 42708 2252 42760 2261
rect 43076 2295 43128 2304
rect 43076 2261 43085 2295
rect 43085 2261 43119 2295
rect 43119 2261 43128 2295
rect 43076 2252 43128 2261
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 1124 2048 1176 2100
rect 22836 2048 22888 2100
rect 20352 348 20404 400
rect 38660 348 38712 400
rect 14004 280 14056 332
rect 34704 280 34756 332
rect 18236 212 18288 264
rect 40868 212 40920 264
rect 1308 144 1360 196
rect 3424 144 3476 196
rect 26424 144 26476 196
rect 16212 76 16264 128
rect 39580 76 39632 128
rect 31760 8 31812 60
<< metal2 >>
rect 5354 11194 5410 11250
rect 5630 11194 5686 11250
rect 5906 11194 5962 11250
rect 6182 11194 6238 11250
rect 6458 11194 6514 11250
rect 6734 11194 6790 11250
rect 7010 11194 7066 11250
rect 7286 11194 7342 11250
rect 7562 11194 7618 11250
rect 7656 11212 7708 11218
rect 1306 9480 1362 9489
rect 1306 9415 1362 9424
rect 1214 7984 1270 7993
rect 1214 7919 1270 7928
rect 1122 7712 1178 7721
rect 1122 7647 1178 7656
rect 1136 2106 1164 7647
rect 1228 6390 1256 7919
rect 1320 7449 1348 9415
rect 2870 9208 2926 9217
rect 2870 9143 2926 9152
rect 2884 8809 2912 9143
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 5368 8634 5396 11194
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 3422 7848 3478 7857
rect 3422 7783 3478 7792
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 1306 7440 1362 7449
rect 1306 7375 1362 7384
rect 3436 7313 3464 7783
rect 3422 7304 3478 7313
rect 3422 7239 3478 7248
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1766 6760 1822 6769
rect 1766 6695 1822 6704
rect 1216 6384 1268 6390
rect 1216 6326 1268 6332
rect 1780 6089 1808 6695
rect 4080 6662 4108 8366
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7546 4384 7822
rect 5184 7546 5212 8434
rect 5644 8090 5672 11194
rect 5920 8634 5948 11194
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5920 7546 5948 8434
rect 6196 8090 6224 11194
rect 6472 8634 6500 11194
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 4068 6656 4120 6662
rect 2870 6624 2926 6633
rect 4068 6598 4120 6604
rect 2870 6559 2926 6568
rect 1766 6080 1822 6089
rect 1766 6015 1822 6024
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2884 5681 2912 6559
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 2870 5672 2926 5681
rect 2870 5607 2926 5616
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2686 5264 2742 5273
rect 2686 5199 2742 5208
rect 2700 5001 2728 5199
rect 2686 4992 2742 5001
rect 1950 4924 2258 4933
rect 2686 4927 2742 4936
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 5538 2952 5594 2961
rect 5538 2887 5594 2896
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 5552 2310 5580 2887
rect 5540 2304 5592 2310
rect 2870 2272 2926 2281
rect 5540 2246 5592 2252
rect 2870 2207 2926 2216
rect 1124 2100 1176 2106
rect 1124 2042 1176 2048
rect 2884 1873 2912 2207
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 5644 2122 5672 6190
rect 6288 5914 6316 7822
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 5914 6500 6734
rect 6564 6662 6592 8434
rect 6748 8090 6776 11194
rect 7024 8634 7052 11194
rect 7300 8634 7328 11194
rect 7576 8634 7604 11194
rect 7838 11194 7894 11250
rect 8114 11194 8170 11250
rect 8390 11194 8446 11250
rect 8666 11194 8722 11250
rect 8942 11194 8998 11250
rect 9218 11194 9274 11250
rect 9494 11194 9550 11250
rect 9770 11194 9826 11250
rect 10046 11194 10102 11250
rect 10322 11194 10378 11250
rect 10598 11194 10654 11250
rect 10874 11194 10930 11250
rect 11150 11194 11206 11250
rect 11426 11194 11482 11250
rect 11702 11194 11758 11250
rect 11978 11194 12034 11250
rect 12254 11194 12310 11250
rect 12530 11194 12586 11250
rect 12806 11194 12862 11250
rect 13082 11194 13138 11250
rect 13358 11194 13414 11250
rect 13634 11194 13690 11250
rect 13910 11194 13966 11250
rect 14186 11194 14242 11250
rect 14462 11194 14518 11250
rect 14738 11194 14794 11250
rect 15014 11194 15070 11250
rect 15290 11194 15346 11250
rect 15566 11194 15622 11250
rect 15842 11194 15898 11250
rect 16118 11194 16174 11250
rect 16394 11194 16450 11250
rect 16670 11194 16726 11250
rect 16946 11194 17002 11250
rect 17222 11194 17278 11250
rect 17498 11194 17554 11250
rect 17774 11194 17830 11250
rect 18050 11194 18106 11250
rect 18326 11194 18382 11250
rect 18602 11194 18658 11250
rect 18878 11194 18934 11250
rect 19154 11194 19210 11250
rect 19430 11194 19486 11250
rect 19706 11194 19762 11250
rect 19982 11194 20038 11250
rect 20258 11194 20314 11250
rect 20534 11194 20590 11250
rect 20810 11194 20866 11250
rect 21086 11194 21142 11250
rect 21362 11194 21418 11250
rect 21638 11194 21694 11250
rect 21914 11194 21970 11250
rect 22190 11194 22246 11250
rect 22466 11194 22522 11250
rect 22742 11194 22798 11250
rect 23018 11194 23074 11250
rect 23294 11194 23350 11250
rect 23570 11194 23626 11250
rect 23846 11194 23902 11250
rect 24122 11194 24178 11250
rect 24398 11194 24454 11250
rect 24674 11194 24730 11250
rect 24950 11212 25006 11250
rect 24950 11194 24952 11212
rect 7656 11154 7708 11160
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7002 6868 7822
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7024 6662 7052 8434
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7392 6934 7420 8298
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 7208 5778 7236 6734
rect 7484 6118 7512 8366
rect 7668 8072 7696 11154
rect 7852 8616 7880 11194
rect 8128 8634 8156 11194
rect 7760 8588 7880 8616
rect 8116 8628 8168 8634
rect 7760 8090 7788 8588
rect 8116 8570 8168 8576
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7576 8044 7696 8072
rect 7748 8084 7800 8090
rect 7576 7868 7604 8044
rect 7748 8026 7800 8032
rect 7576 7840 7788 7868
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 6458 7696 6870
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7760 6322 7788 7840
rect 7852 7002 7880 8434
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8404 8090 8432 11194
rect 8680 8634 8708 11194
rect 8956 8820 8984 11194
rect 9232 9466 9260 11194
rect 9232 9438 9444 9466
rect 8864 8792 8984 8820
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8680 7002 8708 7822
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8772 6458 8800 8434
rect 8864 8362 8892 8792
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 9416 8090 9444 9438
rect 9508 8634 9536 11194
rect 9784 8634 9812 11194
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 6934 8892 7822
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 8864 5302 8892 6326
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5574 9168 6258
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 8852 5296 8904 5302
rect 7838 5264 7894 5273
rect 8852 5238 8904 5244
rect 7838 5199 7894 5208
rect 7010 4992 7066 5001
rect 7010 4927 7066 4936
rect 7024 3058 7052 4927
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 5552 2094 5672 2122
rect 2870 1864 2926 1873
rect 2870 1799 2926 1808
rect 1308 196 1360 202
rect 1308 138 1360 144
rect 3424 196 3476 202
rect 3424 138 3476 144
rect 1320 56 1348 138
rect 3436 56 3464 138
rect 5552 56 5580 2094
rect 7668 56 7696 3538
rect 7852 3194 7880 5199
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 9416 4826 9444 7890
rect 9508 6186 9536 8434
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9600 6458 9628 7822
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9692 5642 9720 6734
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9494 4040 9550 4049
rect 9494 3975 9550 3984
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 9508 2990 9536 3975
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 1465 9444 2858
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9508 1737 9536 2790
rect 9600 2553 9628 3334
rect 9586 2544 9642 2553
rect 9586 2479 9642 2488
rect 9494 1728 9550 1737
rect 9494 1663 9550 1672
rect 9402 1456 9458 1465
rect 9402 1391 9458 1400
rect 9784 56 9812 7822
rect 9876 5914 9904 8434
rect 10060 8090 10088 11194
rect 10138 10840 10194 10849
rect 10138 10775 10194 10784
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 9956 8016 10008 8022
rect 9954 7984 9956 7993
rect 10008 7984 10010 7993
rect 9954 7919 10010 7928
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6390 10088 6734
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10152 6322 10180 10775
rect 10336 8634 10364 11194
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10520 8498 10548 8774
rect 10612 8634 10640 11194
rect 10784 9240 10836 9246
rect 10784 9182 10836 9188
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10796 8514 10824 9182
rect 10888 8634 10916 11194
rect 10968 9444 11020 9450
rect 10968 9386 11020 9392
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10508 8492 10560 8498
rect 10796 8486 10916 8514
rect 10980 8498 11008 9386
rect 10508 8434 10560 8440
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10336 5370 10364 8298
rect 10704 6458 10732 8366
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10506 6352 10562 6361
rect 10506 6287 10508 6296
rect 10560 6287 10562 6296
rect 10508 6258 10560 6264
rect 10888 5710 10916 8486
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11164 8090 11192 11194
rect 11440 8634 11468 11194
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11532 6914 11560 11086
rect 11716 8090 11744 11194
rect 11992 8634 12020 11194
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12268 8090 12296 11194
rect 12544 8634 12572 11194
rect 12820 8634 12848 11194
rect 13096 8634 13124 11194
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11624 7274 11652 7414
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11716 7206 11744 7346
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11532 6886 11652 6914
rect 10966 6760 11022 6769
rect 10966 6695 11022 6704
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10980 4826 11008 6695
rect 11624 6458 11652 6886
rect 12360 6458 12388 7822
rect 12452 7546 12480 8434
rect 12820 8090 12848 8434
rect 13372 8090 13400 11194
rect 13648 8634 13676 11194
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 7206 12480 7346
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12912 5370 12940 7686
rect 13096 7478 13124 7686
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13372 7002 13400 7375
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13464 6458 13492 8502
rect 13924 8378 13952 11194
rect 14200 8634 14228 11194
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 13832 8350 13952 8378
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7886 13676 8230
rect 13832 8090 13860 8350
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14476 8090 14504 11194
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14660 8498 14688 9454
rect 14752 8634 14780 11194
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14738 8120 14794 8129
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14464 8084 14516 8090
rect 14738 8055 14794 8064
rect 14464 8026 14516 8032
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 12900 5364 12952 5370
rect 12900 5306 12952 5312
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 13556 3942 13584 7754
rect 14384 7546 14412 7822
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14660 7177 14688 7210
rect 14752 7206 14780 8055
rect 14844 8022 14872 11018
rect 15028 8922 15056 11194
rect 14936 8894 15056 8922
rect 15304 8922 15332 11194
rect 15304 8894 15424 8922
rect 14936 8634 14964 8894
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 8894
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14936 8498 15056 8514
rect 14924 8492 15056 8498
rect 14976 8486 15056 8492
rect 14924 8434 14976 8440
rect 15028 8362 15056 8486
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14844 7206 14872 7346
rect 14936 7274 14964 8298
rect 15304 8090 15332 8366
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15396 7857 15424 8434
rect 15580 8090 15608 11194
rect 15750 10568 15806 10577
rect 15750 10503 15806 10512
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15764 8022 15792 10503
rect 15856 8634 15884 11194
rect 16026 10976 16082 10985
rect 16026 10911 16082 10920
rect 15934 9752 15990 9761
rect 15934 9687 15990 9696
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15198 7848 15254 7857
rect 15198 7783 15254 7792
rect 15382 7848 15438 7857
rect 15382 7783 15438 7792
rect 15212 7750 15240 7783
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14740 7200 14792 7206
rect 14646 7168 14702 7177
rect 14740 7142 14792 7148
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 13950 7100 14258 7109
rect 14646 7103 14702 7112
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 15212 7002 15240 7346
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13726 5672 13782 5681
rect 13726 5607 13782 5616
rect 13740 5234 13768 5607
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9876 3058 9904 3606
rect 15396 3466 15424 7686
rect 15948 6662 15976 9687
rect 16040 7410 16068 10911
rect 16132 8634 16160 11194
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 8634 16344 8774
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16132 6769 16160 8434
rect 16408 8090 16436 11194
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16486 8936 16542 8945
rect 16486 8871 16542 8880
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16500 7886 16528 8871
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16316 7342 16344 7822
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16118 6760 16174 6769
rect 16118 6695 16174 6704
rect 16592 6662 16620 8978
rect 16684 8838 16712 11194
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16776 8566 16804 9318
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16960 8090 16988 11194
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17040 9240 17092 9246
rect 17040 9182 17092 9188
rect 17052 8498 17080 9182
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 15566 6216 15622 6225
rect 15566 6151 15622 6160
rect 15580 4282 15608 6151
rect 16776 6118 16804 7822
rect 17144 7206 17172 9522
rect 17236 8634 17264 11194
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17328 6254 17356 9658
rect 17512 8634 17540 11194
rect 17682 10704 17738 10713
rect 17682 10639 17738 10648
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17604 8498 17632 8774
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17420 8090 17448 8298
rect 17696 8294 17724 10639
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17788 8090 17816 11194
rect 18064 8634 18092 11194
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17868 8424 17920 8430
rect 17920 8384 18000 8412
rect 17868 8366 17920 8372
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17972 6186 18000 8384
rect 18050 8256 18106 8265
rect 18050 8191 18106 8200
rect 18064 7886 18092 8191
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18156 7410 18184 8978
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8566 18276 8910
rect 18340 8634 18368 11194
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18432 6730 18460 9590
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16486 5808 16542 5817
rect 16486 5743 16542 5752
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 14016 3126 14044 3334
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 16500 3126 16528 5743
rect 18524 5574 18552 9046
rect 18616 8634 18644 11194
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18708 8022 18736 8434
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18602 6896 18658 6905
rect 18602 6831 18658 6840
rect 18616 5914 18644 6831
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18604 5704 18656 5710
rect 18800 5692 18828 10678
rect 18892 8634 18920 11194
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 19076 7886 19104 10950
rect 19168 8362 19196 11194
rect 19444 8634 19472 11194
rect 19720 9450 19748 11194
rect 19996 9761 20024 11194
rect 19982 9752 20038 9761
rect 19982 9687 20038 9696
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19708 9308 19760 9314
rect 19708 9250 19760 9256
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19260 7018 19288 8230
rect 19536 7478 19564 8434
rect 19628 8090 19656 8434
rect 19720 8129 19748 9250
rect 19706 8120 19762 8129
rect 19616 8084 19668 8090
rect 19812 8090 19840 9454
rect 20272 9314 20300 11194
rect 20260 9308 20312 9314
rect 20260 9250 20312 9256
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 19706 8055 19762 8064
rect 19800 8084 19852 8090
rect 19616 8026 19668 8032
rect 19800 8026 19852 8032
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19524 7472 19576 7478
rect 19720 7449 19748 7754
rect 19798 7712 19854 7721
rect 19798 7647 19854 7656
rect 19524 7414 19576 7420
rect 19706 7440 19762 7449
rect 19706 7375 19762 7384
rect 19812 7177 19840 7647
rect 20272 7478 20300 7822
rect 20364 7750 20392 8434
rect 20442 8120 20498 8129
rect 20442 8055 20498 8064
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20456 7585 20484 8055
rect 20548 7721 20576 11194
rect 20718 9344 20774 9353
rect 20718 9279 20774 9288
rect 20732 8090 20760 9279
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20534 7712 20590 7721
rect 20534 7647 20590 7656
rect 20442 7576 20498 7585
rect 20442 7511 20498 7520
rect 20260 7472 20312 7478
rect 20260 7414 20312 7420
rect 19798 7168 19854 7177
rect 19798 7103 19854 7112
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 19260 6990 19380 7018
rect 19352 6934 19380 6990
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19982 6896 20038 6905
rect 19260 6458 19288 6870
rect 19982 6831 20038 6840
rect 19996 6798 20024 6831
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 20824 6322 20852 11194
rect 21100 8922 21128 11194
rect 21376 9058 21404 11194
rect 21376 9030 21496 9058
rect 21100 8894 21404 8922
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 19076 6225 19104 6258
rect 19062 6216 19118 6225
rect 19062 6151 19118 6160
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 18656 5664 18828 5692
rect 18604 5646 18656 5652
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17052 5098 17080 5306
rect 17222 5128 17278 5137
rect 17040 5092 17092 5098
rect 17222 5063 17278 5072
rect 18510 5128 18566 5137
rect 18510 5063 18566 5072
rect 17040 5034 17092 5040
rect 17236 3738 17264 5063
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 18248 3602 18276 3946
rect 18524 3738 18552 5063
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20640 4758 20668 4966
rect 20628 4752 20680 4758
rect 19430 4720 19486 4729
rect 20628 4694 20680 4700
rect 19430 4655 19486 4664
rect 19338 4584 19394 4593
rect 19338 4519 19340 4528
rect 19392 4519 19394 4528
rect 19340 4490 19392 4496
rect 19444 4146 19472 4655
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 20732 4078 20760 5850
rect 20916 4185 20944 6394
rect 21376 6390 21404 8894
rect 21468 6905 21496 9030
rect 21454 6896 21510 6905
rect 21454 6831 21510 6840
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21652 5710 21680 11194
rect 21928 8514 21956 11194
rect 22098 9616 22154 9625
rect 22098 9551 22154 9560
rect 21744 8486 21956 8514
rect 21744 5778 21772 8486
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 7546 21864 8366
rect 22112 8090 22140 9551
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21928 7206 21956 7686
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 22204 6866 22232 11194
rect 22480 9058 22508 11194
rect 22756 9586 22784 11194
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22388 9030 22508 9058
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22296 7478 22324 8230
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22388 5778 22416 9030
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22480 8090 22508 8910
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22572 7478 22600 7890
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 23032 6866 23060 11194
rect 23110 6896 23166 6905
rect 23020 6860 23072 6866
rect 23110 6831 23166 6840
rect 23020 6802 23072 6808
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 21732 5772 21784 5778
rect 21732 5714 21784 5720
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20902 4176 20958 4185
rect 20902 4111 20958 4120
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 21836 4010 21864 5510
rect 21824 4004 21876 4010
rect 21824 3946 21876 3952
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 14004 3120 14056 3126
rect 10966 3088 11022 3097
rect 9864 3052 9916 3058
rect 14004 3062 14056 3068
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 19996 3058 20024 3674
rect 21928 3602 21956 3878
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 10966 3023 11022 3032
rect 19984 3052 20036 3058
rect 9864 2994 9916 3000
rect 10980 2378 11008 3023
rect 19984 2994 20036 3000
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20166 2952 20222 2961
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 14372 2916 14424 2922
rect 20166 2887 20168 2896
rect 14372 2858 14424 2864
rect 20220 2887 20222 2896
rect 20168 2858 20220 2864
rect 12176 2446 12204 2858
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14384 2514 14412 2858
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18156 2582 18184 2790
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 12164 2440 12216 2446
rect 11886 2408 11942 2417
rect 10968 2372 11020 2378
rect 12164 2382 12216 2388
rect 11886 2343 11942 2352
rect 10968 2314 11020 2320
rect 11900 56 11928 2343
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 20364 1873 20392 2994
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 2650 20668 2790
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20732 2009 20760 2994
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 20718 2000 20774 2009
rect 20718 1935 20774 1944
rect 20350 1864 20406 1873
rect 20350 1799 20406 1808
rect 20352 400 20404 406
rect 20352 342 20404 348
rect 14004 332 14056 338
rect 14004 274 14056 280
rect 14016 56 14044 274
rect 18236 264 18288 270
rect 16132 190 16252 218
rect 18236 206 18288 212
rect 16132 56 16160 190
rect 16224 134 16252 190
rect 16212 128 16264 134
rect 16212 70 16264 76
rect 18248 56 18276 206
rect 20364 56 20392 342
rect 22480 56 22508 6258
rect 23018 5264 23074 5273
rect 23018 5199 23074 5208
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22848 4282 22876 4422
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22756 3738 22784 3878
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22848 2106 22876 4082
rect 23032 4010 23060 5199
rect 23020 4004 23072 4010
rect 23020 3946 23072 3952
rect 23124 3534 23152 6831
rect 23308 6225 23336 11194
rect 23386 9888 23442 9897
rect 23386 9823 23442 9832
rect 23400 8430 23428 9823
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23386 7168 23442 7177
rect 23386 7103 23442 7112
rect 23400 7002 23428 7103
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23294 6216 23350 6225
rect 23294 6151 23350 6160
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23308 3194 23336 5714
rect 23584 5166 23612 11194
rect 23860 10742 23888 11194
rect 24136 10849 24164 11194
rect 24122 10840 24178 10849
rect 24122 10775 24178 10784
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 24412 9722 24440 11194
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24216 9444 24268 9450
rect 24216 9386 24268 9392
rect 23846 9208 23902 9217
rect 23846 9143 23902 9152
rect 23860 8090 23888 9143
rect 24228 8090 24256 9386
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24398 9072 24454 9081
rect 24398 9007 24454 9016
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 24412 7886 24440 9007
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24504 7546 24532 9114
rect 24688 9110 24716 11194
rect 25004 11194 25006 11212
rect 25226 11194 25282 11250
rect 25502 11194 25558 11250
rect 25778 11194 25834 11250
rect 26054 11194 26110 11250
rect 26330 11194 26386 11250
rect 26606 11194 26662 11250
rect 26882 11194 26938 11250
rect 27158 11194 27214 11250
rect 27434 11194 27490 11250
rect 27710 11194 27766 11250
rect 27986 11194 28042 11250
rect 28262 11194 28318 11250
rect 28538 11194 28594 11250
rect 28814 11194 28870 11250
rect 29090 11194 29146 11250
rect 29366 11194 29422 11250
rect 29642 11194 29698 11250
rect 29918 11194 29974 11250
rect 30194 11194 30250 11250
rect 30470 11194 30526 11250
rect 30746 11194 30802 11250
rect 31022 11194 31078 11250
rect 31298 11194 31354 11250
rect 31574 11194 31630 11250
rect 31850 11194 31906 11250
rect 32126 11194 32182 11250
rect 32402 11194 32458 11250
rect 32678 11194 32734 11250
rect 32954 11194 33010 11250
rect 33230 11194 33286 11250
rect 33506 11194 33562 11250
rect 33782 11194 33838 11250
rect 34058 11194 34114 11250
rect 34334 11194 34390 11250
rect 34610 11194 34666 11250
rect 34886 11194 34942 11250
rect 35162 11194 35218 11250
rect 35438 11194 35494 11250
rect 35714 11194 35770 11250
rect 35990 11194 36046 11250
rect 36266 11194 36322 11250
rect 36542 11194 36598 11250
rect 36818 11194 36874 11250
rect 37094 11194 37150 11250
rect 37370 11194 37426 11250
rect 37646 11194 37702 11250
rect 37922 11194 37978 11250
rect 38198 11194 38254 11250
rect 38474 11194 38530 11250
rect 38750 11194 38806 11250
rect 39026 11194 39082 11250
rect 39302 11194 39358 11250
rect 39578 11194 39634 11250
rect 24952 11154 25004 11160
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24688 8129 24716 8502
rect 24674 8120 24730 8129
rect 24674 8055 24730 8064
rect 25240 7954 25268 11194
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 24596 7546 24624 7686
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24858 7304 24914 7313
rect 24858 7239 24860 7248
rect 24912 7239 24914 7248
rect 24860 7210 24912 7216
rect 25332 7206 25360 8978
rect 25516 8294 25544 11194
rect 25792 8945 25820 11194
rect 25778 8936 25834 8945
rect 25778 8871 25834 8880
rect 26068 8786 26096 11194
rect 26344 10985 26372 11194
rect 26330 10976 26386 10985
rect 26330 10911 26386 10920
rect 26620 10577 26648 11194
rect 26606 10568 26662 10577
rect 26606 10503 26662 10512
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 25792 8758 26096 8786
rect 25504 8288 25556 8294
rect 25792 8265 25820 8758
rect 26330 8528 26386 8537
rect 25872 8492 25924 8498
rect 26330 8463 26386 8472
rect 25872 8434 25924 8440
rect 25504 8230 25556 8236
rect 25778 8256 25834 8265
rect 25778 8191 25834 8200
rect 25884 8090 25912 8434
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26344 6866 26372 8463
rect 26424 8288 26476 8294
rect 26424 8230 26476 8236
rect 26436 7886 26464 8230
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24412 6458 24440 6734
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24596 6458 24624 6598
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24584 6452 24636 6458
rect 24584 6394 24636 6400
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26424 5704 26476 5710
rect 26424 5646 26476 5652
rect 23572 5160 23624 5166
rect 23572 5102 23624 5108
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 23386 3496 23442 3505
rect 23386 3431 23442 3440
rect 23400 3194 23428 3431
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 24596 56 24624 4082
rect 24858 3632 24914 3641
rect 24858 3567 24860 3576
rect 24912 3567 24914 3576
rect 24860 3538 24912 3544
rect 24766 3496 24822 3505
rect 24766 3431 24822 3440
rect 24780 2854 24808 3431
rect 25148 3058 25176 4762
rect 25870 4040 25926 4049
rect 25870 3975 25872 3984
rect 25924 3975 25926 3984
rect 25872 3946 25924 3952
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25424 3398 25452 3538
rect 25412 3392 25464 3398
rect 25412 3334 25464 3340
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 25516 2854 25544 3538
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26146 2544 26202 2553
rect 26146 2479 26148 2488
rect 26200 2479 26202 2488
rect 26148 2450 26200 2456
rect 26436 202 26464 5646
rect 26620 5574 26648 8910
rect 26896 8362 26924 11194
rect 27172 9058 27200 11194
rect 27448 10713 27476 11194
rect 27434 10704 27490 10713
rect 27434 10639 27490 10648
rect 27618 9480 27674 9489
rect 27618 9415 27674 9424
rect 27172 9030 27384 9058
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 26974 8120 27030 8129
rect 26974 8055 27030 8064
rect 26988 7886 27016 8055
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26896 6934 26924 7686
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27356 7313 27384 9030
rect 27632 8514 27660 9415
rect 27724 9110 27752 11194
rect 28000 11150 28028 11194
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 27632 8486 27752 8514
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27632 7993 27660 8298
rect 27618 7984 27674 7993
rect 27618 7919 27674 7928
rect 27342 7304 27398 7313
rect 27342 7239 27398 7248
rect 26884 6928 26936 6934
rect 26884 6870 26936 6876
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26804 6118 26832 6802
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 26792 6112 26844 6118
rect 26792 6054 26844 6060
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26424 196 26476 202
rect 26424 138 26476 144
rect 26712 56 26740 3878
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27620 3120 27672 3126
rect 27620 3062 27672 3068
rect 27632 2854 27660 3062
rect 27724 3058 27752 8486
rect 28276 5370 28304 11194
rect 28446 7984 28502 7993
rect 28446 7919 28502 7928
rect 28460 7886 28488 7919
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28264 5364 28316 5370
rect 28264 5306 28316 5312
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 28092 2854 28120 4626
rect 28552 4622 28580 11194
rect 28724 9308 28776 9314
rect 28724 9250 28776 9256
rect 28632 8424 28684 8430
rect 28632 8366 28684 8372
rect 28644 7954 28672 8366
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28632 7812 28684 7818
rect 28632 7754 28684 7760
rect 28644 7721 28672 7754
rect 28630 7712 28686 7721
rect 28630 7647 28686 7656
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 27068 2848 27120 2854
rect 27068 2790 27120 2796
rect 27620 2848 27672 2854
rect 27620 2790 27672 2796
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27080 2378 27108 2790
rect 27158 2544 27214 2553
rect 27158 2479 27214 2488
rect 27172 2378 27200 2479
rect 28552 2417 28580 2994
rect 28736 2854 28764 9250
rect 28828 6361 28856 11194
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 29012 8090 29040 8842
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 29104 7834 29132 11194
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29182 8120 29238 8129
rect 29182 8055 29184 8064
rect 29236 8055 29238 8064
rect 29184 8026 29236 8032
rect 29012 7806 29132 7834
rect 29184 7812 29236 7818
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 28920 7478 28948 7686
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 29012 6905 29040 7806
rect 29184 7754 29236 7760
rect 29196 7721 29224 7754
rect 29288 7750 29316 8774
rect 29276 7744 29328 7750
rect 29182 7712 29238 7721
rect 29276 7686 29328 7692
rect 29182 7647 29238 7656
rect 28998 6896 29054 6905
rect 28998 6831 29054 6840
rect 29380 6730 29408 11194
rect 29656 11082 29684 11194
rect 29644 11076 29696 11082
rect 29644 11018 29696 11024
rect 29932 11014 29960 11194
rect 29920 11008 29972 11014
rect 29920 10950 29972 10956
rect 30208 9178 30236 11194
rect 30196 9172 30248 9178
rect 30196 9114 30248 9120
rect 30484 8294 30512 11194
rect 30472 8288 30524 8294
rect 30472 8230 30524 8236
rect 30760 8090 30788 11194
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 31036 8022 31064 11194
rect 29460 8016 29512 8022
rect 29458 7984 29460 7993
rect 31024 8016 31076 8022
rect 29512 7984 29514 7993
rect 31024 7958 31076 7964
rect 31312 7954 31340 11194
rect 29458 7919 29514 7928
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 31588 7886 31616 11194
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31206 7440 31262 7449
rect 31772 7410 31800 8230
rect 31864 7478 31892 11194
rect 32140 8294 32168 11194
rect 32416 9330 32444 11194
rect 32416 9302 32536 9330
rect 32312 9240 32364 9246
rect 32312 9182 32364 9188
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31852 7472 31904 7478
rect 31852 7414 31904 7420
rect 31206 7375 31262 7384
rect 31760 7404 31812 7410
rect 31220 7206 31248 7375
rect 31760 7346 31812 7352
rect 32324 7206 32352 9182
rect 32404 8492 32456 8498
rect 32404 8434 32456 8440
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 29368 6724 29420 6730
rect 29368 6666 29420 6672
rect 30380 6384 30432 6390
rect 28814 6352 28870 6361
rect 30380 6326 30432 6332
rect 28814 6287 28870 6296
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 28538 2408 28594 2417
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 27160 2372 27212 2378
rect 28538 2343 28594 2352
rect 27160 2314 27212 2320
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 28828 56 28856 4966
rect 30392 4758 30420 6326
rect 30668 6186 30696 7142
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 30656 6180 30708 6186
rect 30656 6122 30708 6128
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 30380 4752 30432 4758
rect 30380 4694 30432 4700
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 30392 4078 30420 4422
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28920 2854 28948 3130
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 30392 2310 30420 2994
rect 30380 2304 30432 2310
rect 30380 2246 30432 2252
rect 30944 56 30972 5170
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32416 4826 32444 8434
rect 32508 7410 32536 9302
rect 32588 9240 32640 9246
rect 32588 9182 32640 9188
rect 32496 7404 32548 7410
rect 32496 7346 32548 7352
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 31760 4616 31812 4622
rect 31760 4558 31812 4564
rect 31772 66 31800 4558
rect 32600 4049 32628 9182
rect 32692 6798 32720 11194
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32784 5166 32812 9114
rect 32968 9058 32996 11194
rect 33244 9330 33272 11194
rect 33244 9302 33456 9330
rect 32876 9030 32996 9058
rect 32876 6866 32904 9030
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33428 7410 33456 9302
rect 33520 7750 33548 11194
rect 33600 8424 33652 8430
rect 33600 8366 33652 8372
rect 33508 7744 33560 7750
rect 33508 7686 33560 7692
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 33230 6760 33286 6769
rect 33230 6695 33286 6704
rect 33244 6662 33272 6695
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33612 5846 33640 8366
rect 33692 7472 33744 7478
rect 33692 7414 33744 7420
rect 33600 5840 33652 5846
rect 33600 5782 33652 5788
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32772 5160 32824 5166
rect 32772 5102 32824 5108
rect 33704 4826 33732 7414
rect 33796 7002 33824 11194
rect 34072 8634 34100 11194
rect 34348 8634 34376 11194
rect 34428 9376 34480 9382
rect 34428 9318 34480 9324
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34440 7206 34468 9318
rect 34624 9110 34652 11194
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34716 8498 34744 8910
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34428 7200 34480 7206
rect 34428 7142 34480 7148
rect 33784 6996 33836 7002
rect 33784 6938 33836 6944
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 34808 4758 34836 8910
rect 34900 8616 34928 11194
rect 35176 8838 35204 11194
rect 35256 9104 35308 9110
rect 35256 9046 35308 9052
rect 35164 8832 35216 8838
rect 35164 8774 35216 8780
rect 35268 8634 35296 9046
rect 34980 8628 35032 8634
rect 34900 8588 34980 8616
rect 34980 8570 35032 8576
rect 35256 8628 35308 8634
rect 35256 8570 35308 8576
rect 35452 8480 35480 11194
rect 35728 9110 35756 11194
rect 35716 9104 35768 9110
rect 35716 9046 35768 9052
rect 35808 8832 35860 8838
rect 35808 8774 35860 8780
rect 35820 8634 35848 8774
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35532 8492 35584 8498
rect 35452 8452 35532 8480
rect 35532 8434 35584 8440
rect 35808 8288 35860 8294
rect 35808 8230 35860 8236
rect 34796 4752 34848 4758
rect 34796 4694 34848 4700
rect 35164 4616 35216 4622
rect 35164 4558 35216 4564
rect 32772 4548 32824 4554
rect 32772 4490 32824 4496
rect 32586 4040 32642 4049
rect 32586 3975 32642 3984
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31760 60 31812 66
rect 1306 0 1362 56
rect 3422 0 3478 56
rect 5538 0 5594 56
rect 7654 0 7710 56
rect 9770 0 9826 56
rect 11886 0 11942 56
rect 14002 0 14058 56
rect 16118 0 16174 56
rect 18234 0 18290 56
rect 20350 0 20406 56
rect 22466 0 22522 56
rect 24582 0 24638 56
rect 26698 0 26754 56
rect 28814 0 28870 56
rect 30930 0 30986 56
rect 32784 42 32812 4490
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 34716 338 34744 3470
rect 34704 332 34756 338
rect 34704 274 34756 280
rect 32968 56 33088 82
rect 35176 56 35204 4558
rect 35820 3738 35848 8230
rect 36004 8090 36032 11194
rect 36176 9308 36228 9314
rect 36176 9250 36228 9256
rect 36188 8498 36216 9250
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36280 8090 36308 11194
rect 36556 8634 36584 11194
rect 36728 9104 36780 9110
rect 36728 9046 36780 9052
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 36636 8560 36688 8566
rect 36636 8502 36688 8508
rect 35992 8084 36044 8090
rect 35992 8026 36044 8032
rect 36268 8084 36320 8090
rect 36268 8026 36320 8032
rect 36452 7812 36504 7818
rect 36452 7754 36504 7760
rect 36464 7410 36492 7754
rect 36544 7540 36596 7546
rect 36544 7482 36596 7488
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36556 7206 36584 7482
rect 36544 7200 36596 7206
rect 36544 7142 36596 7148
rect 36452 6860 36504 6866
rect 36452 6802 36504 6808
rect 36464 6390 36492 6802
rect 36452 6384 36504 6390
rect 36452 6326 36504 6332
rect 36648 4826 36676 8502
rect 36740 8362 36768 9046
rect 36832 8362 36860 11194
rect 37108 8430 37136 11194
rect 37096 8424 37148 8430
rect 37096 8366 37148 8372
rect 36728 8356 36780 8362
rect 36728 8298 36780 8304
rect 36820 8356 36872 8362
rect 36820 8298 36872 8304
rect 37384 8090 37412 11194
rect 37660 8634 37688 11194
rect 37936 9110 37964 11194
rect 38016 9240 38068 9246
rect 38016 9182 38068 9188
rect 37924 9104 37976 9110
rect 37924 9046 37976 9052
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37648 8628 37700 8634
rect 37648 8570 37700 8576
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 36820 8084 36872 8090
rect 36820 8026 36872 8032
rect 37372 8084 37424 8090
rect 37372 8026 37424 8032
rect 36832 7342 36860 8026
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 36820 7336 36872 7342
rect 36820 7278 36872 7284
rect 36636 4820 36688 4826
rect 36636 4762 36688 4768
rect 37292 4758 37320 7686
rect 37280 4752 37332 4758
rect 37280 4694 37332 4700
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 35808 3732 35860 3738
rect 35808 3674 35860 3680
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 35820 3097 35848 3130
rect 35806 3088 35862 3097
rect 35806 3023 35862 3032
rect 36556 2854 36584 3674
rect 36544 2848 36596 2854
rect 36544 2790 36596 2796
rect 37292 56 37320 4082
rect 37370 3496 37426 3505
rect 37370 3431 37426 3440
rect 37384 3058 37412 3431
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 37476 2961 37504 7822
rect 37568 7546 37596 8434
rect 37556 7540 37608 7546
rect 37556 7482 37608 7488
rect 37660 6458 37688 8434
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 37752 7478 37780 7822
rect 37740 7472 37792 7478
rect 37740 7414 37792 7420
rect 37844 6730 37872 8774
rect 38028 8498 38056 9182
rect 38212 8498 38240 11194
rect 38384 9172 38436 9178
rect 38384 9114 38436 9120
rect 38396 8498 38424 9114
rect 38016 8492 38068 8498
rect 38016 8434 38068 8440
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 38384 8492 38436 8498
rect 38384 8434 38436 8440
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38488 8090 38516 11194
rect 38568 9104 38620 9110
rect 38568 9046 38620 9052
rect 38580 8362 38608 9046
rect 38660 8492 38712 8498
rect 38660 8434 38712 8440
rect 38568 8356 38620 8362
rect 38568 8298 38620 8304
rect 38476 8084 38528 8090
rect 38476 8026 38528 8032
rect 38568 8016 38620 8022
rect 38568 7958 38620 7964
rect 38476 7948 38528 7954
rect 38476 7890 38528 7896
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 37832 6724 37884 6730
rect 37832 6666 37884 6672
rect 38488 6662 38516 7890
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 37648 6452 37700 6458
rect 37648 6394 37700 6400
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 38580 5846 38608 7958
rect 38672 7562 38700 8434
rect 38764 8106 38792 11194
rect 38844 8968 38896 8974
rect 39040 8922 39068 11194
rect 39316 9058 39344 11194
rect 39316 9030 39436 9058
rect 38844 8910 38896 8916
rect 38856 8498 38884 8910
rect 38948 8894 39068 8922
rect 38948 8634 38976 8894
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 38844 8492 38896 8498
rect 38844 8434 38896 8440
rect 39408 8362 39436 9030
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 38764 8090 38884 8106
rect 39592 8090 39620 11194
rect 41786 9888 41842 9897
rect 41786 9823 41842 9832
rect 41696 9444 41748 9450
rect 41696 9386 41748 9392
rect 41604 8900 41656 8906
rect 41604 8842 41656 8848
rect 41616 8498 41644 8842
rect 41708 8498 41736 9386
rect 41800 8634 41828 9823
rect 42338 9616 42394 9625
rect 42338 9551 42394 9560
rect 41880 9036 41932 9042
rect 41880 8978 41932 8984
rect 41892 8922 41920 8978
rect 41892 8894 42104 8922
rect 41972 8832 42024 8838
rect 41972 8774 42024 8780
rect 41788 8628 41840 8634
rect 41788 8570 41840 8576
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 41604 8492 41656 8498
rect 41604 8434 41656 8440
rect 41696 8492 41748 8498
rect 41696 8434 41748 8440
rect 38764 8084 38896 8090
rect 38764 8078 38844 8084
rect 38844 8026 38896 8032
rect 39580 8084 39632 8090
rect 39580 8026 39632 8032
rect 38936 7880 38988 7886
rect 39488 7880 39540 7886
rect 38936 7822 38988 7828
rect 39302 7848 39358 7857
rect 38844 7812 38896 7818
rect 38844 7754 38896 7760
rect 38672 7534 38792 7562
rect 38660 7404 38712 7410
rect 38660 7346 38712 7352
rect 38568 5840 38620 5846
rect 38568 5782 38620 5788
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37462 2952 37518 2961
rect 37462 2887 37518 2896
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38672 406 38700 7346
rect 38764 5370 38792 7534
rect 38856 7478 38884 7754
rect 38844 7472 38896 7478
rect 38844 7414 38896 7420
rect 38752 5364 38804 5370
rect 38752 5306 38804 5312
rect 38948 4010 38976 7822
rect 39488 7822 39540 7828
rect 39302 7783 39358 7792
rect 39316 7750 39344 7783
rect 39304 7744 39356 7750
rect 39304 7686 39356 7692
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39500 7002 39528 7822
rect 39488 6996 39540 7002
rect 39488 6938 39540 6944
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39580 5704 39632 5710
rect 39580 5646 39632 5652
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39396 4684 39448 4690
rect 39396 4626 39448 4632
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 38936 4004 38988 4010
rect 38936 3946 38988 3952
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38660 400 38712 406
rect 38660 342 38712 348
rect 39408 56 39436 4626
rect 39592 134 39620 5646
rect 39960 4826 39988 8434
rect 40316 8424 40368 8430
rect 40316 8366 40368 8372
rect 41984 8378 42012 8774
rect 42076 8566 42104 8894
rect 42154 8800 42210 8809
rect 42154 8735 42210 8744
rect 42168 8634 42196 8735
rect 42156 8628 42208 8634
rect 42156 8570 42208 8576
rect 42064 8560 42116 8566
rect 42064 8502 42116 8508
rect 42156 8492 42208 8498
rect 42156 8434 42208 8440
rect 42168 8378 42196 8434
rect 40132 6316 40184 6322
rect 40132 6258 40184 6264
rect 40040 5228 40092 5234
rect 40040 5170 40092 5176
rect 39948 4820 40000 4826
rect 39948 4762 40000 4768
rect 40052 3398 40080 5170
rect 40144 3602 40172 6258
rect 40328 5098 40356 8366
rect 41984 8350 42196 8378
rect 42352 8090 42380 9551
rect 43166 9344 43222 9353
rect 43166 9279 43222 9288
rect 42614 9072 42670 9081
rect 42614 9007 42670 9016
rect 42628 8090 42656 9007
rect 42708 8628 42760 8634
rect 42708 8570 42760 8576
rect 42720 8537 42748 8570
rect 42706 8528 42762 8537
rect 42706 8463 42762 8472
rect 43076 8356 43128 8362
rect 43076 8298 43128 8304
rect 43088 8265 43116 8298
rect 43074 8256 43130 8265
rect 43074 8191 43130 8200
rect 42340 8084 42392 8090
rect 42340 8026 42392 8032
rect 42616 8084 42668 8090
rect 42616 8026 42668 8032
rect 40684 7880 40736 7886
rect 40684 7822 40736 7828
rect 42524 7880 42576 7886
rect 42524 7822 42576 7828
rect 40316 5092 40368 5098
rect 40316 5034 40368 5040
rect 40696 4010 40724 7822
rect 41788 7336 41840 7342
rect 41788 7278 41840 7284
rect 40868 6792 40920 6798
rect 40868 6734 40920 6740
rect 40684 4004 40736 4010
rect 40684 3946 40736 3952
rect 40132 3596 40184 3602
rect 40132 3538 40184 3544
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 40880 270 40908 6734
rect 41800 5137 41828 7278
rect 42536 7206 42564 7822
rect 43076 7744 43128 7750
rect 43076 7686 43128 7692
rect 43088 7449 43116 7686
rect 43180 7546 43208 9279
rect 43444 8356 43496 8362
rect 43444 8298 43496 8304
rect 43456 7993 43484 8298
rect 43442 7984 43498 7993
rect 43442 7919 43498 7928
rect 43260 7880 43312 7886
rect 43260 7822 43312 7828
rect 43168 7540 43220 7546
rect 43168 7482 43220 7488
rect 43074 7440 43130 7449
rect 43074 7375 43130 7384
rect 42524 7200 42576 7206
rect 42524 7142 42576 7148
rect 42984 6792 43036 6798
rect 42984 6734 43036 6740
rect 42996 5642 43024 6734
rect 43076 6656 43128 6662
rect 43074 6624 43076 6633
rect 43128 6624 43130 6633
rect 43074 6559 43130 6568
rect 43168 6248 43220 6254
rect 43168 6190 43220 6196
rect 43076 6112 43128 6118
rect 43074 6080 43076 6089
rect 43128 6080 43130 6089
rect 43074 6015 43130 6024
rect 42984 5636 43036 5642
rect 42984 5578 43036 5584
rect 43076 5568 43128 5574
rect 43074 5536 43076 5545
rect 43128 5536 43130 5545
rect 43074 5471 43130 5480
rect 42340 5160 42392 5166
rect 41786 5128 41842 5137
rect 42340 5102 42392 5108
rect 41786 5063 41842 5072
rect 41512 4616 41564 4622
rect 41512 4558 41564 4564
rect 40960 4140 41012 4146
rect 40960 4082 41012 4088
rect 40972 2922 41000 4082
rect 40960 2916 41012 2922
rect 40960 2858 41012 2864
rect 40868 264 40920 270
rect 40868 206 40920 212
rect 39580 128 39632 134
rect 39580 70 39632 76
rect 41524 56 41552 4558
rect 42352 3670 42380 5102
rect 43076 5024 43128 5030
rect 43074 4992 43076 5001
rect 43128 4992 43130 5001
rect 43074 4927 43130 4936
rect 42892 4616 42944 4622
rect 42892 4558 42944 4564
rect 42904 4282 42932 4558
rect 43076 4480 43128 4486
rect 43074 4448 43076 4457
rect 43128 4448 43130 4457
rect 43074 4383 43130 4392
rect 42892 4276 42944 4282
rect 42892 4218 42944 4224
rect 43180 4146 43208 6190
rect 43272 5273 43300 7822
rect 43444 7744 43496 7750
rect 43442 7712 43444 7721
rect 43496 7712 43498 7721
rect 43442 7647 43498 7656
rect 43444 7200 43496 7206
rect 43442 7168 43444 7177
rect 43496 7168 43498 7177
rect 43442 7103 43498 7112
rect 43442 6896 43498 6905
rect 43442 6831 43498 6840
rect 43456 6662 43484 6831
rect 43444 6656 43496 6662
rect 43444 6598 43496 6604
rect 43444 6452 43496 6458
rect 43444 6394 43496 6400
rect 43456 6361 43484 6394
rect 43442 6352 43498 6361
rect 43442 6287 43498 6296
rect 43444 5840 43496 5846
rect 43442 5808 43444 5817
rect 43496 5808 43498 5817
rect 43442 5743 43498 5752
rect 43352 5704 43404 5710
rect 43352 5646 43404 5652
rect 43258 5264 43314 5273
rect 43258 5199 43314 5208
rect 43168 4140 43220 4146
rect 43168 4082 43220 4088
rect 43076 3936 43128 3942
rect 43074 3904 43076 3913
rect 43128 3904 43130 3913
rect 43074 3839 43130 3848
rect 42340 3664 42392 3670
rect 42340 3606 42392 3612
rect 43076 3392 43128 3398
rect 43074 3360 43076 3369
rect 43128 3360 43130 3369
rect 43074 3295 43130 3304
rect 42890 3088 42946 3097
rect 42890 3023 42892 3032
rect 42944 3023 42946 3032
rect 42892 2994 42944 3000
rect 43364 2990 43392 5646
rect 43444 5364 43496 5370
rect 43444 5306 43496 5312
rect 43456 5273 43484 5306
rect 43442 5264 43498 5273
rect 43442 5199 43498 5208
rect 43444 4752 43496 4758
rect 43442 4720 43444 4729
rect 43496 4720 43498 4729
rect 43442 4655 43498 4664
rect 43442 4176 43498 4185
rect 43442 4111 43498 4120
rect 43456 4010 43484 4111
rect 43628 4072 43680 4078
rect 43628 4014 43680 4020
rect 43444 4004 43496 4010
rect 43444 3946 43496 3952
rect 43444 3664 43496 3670
rect 43442 3632 43444 3641
rect 43496 3632 43498 3641
rect 43442 3567 43498 3576
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 43456 3097 43484 3130
rect 43442 3088 43498 3097
rect 43442 3023 43498 3032
rect 43352 2984 43404 2990
rect 43352 2926 43404 2932
rect 42984 2848 43036 2854
rect 43076 2848 43128 2854
rect 42984 2790 43036 2796
rect 43074 2816 43076 2825
rect 43128 2816 43130 2825
rect 42156 2576 42208 2582
rect 42156 2518 42208 2524
rect 42168 1737 42196 2518
rect 42708 2304 42760 2310
rect 42708 2246 42760 2252
rect 42154 1728 42210 1737
rect 42154 1663 42210 1672
rect 42720 1465 42748 2246
rect 42996 2009 43024 2790
rect 43074 2751 43130 2760
rect 43444 2576 43496 2582
rect 43442 2544 43444 2553
rect 43496 2544 43498 2553
rect 43442 2479 43498 2488
rect 43076 2304 43128 2310
rect 43074 2272 43076 2281
rect 43128 2272 43130 2281
rect 43074 2207 43130 2216
rect 42982 2000 43038 2009
rect 42982 1935 43038 1944
rect 42706 1456 42762 1465
rect 42706 1391 42762 1400
rect 43640 56 43668 4014
rect 32968 54 33102 56
rect 32968 42 32996 54
rect 32784 14 32996 42
rect 31760 2 31812 8
rect 33046 0 33102 54
rect 35162 0 35218 56
rect 37278 0 37334 56
rect 39394 0 39450 56
rect 41510 0 41566 56
rect 43626 0 43682 56
<< via2 >>
rect 1306 9424 1362 9480
rect 1214 7928 1270 7984
rect 1122 7656 1178 7712
rect 2870 9152 2926 9208
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3422 7792 3478 7848
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 1306 7384 1362 7440
rect 3422 7248 3478 7304
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1766 6704 1822 6760
rect 2870 6568 2926 6624
rect 1766 6024 1822 6080
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2870 5616 2926 5672
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2686 5208 2742 5264
rect 2686 4936 2742 4992
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 5538 2896 5594 2952
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2870 2216 2926 2272
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 7838 5208 7894 5264
rect 7010 4936 7066 4992
rect 2870 1808 2926 1864
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9494 3984 9550 4040
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9586 2488 9642 2544
rect 9494 1672 9550 1728
rect 9402 1400 9458 1456
rect 10138 10784 10194 10840
rect 9954 7964 9956 7984
rect 9956 7964 10008 7984
rect 10008 7964 10010 7984
rect 9954 7928 10010 7964
rect 10506 6316 10562 6352
rect 10506 6296 10508 6316
rect 10508 6296 10560 6316
rect 10560 6296 10562 6316
rect 10966 6704 11022 6760
rect 13358 7384 13414 7440
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14738 8064 14794 8120
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 15750 10512 15806 10568
rect 16026 10920 16082 10976
rect 15934 9696 15990 9752
rect 15198 7792 15254 7848
rect 15382 7792 15438 7848
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 14646 7112 14702 7168
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13726 5616 13782 5672
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 16486 8880 16542 8936
rect 16118 6704 16174 6760
rect 15566 6160 15622 6216
rect 17682 10648 17738 10704
rect 18050 8200 18106 8256
rect 16486 5752 16542 5808
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 18602 6840 18658 6896
rect 19982 9696 20038 9752
rect 19706 8064 19762 8120
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 19798 7656 19854 7712
rect 19706 7384 19762 7440
rect 20442 8064 20498 8120
rect 20718 9288 20774 9344
rect 20534 7656 20590 7712
rect 20442 7520 20498 7576
rect 19798 7112 19854 7168
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19982 6840 20038 6896
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 19062 6160 19118 6216
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 17222 5072 17278 5128
rect 18510 5072 18566 5128
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19430 4664 19486 4720
rect 19338 4548 19394 4584
rect 19338 4528 19340 4548
rect 19340 4528 19392 4548
rect 19392 4528 19394 4548
rect 21454 6840 21510 6896
rect 22098 9560 22154 9616
rect 23110 6840 23166 6896
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 20902 4120 20958 4176
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 10966 3032 11022 3088
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20166 2916 20222 2952
rect 20166 2896 20168 2916
rect 20168 2896 20220 2916
rect 20220 2896 20222 2916
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 11886 2352 11942 2408
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 20718 1944 20774 2000
rect 20350 1808 20406 1864
rect 23018 5208 23074 5264
rect 23386 9832 23442 9888
rect 23386 7112 23442 7168
rect 23294 6160 23350 6216
rect 24122 10784 24178 10840
rect 23846 9152 23902 9208
rect 24398 9016 24454 9072
rect 24674 8064 24730 8120
rect 24858 7268 24914 7304
rect 24858 7248 24860 7268
rect 24860 7248 24912 7268
rect 24912 7248 24914 7268
rect 25778 8880 25834 8936
rect 26330 10920 26386 10976
rect 26606 10512 26662 10568
rect 26330 8472 26386 8528
rect 25778 8200 25834 8256
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 23386 3440 23442 3496
rect 24858 3596 24914 3632
rect 24858 3576 24860 3596
rect 24860 3576 24912 3596
rect 24912 3576 24914 3596
rect 24766 3440 24822 3496
rect 25870 4004 25926 4040
rect 25870 3984 25872 4004
rect 25872 3984 25924 4004
rect 25924 3984 25926 4004
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 26146 2508 26202 2544
rect 26146 2488 26148 2508
rect 26148 2488 26200 2508
rect 26200 2488 26202 2508
rect 27434 10648 27490 10704
rect 27618 9424 27674 9480
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 26974 8064 27030 8120
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27618 7928 27674 7984
rect 27342 7248 27398 7304
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 28446 7928 28502 7984
rect 28630 7656 28686 7712
rect 27158 2488 27214 2544
rect 29182 8084 29238 8120
rect 29182 8064 29184 8084
rect 29184 8064 29236 8084
rect 29236 8064 29238 8084
rect 29182 7656 29238 7712
rect 28998 6840 29054 6896
rect 29458 7964 29460 7984
rect 29460 7964 29512 7984
rect 29512 7964 29514 7984
rect 29458 7928 29514 7964
rect 31206 7384 31262 7440
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 28814 6296 28870 6352
rect 28538 2352 28594 2408
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33230 6704 33286 6760
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 32586 3984 32642 4040
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 35806 3032 35862 3088
rect 37370 3440 37426 3496
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 41786 9832 41842 9888
rect 42338 9560 42394 9616
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 37462 2896 37518 2952
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39302 7792 39358 7848
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 42154 8744 42210 8800
rect 43166 9288 43222 9344
rect 42614 9016 42670 9072
rect 42706 8472 42762 8528
rect 43074 8200 43130 8256
rect 43442 7928 43498 7984
rect 43074 7384 43130 7440
rect 43074 6604 43076 6624
rect 43076 6604 43128 6624
rect 43128 6604 43130 6624
rect 43074 6568 43130 6604
rect 43074 6060 43076 6080
rect 43076 6060 43128 6080
rect 43128 6060 43130 6080
rect 43074 6024 43130 6060
rect 43074 5516 43076 5536
rect 43076 5516 43128 5536
rect 43128 5516 43130 5536
rect 43074 5480 43130 5516
rect 41786 5072 41842 5128
rect 43074 4972 43076 4992
rect 43076 4972 43128 4992
rect 43128 4972 43130 4992
rect 43074 4936 43130 4972
rect 43074 4428 43076 4448
rect 43076 4428 43128 4448
rect 43128 4428 43130 4448
rect 43074 4392 43130 4428
rect 43442 7692 43444 7712
rect 43444 7692 43496 7712
rect 43496 7692 43498 7712
rect 43442 7656 43498 7692
rect 43442 7148 43444 7168
rect 43444 7148 43496 7168
rect 43496 7148 43498 7168
rect 43442 7112 43498 7148
rect 43442 6840 43498 6896
rect 43442 6296 43498 6352
rect 43442 5788 43444 5808
rect 43444 5788 43496 5808
rect 43496 5788 43498 5808
rect 43442 5752 43498 5788
rect 43258 5208 43314 5264
rect 43074 3884 43076 3904
rect 43076 3884 43128 3904
rect 43128 3884 43130 3904
rect 43074 3848 43130 3884
rect 43074 3340 43076 3360
rect 43076 3340 43128 3360
rect 43128 3340 43130 3360
rect 43074 3304 43130 3340
rect 42890 3052 42946 3088
rect 42890 3032 42892 3052
rect 42892 3032 42944 3052
rect 42944 3032 42946 3052
rect 43442 5208 43498 5264
rect 43442 4700 43444 4720
rect 43444 4700 43496 4720
rect 43496 4700 43498 4720
rect 43442 4664 43498 4700
rect 43442 4120 43498 4176
rect 43442 3612 43444 3632
rect 43444 3612 43496 3632
rect 43496 3612 43498 3632
rect 43442 3576 43498 3612
rect 43442 3032 43498 3088
rect 43074 2796 43076 2816
rect 43076 2796 43128 2816
rect 43128 2796 43130 2816
rect 42154 1672 42210 1728
rect 43074 2760 43130 2796
rect 43442 2524 43444 2544
rect 43444 2524 43496 2544
rect 43496 2524 43498 2544
rect 43442 2488 43498 2524
rect 43074 2252 43076 2272
rect 43076 2252 43128 2272
rect 43128 2252 43130 2272
rect 43074 2216 43130 2252
rect 42982 1944 43038 2000
rect 42706 1400 42762 1456
<< metal3 >>
rect 16021 10978 16087 10981
rect 26325 10978 26391 10981
rect 16021 10976 26391 10978
rect 16021 10920 16026 10976
rect 16082 10920 26330 10976
rect 26386 10920 26391 10976
rect 16021 10918 26391 10920
rect 16021 10915 16087 10918
rect 26325 10915 26391 10918
rect 10133 10842 10199 10845
rect 24117 10842 24183 10845
rect 10133 10840 24183 10842
rect 10133 10784 10138 10840
rect 10194 10784 24122 10840
rect 24178 10784 24183 10840
rect 10133 10782 24183 10784
rect 10133 10779 10199 10782
rect 24117 10779 24183 10782
rect 17677 10706 17743 10709
rect 27429 10706 27495 10709
rect 17677 10704 27495 10706
rect 17677 10648 17682 10704
rect 17738 10648 27434 10704
rect 27490 10648 27495 10704
rect 17677 10646 27495 10648
rect 17677 10643 17743 10646
rect 27429 10643 27495 10646
rect 15745 10570 15811 10573
rect 26601 10570 26667 10573
rect 15745 10568 26667 10570
rect 15745 10512 15750 10568
rect 15806 10512 26606 10568
rect 26662 10512 26667 10568
rect 15745 10510 26667 10512
rect 15745 10507 15811 10510
rect 26601 10507 26667 10510
rect 0 9890 120 9920
rect 23381 9890 23447 9893
rect 0 9888 23447 9890
rect 0 9832 23386 9888
rect 23442 9832 23447 9888
rect 0 9830 23447 9832
rect 0 9800 120 9830
rect 23381 9827 23447 9830
rect 41781 9890 41847 9893
rect 44880 9890 45000 9920
rect 41781 9888 45000 9890
rect 41781 9832 41786 9888
rect 41842 9832 45000 9888
rect 41781 9830 45000 9832
rect 41781 9827 41847 9830
rect 44880 9800 45000 9830
rect 15929 9754 15995 9757
rect 19977 9754 20043 9757
rect 15929 9752 20043 9754
rect 15929 9696 15934 9752
rect 15990 9696 19982 9752
rect 20038 9696 20043 9752
rect 15929 9694 20043 9696
rect 15929 9691 15995 9694
rect 19977 9691 20043 9694
rect 0 9618 120 9648
rect 22093 9618 22159 9621
rect 0 9616 22159 9618
rect 0 9560 22098 9616
rect 22154 9560 22159 9616
rect 0 9558 22159 9560
rect 0 9528 120 9558
rect 22093 9555 22159 9558
rect 42333 9618 42399 9621
rect 44880 9618 45000 9648
rect 42333 9616 45000 9618
rect 42333 9560 42338 9616
rect 42394 9560 45000 9616
rect 42333 9558 45000 9560
rect 42333 9555 42399 9558
rect 44880 9528 45000 9558
rect 1301 9482 1367 9485
rect 27613 9482 27679 9485
rect 1301 9480 27679 9482
rect 1301 9424 1306 9480
rect 1362 9424 27618 9480
rect 27674 9424 27679 9480
rect 1301 9422 27679 9424
rect 1301 9419 1367 9422
rect 27613 9419 27679 9422
rect 0 9346 120 9376
rect 20713 9346 20779 9349
rect 0 9344 20779 9346
rect 0 9288 20718 9344
rect 20774 9288 20779 9344
rect 0 9286 20779 9288
rect 0 9256 120 9286
rect 20713 9283 20779 9286
rect 43161 9346 43227 9349
rect 44880 9346 45000 9376
rect 43161 9344 45000 9346
rect 43161 9288 43166 9344
rect 43222 9288 45000 9344
rect 43161 9286 45000 9288
rect 43161 9283 43227 9286
rect 44880 9256 45000 9286
rect 2865 9210 2931 9213
rect 23841 9210 23907 9213
rect 2865 9208 23907 9210
rect 2865 9152 2870 9208
rect 2926 9152 23846 9208
rect 23902 9152 23907 9208
rect 2865 9150 23907 9152
rect 2865 9147 2931 9150
rect 23841 9147 23907 9150
rect 0 9074 120 9104
rect 24393 9074 24459 9077
rect 0 9072 24459 9074
rect 0 9016 24398 9072
rect 24454 9016 24459 9072
rect 0 9014 24459 9016
rect 0 8984 120 9014
rect 24393 9011 24459 9014
rect 42609 9074 42675 9077
rect 44880 9074 45000 9104
rect 42609 9072 45000 9074
rect 42609 9016 42614 9072
rect 42670 9016 45000 9072
rect 42609 9014 45000 9016
rect 42609 9011 42675 9014
rect 44880 8984 45000 9014
rect 16481 8938 16547 8941
rect 25773 8938 25839 8941
rect 16481 8936 25839 8938
rect 16481 8880 16486 8936
rect 16542 8880 25778 8936
rect 25834 8880 25839 8936
rect 16481 8878 25839 8880
rect 16481 8875 16547 8878
rect 25773 8875 25839 8878
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 42149 8802 42215 8805
rect 44880 8802 45000 8832
rect 42149 8800 45000 8802
rect 42149 8744 42154 8800
rect 42210 8744 45000 8800
rect 42149 8742 45000 8744
rect 42149 8739 42215 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 44880 8712 45000 8742
rect 39006 8671 39322 8672
rect 0 8530 120 8560
rect 26325 8530 26391 8533
rect 0 8528 26391 8530
rect 0 8472 26330 8528
rect 26386 8472 26391 8528
rect 0 8470 26391 8472
rect 0 8440 120 8470
rect 26325 8467 26391 8470
rect 42701 8530 42767 8533
rect 44880 8530 45000 8560
rect 42701 8528 45000 8530
rect 42701 8472 42706 8528
rect 42762 8472 45000 8528
rect 42701 8470 45000 8472
rect 42701 8467 42767 8470
rect 44880 8440 45000 8470
rect 19750 8334 20546 8394
rect 0 8258 120 8288
rect 18045 8258 18111 8261
rect 19750 8258 19810 8334
rect 0 8198 1824 8258
rect 0 8168 120 8198
rect 0 7986 120 8016
rect 1209 7986 1275 7989
rect 0 7984 1275 7986
rect 0 7928 1214 7984
rect 1270 7928 1275 7984
rect 0 7926 1275 7928
rect 0 7896 120 7926
rect 1209 7923 1275 7926
rect 0 7714 120 7744
rect 1117 7714 1183 7717
rect 0 7712 1183 7714
rect 0 7656 1122 7712
rect 1178 7656 1183 7712
rect 0 7654 1183 7656
rect 0 7624 120 7654
rect 1117 7651 1183 7654
rect 0 7442 120 7472
rect 1301 7442 1367 7445
rect 0 7440 1367 7442
rect 0 7384 1306 7440
rect 1362 7384 1367 7440
rect 0 7382 1367 7384
rect 1764 7442 1824 8198
rect 18045 8256 19810 8258
rect 18045 8200 18050 8256
rect 18106 8200 19810 8256
rect 18045 8198 19810 8200
rect 20486 8258 20546 8334
rect 25773 8258 25839 8261
rect 20486 8256 25839 8258
rect 20486 8200 25778 8256
rect 25834 8200 25839 8256
rect 20486 8198 25839 8200
rect 18045 8195 18111 8198
rect 25773 8195 25839 8198
rect 43069 8258 43135 8261
rect 44880 8258 45000 8288
rect 43069 8256 45000 8258
rect 43069 8200 43074 8256
rect 43130 8200 45000 8256
rect 43069 8198 45000 8200
rect 43069 8195 43135 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 44880 8168 45000 8198
rect 37946 8127 38262 8128
rect 14733 8122 14799 8125
rect 19701 8122 19767 8125
rect 14733 8120 19767 8122
rect 14733 8064 14738 8120
rect 14794 8064 19706 8120
rect 19762 8064 19767 8120
rect 14733 8062 19767 8064
rect 14733 8059 14799 8062
rect 19701 8059 19767 8062
rect 20437 8122 20503 8125
rect 24669 8122 24735 8125
rect 20437 8120 24735 8122
rect 20437 8064 20442 8120
rect 20498 8064 24674 8120
rect 24730 8064 24735 8120
rect 20437 8062 24735 8064
rect 20437 8059 20503 8062
rect 24669 8059 24735 8062
rect 26969 8122 27035 8125
rect 29177 8122 29243 8125
rect 26969 8120 29243 8122
rect 26969 8064 26974 8120
rect 27030 8064 29182 8120
rect 29238 8064 29243 8120
rect 26969 8062 29243 8064
rect 26969 8059 27035 8062
rect 29177 8059 29243 8062
rect 9949 7986 10015 7989
rect 27613 7986 27679 7989
rect 9949 7984 27679 7986
rect 9949 7928 9954 7984
rect 10010 7928 27618 7984
rect 27674 7928 27679 7984
rect 9949 7926 27679 7928
rect 9949 7923 10015 7926
rect 27613 7923 27679 7926
rect 28441 7986 28507 7989
rect 29453 7986 29519 7989
rect 28441 7984 29519 7986
rect 28441 7928 28446 7984
rect 28502 7928 29458 7984
rect 29514 7928 29519 7984
rect 28441 7926 29519 7928
rect 28441 7923 28507 7926
rect 29453 7923 29519 7926
rect 43437 7986 43503 7989
rect 44880 7986 45000 8016
rect 43437 7984 45000 7986
rect 43437 7928 43442 7984
rect 43498 7928 45000 7984
rect 43437 7926 45000 7928
rect 43437 7923 43503 7926
rect 44880 7896 45000 7926
rect 3417 7850 3483 7853
rect 15193 7850 15259 7853
rect 3417 7848 11714 7850
rect 3417 7792 3422 7848
rect 3478 7792 11714 7848
rect 3417 7790 11714 7792
rect 3417 7787 3483 7790
rect 11654 7714 11714 7790
rect 12390 7848 15259 7850
rect 12390 7792 15198 7848
rect 15254 7792 15259 7848
rect 12390 7790 15259 7792
rect 12390 7714 12450 7790
rect 15193 7787 15259 7790
rect 15377 7850 15443 7853
rect 39297 7850 39363 7853
rect 15377 7848 39363 7850
rect 15377 7792 15382 7848
rect 15438 7792 39302 7848
rect 39358 7792 39363 7848
rect 15377 7790 39363 7792
rect 15377 7787 15443 7790
rect 39297 7787 39363 7790
rect 11654 7654 12450 7714
rect 19793 7714 19859 7717
rect 20529 7714 20595 7717
rect 19793 7712 20595 7714
rect 19793 7656 19798 7712
rect 19854 7656 20534 7712
rect 20590 7656 20595 7712
rect 19793 7654 20595 7656
rect 19793 7651 19859 7654
rect 20529 7651 20595 7654
rect 28625 7714 28691 7717
rect 29177 7714 29243 7717
rect 28625 7712 29243 7714
rect 28625 7656 28630 7712
rect 28686 7656 29182 7712
rect 29238 7656 29243 7712
rect 28625 7654 29243 7656
rect 28625 7651 28691 7654
rect 29177 7651 29243 7654
rect 43437 7714 43503 7717
rect 44880 7714 45000 7744
rect 43437 7712 45000 7714
rect 43437 7656 43442 7712
rect 43498 7656 45000 7712
rect 43437 7654 45000 7656
rect 43437 7651 43503 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 44880 7624 45000 7654
rect 39006 7583 39322 7584
rect 20437 7578 20503 7581
rect 15518 7576 20503 7578
rect 15518 7520 20442 7576
rect 20498 7520 20503 7576
rect 15518 7518 20503 7520
rect 13353 7442 13419 7445
rect 15518 7442 15578 7518
rect 20437 7515 20503 7518
rect 1764 7382 6930 7442
rect 0 7352 120 7382
rect 1301 7379 1367 7382
rect 3417 7306 3483 7309
rect 1764 7304 3483 7306
rect 1764 7248 3422 7304
rect 3478 7248 3483 7304
rect 1764 7246 3483 7248
rect 6870 7306 6930 7382
rect 13353 7440 15578 7442
rect 13353 7384 13358 7440
rect 13414 7384 15578 7440
rect 13353 7382 15578 7384
rect 19701 7442 19767 7445
rect 31201 7442 31267 7445
rect 19701 7440 31267 7442
rect 19701 7384 19706 7440
rect 19762 7384 31206 7440
rect 31262 7384 31267 7440
rect 19701 7382 31267 7384
rect 13353 7379 13419 7382
rect 19701 7379 19767 7382
rect 31201 7379 31267 7382
rect 43069 7442 43135 7445
rect 44880 7442 45000 7472
rect 43069 7440 45000 7442
rect 43069 7384 43074 7440
rect 43130 7384 45000 7440
rect 43069 7382 45000 7384
rect 43069 7379 43135 7382
rect 44880 7352 45000 7382
rect 24853 7306 24919 7309
rect 27337 7306 27403 7309
rect 6870 7304 24919 7306
rect 6870 7248 24858 7304
rect 24914 7248 24919 7304
rect 6870 7246 24919 7248
rect 0 7170 120 7200
rect 1764 7170 1824 7246
rect 3417 7243 3483 7246
rect 24853 7243 24919 7246
rect 25822 7304 27403 7306
rect 25822 7248 27342 7304
rect 27398 7248 27403 7304
rect 25822 7246 27403 7248
rect 0 7110 1824 7170
rect 14641 7170 14707 7173
rect 19793 7170 19859 7173
rect 14641 7168 19859 7170
rect 14641 7112 14646 7168
rect 14702 7112 19798 7168
rect 19854 7112 19859 7168
rect 14641 7110 19859 7112
rect 0 7080 120 7110
rect 14641 7107 14707 7110
rect 19793 7107 19859 7110
rect 23381 7170 23447 7173
rect 25822 7170 25882 7246
rect 27337 7243 27403 7246
rect 23381 7168 25882 7170
rect 23381 7112 23386 7168
rect 23442 7112 25882 7168
rect 23381 7110 25882 7112
rect 43437 7170 43503 7173
rect 44880 7170 45000 7200
rect 43437 7168 45000 7170
rect 43437 7112 43442 7168
rect 43498 7112 45000 7168
rect 43437 7110 45000 7112
rect 23381 7107 23447 7110
rect 43437 7107 43503 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 44880 7080 45000 7110
rect 37946 7039 38262 7040
rect 0 6898 120 6928
rect 18597 6898 18663 6901
rect 0 6896 18663 6898
rect 0 6840 18602 6896
rect 18658 6840 18663 6896
rect 0 6838 18663 6840
rect 0 6808 120 6838
rect 18597 6835 18663 6838
rect 19977 6898 20043 6901
rect 21449 6898 21515 6901
rect 19977 6896 21515 6898
rect 19977 6840 19982 6896
rect 20038 6840 21454 6896
rect 21510 6840 21515 6896
rect 19977 6838 21515 6840
rect 19977 6835 20043 6838
rect 21449 6835 21515 6838
rect 23105 6898 23171 6901
rect 28993 6898 29059 6901
rect 23105 6896 29059 6898
rect 23105 6840 23110 6896
rect 23166 6840 28998 6896
rect 29054 6840 29059 6896
rect 23105 6838 29059 6840
rect 23105 6835 23171 6838
rect 28993 6835 29059 6838
rect 43437 6898 43503 6901
rect 44880 6898 45000 6928
rect 43437 6896 45000 6898
rect 43437 6840 43442 6896
rect 43498 6840 45000 6896
rect 43437 6838 45000 6840
rect 43437 6835 43503 6838
rect 44880 6808 45000 6838
rect 1761 6762 1827 6765
rect 10961 6762 11027 6765
rect 1761 6760 11027 6762
rect 1761 6704 1766 6760
rect 1822 6704 10966 6760
rect 11022 6704 11027 6760
rect 1761 6702 11027 6704
rect 1761 6699 1827 6702
rect 10961 6699 11027 6702
rect 16113 6762 16179 6765
rect 33225 6762 33291 6765
rect 16113 6760 33291 6762
rect 16113 6704 16118 6760
rect 16174 6704 33230 6760
rect 33286 6704 33291 6760
rect 16113 6702 33291 6704
rect 16113 6699 16179 6702
rect 33225 6699 33291 6702
rect 0 6626 120 6656
rect 2865 6626 2931 6629
rect 0 6624 2931 6626
rect 0 6568 2870 6624
rect 2926 6568 2931 6624
rect 0 6566 2931 6568
rect 0 6536 120 6566
rect 2865 6563 2931 6566
rect 43069 6626 43135 6629
rect 44880 6626 45000 6656
rect 43069 6624 45000 6626
rect 43069 6568 43074 6624
rect 43130 6568 45000 6624
rect 43069 6566 45000 6568
rect 43069 6563 43135 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 44880 6536 45000 6566
rect 39006 6495 39322 6496
rect 0 6354 120 6384
rect 10501 6354 10567 6357
rect 28809 6354 28875 6357
rect 0 6294 6930 6354
rect 0 6264 120 6294
rect 6870 6218 6930 6294
rect 10501 6352 28875 6354
rect 10501 6296 10506 6352
rect 10562 6296 28814 6352
rect 28870 6296 28875 6352
rect 10501 6294 28875 6296
rect 10501 6291 10567 6294
rect 28809 6291 28875 6294
rect 43437 6354 43503 6357
rect 44880 6354 45000 6384
rect 43437 6352 45000 6354
rect 43437 6296 43442 6352
rect 43498 6296 45000 6352
rect 43437 6294 45000 6296
rect 43437 6291 43503 6294
rect 44880 6264 45000 6294
rect 15561 6218 15627 6221
rect 6870 6216 15627 6218
rect 6870 6160 15566 6216
rect 15622 6160 15627 6216
rect 6870 6158 15627 6160
rect 15561 6155 15627 6158
rect 19057 6218 19123 6221
rect 23289 6218 23355 6221
rect 19057 6216 23355 6218
rect 19057 6160 19062 6216
rect 19118 6160 23294 6216
rect 23350 6160 23355 6216
rect 19057 6158 23355 6160
rect 19057 6155 19123 6158
rect 23289 6155 23355 6158
rect 0 6082 120 6112
rect 1761 6082 1827 6085
rect 0 6080 1827 6082
rect 0 6024 1766 6080
rect 1822 6024 1827 6080
rect 0 6022 1827 6024
rect 0 5992 120 6022
rect 1761 6019 1827 6022
rect 43069 6082 43135 6085
rect 44880 6082 45000 6112
rect 43069 6080 45000 6082
rect 43069 6024 43074 6080
rect 43130 6024 45000 6080
rect 43069 6022 45000 6024
rect 43069 6019 43135 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 44880 5992 45000 6022
rect 37946 5951 38262 5952
rect 0 5810 120 5840
rect 16481 5810 16547 5813
rect 0 5808 16547 5810
rect 0 5752 16486 5808
rect 16542 5752 16547 5808
rect 0 5750 16547 5752
rect 0 5720 120 5750
rect 16481 5747 16547 5750
rect 43437 5810 43503 5813
rect 44880 5810 45000 5840
rect 43437 5808 45000 5810
rect 43437 5752 43442 5808
rect 43498 5752 45000 5808
rect 43437 5750 45000 5752
rect 43437 5747 43503 5750
rect 44880 5720 45000 5750
rect 2865 5674 2931 5677
rect 13721 5674 13787 5677
rect 2865 5672 13787 5674
rect 2865 5616 2870 5672
rect 2926 5616 13726 5672
rect 13782 5616 13787 5672
rect 2865 5614 13787 5616
rect 2865 5611 2931 5614
rect 13721 5611 13787 5614
rect 0 5538 120 5568
rect 43069 5538 43135 5541
rect 44880 5538 45000 5568
rect 0 5478 2882 5538
rect 0 5448 120 5478
rect 0 5266 120 5296
rect 2681 5266 2747 5269
rect 0 5264 2747 5266
rect 0 5208 2686 5264
rect 2742 5208 2747 5264
rect 0 5206 2747 5208
rect 2822 5266 2882 5478
rect 43069 5536 45000 5538
rect 43069 5480 43074 5536
rect 43130 5480 45000 5536
rect 43069 5478 45000 5480
rect 43069 5475 43135 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 44880 5448 45000 5478
rect 39006 5407 39322 5408
rect 7833 5266 7899 5269
rect 2822 5264 7899 5266
rect 2822 5208 7838 5264
rect 7894 5208 7899 5264
rect 2822 5206 7899 5208
rect 0 5176 120 5206
rect 2681 5203 2747 5206
rect 7833 5203 7899 5206
rect 23013 5266 23079 5269
rect 43253 5266 43319 5269
rect 23013 5264 43319 5266
rect 23013 5208 23018 5264
rect 23074 5208 43258 5264
rect 43314 5208 43319 5264
rect 23013 5206 43319 5208
rect 23013 5203 23079 5206
rect 43253 5203 43319 5206
rect 43437 5266 43503 5269
rect 44880 5266 45000 5296
rect 43437 5264 45000 5266
rect 43437 5208 43442 5264
rect 43498 5208 45000 5264
rect 43437 5206 45000 5208
rect 43437 5203 43503 5206
rect 44880 5176 45000 5206
rect 17217 5130 17283 5133
rect 1718 5128 17283 5130
rect 1718 5072 17222 5128
rect 17278 5072 17283 5128
rect 1718 5070 17283 5072
rect 0 4994 120 5024
rect 1718 4994 1778 5070
rect 17217 5067 17283 5070
rect 18505 5130 18571 5133
rect 41781 5130 41847 5133
rect 18505 5128 41847 5130
rect 18505 5072 18510 5128
rect 18566 5072 41786 5128
rect 41842 5072 41847 5128
rect 18505 5070 41847 5072
rect 18505 5067 18571 5070
rect 41781 5067 41847 5070
rect 0 4934 1778 4994
rect 2681 4994 2747 4997
rect 7005 4994 7071 4997
rect 2681 4992 7071 4994
rect 2681 4936 2686 4992
rect 2742 4936 7010 4992
rect 7066 4936 7071 4992
rect 2681 4934 7071 4936
rect 0 4904 120 4934
rect 2681 4931 2747 4934
rect 7005 4931 7071 4934
rect 43069 4994 43135 4997
rect 44880 4994 45000 5024
rect 43069 4992 45000 4994
rect 43069 4936 43074 4992
rect 43130 4936 45000 4992
rect 43069 4934 45000 4936
rect 43069 4931 43135 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 44880 4904 45000 4934
rect 37946 4863 38262 4864
rect 0 4722 120 4752
rect 19425 4722 19491 4725
rect 0 4720 19491 4722
rect 0 4664 19430 4720
rect 19486 4664 19491 4720
rect 0 4662 19491 4664
rect 0 4632 120 4662
rect 19425 4659 19491 4662
rect 43437 4722 43503 4725
rect 44880 4722 45000 4752
rect 43437 4720 45000 4722
rect 43437 4664 43442 4720
rect 43498 4664 45000 4720
rect 43437 4662 45000 4664
rect 43437 4659 43503 4662
rect 44880 4632 45000 4662
rect 19333 4586 19399 4589
rect 2822 4584 19399 4586
rect 2822 4528 19338 4584
rect 19394 4528 19399 4584
rect 2822 4526 19399 4528
rect 0 4450 120 4480
rect 2822 4450 2882 4526
rect 19333 4523 19399 4526
rect 0 4390 2882 4450
rect 43069 4450 43135 4453
rect 44880 4450 45000 4480
rect 43069 4448 45000 4450
rect 43069 4392 43074 4448
rect 43130 4392 45000 4448
rect 43069 4390 45000 4392
rect 0 4360 120 4390
rect 43069 4387 43135 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 44880 4360 45000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 20897 4178 20963 4181
rect 0 4176 20963 4178
rect 0 4120 20902 4176
rect 20958 4120 20963 4176
rect 0 4118 20963 4120
rect 0 4088 120 4118
rect 20897 4115 20963 4118
rect 43437 4178 43503 4181
rect 44880 4178 45000 4208
rect 43437 4176 45000 4178
rect 43437 4120 43442 4176
rect 43498 4120 45000 4176
rect 43437 4118 45000 4120
rect 43437 4115 43503 4118
rect 44880 4088 45000 4118
rect 9489 4042 9555 4045
rect 1718 4040 9555 4042
rect 1718 3984 9494 4040
rect 9550 3984 9555 4040
rect 1718 3982 9555 3984
rect 0 3906 120 3936
rect 1718 3906 1778 3982
rect 9489 3979 9555 3982
rect 25865 4042 25931 4045
rect 32581 4042 32647 4045
rect 25865 4040 32647 4042
rect 25865 3984 25870 4040
rect 25926 3984 32586 4040
rect 32642 3984 32647 4040
rect 25865 3982 32647 3984
rect 25865 3979 25931 3982
rect 32581 3979 32647 3982
rect 0 3846 1778 3906
rect 43069 3906 43135 3909
rect 44880 3906 45000 3936
rect 43069 3904 45000 3906
rect 43069 3848 43074 3904
rect 43130 3848 45000 3904
rect 43069 3846 45000 3848
rect 0 3816 120 3846
rect 43069 3843 43135 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 44880 3816 45000 3846
rect 37946 3775 38262 3776
rect 0 3634 120 3664
rect 24853 3634 24919 3637
rect 0 3632 24919 3634
rect 0 3576 24858 3632
rect 24914 3576 24919 3632
rect 0 3574 24919 3576
rect 0 3544 120 3574
rect 24853 3571 24919 3574
rect 43437 3634 43503 3637
rect 44880 3634 45000 3664
rect 43437 3632 45000 3634
rect 43437 3576 43442 3632
rect 43498 3576 45000 3632
rect 43437 3574 45000 3576
rect 43437 3571 43503 3574
rect 44880 3544 45000 3574
rect 23381 3498 23447 3501
rect 2822 3496 23447 3498
rect 2822 3440 23386 3496
rect 23442 3440 23447 3496
rect 2822 3438 23447 3440
rect 0 3362 120 3392
rect 2822 3362 2882 3438
rect 23381 3435 23447 3438
rect 24761 3498 24827 3501
rect 37365 3498 37431 3501
rect 24761 3496 37431 3498
rect 24761 3440 24766 3496
rect 24822 3440 37370 3496
rect 37426 3440 37431 3496
rect 24761 3438 37431 3440
rect 24761 3435 24827 3438
rect 37365 3435 37431 3438
rect 0 3302 2882 3362
rect 43069 3362 43135 3365
rect 44880 3362 45000 3392
rect 43069 3360 45000 3362
rect 43069 3304 43074 3360
rect 43130 3304 45000 3360
rect 43069 3302 45000 3304
rect 0 3272 120 3302
rect 43069 3299 43135 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 44880 3272 45000 3302
rect 39006 3231 39322 3232
rect 0 3090 120 3120
rect 10961 3090 11027 3093
rect 0 3088 11027 3090
rect 0 3032 10966 3088
rect 11022 3032 11027 3088
rect 0 3030 11027 3032
rect 0 3000 120 3030
rect 10961 3027 11027 3030
rect 35801 3090 35867 3093
rect 42885 3090 42951 3093
rect 35801 3088 42951 3090
rect 35801 3032 35806 3088
rect 35862 3032 42890 3088
rect 42946 3032 42951 3088
rect 35801 3030 42951 3032
rect 35801 3027 35867 3030
rect 42885 3027 42951 3030
rect 43437 3090 43503 3093
rect 44880 3090 45000 3120
rect 43437 3088 45000 3090
rect 43437 3032 43442 3088
rect 43498 3032 45000 3088
rect 43437 3030 45000 3032
rect 43437 3027 43503 3030
rect 44880 3000 45000 3030
rect 5533 2954 5599 2957
rect 1718 2952 5599 2954
rect 1718 2896 5538 2952
rect 5594 2896 5599 2952
rect 1718 2894 5599 2896
rect 0 2818 120 2848
rect 1718 2818 1778 2894
rect 5533 2891 5599 2894
rect 20161 2954 20227 2957
rect 37457 2954 37523 2957
rect 20161 2952 37523 2954
rect 20161 2896 20166 2952
rect 20222 2896 37462 2952
rect 37518 2896 37523 2952
rect 20161 2894 37523 2896
rect 20161 2891 20227 2894
rect 37457 2891 37523 2894
rect 0 2758 1778 2818
rect 43069 2818 43135 2821
rect 44880 2818 45000 2848
rect 43069 2816 45000 2818
rect 43069 2760 43074 2816
rect 43130 2760 45000 2816
rect 43069 2758 45000 2760
rect 0 2728 120 2758
rect 43069 2755 43135 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 44880 2728 45000 2758
rect 37946 2687 38262 2688
rect 0 2546 120 2576
rect 9581 2546 9647 2549
rect 0 2544 9647 2546
rect 0 2488 9586 2544
rect 9642 2488 9647 2544
rect 0 2486 9647 2488
rect 0 2456 120 2486
rect 9581 2483 9647 2486
rect 26141 2546 26207 2549
rect 27153 2546 27219 2549
rect 26141 2544 27219 2546
rect 26141 2488 26146 2544
rect 26202 2488 27158 2544
rect 27214 2488 27219 2544
rect 26141 2486 27219 2488
rect 26141 2483 26207 2486
rect 27153 2483 27219 2486
rect 43437 2546 43503 2549
rect 44880 2546 45000 2576
rect 43437 2544 45000 2546
rect 43437 2488 43442 2544
rect 43498 2488 45000 2544
rect 43437 2486 45000 2488
rect 43437 2483 43503 2486
rect 44880 2456 45000 2486
rect 11881 2410 11947 2413
rect 28533 2410 28599 2413
rect 11881 2408 28599 2410
rect 11881 2352 11886 2408
rect 11942 2352 28538 2408
rect 28594 2352 28599 2408
rect 11881 2350 28599 2352
rect 11881 2347 11947 2350
rect 28533 2347 28599 2350
rect 0 2274 120 2304
rect 2865 2274 2931 2277
rect 0 2272 2931 2274
rect 0 2216 2870 2272
rect 2926 2216 2931 2272
rect 0 2214 2931 2216
rect 0 2184 120 2214
rect 2865 2211 2931 2214
rect 43069 2274 43135 2277
rect 44880 2274 45000 2304
rect 43069 2272 45000 2274
rect 43069 2216 43074 2272
rect 43130 2216 45000 2272
rect 43069 2214 45000 2216
rect 43069 2211 43135 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 44880 2184 45000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 20713 2002 20779 2005
rect 0 2000 20779 2002
rect 0 1944 20718 2000
rect 20774 1944 20779 2000
rect 0 1942 20779 1944
rect 0 1912 120 1942
rect 20713 1939 20779 1942
rect 42977 2002 43043 2005
rect 44880 2002 45000 2032
rect 42977 2000 45000 2002
rect 42977 1944 42982 2000
rect 43038 1944 45000 2000
rect 42977 1942 45000 1944
rect 42977 1939 43043 1942
rect 44880 1912 45000 1942
rect 2865 1866 2931 1869
rect 20345 1866 20411 1869
rect 2865 1864 20411 1866
rect 2865 1808 2870 1864
rect 2926 1808 20350 1864
rect 20406 1808 20411 1864
rect 2865 1806 20411 1808
rect 2865 1803 2931 1806
rect 20345 1803 20411 1806
rect 0 1730 120 1760
rect 9489 1730 9555 1733
rect 0 1728 9555 1730
rect 0 1672 9494 1728
rect 9550 1672 9555 1728
rect 0 1670 9555 1672
rect 0 1640 120 1670
rect 9489 1667 9555 1670
rect 42149 1730 42215 1733
rect 44880 1730 45000 1760
rect 42149 1728 45000 1730
rect 42149 1672 42154 1728
rect 42210 1672 45000 1728
rect 42149 1670 45000 1672
rect 42149 1667 42215 1670
rect 44880 1640 45000 1670
rect 0 1458 120 1488
rect 9397 1458 9463 1461
rect 0 1456 9463 1458
rect 0 1400 9402 1456
rect 9458 1400 9463 1456
rect 0 1398 9463 1400
rect 0 1368 120 1398
rect 9397 1395 9463 1398
rect 42701 1458 42767 1461
rect 44880 1458 45000 1488
rect 42701 1456 45000 1458
rect 42701 1400 42706 1456
rect 42762 1400 45000 1456
rect 42701 1398 45000 1400
rect 42701 1395 42767 1398
rect 44880 1368 45000 1398
<< via3 >>
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__clkbuf_2  _000_
timestamp -3599
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _001_
timestamp -3599
transform 1 0 17940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp -3599
transform -1 0 20976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp -3599
transform -1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _004_
timestamp -3599
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _005_
timestamp -3599
transform 1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _006_
timestamp -3599
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _007_
timestamp -3599
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _008_
timestamp -3599
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _009_
timestamp -3599
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _010_
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _011_
timestamp -3599
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _012_
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _013_
timestamp -3599
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _014_
timestamp -3599
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _015_
timestamp -3599
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _016_
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _017_
timestamp -3599
transform 1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _018_
timestamp -3599
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _019_
timestamp -3599
transform 1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _020_
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _021_
timestamp -3599
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _022_
timestamp -3599
transform 1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp -3599
transform -1 0 23092 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _024_
timestamp -3599
transform 1 0 27048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _025_
timestamp -3599
transform 1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _026_
timestamp -3599
transform 1 0 26588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _027_
timestamp -3599
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _028_
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _029_
timestamp -3599
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _030_
timestamp -3599
transform 1 0 22172 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _031_
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp -3599
transform -1 0 26680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _033_
timestamp -3599
transform 1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _034_
timestamp -3599
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _035_
timestamp -3599
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _036_
timestamp -3599
transform 1 0 28520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp -3599
transform -1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp -3599
transform 1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp -3599
transform 1 0 40664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp -3599
transform 1 0 38548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp -3599
transform -1 0 36800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp -3599
transform 1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _043_
timestamp -3599
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _044_
timestamp -3599
transform 1 0 24472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp -3599
transform -1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp -3599
transform -1 0 31556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp -3599
transform -1 0 33764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp -3599
transform -1 0 35328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp -3599
transform -1 0 36708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp -3599
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp -3599
transform 1 0 40664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp -3599
transform -1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp -3599
transform -1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp -3599
transform -1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp -3599
transform -1 0 5060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp -3599
transform -1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp -3599
transform -1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp -3599
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp -3599
transform 1 0 6992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp -3599
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp -3599
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp -3599
transform 1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp -3599
transform -1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp -3599
transform -1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp -3599
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp -3599
transform 1 0 9476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp -3599
transform 1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp -3599
transform 1 0 15824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp -3599
transform 1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _072_
timestamp -3599
transform -1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _073_
timestamp -3599
transform -1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp -3599
transform -1 0 10764 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform -1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp -3599
transform -1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp -3599
transform 1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp -3599
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp -3599
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp -3599
transform 1 0 15364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp -3599
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp -3599
transform 1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp -3599
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp -3599
transform 1 0 22448 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp -3599
transform 1 0 39284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp -3599
transform -1 0 37076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp -3599
transform -1 0 35420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp -3599
transform -1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp -3599
transform -1 0 33304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _093_
timestamp -3599
transform -1 0 32660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _094_
timestamp -3599
transform -1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _095_
timestamp -3599
transform -1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform -1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform -1 0 29348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp -3599
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp -3599
transform 1 0 26772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform 1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp -3599
transform -1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp -3599
transform -1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp -3599
transform 1 0 32200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform 1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 24840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 22632 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 22264 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform 1 0 17204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 17204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 25300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 20424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 18124 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 27876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 26404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform 1 0 23828 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 24840 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform -1 0 21160 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 21988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp -3599
transform 1 0 28612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp -3599
transform 1 0 20240 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp -3599
transform -1 0 27416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp -3599
transform -1 0 23920 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp -3599
transform 1 0 24840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp -3599
transform -1 0 21988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp -3599
transform -1 0 4784 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp -3599
transform 1 0 4140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp -3599
transform -1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp -3599
transform -1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp -3599
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp -3599
transform -1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp -3599
transform -1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp -3599
transform -1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636964856
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636964856
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636964856
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636964856
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp -3599
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636964856
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp -3599
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_441
timestamp -3599
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_449
timestamp -3599
transform 1 0 42412 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp -3599
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_89
timestamp -3599
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_96
timestamp 1636964856
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp -3599
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_137
timestamp -3599
transform 1 0 13708 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1636964856
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp -3599
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_175
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_186
timestamp 1636964856
transform 1 0 18216 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_198
timestamp -3599
transform 1 0 19320 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_204
timestamp -3599
transform 1 0 19872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp -3599
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636964856
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_237
timestamp -3599
transform 1 0 22908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_245
timestamp -3599
transform 1 0 23644 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_251
timestamp -3599
transform 1 0 24196 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_259
timestamp -3599
transform 1 0 24932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_266
timestamp 1636964856
transform 1 0 25576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp -3599
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_294
timestamp -3599
transform 1 0 28152 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_301
timestamp 1636964856
transform 1 0 28796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_313
timestamp -3599
transform 1 0 29900 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_321
timestamp -3599
transform 1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp -3599
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636964856
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636964856
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636964856
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636964856
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636964856
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636964856
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp -3599
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp -3599
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_449
timestamp -3599
transform 1 0 42412 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636964856
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_165
timestamp -3599
transform 1 0 16284 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp -3599
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp -3599
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp -3599
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp -3599
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636964856
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636964856
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636964856
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_233
timestamp -3599
transform 1 0 22540 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_240
timestamp 1636964856
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp -3599
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_263
timestamp 1636964856
transform 1 0 25300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_275
timestamp 1636964856
transform 1 0 26404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_287
timestamp 1636964856
transform 1 0 27508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp -3599
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -3599
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636964856
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636964856
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636964856
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636964856
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_368
timestamp 1636964856
transform 1 0 34960 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_380
timestamp 1636964856
transform 1 0 36064 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_392
timestamp 1636964856
transform 1 0 37168 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_404
timestamp 1636964856
transform 1 0 38272 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp -3599
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636964856
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636964856
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_445
timestamp -3599
transform 1 0 42044 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_453
timestamp -3599
transform 1 0 42780 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636964856
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp -3599
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636964856
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636964856
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636964856
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636964856
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp -3599
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_230
timestamp -3599
transform 1 0 22264 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_239
timestamp 1636964856
transform 1 0 23092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1636964856
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp -3599
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_270
timestamp -3599
transform 1 0 25944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp -3599
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636964856
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636964856
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp -3599
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_361
timestamp -3599
transform 1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_372
timestamp 1636964856
transform 1 0 35328 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_384
timestamp -3599
transform 1 0 36432 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636964856
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636964856
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_429
timestamp -3599
transform 1 0 40572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_433
timestamp 1636964856
transform 1 0 40940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_445
timestamp -3599
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp -3599
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_453
timestamp -3599
transform 1 0 42780 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_88
timestamp 1636964856
transform 1 0 9200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_100
timestamp 1636964856
transform 1 0 10304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_112
timestamp 1636964856
transform 1 0 11408 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_124
timestamp 1636964856
transform 1 0 12512 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp -3599
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636964856
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636964856
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636964856
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_229
timestamp -3599
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_237
timestamp 1636964856
transform 1 0 22908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp -3599
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636964856
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636964856
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636964856
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp -3599
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636964856
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp -3599
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_327
timestamp -3599
transform 1 0 31188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_331
timestamp -3599
transform 1 0 31556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_337
timestamp -3599
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_342
timestamp -3599
transform 1 0 32568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_350
timestamp -3599
transform 1 0 33304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp -3599
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp -3599
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_377
timestamp -3599
transform 1 0 35788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_383
timestamp -3599
transform 1 0 36340 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_387
timestamp 1636964856
transform 1 0 36708 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_399
timestamp -3599
transform 1 0 37812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_410
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp -3599
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636964856
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636964856
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_445
timestamp -3599
transform 1 0 42044 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_453
timestamp -3599
transform 1 0 42780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636964856
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636964856
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp -3599
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_100
timestamp 1636964856
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp -3599
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1636964856
transform 1 0 13156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_143
timestamp 1636964856
transform 1 0 14260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1636964856
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636964856
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp -3599
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp -3599
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636964856
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp -3599
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_253
timestamp -3599
transform 1 0 24380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_257
timestamp 1636964856
transform 1 0 24748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp -3599
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp -3599
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_285
timestamp 1636964856
transform 1 0 27324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_297
timestamp -3599
transform 1 0 28428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp -3599
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_311
timestamp 1636964856
transform 1 0 29716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_323
timestamp 1636964856
transform 1 0 30820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636964856
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636964856
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636964856
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp -3599
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp -3599
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp -3599
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_453
timestamp -3599
transform 1 0 42780 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_37
timestamp -3599
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_43
timestamp 1636964856
transform 1 0 5060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_55
timestamp 1636964856
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_67
timestamp 1636964856
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp -3599
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636964856
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_112
timestamp 1636964856
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_124
timestamp 1636964856
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636964856
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636964856
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636964856
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636964856
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636964856
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636964856
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_230
timestamp 1636964856
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_242
timestamp -3599
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp -3599
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636964856
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp -3599
transform 1 0 26220 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_278
timestamp 1636964856
transform 1 0 26680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_290
timestamp 1636964856
transform 1 0 27784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp -3599
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636964856
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636964856
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636964856
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636964856
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636964856
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636964856
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_413
timestamp -3599
transform 1 0 39100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp -3599
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636964856
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636964856
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_445
timestamp -3599
transform 1 0 42044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_453
timestamp -3599
transform 1 0 42780 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636964856
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636964856
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636964856
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636964856
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_83
timestamp -3599
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_88
timestamp -3599
transform 1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_94
timestamp -3599
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp -3599
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_128
timestamp 1636964856
transform 1 0 12880 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_140
timestamp 1636964856
transform 1 0 13984 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_152
timestamp -3599
transform 1 0 15088 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp -3599
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636964856
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp -3599
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_200
timestamp 1636964856
transform 1 0 19504 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1636964856
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636964856
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636964856
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636964856
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636964856
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636964856
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636964856
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636964856
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp -3599
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636964856
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636964856
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636964856
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636964856
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp -3599
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp -3599
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_449
timestamp -3599
transform 1 0 42412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_453
timestamp -3599
transform 1 0 42780 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_35
timestamp 1636964856
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_47
timestamp -3599
transform 1 0 5428 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_53
timestamp -3599
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp -3599
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_67
timestamp -3599
transform 1 0 7268 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp -3599
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_95
timestamp 1636964856
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_107
timestamp 1636964856
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_119
timestamp 1636964856
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp -3599
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636964856
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636964856
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636964856
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp -3599
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_207
timestamp 1636964856
transform 1 0 20148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_219
timestamp -3599
transform 1 0 21252 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_227
timestamp -3599
transform 1 0 21988 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_232
timestamp 1636964856
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp -3599
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_258
timestamp 1636964856
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp -3599
transform 1 0 25944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp -3599
transform 1 0 26312 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_280
timestamp 1636964856
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_292
timestamp 1636964856
transform 1 0 27968 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636964856
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636964856
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_345
timestamp -3599
transform 1 0 32844 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_350
timestamp 1636964856
transform 1 0 33304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp -3599
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_368
timestamp 1636964856
transform 1 0 34960 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_380
timestamp 1636964856
transform 1 0 36064 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_392
timestamp 1636964856
transform 1 0 37168 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_404
timestamp 1636964856
transform 1 0 38272 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp -3599
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_421
timestamp -3599
transform 1 0 39836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_429
timestamp -3599
transform 1 0 40572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636964856
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_445
timestamp -3599
transform 1 0 42044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_453
timestamp -3599
transform 1 0 42780 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636964856
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_27
timestamp -3599
transform 1 0 3588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_39
timestamp -3599
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_47
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp -3599
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636964856
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636964856
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636964856
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp -3599
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp -3599
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_128
timestamp 1636964856
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_140
timestamp -3599
transform 1 0 13984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_148
timestamp -3599
transform 1 0 14720 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp -3599
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp -3599
transform 1 0 15640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp -3599
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636964856
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636964856
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636964856
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp -3599
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_228
timestamp 1636964856
transform 1 0 22080 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1636964856
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_252
timestamp -3599
transform 1 0 24288 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_263
timestamp 1636964856
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_324
timestamp -3599
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_330
timestamp -3599
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_337
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_343
timestamp 1636964856
transform 1 0 32660 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_355
timestamp 1636964856
transform 1 0 33764 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_367
timestamp -3599
transform 1 0 34868 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636964856
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636964856
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp -3599
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_410
timestamp 1636964856
transform 1 0 38824 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_422
timestamp 1636964856
transform 1 0 39928 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_434
timestamp 1636964856
transform 1 0 41032 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp -3599
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_449
timestamp -3599
transform 1 0 42412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_453
timestamp -3599
transform 1 0 42780 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636964856
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636964856
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636964856
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_54
timestamp -3599
transform 1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp -3599
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_66
timestamp -3599
transform 1 0 7176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp -3599
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_102
timestamp -3599
transform 1 0 10488 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_114
timestamp -3599
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp -3599
transform 1 0 12144 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp -3599
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp -3599
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp -3599
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp -3599
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_180
timestamp -3599
transform 1 0 17664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_205
timestamp -3599
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_218
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_226
timestamp -3599
transform 1 0 21896 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_235
timestamp 1636964856
transform 1 0 22724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_258
timestamp 1636964856
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_270
timestamp -3599
transform 1 0 25944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_276
timestamp -3599
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_282
timestamp -3599
transform 1 0 27048 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_286
timestamp 1636964856
transform 1 0 27416 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp -3599
transform 1 0 28520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_309
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_313
timestamp -3599
transform 1 0 29900 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_317
timestamp 1636964856
transform 1 0 30268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_329
timestamp 1636964856
transform 1 0 31372 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_341
timestamp 1636964856
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp -3599
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp -3599
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1636964856
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_377
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_399
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp -3599
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_425
timestamp 1636964856
transform 1 0 40204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_437
timestamp -3599
transform 1 0 41308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_445
timestamp -3599
transform 1 0 42044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636964856
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636964856
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_29
timestamp 1636964856
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_41
timestamp -3599
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_208
timestamp 1636964856
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp -3599
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636964856
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636964856
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_249
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_253
timestamp 1636964856
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_265
timestamp 1636964856
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp -3599
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636964856
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1636964856
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_305
timestamp -3599
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_309
timestamp 1636964856
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_321
timestamp 1636964856
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp -3599
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1636964856
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_349
timestamp -3599
transform 1 0 33212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_357
timestamp -3599
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_417
timestamp -3599
transform 1 0 39468 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_429
timestamp -3599
transform 1 0 40572 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_437
timestamp -3599
transform 1 0 41308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_449
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output1
timestamp -3599
transform 1 0 42504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp -3599
transform 1 0 43240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp -3599
transform 1 0 42872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform 1 0 43240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform 1 0 42872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 43240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 42872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 43240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 42872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 43240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform 1 0 42872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp -3599
transform 1 0 43240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -3599
transform 1 0 43240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -3599
transform 1 0 42872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -3599
transform 1 0 43240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -3599
transform 1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -3599
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -3599
transform 1 0 42504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -3599
transform 1 0 41952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -3599
transform 1 0 42504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -3599
transform 1 0 42872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp -3599
transform 1 0 42504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp -3599
transform 1 0 42136 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp -3599
transform 1 0 41584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp -3599
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp -3599
transform 1 0 43240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp -3599
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp -3599
transform 1 0 43240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp -3599
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp -3599
transform 1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp -3599
transform 1 0 42872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp -3599
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp -3599
transform 1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp -3599
transform 1 0 39100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp -3599
transform 1 0 38548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp -3599
transform 1 0 38916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp -3599
transform 1 0 39836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp -3599
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp -3599
transform -1 0 40204 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp -3599
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp -3599
transform 1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp -3599
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp -3599
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp -3599
transform -1 0 36432 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp -3599
transform -1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp -3599
transform -1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp -3599
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp -3599
transform 1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform 1 0 5704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 6624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform -1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform -1 0 8832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform -1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform -1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform -1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform -1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform -1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform -1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 13800 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 18400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform -1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output105
timestamp -3599
transform -1 0 34408 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_59
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_73
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_86
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_91
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_92
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_93
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_94
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_95
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_96
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_97
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_98
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_106
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_110
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_130
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_131
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 44880 1368 45000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 44880 4088 45000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 44880 4360 45000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 44880 4632 45000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 44880 4904 45000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 44880 5176 45000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 44880 5448 45000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 44880 5720 45000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 44880 5992 45000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 44880 6264 45000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 44880 6536 45000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 44880 1640 45000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 44880 6808 45000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 44880 7080 45000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 44880 7352 45000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 44880 7624 45000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 44880 7896 45000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 44880 8168 45000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 44880 8440 45000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 44880 8712 45000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 44880 8984 45000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 44880 9256 45000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 44880 1912 45000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 44880 9528 45000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 44880 9800 45000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 44880 2184 45000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 44880 2456 45000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 44880 2728 45000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 44880 3000 45000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 44880 3272 45000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 44880 3544 45000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 44880 3816 45000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 3422 0 3478 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 24582 0 24638 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 26698 0 26754 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 28814 0 28870 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 30930 0 30986 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 33046 0 33102 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 35162 0 35218 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 37278 0 37334 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 39394 0 39450 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 41510 0 41566 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 43626 0 43682 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 5538 0 5594 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 7654 0 7710 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 9770 0 9826 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 11886 0 11942 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 14002 0 14058 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 16118 0 16174 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 18234 0 18290 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 20350 0 20406 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 22466 0 22522 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 34334 11194 34390 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 37094 11194 37150 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 37370 11194 37426 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 37646 11194 37702 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 37922 11194 37978 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 38198 11194 38254 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 38474 11194 38530 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 38750 11194 38806 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 39026 11194 39082 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 39302 11194 39358 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 39578 11194 39634 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 34610 11194 34666 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 34886 11194 34942 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 35162 11194 35218 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 35438 11194 35494 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 35714 11194 35770 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 35990 11194 36046 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 36266 11194 36322 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 36542 11194 36598 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 36818 11194 36874 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 5354 11194 5410 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 5630 11194 5686 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 5906 11194 5962 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 6182 11194 6238 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 6458 11194 6514 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 6734 11194 6790 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 7010 11194 7066 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 7286 11194 7342 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 7562 11194 7618 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 7838 11194 7894 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 8114 11194 8170 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 8390 11194 8446 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 8666 11194 8722 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 8942 11194 8998 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 9218 11194 9274 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 9494 11194 9550 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 9770 11194 9826 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 10046 11194 10102 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 10322 11194 10378 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 10598 11194 10654 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 10874 11194 10930 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 13634 11194 13690 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 13910 11194 13966 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 14186 11194 14242 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 14462 11194 14518 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 14738 11194 14794 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 15014 11194 15070 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 11150 11194 11206 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 11426 11194 11482 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 11702 11194 11758 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 11978 11194 12034 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 12254 11194 12310 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 12530 11194 12586 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 12806 11194 12862 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 13082 11194 13138 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 13358 11194 13414 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 15290 11194 15346 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 18050 11194 18106 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 18326 11194 18382 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 18602 11194 18658 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 18878 11194 18934 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 19154 11194 19210 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 19430 11194 19486 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 15566 11194 15622 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 15842 11194 15898 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 16118 11194 16174 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 16394 11194 16450 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 16670 11194 16726 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 16946 11194 17002 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 17222 11194 17278 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 17498 11194 17554 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 17774 11194 17830 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 19706 11194 19762 11250 0 FreeSans 224 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 19982 11194 20038 11250 0 FreeSans 224 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 20258 11194 20314 11250 0 FreeSans 224 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 20534 11194 20590 11250 0 FreeSans 224 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 23018 11194 23074 11250 0 FreeSans 224 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 23294 11194 23350 11250 0 FreeSans 224 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 23570 11194 23626 11250 0 FreeSans 224 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 23846 11194 23902 11250 0 FreeSans 224 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 24122 11194 24178 11250 0 FreeSans 224 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 24398 11194 24454 11250 0 FreeSans 224 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 24674 11194 24730 11250 0 FreeSans 224 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 24950 11194 25006 11250 0 FreeSans 224 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 20810 11194 20866 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 21086 11194 21142 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 21362 11194 21418 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 21638 11194 21694 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 21914 11194 21970 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 22190 11194 22246 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 22466 11194 22522 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 22742 11194 22798 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 25226 11194 25282 11250 0 FreeSans 224 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 27986 11194 28042 11250 0 FreeSans 224 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 28262 11194 28318 11250 0 FreeSans 224 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 28538 11194 28594 11250 0 FreeSans 224 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 28814 11194 28870 11250 0 FreeSans 224 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 29090 11194 29146 11250 0 FreeSans 224 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 29366 11194 29422 11250 0 FreeSans 224 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 25502 11194 25558 11250 0 FreeSans 224 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 25778 11194 25834 11250 0 FreeSans 224 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 26054 11194 26110 11250 0 FreeSans 224 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 26330 11194 26386 11250 0 FreeSans 224 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 26606 11194 26662 11250 0 FreeSans 224 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 26882 11194 26938 11250 0 FreeSans 224 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 27158 11194 27214 11250 0 FreeSans 224 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 27434 11194 27490 11250 0 FreeSans 224 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 27710 11194 27766 11250 0 FreeSans 224 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 29642 11194 29698 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 32402 11194 32458 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 32678 11194 32734 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 32954 11194 33010 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 33230 11194 33286 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 33506 11194 33562 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 33782 11194 33838 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 29918 11194 29974 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 30194 11194 30250 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 30470 11194 30526 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 30746 11194 30802 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 31022 11194 31078 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 31298 11194 31354 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 31574 11194 31630 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 31850 11194 31906 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 32126 11194 32182 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1306 0 1362 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 34058 11194 34114 11250 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 210 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 211 nsew power bidirectional
rlabel metal1 22494 8704 22494 8704 0 VGND
rlabel metal1 22494 8160 22494 8160 0 VPWR
rlabel metal1 10580 2890 10580 2890 0 FrameData[0]
rlabel metal2 20930 5287 20930 5287 0 FrameData[10]
rlabel metal3 1471 4420 1471 4420 0 FrameData[11]
rlabel metal2 19458 4403 19458 4403 0 FrameData[12]
rlabel metal3 919 4964 919 4964 0 FrameData[13]
rlabel metal3 1402 5236 1402 5236 0 FrameData[14]
rlabel metal3 1471 5508 1471 5508 0 FrameData[15]
rlabel metal1 16652 3094 16652 3094 0 FrameData[16]
rlabel metal3 942 6052 942 6052 0 FrameData[17]
rlabel metal3 3495 6324 3495 6324 0 FrameData[18]
rlabel metal3 1494 6596 1494 6596 0 FrameData[19]
rlabel metal2 9522 2261 9522 2261 0 FrameData[1]
rlabel metal2 18630 6375 18630 6375 0 FrameData[20]
rlabel metal3 942 7140 942 7140 0 FrameData[21]
rlabel metal3 712 7412 712 7412 0 FrameData[22]
rlabel metal3 620 7684 620 7684 0 FrameData[23]
rlabel metal3 666 7956 666 7956 0 FrameData[24]
rlabel metal3 942 8228 942 8228 0 FrameData[25]
rlabel metal1 26404 6834 26404 6834 0 FrameData[26]
rlabel metal3 1494 8772 1494 8772 0 FrameData[27]
rlabel metal2 24426 8449 24426 8449 0 FrameData[28]
rlabel metal2 20746 8687 20746 8687 0 FrameData[29]
rlabel metal3 10418 1972 10418 1972 0 FrameData[2]
rlabel metal2 22126 8823 22126 8823 0 FrameData[30]
rlabel metal2 28658 8160 28658 8160 0 FrameData[31]
rlabel metal3 1494 2244 1494 2244 0 FrameData[3]
rlabel metal2 9614 2941 9614 2941 0 FrameData[4]
rlabel metal3 919 2788 919 2788 0 FrameData[5]
rlabel metal2 10994 2703 10994 2703 0 FrameData[6]
rlabel metal3 1471 3332 1471 3332 0 FrameData[7]
rlabel via2 24886 3587 24886 3587 0 FrameData[8]
rlabel metal3 919 3876 919 3876 0 FrameData[9]
rlabel metal3 43822 1428 43822 1428 0 FrameData_O[0]
rlabel metal3 44190 4148 44190 4148 0 FrameData_O[10]
rlabel metal3 44006 4420 44006 4420 0 FrameData_O[11]
rlabel metal3 44190 4692 44190 4692 0 FrameData_O[12]
rlabel metal3 44006 4964 44006 4964 0 FrameData_O[13]
rlabel metal3 44190 5236 44190 5236 0 FrameData_O[14]
rlabel metal3 44006 5508 44006 5508 0 FrameData_O[15]
rlabel metal3 44190 5780 44190 5780 0 FrameData_O[16]
rlabel metal3 44006 6052 44006 6052 0 FrameData_O[17]
rlabel metal3 44190 6324 44190 6324 0 FrameData_O[18]
rlabel metal3 44006 6596 44006 6596 0 FrameData_O[19]
rlabel metal3 43546 1700 43546 1700 0 FrameData_O[1]
rlabel metal3 44190 6868 44190 6868 0 FrameData_O[20]
rlabel metal3 44190 7140 44190 7140 0 FrameData_O[21]
rlabel metal3 44006 7412 44006 7412 0 FrameData_O[22]
rlabel metal3 44190 7684 44190 7684 0 FrameData_O[23]
rlabel metal3 44190 7956 44190 7956 0 FrameData_O[24]
rlabel metal3 44006 8228 44006 8228 0 FrameData_O[25]
rlabel metal3 43822 8500 43822 8500 0 FrameData_O[26]
rlabel metal2 42182 8687 42182 8687 0 FrameData_O[27]
rlabel metal1 42688 8058 42688 8058 0 FrameData_O[28]
rlabel metal1 43148 7514 43148 7514 0 FrameData_O[29]
rlabel metal3 43960 1972 43960 1972 0 FrameData_O[2]
rlabel metal2 42366 8823 42366 8823 0 FrameData_O[30]
rlabel metal2 41814 9231 41814 9231 0 FrameData_O[31]
rlabel metal3 44006 2244 44006 2244 0 FrameData_O[3]
rlabel metal3 44190 2516 44190 2516 0 FrameData_O[4]
rlabel metal3 44006 2788 44006 2788 0 FrameData_O[5]
rlabel metal3 44190 3060 44190 3060 0 FrameData_O[6]
rlabel metal3 44006 3332 44006 3332 0 FrameData_O[7]
rlabel metal3 44190 3604 44190 3604 0 FrameData_O[8]
rlabel metal3 44006 3876 44006 3876 0 FrameData_O[9]
rlabel metal2 3450 106 3450 106 0 FrameStrobe[0]
rlabel metal1 25162 4114 25162 4114 0 FrameStrobe[10]
rlabel metal2 20010 3366 20010 3366 0 FrameStrobe[11]
rlabel metal1 26680 4998 26680 4998 0 FrameStrobe[12]
rlabel metal1 30222 5202 30222 5202 0 FrameStrobe[13]
rlabel metal2 33074 55 33074 55 0 FrameStrobe[14]
rlabel metal1 34362 4590 34362 4590 0 FrameStrobe[15]
rlabel metal1 36202 4114 36202 4114 0 FrameStrobe[16]
rlabel metal1 37950 4658 37950 4658 0 FrameStrobe[17]
rlabel metal1 40066 4590 40066 4590 0 FrameStrobe[18]
rlabel metal1 40894 4080 40894 4080 0 FrameStrobe[19]
rlabel metal2 5566 1075 5566 1075 0 FrameStrobe[1]
rlabel metal2 7682 1806 7682 1806 0 FrameStrobe[2]
rlabel metal1 9752 7854 9752 7854 0 FrameStrobe[3]
rlabel metal2 11914 1211 11914 1211 0 FrameStrobe[4]
rlabel metal2 14030 174 14030 174 0 FrameStrobe[5]
rlabel metal2 16146 123 16146 123 0 FrameStrobe[6]
rlabel metal2 18262 140 18262 140 0 FrameStrobe[7]
rlabel metal2 20378 208 20378 208 0 FrameStrobe[8]
rlabel metal2 22494 3166 22494 3166 0 FrameStrobe[9]
rlabel metal1 34638 8602 34638 8602 0 FrameStrobe_O[0]
rlabel metal1 38226 8364 38226 8364 0 FrameStrobe_O[10]
rlabel metal1 37536 8058 37536 8058 0 FrameStrobe_O[11]
rlabel metal1 38134 8602 38134 8602 0 FrameStrobe_O[12]
rlabel metal1 38778 8330 38778 8330 0 FrameStrobe_O[13]
rlabel metal1 39330 8364 39330 8364 0 FrameStrobe_O[14]
rlabel metal1 38640 8058 38640 8058 0 FrameStrobe_O[15]
rlabel metal1 39008 8058 39008 8058 0 FrameStrobe_O[16]
rlabel metal1 39514 8602 39514 8602 0 FrameStrobe_O[17]
rlabel metal1 39928 8330 39928 8330 0 FrameStrobe_O[18]
rlabel metal1 39790 8058 39790 8058 0 FrameStrobe_O[19]
rlabel metal2 35282 8840 35282 8840 0 FrameStrobe_O[1]
rlabel metal1 35650 8568 35650 8568 0 FrameStrobe_O[2]
rlabel metal1 35926 8602 35926 8602 0 FrameStrobe_O[3]
rlabel metal1 36386 8568 36386 8568 0 FrameStrobe_O[4]
rlabel metal2 36754 8704 36754 8704 0 FrameStrobe_O[5]
rlabel metal1 36110 8058 36110 8058 0 FrameStrobe_O[6]
rlabel metal1 36432 8058 36432 8058 0 FrameStrobe_O[7]
rlabel metal1 36984 8602 36984 8602 0 FrameStrobe_O[8]
rlabel metal1 37352 8330 37352 8330 0 FrameStrobe_O[9]
rlabel metal2 5382 9904 5382 9904 0 N1BEG[0]
rlabel metal1 5796 8058 5796 8058 0 N1BEG[1]
rlabel metal1 5842 8602 5842 8602 0 N1BEG[2]
rlabel metal1 6348 8058 6348 8058 0 N1BEG[3]
rlabel metal1 6302 8602 6302 8602 0 N2BEG[0]
rlabel metal2 6762 9632 6762 9632 0 N2BEG[1]
rlabel metal2 7038 9904 7038 9904 0 N2BEG[2]
rlabel metal1 7268 8602 7268 8602 0 N2BEG[3]
rlabel metal1 7544 8602 7544 8602 0 N2BEG[4]
rlabel metal1 7912 8058 7912 8058 0 N2BEG[5]
rlabel metal1 8004 8602 8004 8602 0 N2BEG[6]
rlabel metal1 8510 8058 8510 8058 0 N2BEG[7]
rlabel metal1 8510 8602 8510 8602 0 N2BEGb[0]
rlabel metal1 8740 8330 8740 8330 0 N2BEGb[1]
rlabel metal2 9430 8755 9430 8755 0 N2BEGb[2]
rlabel metal1 9430 8602 9430 8602 0 N2BEGb[3]
rlabel metal1 9752 8602 9752 8602 0 N2BEGb[4]
rlabel metal1 10166 8058 10166 8058 0 N2BEGb[5]
rlabel metal1 10212 8602 10212 8602 0 N2BEGb[6]
rlabel metal1 10534 8602 10534 8602 0 N2BEGb[7]
rlabel metal1 10856 8602 10856 8602 0 N4BEG[0]
rlabel metal1 13524 8602 13524 8602 0 N4BEG[10]
rlabel metal1 14030 8058 14030 8058 0 N4BEG[11]
rlabel metal1 13984 8602 13984 8602 0 N4BEG[12]
rlabel metal1 14582 8058 14582 8058 0 N4BEG[13]
rlabel metal1 14628 8602 14628 8602 0 N4BEG[14]
rlabel metal1 14904 8602 14904 8602 0 N4BEG[15]
rlabel metal1 11270 8058 11270 8058 0 N4BEG[1]
rlabel metal1 11362 8602 11362 8602 0 N4BEG[2]
rlabel metal1 11868 8058 11868 8058 0 N4BEG[3]
rlabel metal2 12006 9904 12006 9904 0 N4BEG[4]
rlabel metal2 12282 9632 12282 9632 0 N4BEG[5]
rlabel metal2 12558 9904 12558 9904 0 N4BEG[6]
rlabel metal1 12742 8602 12742 8602 0 N4BEG[7]
rlabel metal1 13064 8602 13064 8602 0 N4BEG[8]
rlabel metal1 13478 8058 13478 8058 0 N4BEG[9]
rlabel metal1 15318 8602 15318 8602 0 NN4BEG[0]
rlabel metal1 17940 8602 17940 8602 0 NN4BEG[10]
rlabel metal1 18262 8602 18262 8602 0 NN4BEG[11]
rlabel metal1 18584 8602 18584 8602 0 NN4BEG[12]
rlabel metal2 18906 9904 18906 9904 0 NN4BEG[13]
rlabel metal1 19642 8330 19642 8330 0 NN4BEG[14]
rlabel metal1 19596 8602 19596 8602 0 NN4BEG[15]
rlabel metal1 15778 8058 15778 8058 0 NN4BEG[1]
rlabel metal1 15732 8602 15732 8602 0 NN4BEG[2]
rlabel metal1 16054 8602 16054 8602 0 NN4BEG[3]
rlabel metal1 16514 8058 16514 8058 0 NN4BEG[4]
rlabel metal2 16330 8704 16330 8704 0 NN4BEG[5]
rlabel metal1 17066 8058 17066 8058 0 NN4BEG[6]
rlabel metal1 17158 8602 17158 8602 0 NN4BEG[7]
rlabel metal1 17480 8602 17480 8602 0 NN4BEG[8]
rlabel metal1 17894 8058 17894 8058 0 NN4BEG[9]
rlabel metal1 4784 5678 4784 5678 0 S1END[0]
rlabel metal1 4048 6766 4048 6766 0 S1END[1]
rlabel metal1 4186 7412 4186 7412 0 S1END[2]
rlabel metal1 4462 7344 4462 7344 0 S1END[3]
rlabel metal2 23046 9020 23046 9020 0 S2END[0]
rlabel metal2 19090 6239 19090 6239 0 S2END[1]
rlabel metal1 13110 5168 13110 5168 0 S2END[2]
rlabel metal2 18722 5678 18722 5678 0 S2END[3]
rlabel metal2 10166 8551 10166 8551 0 S2END[4]
rlabel metal1 9706 6256 9706 6256 0 S2END[5]
rlabel metal2 9154 5916 9154 5916 0 S2END[6]
rlabel metal2 7682 7854 7682 7854 0 S2END[7]
rlabel metal2 20838 8748 20838 8748 0 S2MID[0]
rlabel metal2 21114 10057 21114 10057 0 S2MID[1]
rlabel metal1 9798 6732 9798 6732 0 S2MID[2]
rlabel metal2 9706 6188 9706 6188 0 S2MID[3]
rlabel metal2 7222 6256 7222 6256 0 S2MID[4]
rlabel metal1 6831 6766 6831 6766 0 S2MID[5]
rlabel metal2 6486 6324 6486 6324 0 S2MID[6]
rlabel metal2 11730 7276 11730 7276 0 S2MID[7]
rlabel metal2 25254 9564 25254 9564 0 S4END[0]
rlabel metal1 11776 6290 11776 6290 0 S4END[10]
rlabel metal1 10074 5134 10074 5134 0 S4END[11]
rlabel metal1 10695 4590 10695 4590 0 S4END[12]
rlabel via2 10534 6307 10534 6307 0 S4END[13]
rlabel metal2 29118 9513 29118 9513 0 S4END[14]
rlabel metal2 29394 8952 29394 8952 0 S4END[15]
rlabel metal2 20286 7650 20286 7650 0 S4END[1]
rlabel metal2 16514 8381 16514 8381 0 S4END[2]
rlabel metal3 20516 8296 20516 8296 0 S4END[3]
rlabel metal1 16100 7378 16100 7378 0 S4END[4]
rlabel metal2 15778 9265 15778 9265 0 S4END[5]
rlabel metal1 15318 7888 15318 7888 0 S4END[6]
rlabel metal2 15226 7174 15226 7174 0 S4END[7]
rlabel metal2 17710 9469 17710 9469 0 S4END[8]
rlabel metal1 12834 7344 12834 7344 0 S4END[9]
rlabel metal2 14858 9520 14858 9520 0 SS4END[0]
rlabel metal2 32430 10261 32430 10261 0 SS4END[10]
rlabel metal2 32706 8986 32706 8986 0 SS4END[11]
rlabel metal2 32982 10125 32982 10125 0 SS4END[12]
rlabel metal2 33258 10261 33258 10261 0 SS4END[13]
rlabel metal2 33534 9462 33534 9462 0 SS4END[14]
rlabel metal2 33810 9088 33810 9088 0 SS4END[15]
rlabel metal2 19090 9418 19090 9418 0 SS4END[1]
rlabel metal2 30222 10176 30222 10176 0 SS4END[2]
rlabel metal2 30498 9734 30498 9734 0 SS4END[3]
rlabel metal2 30774 9632 30774 9632 0 SS4END[4]
rlabel metal2 31050 9598 31050 9598 0 SS4END[5]
rlabel metal2 31326 9564 31326 9564 0 SS4END[6]
rlabel metal2 31602 9530 31602 9530 0 SS4END[7]
rlabel metal2 31878 9326 31878 9326 0 SS4END[8]
rlabel metal2 32154 9734 32154 9734 0 SS4END[9]
rlabel metal2 1334 106 1334 106 0 UserCLK
rlabel metal1 34132 8602 34132 8602 0 UserCLKo
rlabel metal1 42550 2380 42550 2380 0 net1
rlabel metal1 18400 4046 18400 4046 0 net10
rlabel metal1 32384 7174 32384 7174 0 net100
rlabel metal2 19734 7599 19734 7599 0 net101
rlabel metal2 17986 7276 17986 7276 0 net102
rlabel metal2 17618 8636 17618 8636 0 net103
rlabel metal1 18170 7888 18170 7888 0 net104
rlabel metal2 32430 6630 32430 6630 0 net105
rlabel metal2 20654 4862 20654 4862 0 net11
rlabel metal1 41906 2482 41906 2482 0 net12
rlabel metal1 18998 5576 18998 5576 0 net13
rlabel metal2 18538 4403 18538 4403 0 net14
rlabel metal1 36386 4692 36386 4692 0 net15
rlabel metal2 23046 4607 23046 4607 0 net16
rlabel metal2 40342 6732 40342 6732 0 net17
rlabel metal1 25300 7174 25300 7174 0 net18
rlabel metal1 33166 6664 33166 6664 0 net19
rlabel metal1 36662 6324 36662 6324 0 net2
rlabel metal2 24242 8738 24242 8738 0 net20
rlabel metal2 36570 7344 36570 7344 0 net21
rlabel metal2 21942 7446 21942 7446 0 net22
rlabel metal1 21758 2856 21758 2856 0 net23
rlabel metal2 36478 7582 36478 7582 0 net24
rlabel metal2 41630 8670 41630 8670 0 net25
rlabel metal1 42734 2516 42734 2516 0 net26
rlabel metal1 42642 2312 42642 2312 0 net27
rlabel metal2 35834 3111 35834 3111 0 net28
rlabel metal2 27646 2958 27646 2958 0 net29
rlabel metal2 22862 4352 22862 4352 0 net3
rlabel metal2 36570 3264 36570 3264 0 net30
rlabel metal1 34638 3468 34638 3468 0 net31
rlabel metal1 21850 2924 21850 2924 0 net32
rlabel metal2 34730 8704 34730 8704 0 net33
rlabel metal2 32614 6613 32614 6613 0 net34
rlabel via2 20194 2907 20194 2907 0 net35
rlabel metal2 32798 7140 32798 7140 0 net36
rlabel metal2 38778 6443 38778 6443 0 net37
rlabel metal2 34822 6834 34822 6834 0 net38
rlabel metal2 33718 6120 33718 6120 0 net39
rlabel metal1 22034 4012 22034 4012 0 net4
rlabel metal1 37122 3978 37122 3978 0 net40
rlabel metal2 36662 6664 36662 6664 0 net41
rlabel metal1 39376 4794 39376 4794 0 net42
rlabel metal2 40710 5916 40710 5916 0 net43
rlabel metal2 13386 7191 13386 7191 0 net44
rlabel metal2 33626 7106 33626 7106 0 net45
rlabel metal1 9936 7990 9936 7990 0 net46
rlabel metal2 36202 8874 36202 8874 0 net47
rlabel metal1 35374 3706 35374 3706 0 net48
rlabel metal1 39008 5814 39008 5814 0 net49
rlabel metal1 17618 3400 17618 3400 0 net5
rlabel metal1 39606 6630 39606 6630 0 net50
rlabel metal1 38088 7514 38088 7514 0 net51
rlabel metal1 37214 6426 37214 6426 0 net52
rlabel metal1 4922 7514 4922 7514 0 net53
rlabel metal2 4370 7684 4370 7684 0 net54
rlabel metal1 4830 8398 4830 8398 0 net55
rlabel metal1 5658 5882 5658 5882 0 net56
rlabel metal2 5934 7990 5934 7990 0 net57
rlabel metal1 6578 6970 6578 6970 0 net58
rlabel metal1 6624 8466 6624 8466 0 net59
rlabel metal2 9890 3332 9890 3332 0 net6
rlabel metal2 7038 7548 7038 7548 0 net60
rlabel metal2 7866 7718 7866 7718 0 net61
rlabel metal1 9154 6970 9154 6970 0 net62
rlabel metal1 7774 8398 7774 8398 0 net63
rlabel metal2 8878 7378 8878 7378 0 net64
rlabel metal1 7820 6426 7820 6426 0 net65
rlabel metal1 8878 6426 8878 6426 0 net66
rlabel metal1 9568 6426 9568 6426 0 net67
rlabel metal1 9752 6154 9752 6154 0 net68
rlabel metal1 10534 5882 10534 5882 0 net69
rlabel metal1 32522 5712 32522 5712 0 net7
rlabel metal1 10442 7786 10442 7786 0 net70
rlabel metal1 10258 8500 10258 8500 0 net71
rlabel metal2 10534 8636 10534 8636 0 net72
rlabel metal2 10994 8942 10994 8942 0 net73
rlabel metal1 15364 8058 15364 8058 0 net74
rlabel metal1 15180 7514 15180 7514 0 net75
rlabel metal2 17434 8194 17434 8194 0 net76
rlabel metal1 14858 7820 14858 7820 0 net77
rlabel metal1 19964 8058 19964 8058 0 net78
rlabel metal2 22494 8500 22494 8500 0 net79
rlabel metal1 19527 3094 19527 3094 0 net8
rlabel metal1 11546 7820 11546 7820 0 net80
rlabel metal1 10902 8398 10902 8398 0 net81
rlabel metal1 9292 4794 9292 4794 0 net82
rlabel metal1 10304 5338 10304 5338 0 net83
rlabel metal1 12190 6426 12190 6426 0 net84
rlabel metal1 12558 7514 12558 7514 0 net85
rlabel metal1 13018 8058 13018 8058 0 net86
rlabel metal1 14996 7242 14996 7242 0 net87
rlabel metal1 13754 7888 13754 7888 0 net88
rlabel metal2 15410 8143 15410 8143 0 net89
rlabel metal2 40158 4930 40158 4930 0 net9
rlabel metal2 19366 6953 19366 6953 0 net90
rlabel metal1 18354 8500 18354 8500 0 net91
rlabel metal2 18722 8228 18722 8228 0 net92
rlabel metal2 21850 7956 21850 7956 0 net93
rlabel metal1 19044 8058 19044 8058 0 net94
rlabel metal2 13110 7582 13110 7582 0 net95
rlabel metal2 16330 7582 16330 7582 0 net96
rlabel metal1 34822 7174 34822 7174 0 net97
rlabel metal2 16146 7599 16146 7599 0 net98
rlabel metal2 16790 6970 16790 6970 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 11250
<< end >>
