* NGSPICE file created from S_term_DSP.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

.subckt S_term_DSP FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_5_343 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_4
XFILLER_3_89 VPWR VGND sg13g2_fill_2
XFILLER_2_324 VPWR VGND sg13g2_decap_8
X_062_ S2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_110 VPWR VGND sg13g2_decap_8
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_7_279 VPWR VGND sg13g2_decap_8
X_045_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
XFILLER_4_205 VPWR VGND sg13g2_decap_8
X_028_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput97 net97 NN4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput75 net75 N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput86 net86 N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput64 net64 N2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput53 net53 N1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_5_322 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_8_182 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_decap_8
XFILLER_2_303 VPWR VGND sg13g2_decap_8
XFILLER_5_141 VPWR VGND sg13g2_fill_2
XFILLER_9_67 VPWR VGND sg13g2_fill_2
XFILLER_9_56 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_188 VPWR VGND sg13g2_fill_2
X_061_ S2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_7_258 VPWR VGND sg13g2_decap_8
XFILLER_7_247 VPWR VGND sg13g2_decap_8
X_044_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
X_027_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XFILLER_6_35 VPWR VGND sg13g2_decap_8
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput98 net98 NN4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput76 net76 N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput87 net87 N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput65 net65 N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput54 net54 N1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_8_320 VPWR VGND sg13g2_fill_2
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_0_231 VPWR VGND sg13g2_decap_8
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_8_375 VPWR VGND sg13g2_fill_2
XFILLER_5_301 VPWR VGND sg13g2_decap_8
XFILLER_8_161 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_fill_2
XFILLER_2_359 VPWR VGND sg13g2_decap_8
XFILLER_5_120 VPWR VGND sg13g2_decap_8
XFILLER_5_197 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_2_145 VPWR VGND sg13g2_decap_4
X_060_ S2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_7_226 VPWR VGND sg13g2_decap_8
X_043_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
X_026_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_3_273 VPWR VGND sg13g2_decap_8
XFILLER_3_295 VPWR VGND sg13g2_decap_8
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput99 net99 NN4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput77 net77 N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput88 net88 N4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput66 net66 N2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput55 net55 N1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
X_009_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
XFILLER_8_140 VPWR VGND sg13g2_decap_8
XFILLER_5_357 VPWR VGND sg13g2_decap_8
XFILLER_2_338 VPWR VGND sg13g2_decap_8
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_5_143 VPWR VGND sg13g2_fill_1
XFILLER_5_176 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_2_124 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_fill_1
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_7_205 VPWR VGND sg13g2_fill_2
X_042_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_6_293 VPWR VGND sg13g2_fill_1
XFILLER_6_282 VPWR VGND sg13g2_decap_8
XFILLER_1_92 VPWR VGND sg13g2_decap_8
XFILLER_4_219 VPWR VGND sg13g2_decap_8
X_025_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XFILLER_3_252 VPWR VGND sg13g2_decap_8
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput89 net89 NN4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput78 net78 N4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput67 net67 N2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput56 net56 N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_8_333 VPWR VGND sg13g2_decap_8
X_008_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_5_336 VPWR VGND sg13g2_decap_8
XFILLER_3_27 VPWR VGND sg13g2_fill_1
XFILLER_2_317 VPWR VGND sg13g2_decap_8
XFILLER_1_361 VPWR VGND sg13g2_decap_8
XFILLER_1_372 VPWR VGND sg13g2_fill_1
XFILLER_2_103 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_9_280 VPWR VGND sg13g2_decap_4
X_041_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_6_261 VPWR VGND sg13g2_decap_8
X_024_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XFILLER_6_49 VPWR VGND sg13g2_decap_8
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput57 net57 N2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput79 net79 N4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput68 net68 N2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_0_245 VPWR VGND sg13g2_decap_8
X_007_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_5_315 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_8_175 VPWR VGND sg13g2_decap_8
XFILLER_4_370 VPWR VGND sg13g2_decap_8
XFILLER_1_340 VPWR VGND sg13g2_decap_8
XFILLER_5_134 VPWR VGND sg13g2_decap_8
XFILLER_9_49 VPWR VGND sg13g2_decap_8
XFILLER_7_207 VPWR VGND sg13g2_fill_1
X_040_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_6_240 VPWR VGND sg13g2_decap_8
X_023_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_3_232 VPWR VGND sg13g2_decap_8
XFILLER_3_287 VPWR VGND sg13g2_decap_4
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput69 net69 N2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput58 net58 N2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_8_368 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
X_006_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
XFILLER_8_154 VPWR VGND sg13g2_decap_8
XFILLER_5_113 VPWR VGND sg13g2_decap_8
XFILLER_4_94 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_2_138 VPWR VGND sg13g2_decap_8
XFILLER_2_149 VPWR VGND sg13g2_fill_1
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_1_193 VPWR VGND sg13g2_decap_8
XFILLER_7_219 VPWR VGND sg13g2_decap_8
X_099_ SS4END[4] net91 VPWR VGND sg13g2_buf_1
XFILLER_10_60 VPWR VGND sg13g2_fill_1
X_022_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
XFILLER_3_211 VPWR VGND sg13g2_decap_8
XFILLER_3_266 VPWR VGND sg13g2_decap_8
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput59 net59 N2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_8_347 VPWR VGND sg13g2_decap_8
X_005_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
XFILLER_8_133 VPWR VGND sg13g2_decap_8
XFILLER_4_191 VPWR VGND sg13g2_decap_8
XFILLER_2_117 VPWR VGND sg13g2_decap_8
XFILLER_1_172 VPWR VGND sg13g2_decap_8
X_098_ SS4END[5] net90 VPWR VGND sg13g2_buf_1
XFILLER_6_275 VPWR VGND sg13g2_decap_8
XFILLER_1_85 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_3_245 VPWR VGND sg13g2_decap_8
X_021_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_326 VPWR VGND sg13g2_decap_8
X_004_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_8_189 VPWR VGND sg13g2_fill_2
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_5_329 VPWR VGND sg13g2_decap_8
XFILLER_1_354 VPWR VGND sg13g2_decap_8
XFILLER_4_52 VPWR VGND sg13g2_decap_8
XFILLER_4_170 VPWR VGND sg13g2_decap_8
XFILLER_9_284 VPWR VGND sg13g2_fill_1
XFILLER_9_273 VPWR VGND sg13g2_decap_8
XFILLER_10_261 VPWR VGND sg13g2_decap_8
X_097_ SS4END[6] net104 VPWR VGND sg13g2_buf_1
XFILLER_6_254 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_020_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_8_316 VPWR VGND sg13g2_decap_4
X_003_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_7_371 VPWR VGND sg13g2_decap_4
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_5_308 VPWR VGND sg13g2_decap_8
XFILLER_8_168 VPWR VGND sg13g2_decap_8
XFILLER_4_363 VPWR VGND sg13g2_decap_8
XFILLER_5_127 VPWR VGND sg13g2_decap_8
XFILLER_1_333 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_4
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_1_163 VPWR VGND sg13g2_decap_4
XFILLER_1_130 VPWR VGND sg13g2_decap_8
XFILLER_9_252 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_10_240 VPWR VGND sg13g2_decap_8
X_096_ SS4END[7] net103 VPWR VGND sg13g2_buf_1
XFILLER_6_233 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_3_225 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
X_079_ S4END[8] net86 VPWR VGND sg13g2_buf_1
X_002_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_7_350 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_decap_8
XFILLER_4_342 VPWR VGND sg13g2_decap_8
XFILLER_1_312 VPWR VGND sg13g2_decap_8
XFILLER_5_106 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_4_87 VPWR VGND sg13g2_decap_8
XFILLER_4_150 VPWR VGND sg13g2_decap_8
XFILLER_4_161 VPWR VGND sg13g2_fill_1
XFILLER_9_231 VPWR VGND sg13g2_decap_8
XFILLER_1_186 VPWR VGND sg13g2_decap_8
X_095_ SS4END[8] net102 VPWR VGND sg13g2_buf_1
XFILLER_6_289 VPWR VGND sg13g2_decap_4
XFILLER_6_212 VPWR VGND sg13g2_decap_8
XFILLER_1_99 VPWR VGND sg13g2_decap_8
XFILLER_10_42 VPWR VGND sg13g2_decap_8
XFILLER_3_204 VPWR VGND sg13g2_decap_8
XFILLER_3_259 VPWR VGND sg13g2_decap_8
X_078_ S4END[9] net85 VPWR VGND sg13g2_buf_1
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
X_001_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_4_321 VPWR VGND sg13g2_decap_8
XFILLER_1_368 VPWR VGND sg13g2_decap_4
XFILLER_4_184 VPWR VGND sg13g2_decap_8
XFILLER_9_210 VPWR VGND sg13g2_decap_8
X_094_ SS4END[9] net101 VPWR VGND sg13g2_buf_1
XFILLER_6_268 VPWR VGND sg13g2_decap_8
XFILLER_1_78 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_10_21 VPWR VGND sg13g2_decap_8
X_077_ S4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_7_77 VPWR VGND sg13g2_decap_8
X_000_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_4_300 VPWR VGND sg13g2_decap_8
XFILLER_1_347 VPWR VGND sg13g2_decap_8
XFILLER_9_266 VPWR VGND sg13g2_decap_8
XFILLER_1_111 VPWR VGND sg13g2_decap_8
XFILLER_10_254 VPWR VGND sg13g2_decap_8
X_093_ SS4END[10] net100 VPWR VGND sg13g2_buf_1
XFILLER_6_247 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_3_239 VPWR VGND sg13g2_fill_2
XFILLER_2_272 VPWR VGND sg13g2_decap_8
XFILLER_2_283 VPWR VGND sg13g2_fill_2
X_076_ S4END[11] net83 VPWR VGND sg13g2_buf_1
XFILLER_7_375 VPWR VGND sg13g2_fill_2
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
X_059_ S2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_4_356 VPWR VGND sg13g2_decap_8
XFILLER_1_304 VPWR VGND sg13g2_decap_4
XFILLER_1_326 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_fill_2
XFILLER_1_167 VPWR VGND sg13g2_fill_1
XFILLER_1_156 VPWR VGND sg13g2_decap_8
XFILLER_1_145 VPWR VGND sg13g2_fill_2
XFILLER_9_245 VPWR VGND sg13g2_decap_8
XFILLER_10_233 VPWR VGND sg13g2_decap_8
XFILLER_6_226 VPWR VGND sg13g2_decap_8
X_092_ SS4END[11] net99 VPWR VGND sg13g2_buf_1
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_10_56 VPWR VGND sg13g2_decap_4
XFILLER_5_281 VPWR VGND sg13g2_decap_8
XFILLER_3_218 VPWR VGND sg13g2_decap_8
X_075_ S4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_7_343 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_058_ S2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_4_335 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_143 VPWR VGND sg13g2_decap_8
XFILLER_4_198 VPWR VGND sg13g2_decap_8
XFILLER_1_179 VPWR VGND sg13g2_decap_8
XFILLER_9_224 VPWR VGND sg13g2_decap_8
XFILLER_10_212 VPWR VGND sg13g2_decap_8
X_091_ SS4END[12] net98 VPWR VGND sg13g2_buf_1
XFILLER_6_205 VPWR VGND sg13g2_decap_8
XFILLER_5_260 VPWR VGND sg13g2_decap_8
XFILLER_10_35 VPWR VGND sg13g2_decap_8
X_074_ S4END[13] net81 VPWR VGND sg13g2_buf_1
XFILLER_2_252 VPWR VGND sg13g2_decap_8
XFILLER_2_296 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_057_ S2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_4_314 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_4_177 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_fill_1
XFILLER_1_125 VPWR VGND sg13g2_fill_1
XFILLER_9_203 VPWR VGND sg13g2_decap_8
XFILLER_10_268 VPWR VGND sg13g2_decap_8
X_090_ SS4END[13] net97 VPWR VGND sg13g2_buf_1
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_5_294 VPWR VGND sg13g2_decap_8
XFILLER_10_14 VPWR VGND sg13g2_decap_8
XFILLER_2_231 VPWR VGND sg13g2_decap_8
X_073_ S4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_4_0 VPWR VGND sg13g2_decap_8
X_056_ S2MID[7] net57 VPWR VGND sg13g2_buf_1
XFILLER_7_175 VPWR VGND sg13g2_decap_4
X_039_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_8_91 VPWR VGND sg13g2_decap_8
XFILLER_4_101 VPWR VGND sg13g2_decap_8
XFILLER_4_134 VPWR VGND sg13g2_decap_4
XFILLER_9_259 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_5_92 VPWR VGND sg13g2_decap_8
XFILLER_10_247 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_2_265 VPWR VGND sg13g2_decap_8
X_072_ S4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_2_82 VPWR VGND sg13g2_decap_8
XFILLER_7_357 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
X_055_ S1END[0] net56 VPWR VGND sg13g2_buf_1
XFILLER_4_349 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
X_038_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_1_319 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_157 VPWR VGND sg13g2_decap_4
XFILLER_3_190 VPWR VGND sg13g2_decap_8
XFILLER_9_238 VPWR VGND sg13g2_decap_8
XFILLER_8_293 VPWR VGND sg13g2_fill_2
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_10_226 VPWR VGND sg13g2_decap_8
XFILLER_6_219 VPWR VGND sg13g2_decap_8
XFILLER_5_71 VPWR VGND sg13g2_decap_8
XFILLER_5_274 VPWR VGND sg13g2_decap_8
XFILLER_10_49 VPWR VGND sg13g2_decap_8
X_071_ S2END[0] net72 VPWR VGND sg13g2_buf_1
XFILLER_2_61 VPWR VGND sg13g2_decap_8
XFILLER_7_336 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_054_ S1END[1] net55 VPWR VGND sg13g2_buf_1
XFILLER_4_328 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
X_037_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_3_372 VPWR VGND sg13g2_decap_4
XFILLER_0_364 VPWR VGND sg13g2_fill_1
XFILLER_1_106 VPWR VGND sg13g2_fill_1
XFILLER_9_217 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_10_205 VPWR VGND sg13g2_decap_8
XFILLER_8_250 VPWR VGND sg13g2_fill_1
XFILLER_5_253 VPWR VGND sg13g2_decap_8
XFILLER_10_28 VPWR VGND sg13g2_decap_8
XFILLER_2_245 VPWR VGND sg13g2_decap_8
XFILLER_2_289 VPWR VGND sg13g2_decap_8
X_070_ S2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_7_304 VPWR VGND sg13g2_decap_8
XFILLER_2_0 VPWR VGND sg13g2_decap_8
X_053_ S1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_6_370 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_4_307 VPWR VGND sg13g2_decap_8
X_036_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_3_351 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
X_019_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_1_118 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_8_295 VPWR VGND sg13g2_fill_1
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_5_232 VPWR VGND sg13g2_decap_8
XFILLER_2_224 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_decap_4
XFILLER_2_96 VPWR VGND sg13g2_decap_8
X_052_ S1END[3] net53 VPWR VGND sg13g2_buf_1
XFILLER_7_179 VPWR VGND sg13g2_fill_2
XFILLER_7_168 VPWR VGND sg13g2_decap_8
X_035_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
X_104_ UserCLK net105 VPWR VGND sg13g2_buf_1
XFILLER_3_330 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
X_018_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_4_138 VPWR VGND sg13g2_fill_1
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
XFILLER_8_241 VPWR VGND sg13g2_decap_8
XFILLER_5_85 VPWR VGND sg13g2_decap_8
XFILLER_5_288 VPWR VGND sg13g2_fill_2
XFILLER_5_211 VPWR VGND sg13g2_decap_8
XFILLER_2_42 VPWR VGND sg13g2_fill_1
XFILLER_2_75 VPWR VGND sg13g2_decap_8
X_051_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
X_103_ SS4END[0] net95 VPWR VGND sg13g2_buf_1
XFILLER_7_147 VPWR VGND sg13g2_decap_8
X_034_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_6_180 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
X_017_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_3_183 VPWR VGND sg13g2_decap_8
XFILLER_8_286 VPWR VGND sg13g2_decap_8
XFILLER_8_220 VPWR VGND sg13g2_decap_4
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_5_42 VPWR VGND sg13g2_fill_2
XFILLER_5_64 VPWR VGND sg13g2_decap_8
XFILLER_10_219 VPWR VGND sg13g2_decap_8
XFILLER_5_267 VPWR VGND sg13g2_decap_8
XFILLER_2_259 VPWR VGND sg13g2_fill_2
XFILLER_1_281 VPWR VGND sg13g2_decap_8
XFILLER_1_292 VPWR VGND sg13g2_fill_1
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_54 VPWR VGND sg13g2_decap_8
Xoutput100 net100 NN4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_7_329 VPWR VGND sg13g2_decap_8
X_050_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
X_102_ SS4END[1] net94 VPWR VGND sg13g2_buf_1
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
X_033_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_3_365 VPWR VGND sg13g2_decap_8
XFILLER_3_376 VPWR VGND sg13g2_fill_1
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
X_016_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_3_162 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_5_246 VPWR VGND sg13g2_decap_8
XFILLER_2_216 VPWR VGND sg13g2_decap_4
XFILLER_2_238 VPWR VGND sg13g2_decap_8
XFILLER_4_7 VPWR VGND sg13g2_decap_8
Xoutput101 net101 NN4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_6_363 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_decap_8
X_101_ SS4END[2] net93 VPWR VGND sg13g2_buf_1
X_032_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_3_344 VPWR VGND sg13g2_decap_8
XFILLER_8_98 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_4_108 VPWR VGND sg13g2_fill_2
X_015_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_141 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_8_255 VPWR VGND sg13g2_decap_4
XFILLER_5_99 VPWR VGND sg13g2_decap_8
XFILLER_5_225 VPWR VGND sg13g2_decap_8
XFILLER_2_89 VPWR VGND sg13g2_decap_8
Xoutput102 net102 NN4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_6_342 VPWR VGND sg13g2_decap_8
X_031_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
X_100_ SS4END[3] net92 VPWR VGND sg13g2_buf_1
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_6_161 VPWR VGND sg13g2_fill_1
XFILLER_3_323 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
X_014_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_3_120 VPWR VGND sg13g2_decap_8
XFILLER_3_197 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_5_78 VPWR VGND sg13g2_decap_8
XFILLER_5_204 VPWR VGND sg13g2_decap_8
XFILLER_2_207 VPWR VGND sg13g2_fill_1
XFILLER_9_351 VPWR VGND sg13g2_decap_8
Xoutput103 net103 NN4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_2_68 VPWR VGND sg13g2_decap_8
XFILLER_6_321 VPWR VGND sg13g2_decap_8
X_030_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_3_302 VPWR VGND sg13g2_decap_8
XFILLER_10_191 VPWR VGND sg13g2_decap_8
XFILLER_6_173 VPWR VGND sg13g2_decap_8
XFILLER_6_140 VPWR VGND sg13g2_decap_8
X_013_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_3_176 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_8_279 VPWR VGND sg13g2_decap_8
XFILLER_8_268 VPWR VGND sg13g2_decap_8
XFILLER_8_224 VPWR VGND sg13g2_fill_1
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_4_293 VPWR VGND sg13g2_decap_8
XFILLER_9_330 VPWR VGND sg13g2_decap_8
Xoutput104 net104 NN4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_1_230 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_2_47 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_9_182 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_3_358 VPWR VGND sg13g2_decap_8
X_089_ SS4END[14] net96 VPWR VGND sg13g2_buf_1
XFILLER_8_35 VPWR VGND sg13g2_decap_8
X_012_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_3_155 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_8_236 VPWR VGND sg13g2_fill_1
XFILLER_8_214 VPWR VGND sg13g2_fill_2
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_5_239 VPWR VGND sg13g2_decap_8
XFILLER_4_283 VPWR VGND sg13g2_decap_4
XFILLER_1_297 VPWR VGND sg13g2_decap_8
Xoutput105 net105 UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_10_341 VPWR VGND sg13g2_decap_8
XFILLER_6_356 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_decap_8
XFILLER_3_91 VPWR VGND sg13g2_fill_1
XFILLER_3_337 VPWR VGND sg13g2_decap_8
X_088_ SS4END[15] net89 VPWR VGND sg13g2_buf_1
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
X_011_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_3_134 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_8_259 VPWR VGND sg13g2_fill_1
XFILLER_8_248 VPWR VGND sg13g2_fill_2
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
XFILLER_5_218 VPWR VGND sg13g2_decap_8
XFILLER_4_262 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_1_265 VPWR VGND sg13g2_decap_4
XFILLER_9_365 VPWR VGND sg13g2_decap_4
XFILLER_6_335 VPWR VGND sg13g2_decap_8
XFILLER_6_302 VPWR VGND sg13g2_decap_8
XFILLER_3_316 VPWR VGND sg13g2_decap_8
XFILLER_6_198 VPWR VGND sg13g2_decap_8
XFILLER_6_187 VPWR VGND sg13g2_decap_8
X_087_ S4END[0] net79 VPWR VGND sg13g2_buf_1
XFILLER_6_154 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_010_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_3_113 VPWR VGND sg13g2_decap_8
XFILLER_2_190 VPWR VGND sg13g2_fill_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_7_293 VPWR VGND sg13g2_fill_2
XFILLER_4_241 VPWR VGND sg13g2_decap_8
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_1_244 VPWR VGND sg13g2_decap_4
XFILLER_1_200 VPWR VGND sg13g2_decap_8
XFILLER_1_288 VPWR VGND sg13g2_decap_4
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_9_344 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_9_196 VPWR VGND sg13g2_decap_8
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_3_71 VPWR VGND sg13g2_fill_2
XFILLER_10_184 VPWR VGND sg13g2_decap_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_6_166 VPWR VGND sg13g2_decap_8
XFILLER_6_133 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
X_086_ S4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_3_103 VPWR VGND sg13g2_decap_4
XFILLER_3_169 VPWR VGND sg13g2_decap_8
X_069_ S2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_7_272 VPWR VGND sg13g2_decap_8
XFILLER_1_223 VPWR VGND sg13g2_decap_8
Xoutput90 net90 NN4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_10_355 VPWR VGND sg13g2_decap_4
XFILLER_9_175 VPWR VGND sg13g2_decap_8
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_2_373 VPWR VGND sg13g2_decap_4
X_085_ S4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_3_148 VPWR VGND sg13g2_decap_8
X_068_ S2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_8_229 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_7_295 VPWR VGND sg13g2_fill_1
XFILLER_7_240 VPWR VGND sg13g2_decap_8
XFILLER_4_276 VPWR VGND sg13g2_decap_8
XFILLER_4_287 VPWR VGND sg13g2_fill_2
XFILLER_9_324 VPWR VGND sg13g2_fill_2
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput91 net91 NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput80 net80 N4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_10_334 VPWR VGND sg13g2_decap_8
XFILLER_6_349 VPWR VGND sg13g2_decap_8
XFILLER_6_316 VPWR VGND sg13g2_fill_1
XFILLER_5_371 VPWR VGND sg13g2_decap_4
XFILLER_3_84 VPWR VGND sg13g2_fill_1
XFILLER_2_352 VPWR VGND sg13g2_decap_8
X_084_ S4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_5_190 VPWR VGND sg13g2_decap_8
XFILLER_3_127 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
X_067_ S2END[4] net68 VPWR VGND sg13g2_buf_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_4_233 VPWR VGND sg13g2_decap_4
XFILLER_4_255 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_9_358 VPWR VGND sg13g2_decap_8
XFILLER_1_258 VPWR VGND sg13g2_decap_8
Xoutput92 net92 NN4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput81 net81 N4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput70 net70 N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_6_328 VPWR VGND sg13g2_decap_8
XFILLER_5_350 VPWR VGND sg13g2_decap_8
XFILLER_3_96 VPWR VGND sg13g2_fill_2
XFILLER_3_309 VPWR VGND sg13g2_decap_8
XFILLER_10_198 VPWR VGND sg13g2_decap_8
XFILLER_6_147 VPWR VGND sg13g2_decap_8
XFILLER_2_331 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
X_083_ S4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_2_161 VPWR VGND sg13g2_decap_8
X_066_ S2END[5] net67 VPWR VGND sg13g2_buf_1
X_049_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
XFILLER_7_286 VPWR VGND sg13g2_decap_8
XFILLER_4_212 VPWR VGND sg13g2_decap_8
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_1_248 VPWR VGND sg13g2_fill_2
XFILLER_1_237 VPWR VGND sg13g2_decap_8
XFILLER_9_337 VPWR VGND sg13g2_decap_8
Xoutput93 net93 NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput82 net82 N4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 N2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput60 net60 N2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_9_189 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_10_177 VPWR VGND sg13g2_decap_8
XFILLER_6_126 VPWR VGND sg13g2_decap_8
XFILLER_2_310 VPWR VGND sg13g2_decap_8
X_082_ S4END[5] net74 VPWR VGND sg13g2_buf_1
XFILLER_3_107 VPWR VGND sg13g2_fill_2
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
X_065_ S2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_9_63 VPWR VGND sg13g2_decap_4
XFILLER_7_265 VPWR VGND sg13g2_decap_8
X_048_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XFILLER_1_216 VPWR VGND sg13g2_decap_8
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput94 net94 NN4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput83 net83 N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 N2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput61 net61 N2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_10_359 VPWR VGND sg13g2_fill_2
XFILLER_10_348 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_fill_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
X_081_ S4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_2_366 VPWR VGND sg13g2_decap_8
X_064_ S2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_7_233 VPWR VGND sg13g2_decap_8
X_047_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_6_98 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_4_269 VPWR VGND sg13g2_decap_8
XFILLER_3_280 VPWR VGND sg13g2_decap_8
XFILLER_9_317 VPWR VGND sg13g2_decap_8
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput95 net95 NN4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput84 net84 N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 N4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput62 net62 N2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_0_294 VPWR VGND sg13g2_decap_8
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_8_361 VPWR VGND sg13g2_decap_8
XFILLER_10_327 VPWR VGND sg13g2_decap_8
XFILLER_6_309 VPWR VGND sg13g2_decap_8
XFILLER_5_375 VPWR VGND sg13g2_fill_2
XFILLER_5_364 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_8_191 VPWR VGND sg13g2_fill_1
X_080_ S4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_2_345 VPWR VGND sg13g2_decap_8
XFILLER_5_183 VPWR VGND sg13g2_decap_8
XFILLER_2_131 VPWR VGND sg13g2_decap_8
XFILLER_2_175 VPWR VGND sg13g2_decap_4
XFILLER_3_0 VPWR VGND sg13g2_decap_8
X_063_ S2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_7_212 VPWR VGND sg13g2_decap_8
X_046_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_4_226 VPWR VGND sg13g2_decap_8
XFILLER_4_248 VPWR VGND sg13g2_decap_8
X_029_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
XFILLER_6_77 VPWR VGND sg13g2_decap_8
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_1_207 VPWR VGND sg13g2_fill_1
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput96 net96 NN4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput74 net74 N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput85 net85 N4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput63 net63 N2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_8_340 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
.ends

