* NGSPICE file created from DSP.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VGND VPWR
Xclkbuf_2_2__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3155_ net1002 net666 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__mux2_1
X_3086_ net1033 net983 net1042 net1053 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _1863_ sky130_fd_sc_hd__mux4_1
X_2106_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q _0978_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__a21oi_2
X_2037_ net1020 net1036 net1032 net983 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ _0913_ sky130_fd_sc_hd__mux4_1
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3988_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q _0652_ _0651_
+ _0073_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__a211o_1
X_2939_ net186 net201 net114 net1048 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_148_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4609_ net1228 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_202 net1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_213 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_224 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_268 net349 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_246 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_257 net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_235 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_279 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4960_ net1203 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_19_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4891_ net1197 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3911_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q _0579_ _0133_
+ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__a21o_1
X_3842_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q _0515_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__o21ai_1
X_5512_ Tile_X0Y1_WW4END[7] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_4
X_3773_ net663 _0448_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a21oi_4
X_2724_ _1396_ _1528_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__xor2_1
X_5443_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net535
+ sky130_fd_sc_hd__buf_8
Xoutput401 net401 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[0] sky130_fd_sc_hd__buf_2
X_2655_ _1121_ _1125_ _1502_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__a21o_1
Xoutput412 net412 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput423 net423 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput434 net434 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[7] sky130_fd_sc_hd__buf_2
X_5374_ Tile_X0Y1_E6END[11] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
XFILLER_99_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4325_ net1232 net1147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput445 net445 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput456 net456 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput478 net478 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput467 net467 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[8] sky130_fd_sc_hd__buf_2
X_2586_ net192 net137 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q
+ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__mux4_2
Xoutput489 net489 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[13] sky130_fd_sc_hd__buf_2
X_4256_ _0615_ _0616_ _0821_ _0820_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a31oi_4
X_4187_ net176 net182 net194 net127 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0838_ sky130_fd_sc_hd__mux4_1
X_3207_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _1950_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3138_ net139 net72 net83 net971 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_82_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3069_ _1845_ _1847_ _1848_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_53_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2440_ net989 net1023 net864 net1008 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q VGND VGND VPWR VPWR
+ _1302_ sky130_fd_sc_hd__mux4_1
X_2371_ net193 net25 net68 net104 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q VGND VGND VPWR VPWR
+ _1238_ sky130_fd_sc_hd__mux4_1
X_4110_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q _0764_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ _0763_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__o211a_1
X_5090_ net1207 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4041_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q _0697_ _0698_
+ _0699_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q VGND VGND VPWR
+ VPWR _0702_ sky130_fd_sc_hd__a221o_1
XFILLER_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4943_ net1187 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4874_ net1216 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3825_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0499_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3756_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q _0436_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a21o_1
X_2707_ _1173_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__xor2_1
XFILLER_118_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5426_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net518
+ sky130_fd_sc_hd__buf_4
X_3687_ net1017 net823 net982 net867 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0374_ sky130_fd_sc_hd__mux4_2
Xoutput253 net253 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[2] sky130_fd_sc_hd__buf_4
X_2638_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q _1486_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__o21a_1
Xoutput286 net286 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[11] sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_99_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5357_ net131 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_2
X_2569_ net189 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net225
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__mux4_2
Xoutput297 net297 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[21] sky130_fd_sc_hd__buf_2
X_4308_ net40 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5288_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_6
X_4239_ _0805_ _0807_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__xor2_2
XFILLER_70_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_122_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone248 net986 VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_88_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4590_ net1239 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3610_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q _0299_ VGND VGND
+ VPWR VPWR _0300_ sky130_fd_sc_hd__nand2b_2
X_3541_ net176 net182 net127 net1222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0234_ sky130_fd_sc_hd__mux4_1
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3472_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\] VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_1
X_5211_ net37 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2423_ net990 net1023 net1004 net1011 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1286_ sky130_fd_sc_hd__mux4_2
XFILLER_130_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2354_ _0110_ _1219_ _1220_ _1221_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a221o_1
X_5142_ net156 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2285_ _0896_ _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nand2_2
XFILLER_96_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5073_ net170 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4024_ _0105_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and2_4
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4926_ net1200 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4857_ net1194 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3808_ net1221 net215 net90 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q VGND VGND VPWR VPWR
+ _0484_ sky130_fd_sc_hd__mux4_1
XFILLER_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4788_ net1192 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3739_ net94 net1225 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XFILLER_4_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5409_ net152 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_1
XFILLER_79_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1231 net52 VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__buf_4
Xfanout1220 net145 VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__buf_4
Xfanout1264 net3 VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__buf_4
Xfanout1242 Tile_X0Y0_FrameData[25] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1253 net34 VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__buf_4
XFILLER_78_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2070_ _0855_ _0883_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_77_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2972_ _1767_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__inv_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4711_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C3 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ net1229 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4573_ net1257 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3524_ net925 net970 net999 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0218_ sky130_fd_sc_hd__mux4_2
X_3455_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR
+ VPWR _0150_ sky130_fd_sc_hd__inv_1
X_2406_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1267_ _1269_
+ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__and3_1
X_3386_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q VGND VGND VPWR
+ VPWR _0081_ sky130_fd_sc_hd__inv_2
X_2337_ net208 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q VGND
+ VGND VPWR VPWR _1206_ sky130_fd_sc_hd__mux2_1
X_5125_ net1211 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2268_ _0945_ _0949_ _0950_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__and3_1
X_5056_ net1203 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4007_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q _0669_ VGND VGND
+ VPWR VPWR _0670_ sky130_fd_sc_hd__nand2b_1
XFILLER_84_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2199_ _0984_ _1049_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__xnor2_2
XFILLER_25_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4909_ net1219 net1108 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3240_ _1974_ _1978_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 sky130_fd_sc_hd__mux2_2
XFILLER_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3171_ net1007 _1400_ _1473_ _0841_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q VGND VGND VPWR VPWR
+ _1920_ sky130_fd_sc_hd__mux4_2
X_2122_ _0991_ _0992_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__xnor2_1
Xfanout1061 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q VGND VGND
+ VPWR VPWR net1061 sky130_fd_sc_hd__clkbuf_8
Xfanout1072 net213 VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__buf_4
Xfanout1083 net1085 VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__clkbuf_2
Xfanout1050 net1052 VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__buf_6
Xfanout1094 net1095 VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__buf_2
Xrebuffer17 net633 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2053_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\] net1059 VGND VGND VPWR VPWR _0927_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_22_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q _0560_ _1760_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q VGND VGND VPWR VPWR
+ _1761_ sky130_fd_sc_hd__a211o_1
X_2886_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _1708_ VGND VGND
+ VPWR VPWR _1709_ sky130_fd_sc_hd__or2_1
X_4625_ net1244 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4556_ net1237 net1079 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3507_ net1053 net1048 net1029 net822 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0202_ sky130_fd_sc_hd__mux4_1
X_4487_ net1236 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3438_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR
+ VPWR _0133_ sky130_fd_sc_hd__inv_2
XFILLER_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3369_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR
+ VPWR _0064_ sky130_fd_sc_hd__inv_1
X_5108_ net167 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5039_ net1187 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput120 Tile_X0Y1_E1END[1] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_4
Xinput131 Tile_X0Y1_E2MID[0] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
Xinput142 Tile_X0Y1_EE4END[1] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput153 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_2
Xinput186 Tile_X0Y1_N2MID[0] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_6
Xinput175 Tile_X0Y1_N1END[1] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_4
Xinput164 Tile_X0Y1_FrameData[2] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_2
Xinput197 Tile_X0Y1_N4END[3] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_2
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ net815 net1036 net1032 net985 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1573_ sky130_fd_sc_hd__mux4_1
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2671_ _1517_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] net1067 VGND VGND VPWR VPWR
+ _1518_ sky130_fd_sc_hd__mux2_4
X_4410_ net1254 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_152_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput616 net616 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[9] sky130_fd_sc_hd__buf_2
X_5390_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR net473
+ sky130_fd_sc_hd__clkbuf_2
Xoutput605 net605 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[13] sky130_fd_sc_hd__buf_4
X_4341_ net1248 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4272_ net1242 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3223_ _1961_ _1964_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 sky130_fd_sc_hd__mux2_1
X_3154_ _1906_ _1908_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__nand2_1
X_3085_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _1861_ VGND VGND
+ VPWR VPWR _1862_ sky130_fd_sc_hd__or2_1
X_2105_ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__inv_2
X_2036_ _0908_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q _0911_
+ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a21o_1
X_3987_ net100 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__mux2_1
X_2938_ net189 net200 net1262 net1053 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2869_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _1690_ _1692_
+ _0177_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__o211a_1
X_4608_ net1227 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4539_ net32 net1089 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 net1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_214 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_236 net186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_258 net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_247 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 net403 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4890_ net1196 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3910_ net74 net211 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__mux2_1
XFILLER_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3841_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_17_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3772_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0449_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o211a_4
XFILLER_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5511_ Tile_X0Y1_WW4END[6] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_4
X_2723_ _1562_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 sky130_fd_sc_hd__mux2_4
X_5442_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR net534
+ sky130_fd_sc_hd__buf_4
Xoutput402 net402 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[1] sky130_fd_sc_hd__buf_2
X_2654_ _0928_ _0981_ net832 _0848_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__o22a_1
Xoutput413 net413 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[2] sky130_fd_sc_hd__buf_2
Xoutput424 net424 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput435 net435 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[8] sky130_fd_sc_hd__buf_2
X_5373_ Tile_X0Y1_E6END[10] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_1
X_2585_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _1436_ VGND VGND
+ VPWR VPWR _1437_ sky130_fd_sc_hd__or2_1
XFILLER_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4324_ net1231 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput446 net446 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput457 net457 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput468 net468 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput479 net479 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[4] sky130_fd_sc_hd__buf_2
X_4255_ _0898_ _0899_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4186_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q _0834_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a21bo_1
X_3206_ _1949_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__inv_1
XFILLER_94_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3137_ net1221 net82 net71 net921 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3068_ net920 net1225 net60 net983 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q VGND VGND VPWR VPWR
+ _1848_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_148_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer290 net874 VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2370_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q _1233_ _1236_
+ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a21o_1
X_4040_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__inv_2
XFILLER_110_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4942_ net173 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4873_ net1215 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3824_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__inv_1
XFILLER_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3755_ net1262 net65 net101 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0436_ sky130_fd_sc_hd__mux4_1
X_2706_ _1533_ _1203_ _1550_ _1551_ _1202_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__a311o_1
X_3686_ _0049_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2_4
XFILLER_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5425_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net517
+ sky130_fd_sc_hd__clkbuf_1
X_2637_ net204 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__mux2_1
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput243 net243 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput265 net265 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[6] sky130_fd_sc_hd__buf_2
X_2568_ _1418_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q _1419_
+ _1420_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q VGND VGND VPWR
+ VPWR _1421_ sky130_fd_sc_hd__a221o_1
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput298 net298 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput287 net287 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[12] sky130_fd_sc_hd__buf_2
X_4307_ net41 net1149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5287_ Tile_X0Y1_NN4END[15] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_4
X_2499_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR VPWR
+ _1356_ sky130_fd_sc_hd__mux2_1
X_4238_ _0855_ _0883_ _0854_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__o21a_1
X_4169_ _0819_ _0808_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__xnor2_4
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone205 net1058 VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_8
Xclone249 net1033 VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__buf_8
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3540_ _0034_ _0232_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o21a_1
X_5210_ net36 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_2
X_3471_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\] VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_1
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2422_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q _1284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_149_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2353_ net71 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__o21a_1
X_5141_ net164 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5072_ net171 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4023_ net1018 net1036 net1032 net983 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0685_ sky130_fd_sc_hd__mux4_2
X_2284_ _1152_ _1153_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__xnor2_2
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4925_ net1199 net1100 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ net1193 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3807_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q _0482_ VGND VGND
+ VPWR VPWR _0483_ sky130_fd_sc_hd__and2b_1
X_4787_ net1191 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3738_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q _0419_ VGND VGND
+ VPWR VPWR _0420_ sky130_fd_sc_hd__or2_1
XFILLER_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3669_ _0348_ _0350_ _0355_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a211o_4
XFILLER_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5408_ net151 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_1
X_5339_ Tile_X0Y0_WW4END[14] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__buf_4
XFILLER_125_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1232 net51 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__buf_4
Xfanout1210 net155 VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__buf_4
Xfanout1221 net140 VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__buf_2
XFILLER_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1243 net1244 VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__buf_4
Xfanout1254 net33 VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2971_ _0199_ net621 _0677_ _0384_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q VGND VGND VPWR VPWR
+ _1767_ sky130_fd_sc_hd__mux4_1
X_4710_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C2 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\] sky130_fd_sc_hd__dfxtp_1
X_4641_ net55 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4572_ net1256 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3523_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q net979 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o21ba_4
XFILLER_143_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3454_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q VGND VGND VPWR
+ VPWR _0149_ sky130_fd_sc_hd__inv_1
XFILLER_130_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2405_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q _1268_ VGND VGND
+ VPWR VPWR _1269_ sky130_fd_sc_hd__nand2_1
X_3385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q VGND VGND VPWR
+ VPWR _0080_ sky130_fd_sc_hd__inv_1
XFILLER_111_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2336_ net79 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__mux2_4
X_5124_ net1210 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2267_ _1041_ _1137_ _1040_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__a21o_4
X_5055_ net1201 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4006_ net1019 net1038 net986 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0669_ sky130_fd_sc_hd__mux4_1
X_2198_ _1052_ _1059_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__xor2_2
XFILLER_25_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4908_ net1218 net1108 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_121_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4839_ net1213 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1040 net1041 VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__buf_8
X_3170_ net175 net211 net120 net996 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q VGND VGND VPWR VPWR
+ _1919_ sky130_fd_sc_hd__mux4_1
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2121_ _0991_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__nand2_1
Xfanout1051 net1052 VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__buf_6
Xfanout1062 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q VGND VGND
+ VPWR VPWR net1062 sky130_fd_sc_hd__clkbuf_4
Xfanout1073 net212 VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__clkbuf_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1095 net1097 VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__buf_2
Xfanout1084 net1085 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__buf_2
X_2052_ _0926_ _0907_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A0 sky130_fd_sc_hd__mux2_4
Xrebuffer18 _0258_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2954_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q net1042 VGND
+ VGND VPWR VPWR _1760_ sky130_fd_sc_hd__nor2_1
X_2885_ net57 net61 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q VGND
+ VGND VPWR VPWR _1708_ sky130_fd_sc_hd__mux2_1
X_4624_ net1242 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4555_ net1235 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3506_ _0097_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__and2_1
X_4486_ net50 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_112_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3437_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR
+ VPWR _0132_ sky130_fd_sc_hd__inv_1
X_3368_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0063_ sky130_fd_sc_hd__inv_2
XFILLER_97_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2319_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q _1183_ _1188_
+ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__o21ba_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5107_ net168 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3299_ net819 _2021_ _2030_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ _0197_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_84_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5038_ net1186 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 Tile_X0Y0_W2MID[5] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput121 Tile_X0Y1_E1END[2] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xinput132 Tile_X0Y1_E2MID[1] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_2
Xinput143 Tile_X0Y1_EE4END[2] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xinput154 Tile_X0Y1_FrameData[18] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xinput187 Tile_X0Y1_N2MID[1] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_4
Xinput176 Tile_X0Y1_N1END[2] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__buf_4
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput165 Tile_X0Y1_FrameData[30] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_4
Xinput198 Tile_X0Y1_N4END[4] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_4
XFILLER_29_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2670_ Tile_X0Y1_DSP_bot.C0 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\] net1065 VGND
+ VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux2_2
XFILLER_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput606 net606 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[14] sky130_fd_sc_hd__buf_2
X_4340_ net1247 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4271_ net43 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3222_ _1963_ _1962_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__mux2_1
X_3153_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q net833 _1907_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q VGND VGND VPWR VPWR
+ _1908_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2104_ net189 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net225
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q
+ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__mux4_2
X_3084_ net1263 net1225 net815 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _1861_ sky130_fd_sc_hd__mux4_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3986_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q _0072_ _0650_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0651_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2937_ net188 net199 net1261 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_99_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2868_ _0176_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__or2_1
X_4607_ net28 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2799_ _1601_ _1623_ _1624_ _1622_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__a31o_1
X_4538_ net33 net1089 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4469_ net1248 net1105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_215 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_204 net1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_237 net186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_248 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_259 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3840_ net198 net1262 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
XFILLER_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3771_ _0051_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or2_1
X_5510_ Tile_X0Y1_WW4END[5] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_4
X_2722_ _1410_ _1527_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__xnor2_2
XFILLER_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net533
+ sky130_fd_sc_hd__buf_1
X_2653_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__inv_6
Xoutput414 net414 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput425 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR
+ Tile_X0Y0_WW4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput403 net403 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[2] sky130_fd_sc_hd__buf_2
X_2584_ net185 net130 net76 net232 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q VGND VGND VPWR VPWR
+ _1436_ sky130_fd_sc_hd__mux4_2
X_5372_ Tile_X0Y1_E6END[9] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_1
XFILLER_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput436 net436 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[9] sky130_fd_sc_hd__buf_2
X_4323_ net1230 net1147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput469 net469 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput447 net447 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput458 net458 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_113_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4254_ _0899_ _0898_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__nor2_8
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4185_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q _0835_ VGND VGND
+ VPWR VPWR _0836_ sky130_fd_sc_hd__and2b_1
X_3205_ net980 net656 net1000 net995 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q VGND VGND VPWR VPWR
+ _1949_ sky130_fd_sc_hd__mux4_1
X_3136_ net1003 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 _0413_ _0405_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3067_ _1846_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__a21bo_1
XFILLER_94_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3969_ _0020_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer291 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND VGND VPWR VPWR net908
+ sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer280 net898 VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4941_ net1219 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_106_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4872_ net1214 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3823_ net868 net70 net14 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q VGND VGND VPWR VPWR
+ _0498_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_50_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3754_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q _0434_ VGND VGND
+ VPWR VPWR _0435_ sky130_fd_sc_hd__and2b_1
X_2705_ _1199_ _1201_ _1548_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__a21oi_1
X_3685_ net1050 net1045 net1026 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0372_ sky130_fd_sc_hd__mux4_2
X_5424_ net1193 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_4
X_2636_ net83 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__mux2_1
Xoutput244 net244 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput266 net266 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[8] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput255 net255 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[7] sky130_fd_sc_hd__buf_2
X_5355_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net447
+ sky130_fd_sc_hd__clkbuf_1
X_2567_ net188 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__o21ba_1
X_5286_ Tile_X0Y1_NN4END[14] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_1
Xoutput299 net299 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[13] sky130_fd_sc_hd__buf_2
X_4306_ net42 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2498_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6
+ _1354_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q VGND VGND VPWR
+ VPWR _1355_ sky130_fd_sc_hd__o211a_1
XFILLER_114_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4237_ _0879_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4168_ _0819_ _0808_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__and2b_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4099_ _0746_ _0745_ _0754_ _0102_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__a221o_1
XFILLER_15_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3119_ net987 _0214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 _0228_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_66_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclone206 net1039 VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__buf_8
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3470_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q VGND VGND VPWR
+ VPWR _0165_ sky130_fd_sc_hd__inv_1
X_2421_ net176 net1224 net184 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _1284_ sky130_fd_sc_hd__mux4_1
X_2352_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q _1216_ VGND VGND
+ VPWR VPWR _1220_ sky130_fd_sc_hd__nand2_1
X_5140_ net167 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_149_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2283_ _1152_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nand2b_4
X_5071_ net1187 net1170 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4022_ _0679_ _0682_ _0683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR
+ _0684_ sky130_fd_sc_hd__o221a_1
XFILLER_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4924_ net1198 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4855_ net1220 net1125 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4786_ net1190 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3806_ net179 net195 net1223 net124 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _0482_ sky130_fd_sc_hd__mux4_1
X_3737_ net60 net68 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q VGND
+ VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
XFILLER_118_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3668_ _0348_ _0350_ _0355_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ sky130_fd_sc_hd__a21o_4
X_3599_ net201 net23 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
X_2619_ net190 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__mux2_4
X_5407_ net150 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_1
X_5338_ Tile_X0Y0_WW4END[13] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_4
X_5269_ Tile_X0Y1_N4END[13] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_1
XFILLER_18_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1222 net139 VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__clkbuf_4
Xfanout1200 net159 VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__buf_4
Xfanout1211 net154 VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__buf_4
XFILLER_78_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1244 Tile_X0Y0_FrameData[24] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__clkbuf_2
Xfanout1233 net50 VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1255 net32 VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2970_ net824 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net641 _0317_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ net56 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_62_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4571_ net1255 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_155_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3522_ _0211_ _0212_ _0213_ _0031_ _0032_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a221o_4
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3453_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q VGND VGND VPWR
+ VPWR _0148_ sky130_fd_sc_hd__inv_2
X_2404_ net89 net232 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__mux2_1
X_3384_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q VGND VGND VPWR
+ VPWR _0079_ sky130_fd_sc_hd__inv_1
X_5123_ net1208 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2335_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q VGND VGND VPWR VPWR
+ _1204_ sky130_fd_sc_hd__mux4_2
XFILLER_111_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2266_ _1067_ _1134_ _1087_ _1066_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__a31o_4
XFILLER_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5054_ net1200 net1173 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4005_ _0667_ _0640_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nor2_8
X_2197_ _1063_ _1062_ _1056_ _1058_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__o211ai_2
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4907_ net1217 net1108 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_80_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4838_ net1212 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4769_ net1206 net1144 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 net236 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1030 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VGND VGND VPWR VPWR
+ net1030 sky130_fd_sc_hd__clkbuf_4
Xfanout1052 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 VGND VGND VPWR VPWR
+ net1052 sky130_fd_sc_hd__buf_8
Xfanout1041 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 VGND VGND VPWR VPWR
+ net1041 sky130_fd_sc_hd__buf_8
X_2120_ _0937_ _0942_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__xor2_2
XFILLER_86_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1063 net1065 VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__clkbuf_4
Xfanout1074 net1075 VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__clkbuf_2
Xfanout1096 net1097 VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__clkbuf_2
Xfanout1085 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__buf_2
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2051_ _0925_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q _0912_
+ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer19 _0334_ VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_137_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2953_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q _0554_ _1758_
+ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_45_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2884_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q _1704_ _1706_
+ _0175_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__o211a_1
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4623_ net1240 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4554_ net1234 net1079 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3505_ net1020 net1036 net1032 net985 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0200_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_112_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4485_ net51 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q VGND VGND VPWR
+ VPWR _0131_ sky130_fd_sc_hd__inv_1
X_3367_ net188 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__inv_1
X_2318_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q _1185_ _1187_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q VGND VGND VPWR VPWR
+ _1188_ sky130_fd_sc_hd__a31o_1
XFILLER_97_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5106_ net169 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3298_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__or2_1
X_5037_ net1219 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2249_ _1113_ _1109_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_84_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput100 Tile_X0Y0_W2END[3] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
Xinput111 Tile_X0Y0_W2MID[6] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_2
XFILLER_88_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput122 Tile_X0Y1_E1END[3] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
Xinput133 Tile_X0Y1_E2MID[2] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xinput144 Tile_X0Y1_EE4END[3] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xinput177 Tile_X0Y1_N1END[3] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_4
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput155 Tile_X0Y1_FrameData[19] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xinput166 Tile_X0Y1_FrameData[31] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_4
Xinput199 Tile_X0Y1_N4END[5] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
Xinput188 Tile_X0Y1_N2MID[2] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_59_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput607 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y1_WW4BEG[15] sky130_fd_sc_hd__buf_6
XFILLER_140_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ net44 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3221_ net1025 _0823_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__mux2_1
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3152_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q net1021 VGND
+ VGND VPWR VPWR _1907_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_145_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2103_ _0974_ _0973_ _0975_ _0145_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a221o_1
X_3083_ _1859_ _1857_ _1860_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o22a_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3985_ net64 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q VGND VGND
+ VPWR VPWR _0650_ sky130_fd_sc_hd__nor2_1
X_2936_ _1746_ _1748_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_154_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2867_ net1 net5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q VGND
+ VGND VPWR VPWR _1691_ sky130_fd_sc_hd__mux2_1
X_4606_ net29 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2798_ _1626_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 sky130_fd_sc_hd__mux2_4
XFILLER_116_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4537_ net34 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4468_ net1247 net1105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3419_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR
+ VPWR _0114_ sky130_fd_sc_hd__inv_2
X_4399_ net1240 net1121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_205 net1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_249 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_238 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_227 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3770_ net989 net1024 net994 net1008 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR VPWR
+ _0450_ sky130_fd_sc_hd__mux4_1
X_2721_ _1561_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5440_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net532
+ sky130_fd_sc_hd__buf_2
X_2652_ _1499_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] net1067 VGND VGND VPWR VPWR
+ _1500_ sky130_fd_sc_hd__mux2_4
Xoutput415 net415 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[4] sky130_fd_sc_hd__buf_2
Xoutput426 net426 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[14] sky130_fd_sc_hd__buf_8
Xoutput404 net404 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[3] sky130_fd_sc_hd__buf_2
X_5371_ Tile_X0Y1_E6END[8] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_1
X_2583_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q _1431_ _1434_
+ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__a21o_1
X_4322_ net1229 net1147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput437 net437 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput448 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 VGND VGND VPWR VPWR
+ Tile_X0Y1_E2BEG[7] sky130_fd_sc_hd__buf_6
Xoutput459 net459 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[11] sky130_fd_sc_hd__buf_6
XFILLER_113_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4253_ _0522_ _0818_ _0817_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__o21ba_4
XFILLER_113_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3204_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q _1947_ VGND
+ VGND VPWR VPWR _1948_ sky130_fd_sc_hd__or2_1
X_4184_ net811 net869 net977 net988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0835_ sky130_fd_sc_hd__mux4_1
X_3135_ _1896_ _1897_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3066_ _0700_ _1535_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__mux2_4
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3968_ net194 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q VGND VGND
+ VPWR VPWR _0634_ sky130_fd_sc_hd__or2_1
XFILLER_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2919_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__inv_2
X_3899_ _0569_ _0567_ _0541_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4
+ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_118_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer292 net927 VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__buf_6
Xrebuffer270 net888 VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer281 net899 VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_154_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4940_ net1218 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4871_ net152 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3822_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0496_ VGND VGND
+ VPWR VPWR _0497_ sky130_fd_sc_hd__or2_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3753_ net637 net198 net190 net9 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q VGND VGND VPWR VPWR
+ _0434_ sky130_fd_sc_hd__mux4_2
X_2704_ _1548_ _1549_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__and2_4
X_3684_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q _0370_ VGND VGND
+ VPWR VPWR _0371_ sky130_fd_sc_hd__nor2_1
X_5423_ net165 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkbuf_2
X_2635_ _1482_ _1481_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__xnor2_4
XFILLER_145_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5354_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net446
+ sky130_fd_sc_hd__clkbuf_1
X_4305_ net1243 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput267 net267 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[9] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[5] sky130_fd_sc_hd__buf_2
X_2566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q _0677_ VGND VGND
+ VPWR VPWR _1419_ sky130_fd_sc_hd__nand2_1
X_5285_ Tile_X0Y1_NN4END[13] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__buf_1
Xoutput289 net289 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput278 net278 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[4] sky130_fd_sc_hd__buf_2
X_2497_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q _1353_ VGND VGND
+ VPWR VPWR _1354_ sky130_fd_sc_hd__nand2_1
X_4236_ _0880_ _0614_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__xnor2_2
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4167_ _0522_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3118_ net1025 net918 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 _0405_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_82_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4098_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net15 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3049_ net93 net1044 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__mux2_1
XFILLER_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone207 net1027 VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__buf_6
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q VGND VGND
+ VPWR VPWR net617 sky130_fd_sc_hd__clkbuf_4
X_2420_ _1281_ _1280_ _1282_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ _0154_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__a221o_1
XFILLER_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2351_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net15 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__mux2_1
XFILLER_150_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2282_ _0810_ _0892_ _0894_ _0891_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__o2bb2ai_1
X_5070_ net1186 net1170 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4021_ net190 net9 net87 net101 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q VGND VGND VPWR VPWR
+ _0683_ sky130_fd_sc_hd__mux4_2
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4923_ net162 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_63_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4854_ net1209 net1125 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4785_ net1189 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3805_ _0479_ _0480_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_4
X_3736_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q _0415_ _0417_
+ _0113_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__o211a_1
XFILLER_146_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3667_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__inv_2
X_3598_ net80 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_4
X_5406_ net149 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_4
X_2618_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q net660 _1467_
+ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__a21o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5337_ Tile_X0Y0_WW4END[12] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_4
X_2549_ _1402_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__inv_1
X_5268_ Tile_X0Y1_N4END[12] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4219_ net995 net1025 net1005 net1012 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0867_ sky130_fd_sc_hd__mux4_1
X_5199_ net54 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1212 net153 VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__buf_4
Xfanout1223 net122 VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__buf_4
Xfanout1201 net1202 VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1234 net49 VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__buf_4
Xfanout1245 net42 VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__buf_4
Xfanout1256 net31 VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__buf_4
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ net1254 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_155_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3521_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__inv_2
X_3452_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q VGND VGND VPWR
+ VPWR _0147_ sky130_fd_sc_hd__inv_1
X_3383_ net115 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2403_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q net630 _1266_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR
+ _1267_ sky130_fd_sc_hd__a211o_1
XFILLER_130_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2334_ _1201_ _1199_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__xor2_2
X_5122_ net1207 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_111_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2265_ _1067_ _1087_ _1134_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__and3_1
X_5053_ net1199 net1170 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2196_ _1042_ _1065_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__xnor2_1
X_4004_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ net1062 _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__o21ai_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4906_ net1216 net1108 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4837_ net154 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4768_ net1204 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4699_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] sky130_fd_sc_hd__dfxtp_1
X_3719_ net1222 net71 net216 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0403_ sky130_fd_sc_hd__mux4_1
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 net244 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1020 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 VGND VGND VPWR VPWR
+ net1020 sky130_fd_sc_hd__buf_8
Xfanout1031 net1033 VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__buf_8
Xfanout1042 net1044 VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__buf_2
Xfanout1053 net1055 VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__buf_2
Xfanout1064 net1065 VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__clkbuf_4
Xfanout1086 net1089 VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__buf_2
Xfanout1075 net1077 VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__buf_2
Xfanout1097 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__clkbuf_2
X_2050_ net192 net228 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_37_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2952_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q VGND VGND VPWR VPWR
+ _1758_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_45_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2883_ _0174_ _1705_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__or2_1
X_4622_ net44 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4553_ net27 net1089 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3504_ net1019 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__inv_1
X_4484_ net52 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3435_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q VGND VGND VPWR
+ VPWR _0130_ sky130_fd_sc_hd__inv_2
XFILLER_131_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3366_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q VGND VGND VPWR
+ VPWR _0061_ sky130_fd_sc_hd__inv_2
X_2317_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q _1186_ VGND VGND
+ VPWR VPWR _1187_ sky130_fd_sc_hd__nand2_1
X_3297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q _2028_ _2024_
+ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__and3b_1
X_5105_ net170 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5036_ net1218 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2248_ _1115_ _1111_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__xnor2_2
XFILLER_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2179_ _0984_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nor2_4
XFILLER_72_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 Tile_X0Y0_W2END[4] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_8_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput112 Tile_X0Y0_W2MID[7] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput134 Tile_X0Y1_E2MID[3] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_2
Xinput123 Tile_X0Y1_E2END[0] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xinput145 Tile_X0Y1_FrameData[0] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
Xinput178 Tile_X0Y1_N2END[0] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_2
Xinput156 Tile_X0Y1_FrameData[1] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_2
Xinput167 Tile_X0Y1_FrameData[3] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
Xinput189 Tile_X0Y1_N2MID[3] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_59_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput608 net608 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_98_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3220_ _0977_ _1380_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__mux2_1
X_3151_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q net662 _1905_
+ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__a21o_1
XFILLER_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2102_ net188 net133 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__mux2_1
X_3082_ _0279_ net94 net58 net1051 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _1860_ sky130_fd_sc_hd__mux4_1
X_3984_ _0646_ _0647_ _0648_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR VPWR
+ _0649_ sky130_fd_sc_hd__a221o_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q _0359_ _1747_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q VGND VGND VPWR VPWR
+ _1748_ sky130_fd_sc_hd__a211o_1
XFILLER_148_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2866_ _0239_ net186 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__mux2_1
XFILLER_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4605_ net30 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2797_ _1623_ _1625_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__xnor2_2
XFILLER_117_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4536_ net1252 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4467_ net41 net1105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4398_ net1239 net1121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3418_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR
+ VPWR _0113_ sky130_fd_sc_hd__inv_2
XFILLER_77_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q VGND VGND VPWR
+ VPWR _0044_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_206 net1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5019_ net1197 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_217 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_239 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_228 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2720_ _1526_ _1430_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__xnor2_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2651_ Tile_X0Y1_DSP_bot.C1 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\] net1063 VGND
+ VGND VPWR VPWR _1499_ sky130_fd_sc_hd__mux2_4
XFILLER_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput416 net416 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput405 net405 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[4] sky130_fd_sc_hd__buf_2
X_5370_ Tile_X0Y1_E6END[7] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_1
X_2582_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q _1433_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q
+ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__o21ai_1
Xoutput427 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y0_WW4BEG[15] sky130_fd_sc_hd__buf_6
X_4321_ net1228 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput449 net449 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput438 net438 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[1] sky130_fd_sc_hd__buf_6
X_4252_ _0896_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__or2_1
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3203_ net1223 net1072 net655 net971 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1947_ sky130_fd_sc_hd__mux4_1
X_4183_ net992 net1021 net1003 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0834_ sky130_fd_sc_hd__mux4_1
XFILLER_67_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3134_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 _1378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__mux2_1
XFILLER_27_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3065_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q _0571_ _1844_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q VGND VGND VPWR VPWR
+ _1845_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_2_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3967_ net81 net818 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q VGND
+ VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux2_1
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2918_ net62 net78 net98 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _1733_ sky130_fd_sc_hd__mux4_1
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3898_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0568_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__o21ba_1
X_2849_ _1653_ _1672_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__nand2_1
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4519_ net1236 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5499_ Tile_X0Y1_W6END[4] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer260 net878 VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer271 net889 VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer282 net900 VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4870_ net153 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3821_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net13 net69 _0495_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q VGND VGND VPWR VPWR
+ _0496_ sky130_fd_sc_hd__mux4_1
X_3752_ _0431_ _0432_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_4
X_2703_ _1545_ _1547_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__or2_1
X_3683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0367_ _0369_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR VPWR
+ _0370_ sky130_fd_sc_hd__o211a_1
XFILLER_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5422_ net163 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_2
X_2634_ _1482_ _1481_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__nand2_2
X_2565_ net224 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q
+ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__mux2_2
X_5353_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net445
+ sky130_fd_sc_hd__buf_1
X_4304_ net1241 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput257 net257 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[10] sky130_fd_sc_hd__buf_8
Xoutput268 net268 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[6] sky130_fd_sc_hd__buf_8
X_5284_ Tile_X0Y1_NN4END[12] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__buf_1
Xoutput279 net279 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[5] sky130_fd_sc_hd__buf_2
X_2496_ _1353_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__inv_2
X_4235_ _0613_ _0799_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__nor2_1
X_4166_ _0809_ _0816_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__xor2_1
XFILLER_101_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3117_ net995 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 net666 _1378_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 sky130_fd_sc_hd__mux4_1
X_4097_ _0748_ _0750_ _0753_ _0100_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ sky130_fd_sc_hd__a22o_4
XFILLER_55_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3048_ _0027_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4999_ net1213 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_139_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2350_ _1204_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q VGND VGND
+ VPWR VPWR _1218_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_149_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2281_ _1150_ _0893_ _1151_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__o21ai_4
X_4020_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q _0681_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4922_ net163 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4853_ net1195 net1125 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4784_ net1188 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3804_ net994 net1023 net1004 net1011 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _0480_ sky130_fd_sc_hd__mux4_2
XFILLER_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3735_ _0112_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or2_1
XFILLER_20_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5405_ net1217 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_2
X_3666_ _0069_ _0351_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o21ai_2
X_3597_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q _0287_ _0283_
+ _0201_ _0203_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ sky130_fd_sc_hd__o32a_4
X_2617_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q _1466_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__o21ai_1
X_5336_ Tile_X0Y0_WW4END[11] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__buf_4
XFILLER_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2548_ net191 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net227
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q
+ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux4_1
X_5267_ Tile_X0Y1_N4END[11] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XFILLER_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2479_ net76 net1072 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__mux2_1
X_4218_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _0865_ VGND VGND
+ VPWR VPWR _0866_ sky130_fd_sc_hd__or2_1
X_5198_ net1230 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4149_ _0710_ _0784_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
XFILLER_137_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1213 net152 VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__buf_4
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1202 Tile_X0Y1_FrameData[24] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__clkbuf_2
Xfanout1235 net48 VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1246 net41 VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__clkbuf_4
Xfanout1224 net121 VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__clkbuf_4
XFILLER_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1257 net30 VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__buf_4
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3520_ net651 _0212_ _0213_ _0031_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_155_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3451_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR
+ VPWR _0146_ sky130_fd_sc_hd__inv_2
X_3382_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q VGND VGND VPWR
+ VPWR _0077_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_114_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2402_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q _0442_ VGND VGND
+ VPWR VPWR _1266_ sky130_fd_sc_hd__nor2_1
XFILLER_69_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2333_ _1199_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nor2_1
X_5121_ net1205 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2264_ _1088_ _1086_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__nor2_4
X_5052_ net1198 net1170 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4003_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] net1062 VGND VGND VPWR VPWR _0666_
+ sky130_fd_sc_hd__nand2b_1
X_2195_ _1065_ _1042_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__and2b_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4905_ net1215 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_23_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4836_ net1210 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_31_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4767_ net1202 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4698_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] sky130_fd_sc_hd__dfxtp_1
X_3718_ net180 net196 net119 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0402_ sky130_fd_sc_hd__mux4_1
X_3649_ net1222 net73 net218 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0338_ sky130_fd_sc_hd__mux4_1
X_5319_ Tile_X0Y0_W6END[4] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_132_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_9 net255 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1021 net1022 VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__buf_2
Xfanout1010 net1012 VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 net1044 VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__buf_2
Xfanout1054 net1055 VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__buf_1
Xfanout1032 net1033 VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__buf_4
Xfanout1065 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q VGND VGND
+ VPWR VPWR net1065 sky130_fd_sc_hd__clkbuf_4
Xfanout1087 net1088 VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__buf_2
Xfanout1098 net1100 VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__clkbuf_4
Xfanout1076 net1077 VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__buf_2
XFILLER_74_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2951_ _1752_ _1754_ _1757_ _0082_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4621_ net45 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2882_ net1 net23 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q VGND
+ VGND VPWR VPWR _1705_ sky130_fd_sc_hd__mux2_1
X_4552_ net38 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4483_ net53 net1106 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3503_ net1045 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__inv_1
XFILLER_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3434_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR
+ VPWR _0129_ sky130_fd_sc_hd__inv_1
X_3365_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q VGND VGND VPWR
+ VPWR _0060_ sky130_fd_sc_hd__inv_2
X_2316_ net70 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__mux2_1
X_3296_ net192 _2021_ _2026_ _2027_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__a211o_1
X_5104_ net171 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5035_ net1217 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2247_ _1116_ _1106_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__xnor2_4
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2178_ _1044_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__xor2_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4819_ net1191 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput102 Tile_X0Y0_W2END[5] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput113 Tile_X0Y0_W6END[0] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_8_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput135 Tile_X0Y1_E2MID[4] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xinput124 Tile_X0Y1_E2END[1] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput168 Tile_X0Y1_FrameData[4] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
Xinput146 Tile_X0Y1_FrameData[10] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xinput157 Tile_X0Y1_FrameData[20] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_2
Xinput179 Tile_X0Y1_N2END[1] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_2
XFILLER_44_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput609 net609 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3150_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q VGND VGND VPWR VPWR
+ _1905_ sky130_fd_sc_hd__o21ai_1
X_3081_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _1858_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__a21bo_1
XFILLER_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2101_ net224 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3983_ net8 net1261 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q VGND
+ VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux2_1
X_2934_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q net1050 VGND
+ VGND VPWR VPWR _1747_ sky130_fd_sc_hd__nor2_1
X_2865_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q _1688_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__a21bo_1
XFILLER_148_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4604_ net31 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4535_ net1251 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2796_ _1601_ _1624_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_68_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4466_ net42 net1105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3417_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR
+ VPWR _0112_ sky130_fd_sc_hd__inv_2
X_4397_ net1238 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3348_ net229 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XFILLER_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3279_ _0712_ _0875_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__mux2_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5018_ net1196 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_26_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_207 net1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_218 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_229 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_86_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_95_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2650_ _1498_ _1496_ _1491_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C1 sky130_fd_sc_hd__a21oi_2
XFILLER_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput417 net417 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput406 net406 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[5] sky130_fd_sc_hd__buf_2
X_2581_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__inv_1
Xoutput428 net428 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[1] sky130_fd_sc_hd__buf_2
X_4320_ net1227 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput439 net439 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4251_ _0811_ _0814_ _0895_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3202_ _1945_ _1944_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q
+ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__mux2_1
X_4182_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__inv_2
XFILLER_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3133_ net1022 net666 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__mux2_1
X_3064_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q net1028 VGND VGND
+ VPWR VPWR _1844_ sky130_fd_sc_hd__nor2_1
XFILLER_82_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3966_ _0629_ _0627_ _0632_ _0124_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__a22o_1
X_2917_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q _1731_ VGND VGND
+ VPWR VPWR _1732_ sky130_fd_sc_hd__or2_4
XFILLER_136_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3897_ net175 net183 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0568_ sky130_fd_sc_hd__mux4_1
X_2848_ _1601_ _1623_ _1624_ _1654_ _1622_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__a311o_1
X_2779_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q _1608_ _1606_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q VGND VGND VPWR VPWR
+ _1609_ sky130_fd_sc_hd__o211a_1
XFILLER_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4518_ net1233 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5498_ Tile_X0Y1_W6END[3] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4449_ net1228 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer283 net901 VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer272 net890 VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer261 net879 VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer294 net913 VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_15_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3751_ net1050 net1045 net824 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0432_ sky130_fd_sc_hd__mux4_2
X_2702_ _1547_ _1545_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__nand2_2
XFILLER_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3682_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q _0368_ VGND VGND
+ VPWR VPWR _0369_ sky130_fd_sc_hd__nand2_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5421_ net162 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkbuf_2
X_2633_ _1127_ _1126_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_117_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2564_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q _1416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ _1415_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__o211a_1
X_5352_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net444
+ sky130_fd_sc_hd__clkbuf_2
X_4303_ net1240 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput258 net258 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[11] sky130_fd_sc_hd__buf_6
Xoutput247 net247 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[0] sky130_fd_sc_hd__buf_2
X_5283_ Tile_X0Y1_NN4END[11] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_1
Xoutput269 net269 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[10] sky130_fd_sc_hd__buf_2
X_2495_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q _1352_ _1350_
+ _1344_ _1345_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__o32a_4
X_4234_ _0478_ _0799_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_1
X_4165_ _0814_ _0809_ _0815_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__and3_1
XFILLER_55_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3116_ _1882_ _1884_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__nand2_1
X_4096_ _0751_ _0752_ _0099_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3047_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q _0239_ VGND
+ VGND VPWR VPWR _1830_ sky130_fd_sc_hd__or2_1
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4998_ net1212 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3949_ _0613_ _0521_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__nor2_4
XFILLER_139_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2280_ _0667_ net618 _0710_ _0521_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__o22ai_2
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4921_ net165 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_32_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4852_ net1192 net1125 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3803_ net969 net978 net998 net989 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _0479_ sky130_fd_sc_hd__mux4_1
XFILLER_60_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4783_ net1187 net1150 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_71_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3734_ net1263 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3665_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q _0352_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o21a_1
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5404_ net147 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_1
X_2616_ net183 net128 net90 net219 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q VGND VGND VPWR VPWR
+ _1466_ sky130_fd_sc_hd__mux4_2
X_3596_ _0096_ _0286_ _0285_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o211a_1
X_5335_ Tile_X0Y0_WW4END[10] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_4
X_2547_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1400_ VGND VGND
+ VPWR VPWR _1401_ sky130_fd_sc_hd__or2_1
X_5266_ Tile_X0Y1_N4END[10] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2478_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1336_ VGND VGND
+ VPWR VPWR _1337_ sky130_fd_sc_hd__and2b_1
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4217_ net923 net971 net981 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0865_ sky130_fd_sc_hd__mux4_1
X_5197_ net52 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__buf_2
X_4148_ _0799_ net622 VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_87_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4079_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__inv_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload1 clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_50_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1214 net151 VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__buf_4
Xfanout1203 net1204 VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__clkbuf_4
Xfanout1225 net96 VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__clkbuf_4
Xfanout1236 net47 VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__buf_4
XFILLER_120_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1247 net40 VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__clkbuf_4
Xfanout1258 net29 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3450_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q VGND VGND VPWR
+ VPWR _0145_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_114_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3381_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q VGND VGND VPWR
+ VPWR _0076_ sky130_fd_sc_hd__inv_2
X_2401_ _1260_ _1262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ _1265_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 sky130_fd_sc_hd__o22a_1
X_2332_ _1200_ _1161_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__or2_4
X_5120_ net1203 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5051_ net1197 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4002_ _0664_ _0107_ _0665_ _0660_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ sky130_fd_sc_hd__a31o_4
X_2263_ _1105_ _1132_ _1104_ _1088_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__a211o_1
X_2194_ _1062_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__and2b_1
XFILLER_65_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4904_ net1214 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_23_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4835_ net1208 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4766_ net1200 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3717_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q _0400_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_31_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4697_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3648_ net182 net1224 net194 net127 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q VGND VGND VPWR VPWR
+ _0337_ sky130_fd_sc_hd__mux4_1
X_3579_ net994 net1023 net1004 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0270_ sky130_fd_sc_hd__mux4_2
X_5318_ Tile_X0Y0_W6END[3] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_132_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5249_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR net341
+ sky130_fd_sc_hd__buf_1
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1022 net1024 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__clkbuf_2
Xfanout1011 net1012 VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__buf_6
Xfanout1000 net1001 VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__clkbuf_4
Xfanout1055 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 VGND VGND VPWR VPWR
+ net1055 sky130_fd_sc_hd__buf_2
Xfanout1044 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 VGND VGND VPWR VPWR
+ net1044 sky130_fd_sc_hd__clkbuf_4
Xfanout1033 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 VGND VGND VPWR VPWR
+ net1033 sky130_fd_sc_hd__buf_8
XFILLER_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1088 net1089 VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__buf_2
Xfanout1077 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1066 net1067 VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__buf_2
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1099 net1100 VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2950_ _1755_ _1756_ _0081_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _0239_ net186 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_106_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4620_ net46 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4551_ net1236 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4482_ net1229 net1106 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3502_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR
+ VPWR _0197_ sky130_fd_sc_hd__inv_2
XFILLER_143_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3433_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR
+ VPWR _0128_ sky130_fd_sc_hd__inv_1
XFILLER_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3364_ net86 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__inv_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5103_ net172 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2315_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q _1184_ VGND VGND
+ VPWR VPWR _1185_ sky130_fd_sc_hd__nand2b_1
X_3295_ net131 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _0196_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR VPWR
+ _2027_ sky130_fd_sc_hd__a31o_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5034_ net1216 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2246_ _1116_ _1106_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_123_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2177_ _1047_ _1005_ _1046_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__a21bo_4
XTAP_TAPCELL_ROW_36_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4818_ net1190 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4749_ net1219 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_133_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput103 Tile_X0Y0_W2END[6] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
Xinput114 Tile_X0Y0_W6END[1] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_4
XFILLER_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput136 Tile_X0Y1_E2MID[5] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_2
Xinput125 Tile_X0Y1_E2END[2] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
Xinput169 Tile_X0Y1_FrameData[5] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
Xinput147 Tile_X0Y1_FrameData[11] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
Xinput158 Tile_X0Y1_FrameData[21] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_2
XFILLER_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3080_ _1616_ _0528_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__mux2_4
X_2100_ _0966_ _0968_ _0141_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_109_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3982_ _0048_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q
+ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2933_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q _0384_ _1745_
+ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__a21o_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2864_ net1043 net1047 net1055 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q VGND VGND VPWR VPWR
+ _1688_ sky130_fd_sc_hd__mux4_1
X_2795_ _1173_ _1552_ _1572_ _1599_ _1172_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__a221o_1
X_4603_ net32 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4534_ net1250 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4465_ net1243 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4396_ net1237 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3416_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q VGND VGND VPWR
+ VPWR _0111_ sky130_fd_sc_hd__inv_1
XFILLER_112_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3347_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR
+ VPWR _0042_ sky130_fd_sc_hd__inv_1
XFILLER_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3278_ _1473_ _1400_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__mux2_1
X_5017_ net1194 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2229_ _1047_ _1093_ _1095_ _1097_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__a31o_1
XANTENNA_219 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_208 net1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput407 net407 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[6] sky130_fd_sc_hd__buf_2
X_2580_ net197 net141 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__mux2_1
Xoutput418 net418 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput429 net429 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4250_ _0811_ _0814_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__a21oi_1
X_4181_ net143 net83 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q VGND
+ VGND VPWR VPWR _0832_ sky130_fd_sc_hd__mux2_1
X_3201_ net1025 net1005 net812 net1009 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1945_ sky130_fd_sc_hd__mux4_1
X_3132_ _1893_ _1895_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__nand2_1
X_3063_ _1843_ _1842_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 sky130_fd_sc_hd__mux2_1
XFILLER_103_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3965_ _0630_ _0631_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q
+ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2916_ _0414_ net6 net187 net1261 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q VGND VGND VPWR VPWR
+ _1731_ sky130_fd_sc_hd__mux4_2
X_3896_ _0565_ _0564_ _0566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ _0091_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a221o_1
X_2847_ _1670_ _1669_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__nor2_8
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2778_ _1607_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__inv_2
X_4517_ net1232 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5497_ Tile_X0Y1_W6END[2] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_2
X_4448_ net1227 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4379_ net1255 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_37_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer240 net858 VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer273 net891 VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer251 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR
+ net868 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer262 net880 VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer295 net911 VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__clkbuf_2
Xrebuffer284 net902 VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_118_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3750_ net1017 net823 net866 net867 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0431_ sky130_fd_sc_hd__mux4_2
X_2701_ _1546_ _1149_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nor2_2
X_3681_ net100 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
X_5420_ net1198 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_2
X_2632_ _1480_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] net1066 VGND VGND VPWR VPWR
+ _1481_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_117_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net443
+ sky130_fd_sc_hd__clkbuf_2
X_2563_ net181 net126 net89 net217 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q VGND VGND VPWR VPWR
+ _1416_ sky130_fd_sc_hd__mux4_1
X_5282_ Tile_X0Y1_NN4END[10] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_1
X_4302_ net1239 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput259 net259 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput237 net237 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4233_ _0521_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__or2_1
X_2494_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1351_ VGND VGND
+ VPWR VPWR _1352_ sky130_fd_sc_hd__nor2_1
XFILLER_4_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4164_ _0814_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nand2_1
X_4095_ net181 net197 net120 net126 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0752_ sky130_fd_sc_hd__mux4_1
XFILLER_55_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3115_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q _0257_ _1883_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q VGND VGND VPWR VPWR
+ _1884_ sky130_fd_sc_hd__a211o_1
XFILLER_67_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3046_ _1827_ _1828_ _1829_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 sky130_fd_sc_hd__o22a_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4997_ net1211 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3948_ _0478_ _0576_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__nor2_1
X_3879_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0550_ VGND VGND
+ VPWR VPWR _0551_ sky130_fd_sc_hd__and2b_1
XFILLER_151_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4920_ net166 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4851_ net1191 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3802_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ net1062 _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o21ai_4
X_4782_ net1186 net1150 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3733_ _0414_ net193 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XFILLER_118_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3664_ net655 net971 net980 net1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ _0352_ sky130_fd_sc_hd__mux4_1
XFILLER_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5403_ net146 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_1
X_2615_ _1464_ _1463_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__xnor2_2
XFILLER_133_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3595_ net94 net1225 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
X_5334_ Tile_X0Y0_WW4END[9] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_4
X_2546_ net135 net226 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__mux4_2
X_5265_ Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
X_2477_ _0563_ _0387_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux2_1
X_5196_ net51 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4216_ net182 net127 net91 net218 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q VGND VGND VPWR VPWR
+ _0864_ sky130_fd_sc_hd__mux4_2
X_4147_ net1059 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ _0798_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__o21ai_4
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4078_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q VGND
+ VGND VPWR VPWR _0736_ sky130_fd_sc_hd__mux2_1
X_3029_ net1034 net984 net1043 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR
+ _1815_ sky130_fd_sc_hd__mux4_1
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload2 clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_59_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput590 net590 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[10] sky130_fd_sc_hd__buf_2
Xfanout1204 Tile_X0Y1_FrameData[23] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__clkbuf_2
Xfanout1237 net46 VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__buf_4
Xfanout1226 net95 VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__clkbuf_4
Xfanout1215 net150 VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__clkbuf_4
Xfanout1259 net28 VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__clkbuf_4
Xfanout1248 net39 VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_77_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2400_ _1264_ _1263_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q
+ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__mux2_4
X_3380_ net209 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_1
XFILLER_130_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2331_ _0905_ _1160_ _1149_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nor3_2
XFILLER_111_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2262_ _1105_ _1132_ _1104_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__a21o_1
X_5050_ net1196 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4001_ _0439_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q VGND VGND
+ VPWR VPWR _0665_ sky130_fd_sc_hd__nand2b_1
XFILLER_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2193_ _1056_ _1058_ _1063_ _1062_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__a211o_4
XFILLER_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4903_ net1213 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_23_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4834_ net1207 net1132 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4765_ net1199 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3716_ net992 net1021 net1002 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0400_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_31_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4696_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3647_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q _0335_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a21bo_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3578_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0268_ VGND VGND
+ VPWR VPWR _0269_ sky130_fd_sc_hd__nand2_2
X_5317_ Tile_X0Y0_W6END[2] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_93_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2529_ net186 net131 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5248_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 VGND VGND VPWR VPWR net340
+ sky130_fd_sc_hd__buf_1
X_5179_ Tile_X0Y0_EE4END[7] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 VGND VGND VPWR VPWR net1001
+ sky130_fd_sc_hd__buf_8
Xfanout1012 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VGND VGND VPWR VPWR net1012
+ sky130_fd_sc_hd__buf_8
Xfanout1056 net1058 VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__buf_8
Xfanout1034 net1035 VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__buf_2
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1045 net1046 VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_8
Xfanout1023 net1024 VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__buf_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1089 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__clkbuf_2
Xfanout1078 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__buf_2
Xfanout1067 net1069 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q _1702_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__a21bo_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4550_ net1233 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4481_ net1228 net1104 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3501_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q VGND VGND VPWR
+ VPWR _0196_ sky130_fd_sc_hd__inv_2
XFILLER_116_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3432_ net226 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_1
XFILLER_131_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3363_ net199 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__inv_1
X_5102_ net173 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2314_ net868 net14 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q
+ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__mux2_2
X_3294_ net137 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__o211a_1
XFILLER_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5033_ net1215 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2245_ _1111_ _1114_ _1107_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__o21ai_2
XFILLER_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2176_ _0611_ _0847_ _0612_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_123_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4817_ net1189 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4748_ net1218 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4679_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0007_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_103_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput104 Tile_X0Y0_W2END[7] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_2
XFILLER_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput115 Tile_X0Y0_WW4END[0] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
Xinput126 Tile_X0Y1_E2END[3] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput137 Tile_X0Y1_E2MID[6] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
Xinput148 Tile_X0Y1_FrameData[12] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
Xinput159 Tile_X0Y1_FrameData[25] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3981_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q _0279_ VGND VGND
+ VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
X_2932_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q VGND VGND VPWR VPWR
+ _1745_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2863_ _0177_ _1686_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__and2_1
X_2794_ _1604_ _1621_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__xor2_1
X_4602_ net33 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_156_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4533_ net1248 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ net1241 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4395_ net48 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3415_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q VGND VGND VPWR
+ VPWR _0110_ sky130_fd_sc_hd__inv_1
X_3346_ net57 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_90_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q _2005_ _2007_
+ _2010_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 sky130_fd_sc_hd__a22o_1
X_5016_ net166 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2228_ _1091_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__nor2_4
XANTENNA_209 net1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2159_ _0521_ net832 VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__nor2_2
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput408 net408 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput419 net419 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4180_ net221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__mux2_2
X_3200_ _0823_ _0977_ _1497_ net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1944_ sky130_fd_sc_hd__mux4_1
X_3131_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q net833 _1894_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR
+ _1895_ sky130_fd_sc_hd__a211o_1
XFILLER_79_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3062_ net637 net59 net1226 net1034 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q VGND VGND VPWR VPWR
+ _1843_ sky130_fd_sc_hd__mux4_1
XFILLER_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3964_ net71 net216 net83 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q VGND VGND VPWR VPWR
+ _0631_ sky130_fd_sc_hd__mux4_1
X_2915_ _0055_ _1726_ _1728_ _1730_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5
+ sky130_fd_sc_hd__o22a_4
XFILLER_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3895_ net211 net1072 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux2_1
X_2846_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q _1572_ _1668_
+ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__a21oi_1
X_2777_ net22 net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q VGND
+ VGND VPWR VPWR _1607_ sky130_fd_sc_hd__mux2_1
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4516_ net1231 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ net229 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkbuf_2
X_4447_ net28 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4378_ net1254 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3329_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q VGND VGND VPWR
+ VPWR _0024_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_129_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer241 net859 VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__clkbuf_2
Xrebuffer230 net848 VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__clkbuf_2
Xrebuffer274 net892 VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer263 net881 VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer296 net914 VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__clkbuf_1
XFILLER_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer285 net903 VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_151_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2700_ _1148_ _1146_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__and2b_1
XFILLER_9_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3680_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__inv_1
X_2631_ Tile_X0Y1_DSP_bot.C2 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\] net1063 VGND
+ VGND VPWR VPWR _1480_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_117_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5350_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net442
+ sky130_fd_sc_hd__buf_1
X_2562_ _1411_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q _1414_
+ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__a21o_1
XFILLER_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5281_ Tile_X0Y1_NN4END[9] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_1
X_4301_ net45 net1149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput249 net249 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput238 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 VGND VGND VPWR VPWR
+ Tile_X0Y0_E1BEG[2] sky130_fd_sc_hd__buf_8
XFILLER_87_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4232_ net1061 Tile_X0Y1_DSP_bot.B2 _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__o21ai_4
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2493_ net177 net185 net1223 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1351_ sky130_fd_sc_hd__mux4_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4163_ _0576_ _0762_ _0813_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__o21ai_1
X_4094_ net140 net72 net217 net233 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0751_ sky130_fd_sc_hd__mux4_1
X_3114_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q net991 VGND VGND
+ VPWR VPWR _1883_ sky130_fd_sc_hd__nor2_1
X_3045_ net920 net1225 net4 net986 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR
+ _1829_ sky130_fd_sc_hd__mux4_1
XFILLER_67_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4996_ net155 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3947_ _0613_ _0576_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nor2_4
XFILLER_23_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3878_ net1261 net62 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__mux2_1
X_2829_ _1654_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_96_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5479_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net571
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ net1190 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3801_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] net1062 VGND VGND VPWR VPWR _0477_
+ sky130_fd_sc_hd__nand2b_1
X_4781_ net1219 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3732_ net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 _0413_ _0405_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux4_2
X_3663_ net991 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 net1005 net1009 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ _0351_ sky130_fd_sc_hd__mux4_2
X_5402_ net1186 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkbuf_2
X_2614_ _1128_ _1129_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__xnor2_2
X_5333_ Tile_X0Y0_WW4END[8] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_4
X_3594_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0284_ VGND VGND
+ VPWR VPWR _0285_ sky130_fd_sc_hd__or2_1
X_2545_ _1398_ _1397_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__mux2_1
X_5264_ Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2476_ _1334_ _0157_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__or2_4
X_5195_ net50 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4215_ net203 net142 net82 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q VGND VGND VPWR VPWR
+ _0863_ sky130_fd_sc_hd__mux4_2
X_4146_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] net1059 VGND VGND VPWR VPWR _0798_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_87_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4077_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0734_ VGND VGND
+ VPWR VPWR _0735_ sky130_fd_sc_hd__nor2_1
X_3028_ net1264 net1019 net1226 net1038 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q VGND VGND VPWR VPWR
+ _1814_ sky130_fd_sc_hd__mux4_1
X_4979_ net1191 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_34_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput580 net580 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[7] sky130_fd_sc_hd__buf_2
Xfanout1205 net1206 VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__buf_4
Xfanout1238 net45 VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__buf_4
Xfanout1227 net56 VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__clkbuf_4
Xfanout1216 net149 VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__clkbuf_4
Xoutput591 net591 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[11] sky130_fd_sc_hd__buf_4
Xfanout1249 net38 VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__buf_4
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2330_ net1068 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] _1198_ _1197_ VGND VGND VPWR
+ VPWR _1199_ sky130_fd_sc_hd__o2bb2a_4
X_2261_ _1131_ _1118_ _1117_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__a21o_1
X_4000_ _0662_ _0661_ _0663_ _0106_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__a221o_1
X_2192_ _1033_ _1061_ _1060_ _1051_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__o211a_1
XFILLER_37_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ net153 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_23_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4833_ net1205 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4764_ net1198 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3715_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q _0398_ VGND VGND
+ VPWR VPWR _0399_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4695_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A3 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_106_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3646_ net992 net1022 net1002 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0335_ sky130_fd_sc_hd__mux4_1
X_3577_ _0046_ _0047_ _0033_ _0267_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q VGND VGND VPWR VPWR
+ _0268_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_93_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2528_ net222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q
+ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__o21a_1
X_5316_ net112 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_2
X_5247_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net339
+ sky130_fd_sc_hd__clkbuf_2
X_2459_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1319_ VGND VGND
+ VPWR VPWR _1320_ sky130_fd_sc_hd__nor2_1
X_5178_ Tile_X0Y0_EE4END[6] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_1
X_4129_ _0776_ _0781_ net1060 _0765_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_143_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1002 net1003 VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__buf_6
Xfanout1013 _1422_ VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__buf_8
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1035 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 VGND VGND VPWR VPWR
+ net1035 sky130_fd_sc_hd__clkbuf_2
Xfanout1046 net1049 VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__buf_8
Xfanout1024 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 VGND VGND VPWR VPWR net1024
+ sky130_fd_sc_hd__buf_2
Xfanout1057 net1058 VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__clkbuf_4
Xfanout1068 net1069 VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__buf_2
Xfanout1079 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3500_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q VGND VGND VPWR
+ VPWR _0195_ sky130_fd_sc_hd__inv_1
XFILLER_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4480_ net1227 net1104 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3431_ net135 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_1
X_3362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR
+ VPWR _0057_ sky130_fd_sc_hd__inv_1
X_2313_ net13 net105 net69 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q VGND VGND VPWR VPWR
+ _1183_ sky130_fd_sc_hd__mux4_2
X_5101_ net146 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _0599_ VGND VGND
+ VPWR VPWR _2025_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_29_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5032_ net1214 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2244_ _1107_ _1114_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__xor2_2
X_2175_ _0725_ _0612_ _0611_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_123_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4816_ net1188 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4747_ net1217 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4678_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0006_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3629_ net1019 net1035 net986 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0319_ sky130_fd_sc_hd__mux4_1
XFILLER_134_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput116 Tile_X0Y0_WW4END[1] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput105 Tile_X0Y0_W2MID[0] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput127 Tile_X0Y1_E2END[4] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_1
XFILLER_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput138 Tile_X0Y1_E2MID[7] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
XFILLER_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput149 Tile_X0Y1_FrameData[13] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
XFILLER_56_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3980_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q _0642_ _0644_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR VPWR
+ _0645_ sky130_fd_sc_hd__o211a_1
X_2931_ _1743_ _1744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 sky130_fd_sc_hd__mux2_4
XFILLER_50_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2862_ net1019 net1038 net1034 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR
+ _1686_ sky130_fd_sc_hd__mux4_1
X_4601_ net34 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2793_ _1604_ _1621_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__nor2_1
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4532_ net1247 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4463_ net1240 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3414_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q VGND VGND VPWR
+ VPWR _0109_ sky130_fd_sc_hd__inv_1
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4394_ net49 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ net186 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_1
X_3276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _2009_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q
+ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__a21oi_1
X_5015_ net145 net1085 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2227_ _1096_ _1092_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__xnor2_4
XFILLER_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2158_ Tile_X0Y1_DSP_bot.B0 net1061 _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ _0561_ _0562_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ _0556_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_140_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput409 net409 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_4_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3130_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q net992 VGND VGND
+ VPWR VPWR _1894_ sky130_fd_sc_hd__nor2_1
XFILLER_79_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3061_ net1049 _0756_ _0788_ _1610_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q VGND VGND VPWR VPWR
+ _1842_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3963_ net174 net180 net125 net1222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0630_ sky130_fd_sc_hd__mux4_1
X_2914_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q _1729_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__a21o_1
X_3894_ _0071_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q
+ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__a21oi_1
X_2845_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q _1668_ _1572_
+ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__and3_4
XFILLER_129_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2776_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q _1605_ VGND VGND
+ VPWR VPWR _1606_ sky130_fd_sc_hd__nand2_1
X_4515_ net53 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5495_ net228 VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_4
X_4446_ net29 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4377_ net1253 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3328_ net101 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_129_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ net1011 _1497_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer231 net849 VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__clkbuf_2
Xrebuffer220 net838 VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__clkbuf_2
Xrebuffer242 net860 VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__clkbuf_2
Xrebuffer264 net882 VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer297 net915 VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__clkbuf_1
Xrebuffer286 net904 VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer275 net893 VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2630_ _1479_ _1468_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C2 sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_117_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2561_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q _1413_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__o21ai_1
X_5280_ Tile_X0Y1_NN4END[8] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_1
X_4300_ net46 net1149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput239 net239 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2492_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1347_ _1349_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR VPWR
+ _1350_ sky130_fd_sc_hd__o211a_1
XFILLER_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4231_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] net1061 VGND VGND VPWR VPWR _0877_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4162_ _0576_ _0762_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__or3_1
XFILLER_67_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4093_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q _0749_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__o21a_1
X_3113_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q net661 _1881_
+ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__a21o_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3044_ _1825_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_66_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4995_ net157 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3946_ _0611_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nand2_1
XFILLER_23_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3877_ _0547_ _0546_ _0548_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR VPWR
+ _0549_ sky130_fd_sc_hd__a221o_1
X_2828_ _1604_ _1652_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__nor2_1
X_2759_ net99 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q
+ _1590_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__o211a_1
XFILLER_155_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5478_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net570
+ sky130_fd_sc_hd__buf_4
XFILLER_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4429_ net1238 net1113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q _0470_ _0472_
+ _0476_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ sky130_fd_sc_hd__a31o_4
X_4780_ net1218 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3731_ net191 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net227
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_71_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3662_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q _0349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o21ba_1
X_3593_ net58 net66 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q VGND
+ VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
X_2613_ net1066 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] _1462_ _1461_ VGND VGND VPWR
+ VPWR _1463_ sky130_fd_sc_hd__a22oi_4
X_5401_ net172 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_1
X_5332_ Tile_X0Y0_WW4END[7] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_4
X_2544_ net203 net128 net74 net219 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q VGND VGND VPWR VPWR
+ _1398_ sky130_fd_sc_hd__mux4_2
XFILLER_114_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2475_ net656 net1005 net995 net653 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q VGND VGND VPWR VPWR
+ _1334_ sky130_fd_sc_hd__mux4_2
X_5263_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net355
+ sky130_fd_sc_hd__buf_2
X_5194_ net47 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_10_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4214_ _0857_ _0859_ _0862_ _0140_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ sky130_fd_sc_hd__a22o_4
X_4145_ _0790_ _0797_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X
+ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_79_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4076_ _0279_ net191 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__mux2_1
X_3027_ _1805_ _1808_ _1813_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 sky130_fd_sc_hd__a22o_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4978_ net1190 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_34_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3929_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q _0597_ VGND VGND
+ VPWR VPWR _0598_ sky130_fd_sc_hd__nor2_1
XFILLER_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput581 net581 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput570 net570 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[1] sky130_fd_sc_hd__buf_8
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_148_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1228 net55 VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout1217 net148 VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__buf_4
Xoutput592 net592 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[1] sky130_fd_sc_hd__buf_2
Xfanout1206 Tile_X0Y1_FrameData[22] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1239 net44 VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__buf_4
XFILLER_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2260_ _1119_ _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__nor2_4
X_2191_ _1051_ _1060_ _1033_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__a211oi_4
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4901_ net1211 net1110 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_190 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4832_ net1203 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4763_ net1197 net1144 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3714_ net973 net977 net997 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0398_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_31_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4694_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3645_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q _0333_ VGND VGND
+ VPWR VPWR _0334_ sky130_fd_sc_hd__and2b_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3576_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR _0267_
+ sky130_fd_sc_hd__inv_4
X_5315_ net111 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_1
X_2527_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q _1353_ VGND VGND
+ VPWR VPWR _1382_ sky130_fd_sc_hd__nand2_2
X_2458_ net176 net1224 net184 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _1319_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2389_ _1253_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] net1069 VGND VGND VPWR VPWR
+ _1254_ sky130_fd_sc_hd__mux2_4
X_5177_ Tile_X0Y0_EE4END[5] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_1
X_4128_ _0776_ _0781_ _0765_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X
+ sky130_fd_sc_hd__a21o_1
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4059_ _0717_ _0718_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q
+ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux2_1
XFILLER_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1003 net1006 VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__buf_6
Xfanout1036 net1039 VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__buf_2
Xfanout1014 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 VGND VGND VPWR VPWR
+ net1014 sky130_fd_sc_hd__buf_8
Xfanout1047 net1049 VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__buf_2
Xfanout1025 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 VGND VGND VPWR VPWR net1025
+ sky130_fd_sc_hd__buf_2
Xfanout1058 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 VGND VGND VPWR VPWR
+ net1058 sky130_fd_sc_hd__buf_8
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1069 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q VGND VGND
+ VPWR VPWR net1069 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3430_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q VGND VGND VPWR
+ VPWR _0125_ sky130_fd_sc_hd__inv_1
X_3361_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR
+ VPWR _0056_ sky130_fd_sc_hd__inv_2
X_2312_ _1182_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__inv_2
XFILLER_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5100_ net147 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3292_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q _2020_ _2023_
+ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__a21o_1
X_5031_ net1213 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2243_ _1109_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__nor2_1
X_2174_ _0478_ _0848_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4815_ net1187 net1134 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4746_ net149 net1180 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4677_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0005_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3628_ _0316_ _0315_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ _0300_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o211ai_4
X_3559_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q _0251_ VGND VGND
+ VPWR VPWR _0252_ sky130_fd_sc_hd__or2_4
Xinput117 Tile_X0Y0_WW4END[2] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
Xinput106 Tile_X0Y0_W2MID[1] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5229_ net1115 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_2
Xinput128 Tile_X0Y1_E2END[5] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_2
Xinput139 Tile_X0Y1_E6END[0] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
XFILLER_44_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_90 Tile_X0Y1_E6END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2930_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 _0317_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__mux2_1
XFILLER_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2861_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q _1675_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q
+ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__o21ai_1
X_4600_ net1252 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2792_ net1069 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\] _1620_ VGND VGND VPWR VPWR
+ _1621_ sky130_fd_sc_hd__a21oi_1
X_4531_ net1246 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4462_ net1239 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3413_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q VGND VGND VPWR
+ VPWR _0108_ sky130_fd_sc_hd__inv_2
X_4393_ net1260 net1129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_90_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q VGND VGND VPWR
+ VPWR _0039_ sky130_fd_sc_hd__inv_2
X_3275_ _2008_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__inv_1
XFILLER_97_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5014_ net156 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2226_ _1092_ _1096_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__and2_1
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2157_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] net1061 VGND VGND VPWR VPWR _1028_
+ sky130_fd_sc_hd__nand2b_1
X_2088_ _0360_ _0361_ _0142_ _0386_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_140_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4729_ net1194 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3060_ _1838_ _1840_ _1841_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 sky130_fd_sc_hd__o22a_1
XFILLER_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3962_ _0123_ _0628_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q
+ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__o21a_1
X_2913_ net59 net67 net93 net1226 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1729_ sky130_fd_sc_hd__mux4_1
X_3893_ _0562_ _0561_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ _0556_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__a211o_1
XFILLER_148_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2844_ _1667_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] net1068 VGND VGND VPWR VPWR
+ _1668_ sky130_fd_sc_hd__mux2_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2775_ net118 net654 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__mux2_1
X_4514_ net1229 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5494_ net227 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_2
X_4445_ net1257 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4376_ net35 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3327_ net190 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_1
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3258_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q _1993_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q
+ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_69_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _1071_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_1_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3189_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q _1934_ VGND
+ VGND VPWR VPWR _1935_ sky130_fd_sc_hd__and2b_1
XFILLER_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer210 _0219_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer221 net839 VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__clkbuf_2
Xrebuffer232 net850 VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer243 net861 VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__clkbuf_2
Xrebuffer265 net883 VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer298 _0340_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__clkbuf_1
Xrebuffer287 net905 VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer276 net894 VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_9_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2560_ _1412_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__inv_2
X_2491_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q _1348_ VGND VGND
+ VPWR VPWR _1349_ sky130_fd_sc_hd__nand2_1
XFILLER_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4230_ _0875_ _0876_ _0864_ _0863_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.B2 sky130_fd_sc_hd__mux4_2
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4161_ _0801_ _0810_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a21o_1
X_4092_ net975 net869 net999 net988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0749_ sky130_fd_sc_hd__mux4_1
X_3112_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q VGND VGND VPWR VPWR
+ _1881_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3043_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q _0571_ _1826_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q VGND VGND VPWR VPWR
+ _1827_ sky130_fd_sc_hd__a211oi_1
XFILLER_82_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ net158 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3945_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] net1061 VGND VGND VPWR VPWR _0612_
+ sky130_fd_sc_hd__nand2b_2
XFILLER_23_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3876_ net199 net24 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q VGND
+ VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux2_1
X_2827_ _1604_ _1652_ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__nand2_4
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2758_ _0744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q VGND VGND
+ VPWR VPWR _1590_ sky130_fd_sc_hd__nand2_2
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5477_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net569
+ sky130_fd_sc_hd__buf_1
XFILLER_132_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2689_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q _1535_ VGND VGND
+ VPWR VPWR _1536_ sky130_fd_sc_hd__or2_1
X_4428_ net1237 net1113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_92_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4359_ net1236 net1138 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout990 net991 VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3730_ _0057_ _0408_ _0410_ _0412_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_71_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ net176 net1224 net184 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _0349_ sky130_fd_sc_hd__mux4_1
X_3592_ _0280_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q _0282_
+ _0097_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__o211a_1
X_5400_ net171 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkbuf_2
X_2612_ net1063 _0168_ net1066 VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__a21oi_1
X_5331_ Tile_X0Y0_WW4END[6] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__buf_4
X_2543_ net1221 net82 net235 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__mux4_1
XFILLER_114_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5262_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net354
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2474_ _1332_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q VGND VGND
+ VPWR VPWR _1333_ sky130_fd_sc_hd__or2_4
X_5193_ net38 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_1
X_4213_ _0860_ _0861_ _0139_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__mux2_1
X_4144_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q _0796_ _0795_
+ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_79_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4075_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0732_ VGND VGND
+ VPWR VPWR _0733_ sky130_fd_sc_hd__nand2_1
X_3026_ _1812_ _1811_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__mux2_2
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4977_ net1189 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_98_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3928_ net207 net1263 net6 net1261 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0597_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_34_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3859_ _0530_ _0531_ _0060_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_4
XFILLER_152_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput571 net571 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput560 net560 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[1] sky130_fd_sc_hd__buf_2
Xfanout1229 net54 VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__clkbuf_4
Xfanout1207 net158 VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__buf_4
Xoutput582 net582 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput593 net593 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[2] sky130_fd_sc_hd__buf_2
Xfanout1218 net147 VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2190_ _1010_ _1011_ _1032_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_76_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4900_ net1210 net1110 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4831_ net1201 net1126 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_180 net609 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4762_ net1196 net1144 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3713_ _0396_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__a21bo_1
X_4693_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A1 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3644_ net909 net970 net977 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0333_ sky130_fd_sc_hd__mux4_2
XFILLER_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3575_ _0261_ _0263_ _0266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 sky130_fd_sc_hd__o22a_4
XTAP_TAPCELL_ROW_132_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5314_ net110 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_2
X_2526_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1380_ _1379_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR VPWR
+ _1381_ sky130_fd_sc_hd__o211a_1
X_2457_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1315_ _1317_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR VPWR
+ _1318_ sky130_fd_sc_hd__o211a_1
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2388_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\] net1065 VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__mux2_4
X_5176_ Tile_X0Y0_EE4END[4] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
X_4127_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q _0780_ VGND VGND
+ VPWR VPWR _0781_ sky130_fd_sc_hd__nor2_1
X_4058_ net83 net91 net216 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0718_ sky130_fd_sc_hd__mux4_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3009_ net1015 net968 _1204_ _0471_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1798_ sky130_fd_sc_hd__mux4_1
XFILLER_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1004 net1006 VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__buf_2
Xfanout1015 net1016 VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1037 net1039 VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__buf_8
Xfanout1026 net1027 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__buf_8
Xoutput390 net390 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[1] sky130_fd_sc_hd__buf_2
Xfanout1048 net1049 VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__buf_2
Xfanout1059 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q VGND VGND
+ VPWR VPWR net1059 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_73_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3360_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q VGND VGND VPWR
+ VPWR _0055_ sky130_fd_sc_hd__inv_2
XFILLER_124_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2311_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q _1175_ _1177_
+ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a31o_1
XFILLER_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3291_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _0196_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2
+ _2022_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__a31o_1
XFILLER_2_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5030_ net1212 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2242_ _1092_ _1110_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a21o_1
X_2173_ _0878_ _0640_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_36_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4814_ net1186 net1134 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4745_ net1215 net1180 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4676_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0004_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3627_ _0315_ _0316_ _0300_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o21ai_4
X_3558_ net1017 net1037 net1031 net982 net617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux4_2
X_2509_ net177 net185 net1223 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ _1366_ sky130_fd_sc_hd__mux4_1
Xinput118 Tile_X0Y0_WW4END[3] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xinput107 Tile_X0Y0_W2MID[2] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
X_3489_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR
+ VPWR _0184_ sky130_fd_sc_hd__inv_1
X_5228_ net1122 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_2
Xinput129 Tile_X0Y1_E2END[6] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_2
X_5159_ net16 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_80 net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 Tile_X0Y1_E6END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2860_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _1182_ _1679_
+ _1683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR
+ VPWR _1684_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_41_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ net1068 _1619_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__and2b_1
XFILLER_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4530_ net1245 net1089 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4461_ net1238 net1105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3412_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q VGND VGND VPWR
+ VPWR _0107_ sky130_fd_sc_hd__inv_1
X_4392_ net1249 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q VGND VGND VPWR
+ VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3274_ net978 net990 net998 net864 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q VGND VGND VPWR VPWR
+ _2008_ sky130_fd_sc_hd__mux4_1
X_2225_ _1095_ _1094_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__xnor2_4
X_5013_ net164 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2156_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q _1018_ _1020_
+ _1024_ _1027_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B0 sky130_fd_sc_hd__a32o_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ _0960_ _0228_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q
+ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2989_ _0173_ _1781_ _1780_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2
+ sky130_fd_sc_hd__o21a_1
X_4728_ net1193 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4659_ net1246 net1157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3961_ net992 net1021 net1002 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0628_ sky130_fd_sc_hd__mux4_1
X_2912_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q _1727_ VGND VGND
+ VPWR VPWR _1728_ sky130_fd_sc_hd__and2b_1
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3892_ _0561_ _0562_ _0556_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__a21o_4
X_2843_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\] net1064 VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__mux2_4
X_2774_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q _1572_ VGND VGND
+ VPWR VPWR _1604_ sky130_fd_sc_hd__nand2_2
X_4513_ net55 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_130_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5493_ net226 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__buf_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4444_ net1256 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4375_ net1251 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3326_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q VGND VGND VPWR
+ VPWR _0021_ sky130_fd_sc_hd__inv_2
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3257_ net210 net989 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _1077_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_1_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ net174 net119 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__mux2_1
X_2139_ _0990_ _1009_ _1008_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a21o_1
XFILLER_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer200 net919 VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__buf_8
Xrebuffer222 net840 VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__clkbuf_2
Xrebuffer244 net862 VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__clkbuf_2
Xrebuffer233 net851 VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer288 net906 VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer266 net884 VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer277 net895 VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2490_ net76 net1072 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__mux2_1
XFILLER_141_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4160_ _0667_ _0784_ _0799_ _0710_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__o22a_1
X_3111_ net1000 _0214_ net619 _0228_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4091_ _0099_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__or2_1
X_3042_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q net1027 VGND
+ VGND VPWR VPWR _1826_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4993_ net1205 net1085 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3944_ _0603_ _0602_ _0610_ net1061 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a211o_4
X_3875_ _0026_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q
+ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__a21oi_1
X_2826_ _1651_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__inv_4
X_2757_ net641 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q VGND VGND
+ VPWR VPWR _1589_ sky130_fd_sc_hd__nand2b_1
X_2688_ net191 net86 net10 net102 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q VGND VGND VPWR VPWR
+ _1535_ sky130_fd_sc_hd__mux4_2
XFILLER_144_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4427_ net1235 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_96_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ net1233 net1138 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4289_ net1228 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3309_ net966 _1558_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__and2b_1
XFILLER_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout991 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VGND VGND VPWR VPWR net991
+ sky130_fd_sc_hd__clkbuf_2
Xfanout980 net981 VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3660_ _0346_ _0345_ _0347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ _0069_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a221o_1
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3591_ _0096_ _0281_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__or2_1
X_2611_ Tile_X0Y1_DSP_bot.C3 net1063 VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__or2_4
X_5330_ Tile_X0Y0_WW4END[5] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_4
X_2542_ _1394_ _1393_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__xor2_2
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5261_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net353
+ sky130_fd_sc_hd__buf_4
X_2473_ net655 net971 net980 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1332_ sky130_fd_sc_hd__mux4_2
X_4212_ net205 net120 net126 net1221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0861_ sky130_fd_sc_hd__mux4_1
XFILLER_141_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5192_ net1260 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_4
X_4143_ net206 net63 net7 net99 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q VGND VGND VPWR VPWR
+ _0796_ sky130_fd_sc_hd__mux4_2
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4074_ net1053 net1048 net1028 net1014 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0732_ sky130_fd_sc_hd__mux4_1
X_3025_ net1047 net1030 net1015 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1812_ sky130_fd_sc_hd__mux4_1
XFILLER_36_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4976_ net1188 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3927_ _0085_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3858_ net1017 net823 net1031 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0531_ sky130_fd_sc_hd__mux4_1
X_2809_ _0119_ _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__or2_1
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3789_ _0461_ _0463_ _0466_ _0084_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput572 net572 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput550 net550 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput561 net561 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[2] sky130_fd_sc_hd__buf_2
X_5459_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net542
+ sky130_fd_sc_hd__buf_1
Xfanout1208 net157 VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__buf_4
Xoutput583 net583 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput594 net594 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[3] sky130_fd_sc_hd__buf_2
Xfanout1219 net146 VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_170 net583 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ net159 net1126 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_192 _0414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_181 net610 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ net1194 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3712_ net1042 net1028 net1053 net822 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR VPWR
+ _0396_ sky130_fd_sc_hd__mux4_2
X_4692_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.A0 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3643_ _0331_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__inv_2
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5313_ net109 VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_2
X_3574_ _0264_ _0265_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
X_2525_ net179 net144 net70 net215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q VGND VGND VPWR VPWR
+ _1380_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_132_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5244_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net336
+ sky130_fd_sc_hd__clkbuf_2
X_2456_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q _1316_ VGND VGND
+ VPWR VPWR _1317_ sky130_fd_sc_hd__nand2_1
X_5175_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 VGND VGND VPWR VPWR net258
+ sky130_fd_sc_hd__buf_6
X_2387_ _1237_ _1239_ _1252_ _1251_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ sky130_fd_sc_hd__a22o_1
X_4126_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q _0777_ _0779_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q VGND VGND VPWR VPWR
+ _0780_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_39_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4057_ net204 net143 net119 net1222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q VGND VGND VPWR VPWR
+ _0717_ sky130_fd_sc_hd__mux4_1
XFILLER_71_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3008_ _1794_ _1795_ _1796_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q VGND VGND VPWR VPWR
+ _1797_ sky130_fd_sc_hd__a221o_1
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4959_ net1201 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput380 net380 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_105_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1016 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 VGND VGND VPWR VPWR
+ net1016 sky130_fd_sc_hd__clkbuf_4
Xfanout1027 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 VGND VGND VPWR VPWR
+ net1027 sky130_fd_sc_hd__buf_12
Xfanout1038 net1039 VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__clkbuf_4
Xoutput391 net391 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[2] sky130_fd_sc_hd__buf_6
Xfanout1005 net1006 VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__clkbuf_4
Xfanout1049 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 VGND VGND VPWR VPWR
+ net1049 sky130_fd_sc_hd__buf_8
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _1180_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q VGND VGND
+ VPWR VPWR _1181_ sky130_fd_sc_hd__nor2_1
X_3290_ net222 _2021_ _0197_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__a21o_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2241_ _0726_ _0981_ net832 _0640_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__o22a_1
X_2172_ _1007_ _1003_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__xor2_2
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4813_ net1219 net1134 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4744_ net151 net1180 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4675_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0003_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3626_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q net97 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q
+ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3557_ net867 net1045 net1050 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ net617 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux4_1
X_2508_ _1362_ _1363_ _1364_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ _0160_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__a221o_1
X_5227_ net1131 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput108 Tile_X0Y0_W2MID[3] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
X_3488_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR
+ VPWR _0183_ sky130_fd_sc_hd__inv_2
Xinput119 Tile_X0Y1_E1END[0] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
X_2439_ net974 net972 net978 net831 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR
+ _1301_ sky130_fd_sc_hd__mux4_1
X_5158_ net15 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4109_ net192 net11 net88 net103 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q VGND VGND VPWR VPWR
+ _0764_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_16_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5089_ net1205 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 net436 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_81 net444 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 Tile_X0Y1_EE4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\] net1065 VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__mux2_1
XFILLER_62_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4460_ net1237 net1105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3411_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q VGND VGND VPWR
+ VPWR _0106_ sky130_fd_sc_hd__inv_1
X_4391_ net1236 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3342_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR
+ VPWR _0037_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_90_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3273_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q _2006_ VGND VGND
+ VPWR VPWR _2007_ sky130_fd_sc_hd__or2_1
X_2224_ _0784_ net832 VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_8
X_5012_ net1192 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2155_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q _1026_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q
+ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a21oi_2
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone194 net926 VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__buf_6
X_2086_ net180 net125 net71 net234 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q VGND VGND VPWR VPWR
+ _0960_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_140_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2988_ net1015 net641 _1204_ _0759_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q VGND VGND VPWR VPWR
+ _1781_ sky130_fd_sc_hd__mux4_1
X_4727_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\] sky130_fd_sc_hd__dfxtp_1
X_4658_ net1245 net1157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput90 Tile_X0Y0_SS4END[5] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3609_ net206 net1262 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q
+ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
X_4589_ net1238 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3960_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q _0626_ VGND VGND
+ VPWR VPWR _0627_ sky130_fd_sc_hd__or2_4
X_2911_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net3 net192 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _1727_ sky130_fd_sc_hd__mux4_2
XFILLER_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3891_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q net1052 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__o21ba_1
X_2842_ _1666_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ sky130_fd_sc_hd__inv_2
XFILLER_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2773_ _1603_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 sky130_fd_sc_hd__mux2_4
X_4512_ net56 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5492_ net225 VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__buf_4
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4443_ net1255 net1113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4374_ net1250 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3325_ net1222 VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
X_3256_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q _1991_ VGND VGND
+ VPWR VPWR _1992_ sky130_fd_sc_hd__and2b_1
X_2207_ _0799_ net832 VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3187_ _0442_ net991 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__mux2_1
X_2138_ _0990_ _1008_ _1009_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_1_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2069_ _0937_ _0942_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nor2_4
XFILLER_14_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer201 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR
+ net818 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer223 net841 VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__clkbuf_2
Xrebuffer212 _1125_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__buf_8
Xrebuffer245 net863 VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__clkbuf_2
Xrebuffer234 net852 VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__clkbuf_2
Xrebuffer267 net885 VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer278 net896 VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer289 net907 VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_118_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ net179 net194 net230 net1004 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A sky130_fd_sc_hd__mux4_1
X_4090_ net993 net1022 net1003 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0747_ sky130_fd_sc_hd__mux4_1
XFILLER_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3041_ _0700_ _1195_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_128_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4992_ net1203 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3943_ _0602_ _0603_ _0610_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B3 sky130_fd_sc_hd__a21o_1
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3874_ net813 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q VGND VGND
+ VPWR VPWR _0546_ sky130_fd_sc_hd__or2_4
X_2825_ _1650_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] net1068 VGND VGND VPWR VPWR
+ _1651_ sky130_fd_sc_hd__mux2_4
XFILLER_129_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2756_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q _1585_ _1587_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q VGND VGND VPWR VPWR
+ _1588_ sky130_fd_sc_hd__a211o_1
XFILLER_117_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2687_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q _0554_ VGND VGND
+ VPWR VPWR _1534_ sky130_fd_sc_hd__nand2_1
X_5475_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net558
+ sky130_fd_sc_hd__buf_1
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4426_ net1234 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_96_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4357_ net1232 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4288_ net1227 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3308_ net966 _1560_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and2b_1
XFILLER_100_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3239_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q _1975_ _1977_
+ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__a21bo_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout970 net972 VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__buf_8
Xfanout992 net993 VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__buf_6
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout981 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 VGND VGND VPWR VPWR net981
+ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_28_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3590_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q VGND
+ VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
X_2610_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q _1453_ _1455_
+ _1460_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C3 sky130_fd_sc_hd__a31o_4
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2541_ _1376_ _1392_ _1394_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5260_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net352
+ sky130_fd_sc_hd__buf_6
X_2472_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4
+ _0156_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__o211a_1
XFILLER_141_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4211_ net72 net217 net84 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR
+ _0860_ sky130_fd_sc_hd__mux4_1
X_5191_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR net274
+ sky130_fd_sc_hd__buf_6
X_4142_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q _0791_ _0794_
+ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21o_1
X_4073_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q _0730_ VGND VGND
+ VPWR VPWR _0731_ sky130_fd_sc_hd__nand2b_4
XFILLER_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3024_ _1810_ _1809_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q
+ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_87_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4975_ net172 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3926_ net62 net78 net98 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0595_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_34_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3857_ net1050 net1045 net1026 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0530_ sky130_fd_sc_hd__mux4_2
X_2808_ net1263 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__mux2_1
XFILLER_137_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3788_ _0464_ _0465_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q
+ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
X_2739_ _1167_ _1571_ _1170_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__or3b_4
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput551 net551 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput540 net540 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput562 net562 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[3] sky130_fd_sc_hd__buf_2
X_5458_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net541
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4409_ net1253 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput584 net584 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput573 net573 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput595 net595 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[4] sky130_fd_sc_hd__buf_2
X_5389_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net472
+ sky130_fd_sc_hd__clkbuf_1
Xfanout1209 net156 VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_160 net552 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_182 net613 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 net584 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 _0599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4760_ net1193 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4691_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0019_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_3711_ _0113_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3642_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q VGND VGND VPWR VPWR
+ _0331_ sky130_fd_sc_hd__o21ai_2
X_5312_ net108 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3573_ net73 net81 net218 net234 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0265_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_93_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2524_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q _1377_ VGND VGND
+ VPWR VPWR _1379_ sky130_fd_sc_hd__nand2_1
X_5243_ Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_1
X_2455_ net210 net1073 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__mux2_1
X_5174_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net257
+ sky130_fd_sc_hd__buf_6
X_2386_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _0560_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4125_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q _0778_ VGND VGND
+ VPWR VPWR _0779_ sky130_fd_sc_hd__nand2_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4056_ _0128_ _0715_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3007_ net57 net1043 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__mux2_1
XFILLER_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4958_ net159 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4889_ net1194 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3909_ _0360_ _0361_ _0386_ _0131_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a211o_1
XFILLER_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput370 net370 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput381 net381 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[3] sky130_fd_sc_hd__buf_2
Xfanout1028 net1030 VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__buf_2
Xoutput392 net392 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_10_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1006 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 VGND VGND VPWR VPWR net1006
+ sky130_fd_sc_hd__buf_8
Xfanout1017 net1018 VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__buf_8
Xfanout1039 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 VGND VGND VPWR VPWR
+ net1039 sky130_fd_sc_hd__buf_12
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_98_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2240_ _1092_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2171_ _1037_ _1038_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__xor2_1
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4812_ net1218 net1134 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4743_ net152 net1181 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4674_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0002_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3625_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q _0313_ _0308_
+ _0304_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR
+ VPWR _0315_ sky130_fd_sc_hd__o311a_4
X_3556_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q _0248_ VGND VGND
+ VPWR VPWR _0249_ sky130_fd_sc_hd__nor2_1
XFILLER_130_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2507_ net211 net1072 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__mux2_1
XFILLER_142_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3487_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q VGND VGND VPWR
+ VPWR _0182_ sky130_fd_sc_hd__inv_1
XFILLER_102_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput109 Tile_X0Y0_W2MID[4] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlymetal6s2s_1
X_5226_ net1141 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__buf_4
X_2438_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q _0453_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__a21oi_1
X_2369_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q _1235_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__o21ai_1
X_5157_ net14 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
X_4108_ _0384_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q VGND VGND
+ VPWR VPWR _0763_ sky130_fd_sc_hd__nand2_2
X_5088_ net1203 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4039_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q _0697_ _0699_
+ _0698_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a22o_4
XFILLER_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_71 Tile_X0Y0_WW4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 net401 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 Tile_X0Y1_EE4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 Tile_X0Y1_E6END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3410_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR
+ VPWR _0105_ sky130_fd_sc_hd__inv_2
X_4390_ net1233 net1129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3341_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR
+ VPWR _0036_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_90_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ net1223 net1072 net974 net969 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _2006_ sky130_fd_sc_hd__mux4_1
X_2223_ _0878_ _0928_ _1047_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__or3b_4
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5011_ net168 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_78_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2154_ _1025_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__inv_2
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2085_ _0940_ _0956_ _0957_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__a22o_1
Xclone195 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 VGND VGND VPWR VPWR net812
+ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_140_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2987_ _1777_ _1778_ _1779_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q VGND VGND VPWR VPWR
+ _1780_ sky130_fd_sc_hd__a221o_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4726_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4657_ net1243 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput91 Tile_X0Y0_SS4END[6] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xinput80 Tile_X0Y0_S4END[3] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_151_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3608_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q _0295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o211a_1
X_4588_ net1237 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3539_ net992 net1022 net1002 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0232_ sky130_fd_sc_hd__mux4_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5209_ net1252 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2910_ _1724_ _1725_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__mux2_1
XFILLER_43_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3890_ _0558_ _0557_ _0559_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ _0088_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a221o_2
X_2841_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q _1661_ _1659_
+ _1663_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__o32a_4
X_2772_ _1602_ _1570_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__xnor2_2
XFILLER_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4511_ net1259 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5491_ net224 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkbuf_2
X_4442_ net1254 net1113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4373_ net1248 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3324_ net967 _1718_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__and2b_1
XFILLER_112_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3255_ net174 _0442_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__mux2_1
X_2206_ _1045_ _1072_ _1074_ _1075_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a22o_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3186_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q _1928_ _1932_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o21a_1
X_2137_ _0987_ _0988_ _0989_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__a21o_1
XFILLER_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2068_ _0941_ _0938_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__xnor2_4
XFILLER_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer202 _0237_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__buf_6
X_4709_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs net676 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xrebuffer224 net842 VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__clkbuf_2
Xrebuffer246 _0243_ VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__clkbuf_2
Xrebuffer235 net853 VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__clkbuf_2
Xrebuffer257 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR
+ net874 sky130_fd_sc_hd__buf_6
Xrebuffer279 net897 VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer268 net886 VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_Tile_X0Y1_UserCLK_regs Tile_X0Y1_UserCLK_regs VGND VGND VPWR VPWR clknet_0_Tile_X0Y1_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3040_ _1824_ _1823_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4991_ net1201 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3942_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0609_ _0608_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR VPWR
+ _0610_ sky130_fd_sc_hd__o211a_1
X_3873_ _0542_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q _0544_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR VPWR
+ _0545_ sky130_fd_sc_hd__o211a_1
X_2824_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\] net1064 VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__mux2_4
X_2755_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q _1586_ VGND VGND
+ VPWR VPWR _1587_ sky130_fd_sc_hd__and2b_1
X_2686_ _1532_ _1231_ _1230_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__a21o_1
X_5474_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net557
+ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_52_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4425_ net1260 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_96_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4356_ net1231 net1138 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3307_ net928 _1555_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__and2b_1
X_4287_ net1259 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3238_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q net633 _1976_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q VGND VGND VPWR VPWR
+ _1977_ sky130_fd_sc_hd__a211o_1
XFILLER_100_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3169_ _1918_ _1917_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_61_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_70_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout982 net986 VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__buf_8
Xfanout993 net996 VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__buf_6
Xfanout971 net972 VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__clkbuf_4
XFILLER_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 _1398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2540_ _1135_ _1133_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__xnor2_4
XFILLER_126_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2471_ _0588_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q VGND VGND
+ VPWR VPWR _1330_ sky130_fd_sc_hd__nand2_2
XFILLER_141_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4210_ _0139_ _0858_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q
+ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__o21a_1
X_5190_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net273
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_118_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4141_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q _0793_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__o21ai_1
X_4072_ net815 net1036 net1032 net983 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0730_ sky130_fd_sc_hd__mux4_2
XFILLER_95_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3023_ _0788_ _0756_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4974_ net173 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_127_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3925_ _0085_ _0593_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_34_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3856_ _0527_ _0524_ _0528_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q VGND VGND VPWR VPWR
+ _0529_ sky130_fd_sc_hd__o221a_4
X_2807_ _0414_ net193 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__mux2_1
X_3787_ net1261 net64 net100 net116 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0465_ sky130_fd_sc_hd__mux4_1
X_2738_ _0893_ _1154_ _1150_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__a21oi_1
X_5457_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net540
+ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_136_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4408_ net35 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput530 net530 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput552 net552 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput541 net541 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput563 net563 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[4] sky130_fd_sc_hd__buf_2
X_2669_ _1516_ _1515_ _1511_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C0 sky130_fd_sc_hd__a21o_1
Xoutput585 net585 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput574 net574 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput596 net596 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[5] sky130_fd_sc_hd__buf_2
X_5388_ Tile_X0Y1_EE4END[15] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_1
X_4339_ net1246 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_74_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_150 Tile_X0Y1_NN4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_161 net553 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 net615 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 net590 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _0599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3710_ net815 net1036 net1032 net985 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR
+ _0394_ sky130_fd_sc_hd__mux4_1
X_4690_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0018_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_3641_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q _0330_ _0326_
+ _0320_ _0322_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__o32a_4
X_3572_ net182 net127 net1224 net1222 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0264_ sky130_fd_sc_hd__mux4_1
X_5311_ net107 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_2
X_2523_ _1377_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__inv_4
XFILLER_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5242_ Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
X_2454_ _0343_ _0068_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__mux2_4
X_5173_ Tile_X0Y0_E6END[11] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
X_2385_ _0109_ _1240_ _1250_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__a211o_1
XFILLER_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4124_ net76 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q VGND
+ VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux2_1
Xinput1 Tile_X0Y0_E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XFILLER_110_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4055_ net992 net1021 net1002 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0715_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_39_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3006_ _0027_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4957_ net1199 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4888_ net1193 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3908_ _0561_ _0562_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ _0556_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__a211o_1
X_3839_ net77 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_144_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5509_ Tile_X0Y1_WW4END[4] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__buf_4
Xoutput360 net360 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput371 net371 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_10_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput382 net382 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[4] sky130_fd_sc_hd__buf_2
Xfanout1018 net1020 VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__buf_8
Xfanout1029 net1030 VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__buf_1
Xoutput393 net393 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1007 net1009 VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_153_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2170_ _1001_ _1039_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__xnor2_4
Xclone311 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr VGND VGND VPWR VPWR net928
+ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4811_ net1217 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4742_ net1212 net1181 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4673_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0001_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3624_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q _0308_ _0313_
+ _0304_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__o31a_4
XFILLER_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3555_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0245_ _0247_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR
+ _0248_ sky130_fd_sc_hd__o211a_1
X_3486_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q VGND VGND VPWR
+ VPWR _0181_ sky130_fd_sc_hd__inv_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2506_ _0053_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__a21oi_1
X_5225_ net1149 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_1
XFILLER_88_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2437_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__or2_1
XFILLER_102_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2368_ _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__inv_2
X_5156_ net13 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_1
XFILLER_96_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2299_ _1162_ _1161_ _1168_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__o21ai_4
X_4107_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ net1061 _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__o21ai_4
X_5087_ net1201 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4038_ _0092_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a21oi_1
XFILLER_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_50 Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 Tile_X0Y0_WW4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net404 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 Tile_X0Y1_E6END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_94 Tile_X0Y1_EE4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3340_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q VGND VGND VPWR
+ VPWR _0035_ sky130_fd_sc_hd__inv_1
XFILLER_97_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _2004_ _2003_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q
+ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__mux2_1
X_5010_ net169 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2222_ _0878_ _0928_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__nor2_4
XFILLER_38_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ net193 net138 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 net229
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q
+ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__mux4_2
XFILLER_78_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone196 net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 net816 net814
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__mux4_2
X_2084_ _0940_ _0956_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__xor2_2
XFILLER_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2986_ net93 net1043 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__mux2_1
X_4725_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\] sky130_fd_sc_hd__dfxtp_1
X_4656_ net1241 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput81 Tile_X0Y0_S4END[4] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
Xinput70 Tile_X0Y0_S2MID[1] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_151_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3607_ _0087_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__or2_4
X_4587_ net1235 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput92 Tile_X0Y0_SS4END[7] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
X_3538_ _0230_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q VGND VGND
+ VPWR VPWR _0231_ sky130_fd_sc_hd__or2_4
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3469_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR
+ VPWR _0164_ sky130_fd_sc_hd__inv_1
X_5208_ net34 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_1
X_5139_ net168 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2840_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q _1664_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__o21ai_1
X_2771_ _1600_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__and2_1
X_4510_ net1258 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5490_ net223 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkbuf_2
X_4441_ net1253 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4372_ net1247 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3323_ net967 _1721_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3254_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q _1986_ _1990_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 sky130_fd_sc_hd__o21a_1
XFILLER_58_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2205_ _1045_ _1072_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__a21boi_2
X_3185_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q _1929_ _1930_
+ _1931_ _0189_ VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__a221o_1
Xfanout1190 net169 VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__buf_4
X_2136_ _1003_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2067_ _0939_ _0881_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__xnor2_4
XFILLER_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer203 _0254_ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__clkbuf_2
X_2969_ _1766_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__inv_1
X_4708_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C0 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer236 net854 VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__clkbuf_2
Xrebuffer225 net843 VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__clkbuf_2
Xrebuffer258 net874 VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__clkbuf_2
Xrebuffer269 net887 VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4639_ net1259 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4990_ net1200 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3941_ net178 net69 net142 net214 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q VGND VGND VPWR VPWR
+ _0609_ sky130_fd_sc_hd__mux4_2
XFILLER_149_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3872_ _0089_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or2_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2823_ _1649_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X
+ sky130_fd_sc_hd__inv_2
X_2754_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 net71 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__mux2_1
X_2685_ _1531_ _1258_ _1257_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__o21ai_4
X_5473_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net556
+ sky130_fd_sc_hd__buf_1
X_4424_ net1249 net1121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4355_ net1230 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3306_ net966 _1722_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2b_1
X_4286_ net1258 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q net653 VGND
+ VGND VPWR VPWR _1976_ sky130_fd_sc_hd__nor2_1
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3168_ net174 net119 net210 net990 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _1918_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_146_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ _0987_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__nand2_1
XFILLER_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3099_ net1264 net1018 net1226 net1039 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q VGND VGND VPWR VPWR
+ _1875_ sky130_fd_sc_hd__mux4_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout983 net985 VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__buf_2
Xfanout994 net996 VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__buf_8
Xfanout972 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 VGND VGND VPWR VPWR net972
+ sky130_fd_sc_hd__buf_8
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_310 net183 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_321 net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ _1326_ _1328_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__and2_4
XFILLER_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4140_ _0792_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__inv_1
X_4071_ _0667_ _0726_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ _1204_ net968 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__mux2_1
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4973_ net146 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_62_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3924_ net1051 net1046 net824 net822 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0593_ sky130_fd_sc_hd__mux4_1
XFILLER_149_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3855_ net190 net65 net23 net101 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q VGND VGND VPWR VPWR
+ _0528_ sky130_fd_sc_hd__mux4_2
X_2806_ _1633_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__a21bo_1
X_3786_ net189 net201 net2 net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0464_ sky130_fd_sc_hd__mux4_1
X_2737_ _1173_ _1552_ _1172_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__a21oi_2
X_5456_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net539
+ sky130_fd_sc_hd__buf_4
Xoutput520 net520 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[3] sky130_fd_sc_hd__buf_2
X_2668_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q _0257_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__a21oi_2
X_4407_ net1251 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput531 net531 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput553 net553 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput542 net542 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput586 net586 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[5] sky130_fd_sc_hd__buf_2
X_2599_ net144 net81 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q
+ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__mux2_1
Xoutput575 net575 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput564 net564 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[5] sky130_fd_sc_hd__buf_2
X_5387_ Tile_X0Y1_EE4END[14] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_1
X_4338_ net1245 net1141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput597 net597 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4269_ net1238 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_151 Tile_X0Y1_NN4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_140 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_184 net616 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 net560 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 net596 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_195 _0864_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3640_ _0066_ _0329_ _0328_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__o211a_1
X_3571_ _0262_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a21bo_1
X_5310_ net106 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_2
X_2522_ _0135_ _0134_ _0020_ _0588_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q VGND VGND VPWR VPWR
+ _1377_ sky130_fd_sc_hd__mux4_2
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5241_ Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_93_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2453_ _1311_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q _1313_
+ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o21ai_4
X_5172_ Tile_X0Y0_E6END[10] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
X_2384_ net111 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ _1249_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__o211a_1
X_4123_ _0453_ _0052_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__mux2_1
Xinput2 Tile_X0Y0_E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_4054_ _0713_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q VGND VGND
+ VPWR VPWR _0714_ sky130_fd_sc_hd__or2_4
XFILLER_56_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3005_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q net626 VGND
+ VGND VPWR VPWR _1794_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4956_ net161 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3907_ net1060 _0574_ _0529_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__o31ai_4
X_4887_ net1220 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3838_ _0064_ _0508_ _0512_ _0504_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__a31o_4
X_5508_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net591
+ sky130_fd_sc_hd__buf_1
X_3769_ net974 net969 net979 net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _0449_ sky130_fd_sc_hd__mux4_1
Xoutput361 net361 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput350 net350 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5439_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net531
+ sky130_fd_sc_hd__buf_1
Xoutput383 net383 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput372 net372 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[0] sky130_fd_sc_hd__buf_2
Xfanout1019 net1020 VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__clkbuf_4
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput394 net394 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[1] sky130_fd_sc_hd__buf_2
Xfanout1008 net1009 VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__buf_4
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4810_ net1216 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_61_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4741_ net1211 net1180 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4672_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs _0000_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3623_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0310_ _0312_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR
+ _0313_ sky130_fd_sc_hd__o211a_1
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3554_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q _0246_ VGND VGND
+ VPWR VPWR _0247_ sky130_fd_sc_hd__nand2_1
X_3485_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q VGND VGND VPWR
+ VPWR _0180_ sky130_fd_sc_hd__inv_1
X_2505_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q _0387_ VGND VGND
+ VPWR VPWR _1362_ sky130_fd_sc_hd__or2_1
X_5224_ net1185 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_2
X_2436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ _1297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR
+ VPWR _1298_ sky130_fd_sc_hd__o211a_1
X_5155_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 VGND VGND VPWR VPWR net247
+ sky130_fd_sc_hd__buf_1
X_2367_ net201 net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q VGND
+ VGND VPWR VPWR _1234_ sky130_fd_sc_hd__mux2_1
X_2298_ _1161_ _1168_ _1162_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__or3_4
X_4106_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] net1062 VGND VGND VPWR VPWR _0761_
+ sky130_fd_sc_hd__nand2b_1
X_5086_ net1200 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4037_ _0569_ _0567_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ _0541_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__a211o_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4939_ net148 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_40 net331 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 net408 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 Tile_X0Y0_S4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 Tile_X0Y1_E6END[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_95 Tile_X0Y1_EE4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3270_ net1023 net1004 net1010 net1008 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _2004_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_90_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _0640_ _0981_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__nor2_8
XFILLER_38_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2152_ _1022_ _1021_ _1023_ _0147_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a221o_1
X_2083_ _0799_ _0878_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__nor2_1
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2985_ _0027_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__a21oi_1
X_4724_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4655_ net1240 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput82 Tile_X0Y0_S4END[5] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput71 Tile_X0Y0_S2MID[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xinput60 Tile_X0Y0_S1END[3] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
X_3606_ net989 net1006 net864 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q VGND VGND VPWR VPWR
+ _0296_ sky130_fd_sc_hd__mux4_2
X_4586_ net1234 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_151_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput93 Tile_X0Y0_W1END[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_12
X_3537_ net811 net970 net664 net656 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0230_ sky130_fd_sc_hd__mux4_2
X_3468_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q VGND VGND VPWR
+ VPWR _0163_ sky130_fd_sc_hd__inv_1
X_5207_ net33 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
X_2419_ net75 net1073 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__mux2_1
X_3399_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q VGND VGND VPWR
+ VPWR _0094_ sky130_fd_sc_hd__inv_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5138_ net169 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5069_ net146 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2770_ _1599_ _1572_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__or2_4
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4440_ net35 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4371_ net1246 net1131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3322_ net967 _1657_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__and2b_1
X_3253_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q _1987_ _1988_
+ _1989_ _0193_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__a221o_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2204_ _0611_ _0612_ _0847_ _1073_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__a31o_1
X_3184_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q net1005 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q
+ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__o21ba_1
X_2135_ _1006_ _1004_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__xnor2_2
Xfanout1191 net168 VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__clkbuf_4
Xfanout1180 net1181 VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2066_ _0611_ _0612_ _0782_ _0783_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__and4_1
XFILLER_81_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer204 _0217_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd1_1
X_2968_ _0198_ _0560_ _0599_ _0554_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q VGND VGND VPWR VPWR
+ _1766_ sky130_fd_sc_hd__mux4_1
X_4707_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer237 net855 VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__clkbuf_2
Xrebuffer226 net844 VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__clkbuf_2
Xrebuffer215 _1029_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__buf_12
X_2899_ _1533_ _1550_ _1548_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__a21boi_1
X_4638_ net1258 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer259 net877 VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__buf_4
X_4569_ net1253 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone52 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 VGND VGND VPWR VPWR
+ net669 sky130_fd_sc_hd__buf_8
XFILLER_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3940_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q _0604_ _0607_
+ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a21o_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3871_ net1050 net1045 net824 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _0543_ sky130_fd_sc_hd__mux4_1
X_2822_ _1648_ _1630_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__mux2_4
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2753_ net107 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__mux2_4
XFILLER_117_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5472_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net555
+ sky130_fd_sc_hd__buf_8
X_2684_ _1530_ _1327_ _1326_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__o21a_4
X_4423_ net47 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4354_ net1229 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3305_ net928 _1557_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__and2b_1
XFILLER_100_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4285_ net30 net1185 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3236_ _1400_ _0637_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q
+ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__mux2_2
X_3167_ net1011 net1013 _1497_ _0960_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q VGND VGND VPWR VPWR
+ _1917_ sky130_fd_sc_hd__mux4_1
X_3098_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q _1873_ _1872_
+ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__o21ba_1
X_2118_ _0987_ _0988_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nand3_2
XFILLER_39_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2049_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q _0924_ _0920_
+ _0914_ _0916_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__o32a_4
XFILLER_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout984 net985 VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__buf_2
Xfanout995 net996 VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__clkbuf_4
Xfanout973 net975 VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__buf_8
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_300 net1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_322 net1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_311 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4070_ _0641_ _0708_ _0709_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_79_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3021_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _1807_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q
+ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4972_ net147 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_62_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3923_ _0591_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q VGND VGND
+ VPWR VPWR _0592_ sky130_fd_sc_hd__nor2_2
X_3854_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q _0526_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__o21ai_1
X_2805_ net1044 net1028 net1054 net669 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _1633_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_98_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3785_ _0083_ _0462_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__o21a_1
X_2736_ _1569_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 sky130_fd_sc_hd__mux2_4
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5455_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net538
+ sky130_fd_sc_hd__buf_4
X_2667_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q _1512_ _1514_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q VGND VGND VPWR VPWR
+ _1515_ sky130_fd_sc_hd__a211o_1
Xoutput510 net510 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[3] sky130_fd_sc_hd__buf_2
X_4406_ net1250 net1121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput521 net521 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput532 net532 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput543 net543 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput554 net554 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_132_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput587 net587 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[6] sky130_fd_sc_hd__buf_2
X_2598_ net233 _0237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q
+ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__mux2_1
Xoutput576 net576 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput565 net565 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[6] sky130_fd_sc_hd__buf_2
X_5386_ Tile_X0Y1_EE4END[13] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_1
X_4337_ net1243 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput598 net598 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[7] sky130_fd_sc_hd__buf_2
X_4268_ net1237 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3219_ net176 net1224 net1073 net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q VGND VGND VPWR VPWR
+ _1961_ sky130_fd_sc_hd__mux4_1
XFILLER_39_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4199_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__clkinv_2
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_141 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 Tile_X0Y1_NN4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 Tile_X0Y1_N4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 net560 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 net598 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 Tile_X0Y1_WW4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_196 _0906_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3570_ net992 net1021 net1002 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0262_ sky130_fd_sc_hd__mux4_1
X_2521_ net1066 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] VGND VGND VPWR VPWR _1376_
+ sky130_fd_sc_hd__nand2_1
X_5240_ Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
XFILLER_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2452_ _0151_ _1312_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__o21a_1
X_5171_ Tile_X0Y0_E6END[9] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
X_2383_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q _1248_ VGND VGND
+ VPWR VPWR _1249_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4122_ _0766_ _0767_ _0775_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q VGND VGND VPWR VPWR
+ _0776_ sky130_fd_sc_hd__a221o_1
X_4053_ net811 net664 net997 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0713_ sky130_fd_sc_hd__mux4_2
XFILLER_83_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3004_ _1790_ _1792_ _1793_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o22a_1
Xinput3 Tile_X0Y0_E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_39_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4955_ net1197 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3906_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] net1060 VGND VGND VPWR VPWR _0575_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_22_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4886_ net1209 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3837_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0511_ _0510_
+ _0063_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a211o_1
X_3768_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q _0447_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q
+ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o21ba_1
XFILLER_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5507_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net590
+ sky130_fd_sc_hd__buf_1
X_2719_ _1560_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 sky130_fd_sc_hd__mux2_4
X_3699_ _0075_ _0078_ _0072_ _0383_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q VGND VGND VPWR VPWR
+ _0384_ sky130_fd_sc_hd__mux4_2
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput362 net362 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput351 net351 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput340 net340 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[0] sky130_fd_sc_hd__buf_2
X_5438_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR net530
+ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput384 net384 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput373 net373 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput395 net395 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[2] sky130_fd_sc_hd__buf_2
X_5369_ Tile_X0Y1_E6END[6] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_58_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1009 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 VGND VGND VPWR VPWR net1009
+ sky130_fd_sc_hd__buf_8
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ net1210 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4671_ net1259 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3622_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q _0311_ VGND VGND
+ VPWR VPWR _0312_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ net93 net1226 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3484_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q VGND VGND VPWR
+ VPWR _0179_ sky130_fd_sc_hd__inv_1
X_2504_ _1358_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1360_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR VPWR
+ _1361_ sky130_fd_sc_hd__o211a_1
X_5223_ net49 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_1
XFILLER_142_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2435_ _1291_ _1293_ _1296_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ _0148_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a221o_1
X_5154_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net246
+ sky130_fd_sc_hd__buf_6
X_2366_ net100 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__mux2_1
X_4105_ _0755_ _0103_ _0757_ _0760_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ sky130_fd_sc_hd__a31o_4
X_2297_ _1165_ _1156_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__a21oi_4
XFILLER_110_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5085_ net160 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4036_ net73 net654 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux2_1
X_4938_ net1216 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_41 net345 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 Tile_X0Y0_FrameData[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ net154 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_63 Tile_X0Y0_W2MID[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_52 Tile_X0Y0_S4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 Tile_X0Y1_EE4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 Tile_X0Y1_E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2220_ _1074_ _1076_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__xnor2_4
XFILLER_87_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2151_ net137 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q
+ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__mux2_1
X_2082_ _0478_ _0640_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__nor2_1
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone198 net1020 VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__buf_6
XFILLER_34_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2984_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q net626 VGND VGND
+ VPWR VPWR _1777_ sky130_fd_sc_hd__or2_1
X_4723_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4654_ net1239 net1158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput72 Tile_X0Y0_S2MID[3] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_4
Xinput61 Tile_X0Y0_S2END[0] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_6
Xinput50 Tile_X0Y0_FrameData[3] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
X_3605_ net974 net969 net978 net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR
+ _0295_ sky130_fd_sc_hd__mux4_1
X_4585_ net1260 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput83 Tile_X0Y0_S4END[6] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput94 Tile_X0Y0_W1END[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
X_3536_ _0225_ _0226_ _0227_ _0039_ _0032_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a221o_2
XFILLER_88_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5206_ net32 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_1
X_3467_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR
+ VPWR _0162_ sky130_fd_sc_hd__inv_1
X_3398_ net109 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_1
X_2418_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q _0442_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__o21ba_4
X_2349_ net189 net8 net64 net116 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q VGND VGND VPWR VPWR
+ _1217_ sky130_fd_sc_hd__mux4_2
X_5137_ net1189 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5068_ net147 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4019_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__inv_2
XFILLER_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4370_ net1245 net1131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3321_ net967 _1626_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__and2b_1
X_3252_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q net1003 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__o21ba_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2203_ net1061 Tile_X0Y1_DSP_bot.B2 _0877_ _0725_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__o211a_4
X_3183_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q _0711_ VGND
+ VGND VPWR VPWR _1930_ sky130_fd_sc_hd__nand2_1
X_2134_ _0955_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__xor2_2
Xfanout1192 net167 VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__buf_4
Xfanout1170 net1173 VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__buf_1
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1181 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2065_ _0784_ _0478_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nor2_4
XFILLER_19_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2967_ net1050 net670 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 _0429_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 sky130_fd_sc_hd__mux4_1
X_2898_ _1718_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 sky130_fd_sc_hd__mux2_4
X_4706_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer216 _0257_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer238 net856 VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__clkbuf_2
Xrebuffer227 net845 VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__clkbuf_2
X_4637_ net30 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4568_ net1252 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4499_ net41 net1097 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3519_ net187 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone20 _1565_ net817 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q
+ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__mux2_4
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3870_ net1037 net1033 net865 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _0542_ sky130_fd_sc_hd__mux4_2
X_2821_ _0121_ _1647_ _1646_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2752_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q _1580_ _1584_
+ _1574_ _1576_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6
+ sky130_fd_sc_hd__o32a_4
XFILLER_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5471_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net554
+ sky130_fd_sc_hd__buf_4
XFILLER_129_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4422_ net1233 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2683_ _1375_ _1529_ _1374_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__a21oi_4
XFILLER_132_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4353_ net1228 net1139 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4284_ net1256 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3304_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q _2031_ _2035_
+ _2029_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr sky130_fd_sc_hd__a31o_4
X_3235_ net175 net211 net120 net995 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q VGND VGND VPWR VPWR
+ _1974_ sky130_fd_sc_hd__mux4_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3166_ _1913_ _1916_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A sky130_fd_sc_hd__mux2_1
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3097_ net1048 net1028 net1014 net1058 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR VPWR
+ _1873_ sky130_fd_sc_hd__mux4_1
X_2117_ _0957_ _0958_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_65_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ _0117_ _0923_ _0922_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q
+ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_105_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3999_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net69 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout985 net986 VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__buf_2
Xfanout974 net975 VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__buf_2
XFILLER_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout996 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 VGND VGND VPWR VPWR net996
+ sky130_fd_sc_hd__buf_8
XANTENNA_301 net1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_312 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_323 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3020_ _1806_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__inv_1
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4971_ net1217 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_62_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3922_ net1037 net1031 net982 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _0591_ sky130_fd_sc_hd__mux4_2
X_3853_ _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__inv_2
X_2804_ _1631_ _0120_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_98_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3784_ net1053 net1048 net1028 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0462_ sky130_fd_sc_hd__mux4_1
X_2735_ _1533_ _1550_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__xor2_2
X_5523_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net606
+ sky130_fd_sc_hd__buf_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net552
+ sky130_fd_sc_hd__buf_4
X_2666_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q _1513_ VGND VGND
+ VPWR VPWR _1514_ sky130_fd_sc_hd__and2b_1
Xoutput511 net511 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[4] sky130_fd_sc_hd__buf_2
Xoutput500 net500 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[23] sky130_fd_sc_hd__buf_2
X_4405_ net39 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput522 net522 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput533 net533 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput544 net544 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[1] sky130_fd_sc_hd__buf_2
X_5385_ Tile_X0Y1_EE4END[12] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_1
X_4336_ net1241 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput577 net577 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput566 net566 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput555 net555 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[11] sky130_fd_sc_hd__buf_8
X_2597_ _1446_ _1445_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_148_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput588 net588 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput599 net599 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[8] sky130_fd_sc_hd__buf_2
X_4267_ net1235 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_105_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4198_ Tile_X0Y1_DSP_bot.A1 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] net1059 VGND
+ VGND VPWR VPWR _0847_ sky130_fd_sc_hd__mux2_4
XFILLER_27_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3218_ _1954_ _1960_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 sky130_fd_sc_hd__mux2_1
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3149_ _1899_ _1901_ _1904_ _0186_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_114_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_120 Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 Tile_X0Y1_N4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 Tile_X0Y1_NN4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 net560 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_175 net599 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_197 _1565_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 Tile_X0Y1_WW4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2520_ _1371_ _1373_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__xor2_4
X_2451_ net989 net1023 net1004 net1008 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1312_ sky130_fd_sc_hd__mux4_1
X_5170_ Tile_X0Y0_E6END[8] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
X_2382_ _1248_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5
+ sky130_fd_sc_hd__inv_1
XFILLER_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4121_ net111 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__mux2_1
XFILLER_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4052_ net190 net135 net226 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q
+ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__mux4_2
X_3003_ _0414_ net1263 net60 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q VGND VGND VPWR VPWR
+ _1793_ sky130_fd_sc_hd__mux4_1
Xinput4 Tile_X0Y0_E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_39_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4954_ net1196 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_102_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3905_ _0529_ _0574_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X
+ sky130_fd_sc_hd__or2_1
XFILLER_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4885_ net1195 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3836_ net99 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3767_ net174 net178 net119 net141 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _0447_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_154_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ _1559_ _1524_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__nor2_2
X_5506_ Tile_X0Y1_W6END[11] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_4
XFILLER_145_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3698_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR _0383_
+ sky130_fd_sc_hd__inv_2
Xoutput330 net330 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[4] sky130_fd_sc_hd__buf_2
Xoutput352 net352 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[4] sky130_fd_sc_hd__buf_6
Xoutput341 net341 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[1] sky130_fd_sc_hd__buf_2
X_5437_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net529
+ sky130_fd_sc_hd__clkbuf_1
X_2649_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1497_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__a21oi_1
Xoutput385 net385 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput374 net374 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[11] sky130_fd_sc_hd__buf_8
Xoutput363 net363 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput396 net396 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5368_ Tile_X0Y1_E6END[5] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_1
X_4319_ net1259 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5299_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net391
+ sky130_fd_sc_hd__buf_6
XFILLER_27_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4670_ net1258 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_41_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3621_ net66 net94 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND
+ VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
X_3552_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__inv_2
X_2503_ _0160_ _1359_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__or2_1
X_3483_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR
+ VPWR _0178_ sky130_fd_sc_hd__inv_1
X_5222_ net48 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__buf_1
X_2434_ _1294_ _1295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q
+ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__mux2_1
X_5153_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net245
+ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2365_ _1230_ _1231_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__nand2b_4
X_4104_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0759_ _0758_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR VPWR
+ _0760_ sky130_fd_sc_hd__o211a_1
XFILLER_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2296_ _0900_ _1158_ _1164_ _1166_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a31o_1
X_5084_ net161 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4035_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q _0692_ _0696_
+ _0686_ _0688_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__o32a_4
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4937_ net1215 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_31 Tile_X0Y0_FrameData[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 Tile_X0Y0_EE4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ net1210 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_42 net347 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 Tile_X0Y0_S4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_75 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3819_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q _0491_ _0493_
+ _0487_ _0489_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__o32a_4
XANTENNA_97 Tile_X0Y1_EE4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 Tile_X0Y1_E6END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ net1202 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_153_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ net228 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q
+ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__o21a_1
X_2081_ _0611_ _0612_ _0641_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__and3_1
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2983_ _1773_ _1775_ _1776_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 sky130_fd_sc_hd__o22a_1
X_4722_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4653_ net45 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 Tile_X0Y0_FrameData[21] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
Xinput62 Tile_X0Y0_S2END[1] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput73 Tile_X0Y0_S2MID[4] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
Xinput51 Tile_X0Y0_FrameData[4] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
X_3604_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q _0293_ VGND VGND
+ VPWR VPWR _0294_ sky130_fd_sc_hd__or2_1
X_4584_ net1249 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput84 Tile_X0Y0_S4END[7] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput95 Tile_X0Y0_W1END[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
X_3535_ net668 _0226_ _0227_ _0039_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a22o_2
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3466_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q VGND VGND VPWR
+ VPWR _0161_ sky130_fd_sc_hd__inv_1
XFILLER_115_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5205_ net31 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_2
X_2417_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q net629 VGND VGND
+ VPWR VPWR _1280_ sky130_fd_sc_hd__nand2_1
X_3397_ net17 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
XFILLER_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2348_ _1216_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5
+ sky130_fd_sc_hd__inv_1
XFILLER_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5136_ net1188 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2279_ _0667_ _0521_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__or2_4
X_5067_ net148 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_4_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4018_ net207 net24 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q
+ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux2_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3320_ net967 _1603_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__and2b_1
XFILLER_152_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3251_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q _0711_ VGND VGND
+ VPWR VPWR _1988_ sky130_fd_sc_hd__nand2_1
X_2202_ _0478_ _0928_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__nor2_1
X_3182_ _0875_ _1510_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__mux2_1
Xfanout1182 net1183 VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__buf_2
X_2133_ _0726_ _0478_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__nor2_4
Xfanout1171 net1173 VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__buf_2
Xfanout1160 net1161 VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__buf_2
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1193 net166 VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__buf_4
X_2064_ net618 _0878_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__or2_1
XFILLER_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2966_ net62 net77 net113 net986 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
X_2897_ _1717_ _1674_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__xnor2_1
X_4705_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer217 _0254_ VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer228 net846 VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__clkbuf_2
X_4636_ net31 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer239 net857 VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__clkbuf_2
X_4567_ net1251 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4498_ net1245 net1097 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3518_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q _0030_ _0031_
+ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a21oi_1
X_3449_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR
+ VPWR _0144_ sky130_fd_sc_hd__inv_2
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5119_ net1201 net1153 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_150_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput230 Tile_X0Y1_W6END[0] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2820_ net868 net70 net14 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q VGND VGND VPWR VPWR
+ _1647_ sky130_fd_sc_hd__mux4_1
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2751_ _0114_ _1583_ _1582_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__o211a_1
XFILLER_129_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5470_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net568
+ sky130_fd_sc_hd__buf_6
X_2682_ _1528_ _1396_ _1395_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__o21bai_4
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4421_ net1232 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4352_ net1227 net1139 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4283_ net1255 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3303_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q _2032_ _2034_
+ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__a21o_1
XFILLER_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3234_ _1973_ _1972_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 sky130_fd_sc_hd__mux2_1
X_3165_ _1915_ _1914_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__mux2_1
XFILLER_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3096_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _1869_ _1871_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q VGND VGND VPWR VPWR
+ _1872_ sky130_fd_sc_hd__o211a_1
X_2116_ _0933_ _0986_ _0985_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__a21o_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2047_ net94 net1225 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3998_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q net105 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q
+ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__o21a_1
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2949_ net187 net199 net1263 net6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _1756_ sky130_fd_sc_hd__mux4_1
XFILLER_108_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4619_ net48 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_123_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout986 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 VGND VGND VPWR VPWR
+ net986 sky130_fd_sc_hd__buf_8
Xfanout975 net976 VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__buf_8
Xfanout997 net999 VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__buf_8
XANTENNA_313 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_302 net1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_324 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4970_ net149 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_62_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3921_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q net222 VGND VGND
+ VPWR VPWR _0590_ sky130_fd_sc_hd__or2_1
X_3852_ net199 net1261 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__mux2_1
X_2803_ net815 net1036 net1032 net983 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1631_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_98_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3783_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q _0460_ VGND VGND
+ VPWR VPWR _0461_ sky130_fd_sc_hd__or2_1
X_5522_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net605
+ sky130_fd_sc_hd__buf_1
X_2734_ _1568_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 sky130_fd_sc_hd__mux2_4
XFILLER_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5453_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net551
+ sky130_fd_sc_hd__buf_4
XFILLER_105_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2665_ net192 net137 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux2_1
Xoutput501 net501 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[24] sky130_fd_sc_hd__buf_2
X_4404_ net40 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput523 net523 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput534 net534 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput545 net545 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[2] sky130_fd_sc_hd__buf_2
X_5384_ Tile_X0Y1_EE4END[11] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_1
Xoutput512 net512 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[5] sky130_fd_sc_hd__buf_2
X_2596_ _1445_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__nand2_1
X_4335_ net1240 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput578 net578 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[5] sky130_fd_sc_hd__buf_8
Xoutput567 net567 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput556 net556 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_148_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput589 net589 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[0] sky130_fd_sc_hd__buf_2
X_4266_ net1234 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3217_ _1957_ _1958_ _1959_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__o22a_1
X_4197_ _0843_ _0846_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A1 sky130_fd_sc_hd__mux2_4
XFILLER_27_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3148_ _1902_ _1903_ _0185_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__mux2_1
XFILLER_131_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3079_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q _1856_ VGND VGND
+ VPWR VPWR _1857_ sky130_fd_sc_hd__and2b_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 Tile_X0Y1_N4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 Tile_X0Y1_NN4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 net560 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 Tile_X0Y1_W6END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 _0237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_198 net1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2450_ net974 net969 net979 net831 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1311_ sky130_fd_sc_hd__mux4_2
X_2381_ _0108_ _1243_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__o21ai_2
X_4120_ _0769_ _0771_ _0774_ _0080_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ sky130_fd_sc_hd__a22o_2
X_4051_ _0022_ _0126_ _0127_ _0267_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q VGND VGND VPWR VPWR
+ _0711_ sky130_fd_sc_hd__mux4_2
X_3002_ _1791_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__a21bo_1
Xinput5 Tile_X0Y0_E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4953_ net165 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_102_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3904_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q _0572_ _0573_
+ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__o21a_2
X_4884_ net1192 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3835_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q _0509_ VGND VGND
+ VPWR VPWR _0510_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_30_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3766_ _0444_ _0443_ _0445_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ _0051_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5505_ Tile_X0Y1_W6END[10] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__buf_4
X_2717_ _1465_ _1483_ _1523_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__and3_1
X_3697_ _0379_ _0377_ _0382_ _0077_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ sky130_fd_sc_hd__a22o_4
X_5436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR net528
+ sky130_fd_sc_hd__buf_1
Xoutput320 net320 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[13] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[5] sky130_fd_sc_hd__buf_2
XFILLER_145_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2648_ net189 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net225
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__mux4_2
Xoutput364 net364 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput375 net375 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[12] sky130_fd_sc_hd__buf_6
Xoutput386 net386 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_120_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5367_ Tile_X0Y1_E6END[4] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_1
X_2579_ net84 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__mux2_1
XFILLER_113_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput397 net397 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[4] sky130_fd_sc_hd__buf_2
X_4318_ net1258 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5298_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net390
+ sky130_fd_sc_hd__buf_1
X_4249_ _0891_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3620_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__inv_2
X_3551_ net57 net61 net617 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
X_2502_ net989 net1004 net994 net1011 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _1359_ sky130_fd_sc_hd__mux4_1
X_3482_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q VGND VGND VPWR
+ VPWR _0177_ sky130_fd_sc_hd__inv_2
XFILLER_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5221_ net1237 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2433_ net990 net1024 net996 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q VGND VGND VPWR VPWR
+ _1295_ sky130_fd_sc_hd__mux4_1
X_2364_ _1227_ _1229_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__nand2b_1
X_5152_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net244
+ sky130_fd_sc_hd__clkbuf_2
X_4103_ net188 net63 net7 net117 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q VGND VGND VPWR VPWR
+ _0759_ sky130_fd_sc_hd__mux4_2
X_2295_ _0896_ _1155_ _1164_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__and3_1
X_5083_ net162 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4034_ _0104_ _0695_ _0694_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_142_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4936_ net1214 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_32 net285 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 Tile_X0Y0_E6END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 Tile_X0Y0_EE4END[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ net1208 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_43 net354 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 net414 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3818_ _0095_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__nor2_1
XFILLER_20_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_98 Tile_X0Y1_EE4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_87 Tile_X0Y1_E6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ net1200 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3749_ _0424_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q _0425_
+ _0427_ _0021_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__a311o_1
X_5419_ net160 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_1
XFILLER_121_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2080_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__inv_2
XFILLER_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2982_ net920 net1225 net1263 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q VGND VGND VPWR VPWR
+ _1776_ sky130_fd_sc_hd__mux4_1
X_4721_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\] sky130_fd_sc_hd__dfxtp_1
X_4652_ net46 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput30 Tile_X0Y0_FrameData[12] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
X_3603_ net193 net68 net12 net115 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q VGND VGND VPWR VPWR
+ _0293_ sky130_fd_sc_hd__mux4_1
Xinput63 Tile_X0Y0_S2END[2] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xinput41 Tile_X0Y0_FrameData[22] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput52 Tile_X0Y0_FrameData[5] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
X_4583_ net1236 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput85 Tile_X0Y0_SS4END[0] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput74 Tile_X0Y0_S2MID[5] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput96 Tile_X0Y0_W1END[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
X_3534_ net196 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q
+ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
XFILLER_115_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3465_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR
+ VPWR _0160_ sky130_fd_sc_hd__inv_2
XFILLER_88_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q net809 _1278_
+ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__o21a_1
X_5204_ net1257 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_4
X_3396_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR
+ VPWR _0091_ sky130_fd_sc_hd__inv_2
X_2347_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q _1209_ _1211_
+ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__a31o_2
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5135_ net1187 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_150_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2278_ _1146_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__and2b_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5066_ net1216 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4017_ net78 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q
+ _0678_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__o211a_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4919_ net145 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_148_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3250_ _0875_ _1466_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__mux2_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2201_ net620 _0612_ _0611_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__and3b_1
X_3181_ net177 net1223 _0387_ net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _1928_ sky130_fd_sc_hd__mux4_1
Xfanout1150 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__buf_4
XFILLER_120_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1183 net1185 VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__buf_2
X_2132_ _0784_ _0878_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__nor2_1
Xfanout1172 net1173 VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1161 net1162 VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net165 VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__buf_4
X_2063_ _0934_ _0935_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_17_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2965_ net61 net114 net80 net1035 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
X_4704_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_2896_ _1604_ _1716_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__xor2_1
Xrebuffer229 net847 VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__clkbuf_2
Xrebuffer218 net836 VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__clkbuf_2
X_4635_ net32 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4566_ net1250 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3517_ _0205_ _0207_ _0210_ _0029_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q
+ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__a221o_2
X_4497_ net1243 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3448_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR
+ VPWR _0143_ sky130_fd_sc_hd__inv_1
X_3379_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q VGND VGND VPWR
+ VPWR _0074_ sky130_fd_sc_hd__inv_1
X_5118_ net1200 net1152 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5049_ net1194 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_27_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput220 Tile_X0Y1_W2END[6] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput231 Tile_X0Y1_W6END[1] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_4
XFILLER_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2750_ net68 net1225 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__mux2_1
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2681_ _1527_ _1409_ _1408_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__a21boi_4
X_4420_ net1231 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4351_ net28 net1139 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4282_ net1254 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3302_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 _2021_ _2033_ VGND VGND
+ VPWR VPWR _2034_ sky130_fd_sc_hd__a21o_1
XFILLER_140_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3233_ net174 net119 net210 net656 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q VGND VGND VPWR VPWR
+ _1973_ sky130_fd_sc_hd__mux4_1
XFILLER_140_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3164_ net1006 _0712_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__mux2_1
XFILLER_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3095_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q _1870_ VGND VGND
+ VPWR VPWR _1871_ sky130_fd_sc_hd__nand2_1
X_2115_ _0933_ _0985_ _0986_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__nand3_2
XFILLER_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2046_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _0921_ VGND VGND
+ VPWR VPWR _0922_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3997_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q _0314_ VGND VGND
+ VPWR VPWR _0661_ sky130_fd_sc_hd__nand2_1
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2948_ net1261 net98 net86 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q VGND VGND VPWR VPWR
+ _1755_ sky130_fd_sc_hd__mux4_1
XFILLER_148_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4618_ net49 net1167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2879_ net1043 net1047 net1055 net669 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q VGND VGND VPWR VPWR
+ _1702_ sky130_fd_sc_hd__mux4_1
XFILLER_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4549_ net51 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout976 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND VGND VPWR VPWR net976
+ sky130_fd_sc_hd__buf_8
XFILLER_38_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout998 net999 VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__buf_2
Xfanout987 net988 VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__buf_6
XANTENNA_303 net1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_314 net191 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_325 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3920_ _0583_ _0581_ _0587_ _0130_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a211o_1
X_3851_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q _0523_ VGND VGND
+ VPWR VPWR _0524_ sky130_fd_sc_hd__and2_1
X_3782_ net1018 net1036 net983 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q VGND VGND VPWR VPWR
+ _0460_ sky130_fd_sc_hd__mux4_1
X_2802_ _1629_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_98_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2733_ _1232_ _1532_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__xnor2_2
XFILLER_145_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5452_ Tile_X0Y0_S4END[15] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__buf_4
X_2664_ net228 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__mux2_4
Xoutput502 net502 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[25] sky130_fd_sc_hd__buf_2
X_4403_ net41 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput524 net524 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput535 net535 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[6] sky130_fd_sc_hd__buf_8
X_5383_ Tile_X0Y1_EE4END[10] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_1
Xoutput513 net513 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[6] sky130_fd_sc_hd__buf_2
X_2595_ _1119_ _1130_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__xor2_2
X_4334_ net1239 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput546 net546 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput557 net557 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput568 net568 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[9] sky130_fd_sc_hd__buf_8
XFILLER_113_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput579 net579 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[6] sky130_fd_sc_hd__buf_8
XFILLER_59_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4265_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q _0910_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__o21ai_1
X_4196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q _0841_ _0845_
+ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o21a_1
X_3216_ net1025 net1005 net812 net1009 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1959_ sky130_fd_sc_hd__mux4_1
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3147_ net203 net1223 net124 net1221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1903_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_19_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3078_ net822 net647 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q
+ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 Tile_X0Y1_EE4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 Tile_X0Y1_N4END[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 Tile_X0Y1_NN4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 net560 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 _0239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_177 net603 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2380_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1246_ _1245_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q VGND VGND VPWR VPWR
+ _1247_ sky130_fd_sc_hd__a211o_1
X_4050_ _0708_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__nand2_2
X_3001_ _0700_ _1238_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__mux2_4
Xinput6 Tile_X0Y0_E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4952_ net166 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3903_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q _0359_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q
+ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a21oi_1
X_4883_ net1191 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3834_ net63 net79 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3765_ net210 net1073 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3696_ _0380_ _0381_ _0076_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
X_2716_ _1558_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 sky130_fd_sc_hd__mux2_4
X_5504_ Tile_X0Y1_W6END[9] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__buf_4
XFILLER_145_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput310 net310 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5435_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR net527
+ sky130_fd_sc_hd__buf_1
X_2647_ _1492_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q _1493_
+ _1495_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q VGND VGND VPWR
+ VPWR _1496_ sky130_fd_sc_hd__a311o_1
Xoutput321 net321 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput343 net343 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput376 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR
+ Tile_X0Y0_NN4BEG[13] sky130_fd_sc_hd__buf_6
Xoutput365 net365 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput387 net387 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[9] sky130_fd_sc_hd__buf_4
X_5366_ Tile_X0Y1_E6END[3] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_1
XFILLER_59_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2578_ _1426_ _1427_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__xor2_2
XFILLER_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput398 net398 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4317_ net1257 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5297_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net389
+ sky130_fd_sc_hd__buf_1
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4248_ _0810_ _0892_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4179_ _0827_ _0825_ _0830_ _0137_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1
+ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_38_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3550_ _0241_ _0240_ _0242_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR VPWR
+ _0243_ sky130_fd_sc_hd__a221o_1
X_2501_ net974 net969 net978 net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR VPWR
+ _1358_ sky130_fd_sc_hd__mux4_2
X_3481_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR
+ VPWR _0176_ sky130_fd_sc_hd__inv_2
XFILLER_142_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5220_ net1238 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2432_ net974 net972 net978 net831 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1294_ sky130_fd_sc_hd__mux4_1
XFILLER_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2363_ _1229_ _1227_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and2b_1
X_5151_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net243
+ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_63_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4102_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q _0428_ VGND VGND
+ VPWR VPWR _0758_ sky130_fd_sc_hd__nand2_1
X_5082_ net163 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2294_ _0900_ _1158_ _1164_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a21oi_4
X_4033_ net94 net1225 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux2_1
XFILLER_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4935_ net1213 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_11 Tile_X0Y0_E6END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 Tile_X0Y0_EE4END[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ net158 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_44 net355 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net286 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4797_ net1199 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3817_ net65 net101 net77 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0492_ sky130_fd_sc_hd__mux4_1
XANTENNA_99 Tile_X0Y1_EE4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_88 Tile_X0Y1_E6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3748_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__inv_2
XFILLER_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3679_ net1261 net64 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
XFILLER_133_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5418_ net1200 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__buf_1
X_5349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net441
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2981_ _1774_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4720_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\] sky130_fd_sc_hd__dfxtp_1
X_4651_ net48 net1157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput31 Tile_X0Y0_FrameData[13] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
X_3602_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q _0288_ _0291_
+ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a21o_1
Xinput20 Tile_X0Y0_E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
Xinput64 Tile_X0Y0_S2END[3] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xinput42 Tile_X0Y0_FrameData[23] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput53 Tile_X0Y0_FrameData[6] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
X_4582_ net1233 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput86 Tile_X0Y0_SS4END[1] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
Xinput75 Tile_X0Y0_S2MID[6] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput97 Tile_X0Y0_W2END[0] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
X_3533_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q net221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__o21a_1
XFILLER_115_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3464_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q VGND VGND VPWR
+ VPWR _0159_ sky130_fd_sc_hd__inv_1
X_5203_ net29 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
X_2415_ _1277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a21oi_2
X_5134_ net1186 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3395_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q VGND VGND VPWR
+ VPWR _0090_ sky130_fd_sc_hd__inv_1
X_2346_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q _1214_ VGND VGND
+ VPWR VPWR _1215_ sky130_fd_sc_hd__nor2_1
XFILLER_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2277_ _0905_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__and2b_1
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5065_ net150 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4016_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q _0677_ VGND VGND
+ VPWR VPWR _0678_ sky130_fd_sc_hd__nand2_1
X_4918_ net156 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4849_ net1189 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_119_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2200_ _0981_ _0784_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__nor2_8
Xfanout1140 net1141 VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__clkbuf_4
X_3180_ _1922_ _1924_ _1927_ _0188_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1173 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__clkbuf_4
X_2131_ _0985_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__or2_1
Xfanout1151 net1152 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__clkbuf_2
Xfanout1162 net1163 VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1184 net1185 VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__buf_2
X_2062_ _0935_ _0934_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__and2b_1
Xfanout1195 net164 VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2964_ net21 net79 net64 net1038 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 sky130_fd_sc_hd__mux4_1
X_4703_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B3 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] sky130_fd_sc_hd__dfxtp_1
X_2895_ _1715_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] net1068 VGND VGND VPWR VPWR
+ _1716_ sky130_fd_sc_hd__mux2_4
Xrebuffer208 net835 VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__clkbuf_2
Xrebuffer219 net837 VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__clkbuf_2
X_4634_ net33 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4565_ net1248 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3516_ _0207_ _0205_ _0210_ _0029_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_4
X_4496_ net1241 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q VGND VGND VPWR
+ VPWR _0142_ sky130_fd_sc_hd__inv_1
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3378_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q VGND VGND VPWR
+ VPWR _0073_ sky130_fd_sc_hd__inv_2
X_2329_ net1064 _0171_ net1068 VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a21o_1
X_5117_ net1199 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5048_ net1193 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput210 Tile_X0Y1_W1END[0] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_4
XFILLER_102_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput232 Tile_X0Y1_WW4END[0] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
Xinput221 Tile_X0Y1_W2END[7] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2680_ _1526_ _1429_ _1428_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__o21ai_4
XFILLER_144_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4350_ net29 net1139 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3301_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q _0196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR VPWR
+ _2033_ sky130_fd_sc_hd__a31o_1
X_4281_ net1253 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3232_ net812 net1013 _1497_ _0609_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q VGND VGND VPWR VPWR
+ _1972_ sky130_fd_sc_hd__mux4_1
X_3163_ _0875_ _1489_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__mux2_1
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2114_ _0930_ _0932_ _0931_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__a21o_1
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3094_ net648 _1616_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__mux2_1
X_2045_ net60 net68 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q VGND
+ VGND VPWR VPWR _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3996_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q _0659_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ _0658_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__o211a_1
XFILLER_22_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2947_ _0081_ _1753_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__o21a_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4617_ net27 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2878_ _0175_ _1700_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__and2_1
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4548_ net1231 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4479_ net1259 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout977 net979 VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__buf_8
Xfanout966 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr VGND VGND VPWR VPWR net966
+ sky130_fd_sc_hd__buf_8
XFILLER_97_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout999 net1001 VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__buf_8
Xfanout988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VGND VGND VPWR VPWR net988
+ sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_304 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_326 net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3850_ net114 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
X_3781_ _0458_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] net1068 VGND VGND VPWR VPWR
+ _0459_ sky130_fd_sc_hd__mux2_4
X_2801_ _0317_ _1628_ _0121_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__mux2_1
X_2732_ _1567_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 sky130_fd_sc_hd__mux2_4
XFILLER_12_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5520_ Tile_X0Y1_WW4END[15] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5451_ Tile_X0Y0_S4END[14] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__buf_1
X_2663_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q _1510_ _1509_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR
+ _1511_ sky130_fd_sc_hd__o211a_1
X_4402_ net42 net1122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput525 net525 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[4] sky130_fd_sc_hd__buf_4
Xoutput536 net536 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[7] sky130_fd_sc_hd__buf_8
X_5382_ Tile_X0Y1_EE4END[9] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_1
Xoutput514 net514 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[7] sky130_fd_sc_hd__buf_2
X_2594_ net1067 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] _1444_ _1443_ VGND VGND VPWR
+ VPWR _1445_ sky130_fd_sc_hd__a22o_4
Xoutput503 net503 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[26] sky130_fd_sc_hd__buf_2
X_4333_ net1238 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput569 net569 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput547 net547 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput558 net558 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[14] sky130_fd_sc_hd__buf_2
X_4264_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_148_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3215_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _1955_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4195_ _0831_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q _0844_
+ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__a21o_1
X_3146_ net70 net82 net215 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1902_ sky130_fd_sc_hd__mux4_1
X_3077_ _0182_ _1855_ _1852_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2
+ sky130_fd_sc_hd__o21a_1
XFILLER_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3979_ _0643_ _0073_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__or2_4
XFILLER_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_134 Tile_X0Y1_N4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 Tile_X0Y1_EE4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 Tile_X0Y1_NN4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 net563 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_178 net606 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_189 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3000_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q _0571_ _1789_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q VGND VGND VPWR VPWR
+ _1790_ sky130_fd_sc_hd__a211oi_1
Xinput7 Tile_X0Y0_E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4951_ net1220 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3902_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 net109 net17 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux4_1
X_4882_ net1190 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3833_ _0505_ _0506_ _0507_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR VPWR
+ _0508_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3764_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q _0050_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_154_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3695_ net188 net1 net200 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q VGND VGND VPWR VPWR
+ _0381_ sky130_fd_sc_hd__mux4_1
X_5503_ Tile_X0Y1_W6END[8] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__buf_2
X_2715_ _1448_ _1525_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__xor2_1
Xoutput300 net300 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[24] sky130_fd_sc_hd__buf_2
X_5434_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR net526
+ sky130_fd_sc_hd__clkbuf_1
X_2646_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q _1494_ VGND VGND
+ VPWR VPWR _1495_ sky130_fd_sc_hd__nor2_1
Xoutput344 net344 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[15] sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput377 net377 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[14] sky130_fd_sc_hd__buf_8
Xoutput366 net366 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[7] sky130_fd_sc_hd__buf_2
XFILLER_113_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5365_ Tile_X0Y1_E6END[2] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_1
X_2577_ _1427_ _1426_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__nor2_4
Xoutput388 net388 VGND VGND VPWR VPWR Tile_X0Y0_UserCLKo sky130_fd_sc_hd__buf_1
XFILLER_141_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput399 net399 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[6] sky130_fd_sc_hd__clkbuf_4
X_5296_ clknet_1_0__leaf_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_2
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4316_ net1256 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4247_ _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__inv_2
X_4178_ _0828_ _0829_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q
+ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3129_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q net662 _1892_
+ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__a21o_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3480_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR
+ VPWR _0175_ sky130_fd_sc_hd__inv_2
XFILLER_127_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2500_ _0156_ _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__and2_1
X_2431_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q _1292_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__o21ba_1
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2362_ _0953_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__xnor2_1
X_5150_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net242
+ sky130_fd_sc_hd__buf_2
X_2293_ _1163_ _1154_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__xnor2_4
X_4101_ _0756_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q VGND VGND
+ VPWR VPWR _0757_ sky130_fd_sc_hd__nand2b_1
X_5081_ net1194 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4032_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0693_ VGND VGND
+ VPWR VPWR _0694_ sky130_fd_sc_hd__or2_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_regs_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK VGND VGND VPWR VPWR Tile_X0Y1_UserCLK_regs
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4934_ net1212 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_23 Tile_X0Y0_EE4END[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 Tile_X0Y0_E6END[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ net1206 net1118 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_45 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net293 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 Tile_X0Y0_S4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3816_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q _0490_ VGND VGND
+ VPWR VPWR _0491_ sky130_fd_sc_hd__nor2_1
X_4796_ net1198 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_67 net424 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q _0424_ _0425_
+ _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__a31oi_4
XANTENNA_89 Tile_X0Y1_E6END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3678_ _0363_ _0362_ _0364_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR VPWR
+ _0365_ sky130_fd_sc_hd__a221o_1
XFILLER_133_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2629_ _1472_ _0169_ _1478_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__a211o_1
X_5417_ net1201 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__buf_1
X_5348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 VGND VGND VPWR VPWR net440
+ sky130_fd_sc_hd__buf_1
XFILLER_153_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5279_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net362
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _0700_ _1217_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q
+ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__mux2_4
X_4650_ net1234 net1157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3601_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q _0290_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q
+ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o21ai_1
Xinput21 Tile_X0Y0_E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput10 Tile_X0Y0_E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput43 Tile_X0Y0_FrameData[26] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput32 Tile_X0Y0_FrameData[14] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput54 Tile_X0Y0_FrameData[7] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
X_4581_ net1232 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput65 Tile_X0Y0_S2END[4] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput76 Tile_X0Y0_S2MID[7] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput87 Tile_X0Y0_SS4END[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput98 Tile_X0Y0_W2END[1] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
X_3532_ _0219_ _0221_ _0224_ _0038_ _0036_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a221o_1
X_3463_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q VGND VGND VPWR
+ VPWR _0158_ sky130_fd_sc_hd__inv_1
X_5202_ net28 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_2
XFILLER_115_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2414_ _1277_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7
+ sky130_fd_sc_hd__inv_1
XFILLER_69_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5133_ net1219 net1152 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3394_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q VGND VGND VPWR
+ VPWR _0089_ sky130_fd_sc_hd__inv_2
X_2345_ _1213_ _1212_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q
+ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__mux2_1
XFILLER_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2276_ _0890_ _0904_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nand2_2
X_5064_ net151 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4015_ _0677_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_108_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4917_ net1195 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4848_ net1188 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4779_ net1217 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_87_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1130 net1132 VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__buf_2
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1174 net1176 VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__buf_2
X_2130_ net622 _0848_ net620 _0710_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__o22a_1
XFILLER_93_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1152 net1153 VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__clkbuf_2
Xfanout1163 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__clkbuf_2
X_2061_ _0850_ _0851_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__xnor2_1
Xfanout1196 net163 VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__buf_4
Xfanout1185 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_17_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2963_ net22 net78 net63 net1019 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 sky130_fd_sc_hd__mux4_1
X_4702_ clknet_2_2__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B2 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2894_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\] net1064 VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__mux2_4
Xrebuffer209 _0229_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd1_1
X_4633_ net34 net1165 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4564_ net1247 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3515_ _0208_ _0209_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q
+ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
X_4495_ net43 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3446_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q VGND VGND VPWR
+ VPWR _0141_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_139_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3377_ net80 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
X_2328_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ net1064 VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__nor2_4
X_5116_ net1198 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5047_ net1220 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_150_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2259_ _1128_ _1129_ _1124_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone24 net642 VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_8
XFILLER_138_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput211 Tile_X0Y1_W1END[1] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_4
Xinput200 Tile_X0Y1_N4END[6] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_4
Xinput233 Tile_X0Y1_WW4END[1] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
Xinput222 Tile_X0Y1_W2MID[0] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3300_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q VGND VGND VPWR VPWR
+ _2032_ sky130_fd_sc_hd__mux2_1
XFILLER_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4280_ net1252 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3231_ _0191_ _1967_ _1971_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1
+ sky130_fd_sc_hd__o21a_1
X_3162_ net177 net1223 net1072 net830 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q VGND VGND VPWR VPWR
+ _1913_ sky130_fd_sc_hd__mux4_1
XFILLER_39_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2113_ _0710_ _0848_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__nor3_1
X_3093_ _0571_ _0701_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__mux2_1
X_2044_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q _0917_ _0919_
+ _0118_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_65_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3995_ net186 net61 net24 net97 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q VGND VGND VPWR VPWR
+ _0659_ sky130_fd_sc_hd__mux4_2
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2946_ net1054 net1048 net1029 net1058 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _1753_ sky130_fd_sc_hd__mux4_1
X_2877_ net1019 net1038 net1034 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR VPWR
+ _1700_ sky130_fd_sc_hd__mux4_1
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4616_ net38 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4547_ net1230 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_147_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4478_ net1258 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR
+ VPWR _0124_ sky130_fd_sc_hd__inv_1
Xfanout967 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr VGND VGND VPWR VPWR net967
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout989 net990 VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__buf_2
Xfanout978 net979 VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_28_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_305 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_156_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_327 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3780_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\] net1064 VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_4
X_2800_ net187 net62 net26 net98 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q VGND VGND VPWR VPWR
+ _1628_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_70_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ _1531_ _1258_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__xor2_1
X_5450_ Tile_X0Y0_S4END[13] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__buf_1
XFILLER_145_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4401_ net1243 net1121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2662_ net185 net143 net76 net221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q VGND VGND VPWR VPWR
+ _1510_ sky130_fd_sc_hd__mux4_1
Xoutput526 net526 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[5] sky130_fd_sc_hd__buf_6
X_5381_ Tile_X0Y1_EE4END[8] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
X_2593_ net1063 _0167_ net1066 VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__a21oi_1
Xoutput515 net515 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput504 net504 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[27] sky130_fd_sc_hd__buf_2
Xoutput548 net548 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput559 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y1_SS4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput537 net537 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[0] sky130_fd_sc_hd__buf_2
X_4332_ net1237 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4263_ net193 net138 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__mux2_1
XFILLER_86_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q _1956_ VGND
+ VGND VPWR VPWR _1957_ sky130_fd_sc_hd__and2b_1
X_4194_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q _0833_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3145_ _0185_ _1900_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__o21a_1
X_3076_ _1853_ _1854_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__mux2_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3978_ net1050 net1045 net824 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0643_ sky130_fd_sc_hd__mux4_2
XFILLER_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2929_ net1042 net638 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__mux2_4
XFILLER_10_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 Tile_X0Y1_FrameData[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 net521 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_179 net608 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 net567 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer370 net1287 VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput8 Tile_X0Y0_E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4950_ net156 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3901_ _0570_ _0093_ _0092_ _0537_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q VGND VGND VPWR VPWR
+ _0571_ sky130_fd_sc_hd__mux4_2
X_4881_ net1189 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3832_ net7 net1262 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q VGND
+ VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_32_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5502_ Tile_X0Y1_W6END[7] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkbuf_2
X_3763_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0430_ _0438_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q _0441_ VGND VGND VPWR
+ VPWR _0443_ sky130_fd_sc_hd__a311o_1
XFILLER_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3694_ net1262 net99 net63 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q VGND VGND VPWR VPWR
+ _0380_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ _1557_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_154_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput301 net301 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[25] sky130_fd_sc_hd__buf_2
X_5433_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR net525
+ sky130_fd_sc_hd__buf_1
X_2645_ net188 net133 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__mux2_1
Xoutput334 net334 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
Xoutput323 net323 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput312 net312 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[6] sky130_fd_sc_hd__buf_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5364_ net138 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_2
Xoutput378 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y0_NN4BEG[15] sky130_fd_sc_hd__buf_6
Xoutput367 net367 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput356 net356 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput345 net345 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2576_ _1426_ _1427_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__nand2_1
X_4315_ net1255 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput389 net389 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[0] sky130_fd_sc_hd__buf_2
X_4246_ _0576_ _0710_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nor2_1
X_4177_ net1222 net71 net216 net235 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0829_ sky130_fd_sc_hd__mux4_1
X_3128_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q VGND VGND VPWR VPWR
+ _1892_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_38_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3059_ _0279_ net94 net2 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q VGND VGND VPWR VPWR
+ _1841_ sky130_fd_sc_hd__mux4_1
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2430_ net174 net178 net119 net123 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1292_ sky130_fd_sc_hd__mux4_1
X_2361_ _1141_ _1144_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__nor2_1
X_4100_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q VGND VGND VPWR VPWR
+ _0756_ sky130_fd_sc_hd__mux4_2
X_2292_ _0892_ _1150_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_102_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5080_ net1193 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_110_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4031_ net58 net66 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q VGND
+ VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4933_ net1211 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_111_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_13 Tile_X0Y0_E6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4864_ net1204 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_46 net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 net307 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 Tile_X0Y0_EE4END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4795_ net1197 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3815_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net9 net190 net1262 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q VGND VGND VPWR VPWR
+ _0490_ sky130_fd_sc_hd__mux4_1
XANTENNA_68 net432 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ net7 _0025_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__o21a_1
XANTENNA_79 net440 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3677_ net201 net8 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q VGND
+ VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux2_1
X_5416_ net1203 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkbuf_2
X_2628_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q _1475_ _1477_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q VGND VGND VPWR VPWR
+ _1478_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_120_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 VGND VGND VPWR VPWR net439
+ sky130_fd_sc_hd__buf_1
X_2559_ net196 net91 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__mux2_1
X_5278_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net361
+ sky130_fd_sc_hd__buf_1
X_4229_ net191 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net227
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q
+ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__mux4_1
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3600_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__inv_2
Xinput22 Tile_X0Y0_E6END[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput11 Tile_X0Y0_E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
X_4580_ net1231 net1078 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
Xinput44 Tile_X0Y0_FrameData[27] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput33 Tile_X0Y0_FrameData[15] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
Xinput55 Tile_X0Y0_FrameData[8] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
X_3531_ net827 _0221_ _0224_ _0038_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2
+ sky130_fd_sc_hd__a22o_4
Xinput88 Tile_X0Y0_SS4END[3] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 Tile_X0Y0_S4END[0] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 Tile_X0Y0_S2END[5] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_155_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput99 Tile_X0Y0_W2END[2] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
X_3462_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR
+ VPWR _0157_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5201_ net1227 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_4
X_2413_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q _1270_ _1272_
+ _1276_ _1274_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__o32a_1
X_3393_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q VGND VGND VPWR
+ VPWR _0088_ sky130_fd_sc_hd__inv_2
X_2344_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net1264 net192 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _1213_ sky130_fd_sc_hd__mux4_1
XFILLER_130_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5132_ net1218 net1152 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2275_ _0954_ _1138_ _1143_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__a31oi_4
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5063_ net1213 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4014_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q _0670_ _0672_
+ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_108_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4916_ net1192 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ net1187 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4778_ net1216 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3729_ _0056_ _0411_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a21o_1
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1131 net1132 VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1120 net1121 VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__clkbuf_2
Xfanout1164 net1165 VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__buf_2
Xfanout1142 net1150 VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__buf_2
Xfanout1153 net1155 VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__clkbuf_2
Xfanout1175 net1176 VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__clkbuf_4
X_2060_ _0930_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__nand2_2
Xfanout1197 net162 VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net173 VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2962_ _1763_ _1765_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4701_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B1 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] sky130_fd_sc_hd__dfxtp_1
X_4632_ net1252 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2893_ _1685_ _1684_ _1714_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ sky130_fd_sc_hd__o21ai_2
XFILLER_8_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4563_ net1246 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4494_ net44 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3514_ net79 net87 net99 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0209_ sky130_fd_sc_hd__mux4_1
X_3445_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q VGND VGND VPWR
+ VPWR _0140_ sky130_fd_sc_hd__inv_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3376_ net74 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
X_2327_ _1196_ _1189_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X
+ sky130_fd_sc_hd__or2_4
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5115_ net1197 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5046_ net1209 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2258_ _1120_ _1123_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__xnor2_2
X_2189_ _1052_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone47 net979 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__buf_8
Xclone36 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 VGND VGND VPWR VPWR net653
+ sky130_fd_sc_hd__buf_8
XFILLER_119_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput201 Tile_X0Y1_N4END[7] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput234 Tile_X0Y1_WW4END[2] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_2
Xinput223 Tile_X0Y1_W2MID[1] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_2
Xinput212 Tile_X0Y1_W1END[2] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_59_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3230_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q _1970_ _1969_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q VGND VGND VPWR VPWR
+ _1971_ sky130_fd_sc_hd__a211o_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3161_ _1911_ _1912_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A sky130_fd_sc_hd__mux2_1
XFILLER_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2112_ net622 net620 VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__or2_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3092_ _1862_ _1865_ _1868_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 sky130_fd_sc_hd__a22o_1
X_2043_ _0117_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3994_ _0654_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q _0657_
+ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__a21o_1
X_2945_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q _1751_ VGND VGND
+ VPWR VPWR _1752_ sky130_fd_sc_hd__or2_1
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2876_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _1216_ _1698_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR VPWR
+ _1699_ sky130_fd_sc_hd__o211a_1
X_4615_ net1236 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4546_ net1229 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_116_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4477_ net30 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3428_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q VGND VGND VPWR
+ VPWR _0123_ sky130_fd_sc_hd__inv_1
Xfanout968 _0340_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__buf_8
X_3359_ net191 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__inv_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout979 net981 VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__buf_12
XANTENNA_306 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5029_ net1211 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2730_ _1565_ _1566_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 sky130_fd_sc_hd__mux2_8
XTAP_TAPCELL_ROW_70_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2661_ _1505_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q _1508_
+ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__a21o_1
X_4400_ net1241 net1121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput527 net527 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[6] sky130_fd_sc_hd__buf_2
X_5380_ Tile_X0Y1_EE4END[7] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_1
Xoutput516 net516 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[9] sky130_fd_sc_hd__buf_2
X_2592_ net1065 Tile_X0Y1_DSP_bot.C4 VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__or2_4
Xoutput505 net505 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[28] sky130_fd_sc_hd__buf_2
XFILLER_113_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput549 net549 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput538 net538 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[10] sky130_fd_sc_hd__buf_2
X_4331_ net1235 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4262_ net875 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q
+ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__mux2_4
XFILLER_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3213_ _0712_ _0875_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__mux2_2
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4193_ _0842_ _0823_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__mux2_1
X_3144_ net992 net1021 net1002 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1900_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_78_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3075_ net641 _0683_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__mux2_1
XFILLER_94_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3977_ net1017 net823 net865 net867 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0642_ sky130_fd_sc_hd__mux4_2
XFILLER_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2928_ _1739_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q _1740_
+ _1742_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 sky130_fd_sc_hd__a31o_4
XFILLER_10_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2859_ _0179_ _1682_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__o21ai_1
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4529_ net1244 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_125 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 Tile_X0Y1_FrameData[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_114 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_136 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 net532 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_169 net572 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer371 net1288 VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__clkbuf_2
Xrebuffer360 net1277 VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 Tile_X0Y0_E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3900_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR _0570_
+ sky130_fd_sc_hd__inv_1
X_4880_ net1188 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_102_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ _0062_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q
+ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a21oi_1
X_3762_ _0430_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q _0438_
+ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__a31o_4
X_5501_ Tile_X0Y1_W6END[6] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkbuf_2
X_3693_ _0076_ _0378_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2713_ _1556_ _1519_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_154_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5432_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR net524
+ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_33_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2644_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q _0677_ VGND VGND
+ VPWR VPWR _1493_ sky130_fd_sc_hd__or2_1
Xoutput324 net324 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput302 net302 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[26] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[7] sky130_fd_sc_hd__buf_2
X_5363_ net137 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_1
X_2575_ _1118_ _1131_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__xor2_4
Xoutput368 net368 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput357 net357 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput346 net346 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[6] sky130_fd_sc_hd__buf_2
X_4314_ net1254 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput379 net379 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[1] sky130_fd_sc_hd__buf_2
X_5294_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net377
+ sky130_fd_sc_hd__buf_4
X_4245_ _0521_ _0762_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__or2_1
XFILLER_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4176_ net174 net180 net196 net125 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0828_ sky130_fd_sc_hd__mux4_1
X_3127_ _1886_ _1888_ _1891_ _0184_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3058_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q _1839_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q
+ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer190 net808 VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_142_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2360_ _1226_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] net1069 VGND VGND VPWR VPWR
+ _1227_ sky130_fd_sc_hd__mux2_4
X_2291_ _0903_ _1158_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__and2_1
X_4030_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q _0689_ _0691_
+ _0105_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4932_ net1210 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_14 Tile_X0Y0_E6END[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4863_ net1202 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_47 net385 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net309 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 Tile_X0Y0_EE4END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ net1196 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3814_ _0488_ _0095_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q
+ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__o21ai_2
XANTENNA_69 net433 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net398 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ net200 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q
+ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3676_ _0048_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a21oi_1
X_5415_ net1205 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkbuf_2
X_2627_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q _1476_ VGND VGND
+ VPWR VPWR _1477_ sky130_fd_sc_hd__nand2_1
X_2558_ net216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__mux2_4
X_5346_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net438
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5277_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net360
+ sky130_fd_sc_hd__buf_1
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2489_ _1346_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__inv_2
X_4228_ net190 net135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q
+ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__mux4_2
XFILLER_101_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4159_ _0801_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__nand2_1
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 Tile_X0Y0_E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
Xinput45 Tile_X0Y0_FrameData[28] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput34 Tile_X0Y0_FrameData[16] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput23 Tile_X0Y0_EE4END[0] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
X_3530_ _0222_ _0223_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
Xinput78 Tile_X0Y0_S4END[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
Xinput89 Tile_X0Y0_SS4END[4] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput67 Tile_X0Y0_S2END[6] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput56 Tile_X0Y0_FrameData[9] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3461_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q VGND VGND VPWR
+ VPWR _0156_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2412_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1275_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q
+ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__o21ai_1
X_3392_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q VGND VGND VPWR
+ VPWR _0087_ sky130_fd_sc_hd__inv_2
X_5200_ net1228 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__buf_4
X_2343_ net57 net59 net67 net1226 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1212_ sky130_fd_sc_hd__mux4_1
XFILLER_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5131_ net1217 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5062_ net1212 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4013_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q _0675_ VGND VGND
+ VPWR VPWR _0676_ sky130_fd_sc_hd__nor2_1
X_2274_ _0951_ _1141_ _0952_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__o21a_1
XFILLER_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4915_ net1191 net1108 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4846_ net1186 net1125 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4777_ net1215 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3728_ net175 net181 net126 net1221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0411_ sky130_fd_sc_hd__mux4_1
X_3659_ net210 net1073 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__mux2_1
X_5329_ Tile_X0Y0_WW4END[4] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_3_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1132 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net1122 VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1110 net1111 VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__clkbuf_2
Xfanout1165 net1167 VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__buf_1
Xfanout1154 net1155 VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__clkbuf_4
Xfanout1143 net1144 VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1176 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__buf_2
Xfanout1198 net161 VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__buf_4
XFILLER_66_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1187 net172 VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2961_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q net621 _1764_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q VGND VGND VPWR VPWR
+ _1765_ sky130_fd_sc_hd__a211o_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4700_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.B0 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] sky130_fd_sc_hd__dfxtp_1
X_4631_ net1251 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2892_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q _1699_ _1713_
+ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__or3_1
XFILLER_8_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
X_4562_ net1245 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3513_ net208 net1 net25 net1262 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0208_ sky130_fd_sc_hd__mux4_1
X_4493_ net1238 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3444_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q VGND VGND VPWR
+ VPWR _0139_ sky130_fd_sc_hd__inv_2
X_3375_ net18 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkinv_2
X_2326_ _1194_ _1191_ _1195_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q VGND VGND VPWR VPWR
+ _1196_ sky130_fd_sc_hd__o221a_1
X_5114_ net1196 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5045_ net1195 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2257_ _1121_ _1125_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ _1057_ _1053_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4829_ net160 net1126 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput202 Tile_X0Y1_NN4END[0] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__buf_1
Xinput235 Tile_X0Y1_WW4END[3] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
Xinput224 Tile_X0Y1_W2MID[2] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
Xinput213 Tile_X0Y1_W1END[3] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_59_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3160_ net1025 _0823_ _0977_ _1416_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ _1912_ sky130_fd_sc_hd__mux4_1
X_3091_ _1867_ _1866_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q
+ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__mux2_4
X_2111_ _0959_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__nand2_4
X_2042_ net1263 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3993_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q _0656_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__o21ai_1
X_2944_ net1036 net1032 net985 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q VGND VGND VPWR VPWR
+ _1751_ sky130_fd_sc_hd__mux4_1
X_2875_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__nand2_1
X_4614_ net1233 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4545_ net1228 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4476_ net1256 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3427_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q VGND VGND VPWR
+ VPWR _0122_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3358_ net76 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__inv_2
X_2309_ _1178_ _1179_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q
+ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__mux2_2
Xfanout969 net972 VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__clkbuf_4
X_3289_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__nor2_1
XANTENNA_307 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5028_ net1210 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_318 Tile_X0Y0_E6END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_79_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2660_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q _1507_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput517 net517 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[0] sky130_fd_sc_hd__buf_2
X_2591_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q _1435_ _1437_
+ _1442_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C4 sky130_fd_sc_hd__a31o_1
Xoutput506 net506 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[29] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_97_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput528 net528 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput539 net539 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[11] sky130_fd_sc_hd__buf_2
X_4330_ net1234 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4261_ _0906_ _0405_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__mux2_1
XFILLER_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3212_ _1473_ _1400_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4192_ net133 net224 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__mux4_1
X_3143_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q _1898_ VGND VGND
+ VPWR VPWR _1899_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3074_ net669 _1204_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__inv_2
X_2927_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q _0560_ _1741_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q VGND VGND VPWR VPWR
+ _1742_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_33_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2858_ _1680_ _1681_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__mux2_1
XFILLER_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2789_ _1609_ _1611_ _1618_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X
+ sky130_fd_sc_hd__o21ai_1
X_4528_ net1241 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4459_ net1235 net1104 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_159 net541 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer361 net1278 VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__clkbuf_2
Xrebuffer372 net1289 VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q _0239_ VGND VGND
+ VPWR VPWR _0505_ sky130_fd_sc_hd__or2_1
X_3761_ _0439_ _0021_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o21a_1
X_5500_ Tile_X0Y1_W6END[5] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_2
X_2712_ _1518_ net829 VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__nor2_4
XFILLER_118_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3692_ net1053 net828 net1028 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0378_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5431_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR net523
+ sky130_fd_sc_hd__clkbuf_1
X_2643_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__nand2_2
Xoutput325 net325 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[18] sky130_fd_sc_hd__buf_2
Xoutput303 net303 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[27] sky130_fd_sc_hd__buf_2
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput314 net314 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[8] sky130_fd_sc_hd__buf_2
XFILLER_126_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5362_ net136 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__buf_1
X_2574_ _1425_ _1424_ net1066 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] VGND VGND VPWR
+ VPWR _1426_ sky130_fd_sc_hd__a2bb2o_4
Xoutput369 net369 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput347 net347 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput336 net336 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_141_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4313_ net1253 net1146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4244_ _0889_ _0822_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nand2_2
XFILLER_113_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4175_ _0136_ _0826_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__o21a_1
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3126_ _1889_ _1890_ _0183_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__mux2_1
XFILLER_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3057_ _1616_ _0518_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3959_ net973 net977 net830 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0626_ sky130_fd_sc_hd__mux4_2
XFILLER_129_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer180 net798 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer191 net810 VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2290_ _0905_ _1149_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__o21a_1
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4931_ net157 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4862_ net1200 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3813_ net1050 net1045 net1026 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0488_ sky130_fd_sc_hd__mux4_2
XANTENNA_37 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 Tile_X0Y0_E6END[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 Tile_X0Y0_EE4END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 Tile_X0Y0_S4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ net1194 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_59 net400 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q net104 VGND VGND
+ VPWR VPWR _0425_ sky130_fd_sc_hd__or2_1
X_3675_ net635 _0259_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ _0278_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a211o_1
XFILLER_118_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5414_ net158 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_2
X_2626_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net227 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__mux2_2
X_5345_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net437
+ sky130_fd_sc_hd__buf_1
X_2557_ _1408_ _1409_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nand2_4
X_5276_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net359
+ sky130_fd_sc_hd__buf_1
X_2488_ _0563_ _0387_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__mux2_4
XFILLER_101_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4227_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q _0866_ _0868_
+ _0872_ _0874_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__a32o_4
X_4158_ _0667_ _0799_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nor2_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4089_ net107 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q
+ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__o21a_1
X_3109_ net178 net197 net231 net1023 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A sky130_fd_sc_hd__mux4_1
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 Tile_X0Y0_E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput46 Tile_X0Y0_FrameData[29] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput35 Tile_X0Y0_FrameData[17] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput24 Tile_X0Y0_EE4END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput79 Tile_X0Y0_S4END[2] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xinput57 Tile_X0Y0_S1END[0] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_6
Xinput68 Tile_X0Y0_S2END[7] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q VGND VGND VPWR
+ VPWR _0155_ sky130_fd_sc_hd__inv_1
X_3391_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q VGND VGND VPWR
+ VPWR _0086_ sky130_fd_sc_hd__inv_1
X_2411_ net975 net972 net979 net831 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR
+ _1275_ sky130_fd_sc_hd__mux4_1
X_2342_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _1210_ VGND VGND
+ VPWR VPWR _1211_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5130_ net149 net1152 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5061_ net1211 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4012_ _0673_ _0674_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q
+ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__mux2_1
X_2273_ _1143_ _1138_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__and2_4
XFILLER_92_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4914_ net1190 net1108 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4845_ net1219 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4776_ net1214 net1142 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3727_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q _0409_ VGND VGND
+ VPWR VPWR _0410_ sky130_fd_sc_hd__and2_1
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3658_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q _0068_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q
+ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a21oi_1
X_3589_ _0279_ net191 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q
+ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_4
X_2609_ _1456_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1459_
+ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__o21a_1
X_5328_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net411
+ sky130_fd_sc_hd__buf_6
X_5259_ net619 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_4
XFILLER_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1122 net1123 VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__clkbuf_4
Xfanout1100 net1101 VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_2
Xfanout1111 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__clkbuf_2
Xfanout1155 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__clkbuf_1
Xfanout1144 net1145 VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__buf_1
Xfanout1133 net1134 VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__buf_2
XFILLER_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1166 net1167 VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__clkbuf_2
Xfanout1177 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__clkbuf_2
Xfanout1188 net171 VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__clkbuf_4
Xfanout1199 net160 VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2960_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q net828 VGND
+ VGND VPWR VPWR _1764_ sky130_fd_sc_hd__nor2_1
X_2891_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q _1248_ _1712_
+ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__o21a_1
X_4630_ net1250 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4561_ net1243 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4492_ net1237 net1097 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3512_ _0028_ _0206_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q
+ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__o21a_1
XFILLER_143_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3443_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q VGND VGND VPWR
+ VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5113_ net1194 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3374_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q VGND VGND VPWR
+ VPWR _0069_ sky130_fd_sc_hd__inv_2
X_2325_ net208 net6 net62 net98 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q VGND VGND VPWR VPWR
+ _1195_ sky130_fd_sc_hd__mux4_2
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5044_ net1192 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2256_ _1093_ _1122_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__xor2_2
XFILLER_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_108_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2187_ _1053_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4828_ net1198 net1126 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_117_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone49 _1422_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__clkbuf_1
Xclone38 net908 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__buf_6
X_4759_ net1220 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput214 Tile_X0Y1_W2END[0] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput225 Tile_X0Y1_W2MID[3] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_2
Xinput203 Tile_X0Y1_NN4END[1] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_126_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3090_ net1048 net1028 net1014 net822 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _1867_ sky130_fd_sc_hd__mux4_1
X_2110_ _0521_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nor2_2
X_2041_ _0414_ net193 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q
+ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__mux2_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3992_ _0655_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__inv_1
X_2943_ _1749_ _1750_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 sky130_fd_sc_hd__mux2_1
X_2874_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q _1693_ _1697_
+ _1687_ _1689_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7
+ sky130_fd_sc_hd__o32a_1
X_4613_ net1232 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4544_ net1227 net1086 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4475_ net1255 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3426_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR
+ VPWR _0121_ sky130_fd_sc_hd__inv_2
X_3357_ net20 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
X_2308_ net57 net59 net67 net1226 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1179_ sky130_fd_sc_hd__mux4_1
X_3288_ net619 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__mux2_4
X_5027_ net1208 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ net832 _0726_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__nor2_4
XANTENNA_308 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_319 _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_143_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput518 net518 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[1] sky130_fd_sc_hd__buf_8
Xoutput507 net507 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[2] sky130_fd_sc_hd__buf_2
X_2590_ _1438_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _1441_
+ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__o21a_1
XFILLER_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput529 net529 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4260_ net184 net129 net92 net220 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q VGND VGND VPWR VPWR
+ _0906_ sky130_fd_sc_hd__mux4_2
XFILLER_86_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4191_ net202 net71 net125 net216 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q VGND VGND VPWR VPWR
+ _0841_ sky130_fd_sc_hd__mux4_1
X_3211_ _1952_ _1953_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q
+ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__mux2_1
X_3142_ net869 net664 net830 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q VGND VGND VPWR VPWR
+ _1898_ sky130_fd_sc_hd__mux4_1
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3073_ _1849_ _1850_ _1851_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q VGND VGND VPWR VPWR
+ _1852_ sky130_fd_sc_hd__a221o_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3975_ net1059 Tile_X0Y1_DSP_bot.A3 _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__o21ai_4
X_2926_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q net983 VGND
+ VGND VPWR VPWR _1741_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2857_ net1043 net1047 net1055 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q VGND VGND VPWR VPWR
+ _1681_ sky130_fd_sc_hd__mux4_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2788_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q _1613_ _1615_
+ _1617_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q VGND VGND VPWR
+ VPWR _1618_ sky130_fd_sc_hd__a311o_1
X_4527_ net1240 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4458_ net1234 net1104 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3409_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR
+ VPWR _0104_ sky130_fd_sc_hd__inv_2
XFILLER_77_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4389_ net1232 net1129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_116 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_105 net497 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer340 net958 VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__clkbuf_2
Xrebuffer373 net1290 VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__clkbuf_2
Xrebuffer362 net1279 VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q net867 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q
+ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o21ba_1
X_2711_ _1555_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 sky130_fd_sc_hd__mux2_4
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3691_ _0376_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q VGND VGND
+ VPWR VPWR _0377_ sky130_fd_sc_hd__or2_4
X_5430_ net665 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_30_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2642_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q _1488_ _1490_
+ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__and3_1
XFILLER_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput326 net326 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[19] sky130_fd_sc_hd__buf_2
Xoutput304 net304 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[9] sky130_fd_sc_hd__buf_2
XFILLER_133_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5361_ net135 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_2
X_2573_ net1063 _0166_ net1066 VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__a21o_1
Xoutput359 net359 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput348 net348 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput337 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 VGND VGND VPWR VPWR
+ Tile_X0Y0_N1BEG[1] sky130_fd_sc_hd__buf_8
X_5292_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net375
+ sky130_fd_sc_hd__clkbuf_2
X_4312_ net1252 net1147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4243_ _0887_ _0888_ _0886_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__a21bo_1
XFILLER_113_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4174_ net992 net1021 net1002 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0826_ sky130_fd_sc_hd__mux4_1
X_3125_ net177 net179 net195 net142 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _1890_ sky130_fd_sc_hd__mux4_1
XFILLER_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3056_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q _1837_ VGND
+ VGND VPWR VPWR _1838_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3958_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0622_ _0624_
+ _0122_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a211o_1
XFILLER_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2909_ net1043 net1030 net1047 net1015 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q VGND VGND VPWR VPWR
+ _1725_ sky130_fd_sc_hd__mux4_1
X_3889_ _0557_ _0558_ _0559_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a22oi_4
XFILLER_104_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer181 net799 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer170 net788 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer192 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 VGND VGND VPWR VPWR
+ net809 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4930_ net158 net1100 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4861_ net1199 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_43_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3812_ _0486_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q VGND VGND
+ VPWR VPWR _0487_ sky130_fd_sc_hd__nor2_2
XANTENNA_38 net315 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 Tile_X0Y0_EE4END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 Tile_X0Y0_E6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4792_ net1193 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3743_ _0371_ _0365_ _0375_ _0025_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__a211o_1
XANTENNA_49 Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3674_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q net1027 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o21ba_1
X_2625_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__inv_1
X_5413_ net157 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2556_ _1406_ _1407_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__or2_1
XFILLER_87_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5275_ Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_4
X_2487_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q _1342_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q
+ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4226_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q _0873_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__o21ba_1
X_4157_ _0668_ _0801_ _0800_ _0802_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3108_ net181 net1222 net196 net993 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A sky130_fd_sc_hd__mux4_1
X_4088_ _0744_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q VGND VGND
+ VPWR VPWR _0745_ sky130_fd_sc_hd__nand2_2
X_3039_ net637 net1264 net95 net1035 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q VGND VGND VPWR VPWR
+ _1824_ sky130_fd_sc_hd__mux4_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 Tile_X0Y0_FrameData[18] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xinput25 Tile_X0Y0_EE4END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 Tile_X0Y0_E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
Xinput69 Tile_X0Y0_S2MID[0] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
Xinput58 Tile_X0Y0_S1END[1] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xinput47 Tile_X0Y0_FrameData[2] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
X_2410_ _1273_ _0149_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__nor2_1
X_3390_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR
+ VPWR _0085_ sky130_fd_sc_hd__inv_2
X_2341_ net1043 net1030 net1047 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _1210_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_110_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2272_ _1142_ _1141_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__nor2_4
XFILLER_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5060_ net155 net1172 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4011_ net64 net100 net80 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q VGND VGND VPWR VPWR
+ _0674_ sky130_fd_sc_hd__mux4_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4913_ net1189 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4844_ net1218 net1125 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4775_ net152 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3726_ net72 net217 net84 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q VGND VGND VPWR VPWR
+ _0409_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_119_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3657_ _0318_ _0332_ _0342_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q
+ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a211o_1
X_2608_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1458_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q
+ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__a21oi_1
X_3588_ net635 _0259_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__a21o_4
X_5327_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net410
+ sky130_fd_sc_hd__buf_6
X_2539_ _1376_ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__nand2_2
X_5258_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net350
+ sky130_fd_sc_hd__buf_4
X_5189_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR net272
+ sky130_fd_sc_hd__buf_6
X_4209_ net993 net1021 net1002 net1010 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0858_ sky130_fd_sc_hd__mux4_1
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1112 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__buf_2
XFILLER_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1101 net1106 VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__clkbuf_4
Xfanout1156 net1158 VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__buf_2
Xfanout1134 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__clkbuf_2
Xfanout1123 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__buf_2
Xfanout1145 net1150 VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__buf_2
Xfanout1167 net1168 VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1189 net170 VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__clkbuf_4
Xfanout1178 net1180 VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__buf_2
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2890_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q VGND VGND VPWR VPWR
+ _1712_ sky130_fd_sc_hd__a21oi_1
X_4560_ net1241 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4491_ net1235 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3511_ net1050 net1045 net1026 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0206_ sky130_fd_sc_hd__mux4_2
XFILLER_143_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3442_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q VGND VGND VPWR
+ VPWR _0137_ sky130_fd_sc_hd__inv_1
XFILLER_143_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3373_ net75 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
X_2324_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q _1193_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q
+ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__o21ai_1
X_5112_ net1193 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5043_ net1191 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2255_ _1121_ net829 VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__nand2_4
X_2186_ _1055_ _1054_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__xnor2_4
XFILLER_84_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4827_ net1197 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclone39 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 VGND VGND VPWR VPWR net656
+ sky130_fd_sc_hd__buf_8
X_4758_ net1209 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4689_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0017_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_108_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3709_ _0391_ _0393_ _0298_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6
+ sky130_fd_sc_hd__a21o_4
XFILLER_104_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput215 Tile_X0Y1_W2END[1] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
Xinput226 Tile_X0Y1_W2MID[4] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
Xinput204 Tile_X0Y1_NN4END[2] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2040_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q _0915_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q
+ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a21bo_1
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3991_ net198 net85 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2942_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 _0429_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q
+ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__mux2_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2873_ _0176_ _1696_ _1695_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__o211a_1
X_4612_ net1231 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4543_ net1259 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4474_ net1254 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3425_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q VGND VGND VPWR
+ VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3356_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q VGND VGND VPWR
+ VPWR _0051_ sky130_fd_sc_hd__inv_2
X_2307_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net1264 net192 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _1178_ sky130_fd_sc_hd__mux4_2
X_3287_ _2019_ _2016_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux2_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5026_ net1207 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2238_ _1094_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ _1039_ _1001_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and2b_1
XANTENNA_309 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput508 net508 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput519 net519 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[2] sky130_fd_sc_hd__buf_2
X_3210_ net980 net656 net1000 net995 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q VGND VGND VPWR VPWR
+ _1953_ sky130_fd_sc_hd__mux4_1
X_4190_ _0837_ _0836_ _0840_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 sky130_fd_sc_hd__o22a_4
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3141_ net993 _0214_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 _0228_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_78_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3072_ net93 net1044 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__mux2_1
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] net1059 VGND VGND VPWR VPWR _0639_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2925_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q _0554_ VGND
+ VGND VPWR VPWR _1740_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2856_ net1020 net1038 net1034 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1680_ sky130_fd_sc_hd__mux4_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2787_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q _1616_ VGND VGND
+ VPWR VPWR _1617_ sky130_fd_sc_hd__nor2_1
X_4526_ net1239 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4457_ net27 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3408_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q VGND VGND VPWR
+ VPWR _0103_ sky130_fd_sc_hd__inv_1
XFILLER_105_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4388_ net52 net1129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_105_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3339_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR
+ VPWR _0034_ sky130_fd_sc_hd__inv_1
XFILLER_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5009_ net170 net1085 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_106 net506 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_128 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer330 net948 VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__clkbuf_2
Xrebuffer341 net959 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer374 net1291 VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__clkbuf_2
Xrebuffer363 net1280 VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__clkbuf_2
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2710_ _1554_ _1523_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__and2_4
X_3690_ net1017 net1031 net982 net1042 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q VGND VGND VPWR VPWR
+ _0376_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_30_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2641_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q _1489_ VGND VGND
+ VPWR VPWR _1490_ sky130_fd_sc_hd__nand2b_1
Xoutput316 net316 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[0] sky130_fd_sc_hd__buf_2
Xoutput305 net305 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[29] sky130_fd_sc_hd__buf_2
X_2572_ Tile_X0Y1_DSP_bot.C5 net1063 VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__nor2_2
X_5360_ net134 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__buf_1
Xoutput327 net327 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput349 net349 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput338 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 VGND VGND VPWR VPWR
+ Tile_X0Y0_N1BEG[2] sky130_fd_sc_hd__buf_8
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4311_ net1251 net1147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5291_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_6
X_4242_ _0884_ _0885_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4173_ _0824_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q VGND VGND
+ VPWR VPWR _0825_ sky130_fd_sc_hd__or2_4
X_3124_ net1221 net215 net70 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q VGND VGND VPWR VPWR
+ _1889_ sky130_fd_sc_hd__mux4_1
X_3055_ net1057 net649 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q
+ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__mux2_4
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3957_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q _0623_ VGND VGND
+ VPWR VPWR _0624_ sky130_fd_sc_hd__and2b_1
X_2908_ net1020 net1038 net1034 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q VGND VGND VPWR VPWR
+ _1724_ sky130_fd_sc_hd__mux4_1
X_3888_ net76 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux2_1
X_2839_ net654 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q
+ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__mux2_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4509_ net1257 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5489_ net222 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer160 net778 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer171 net789 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer182 net800 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_123_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer193 Tile_X0Y1_DSP_bot.C1 VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4860_ net1198 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3811_ net1017 net823 net866 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0486_ sky130_fd_sc_hd__mux4_2
XANTENNA_39 net316 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 Tile_X0Y0_E6END[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 Tile_X0Y0_EE4END[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4791_ net1220 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3742_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 net19 net75 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux4_1
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3673_ _0357_ _0356_ _0358_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ _0086_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a221o_2
X_2624_ net191 net136 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q
+ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__mux2_1
X_5412_ net1210 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__buf_1
X_5343_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net426
+ sky130_fd_sc_hd__buf_6
X_2555_ _1407_ _1406_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__nand2_2
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5274_ Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_4
X_2486_ _0162_ _1343_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__nor2_1
XFILLER_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4225_ net175 net183 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0873_ sky130_fd_sc_hd__mux4_1
X_4156_ _0805_ _0807_ _0804_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o21bai_4
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3107_ net180 net1221 net195 net989 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A sky130_fd_sc_hd__mux4_1
X_4087_ _0744_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4
+ sky130_fd_sc_hd__inv_1
X_3038_ net1049 _0756_ _0788_ _1628_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q VGND VGND VPWR VPWR
+ _1823_ sky130_fd_sc_hd__mux4_1
XFILLER_102_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4989_ net1199 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 Tile_X0Y0_FrameData[19] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput26 Tile_X0Y0_EE4END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 Tile_X0Y0_E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput59 Tile_X0Y0_S1END[2] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_6
Xinput48 Tile_X0Y0_FrameData[30] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
X_2340_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q _1208_ VGND VGND
+ VPWR VPWR _1209_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_110_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2271_ _0998_ _1000_ _1140_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nor3_1
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4010_ net209 net2 net8 net1261 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0673_ sky130_fd_sc_hd__mux4_1
XFILLER_37_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4912_ net1188 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_45_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4843_ net1217 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_20_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4774_ net153 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3725_ _0406_ _0407_ _0056_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
XFILLER_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3656_ net629 VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__inv_6
X_2607_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__inv_2
X_3587_ _0277_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q _0269_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q VGND VGND VPWR VPWR
+ _0278_ sky130_fd_sc_hd__o211a_4
X_5326_ Tile_X0Y0_W6END[11] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_4
X_2538_ net1066 _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__nand2b_4
XFILLER_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5257_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR net349
+ sky130_fd_sc_hd__buf_6
XFILLER_87_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4208_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q _0856_ VGND VGND
+ VPWR VPWR _0857_ sky130_fd_sc_hd__or2_4
X_2469_ _1324_ _1325_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__or2_1
X_5188_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net271
+ sky130_fd_sc_hd__buf_1
X_4139_ net25 net79 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q VGND
+ VGND VPWR VPWR _0792_ sky130_fd_sc_hd__mux2_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout1113 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1102 net1106 VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__clkbuf_2
Xfanout1124 net1126 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__buf_2
Xfanout1135 net1136 VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__clkbuf_2
Xfanout1146 net1150 VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__clkbuf_2
Xfanout1157 net1158 VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__clkbuf_2
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1179 net1180 VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__buf_2
Xfanout1168 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__buf_2
XFILLER_19_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3510_ _0204_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q VGND VGND
+ VPWR VPWR _0205_ sky130_fd_sc_hd__or2_4
XFILLER_155_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4490_ net1234 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3441_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q VGND VGND VPWR
+ VPWR _0136_ sky130_fd_sc_hd__inv_1
XFILLER_143_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3372_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q VGND VGND VPWR
+ VPWR _0067_ sky130_fd_sc_hd__inv_2
X_2323_ _1192_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__inv_2
X_5111_ net1220 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5042_ net1190 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2254_ _0928_ net832 VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__nor2_8
X_2185_ _1054_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4826_ net1196 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4757_ net164 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4688_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0016_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3708_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q _0392_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q
+ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3639_ net99 net118 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q VGND
+ VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
XFILLER_108_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5309_ net105 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_2
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput216 Tile_X0Y1_W2END[2] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_2
Xinput227 Tile_X0Y1_W2MID[5] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput205 Tile_X0Y1_NN4END[3] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3990_ net113 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q
+ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux2_4
XFILLER_74_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2941_ net865 net670 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q
+ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__mux2_1
X_2872_ net85 net115 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__mux2_1
X_4611_ net1230 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4542_ net1258 net1087 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_116_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4473_ net1253 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3424_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR
+ VPWR _0119_ sky130_fd_sc_hd__inv_2
XFILLER_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3355_ net69 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
X_2306_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q _1176_ VGND VGND
+ VPWR VPWR _1177_ sky130_fd_sc_hd__nand2_1
X_3286_ _2017_ _2018_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__mux2_1
X_2237_ _0848_ _0878_ _1072_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__o21bai_1
X_5025_ net1205 net1077 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_127_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _1037_ _1038_ _1036_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__a21oi_4
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2099_ _0968_ _0966_ _0972_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4809_ net1215 net1134 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput509 net509 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[31] sky130_fd_sc_hd__buf_2
XFILLER_153_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3140_ net70 net81 net230 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_66_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3071_ _0041_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q
+ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_61_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3973_ _0621_ _0125_ _0625_ _0638_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A3 sky130_fd_sc_hd__a31o_4
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2924_ _1735_ _1732_ _1738_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q VGND VGND VPWR VPWR
+ _1739_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_75_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2855_ _0178_ _1676_ _1678_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4525_ net45 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2786_ net17 net109 net73 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q VGND VGND VPWR VPWR
+ _1616_ sky130_fd_sc_hd__mux4_2
X_4456_ net1249 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3407_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q VGND VGND VPWR
+ VPWR _0102_ sky130_fd_sc_hd__inv_1
X_4387_ net1230 net1129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_84_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3338_ net218 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3269_ _0823_ _0977_ _1497_ net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q VGND VGND VPWR VPWR
+ _2003_ sky130_fd_sc_hd__mux4_1
XFILLER_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5008_ net171 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_107 net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 Tile_X0Y1_FrameStrobe[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 Tile_X0Y1_N4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer331 net949 VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__clkbuf_2
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer364 net1281 VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__clkbuf_2
Xrebuffer375 net973 VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer342 net1276 VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2640_ net181 net126 net72 net233 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q VGND VGND VPWR VPWR
+ _1489_ sky130_fd_sc_hd__mux4_1
Xoutput317 net317 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput306 net306 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[2] sky130_fd_sc_hd__buf_2
X_2571_ _1421_ _0165_ _1423_ _1417_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C5 sky130_fd_sc_hd__a31o_1
Xoutput328 net328 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4310_ net1250 net1147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_99_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5290_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__buf_4
X_4241_ _0614_ _0880_ _0882_ _0879_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__o2bb2ai_1
X_4172_ net811 net664 net997 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0824_ sky130_fd_sc_hd__mux4_2
XFILLER_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3123_ _0183_ _1887_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q
+ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__o21a_1
X_3054_ _0181_ _1836_ _1833_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_38_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3956_ net187 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__mux2_1
X_2907_ _1723_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 sky130_fd_sc_hd__mux2_4
XFILLER_136_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3887_ _0052_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a21oi_2
X_2838_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q _0314_ _1662_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _1663_ sky130_fd_sc_hd__o211a_1
X_2769_ _1572_ _1599_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__nand2_1
X_4508_ net31 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5488_ net221 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__buf_1
X_4439_ net1251 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer150 net768 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_153_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer172 net790 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer161 net779 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer183 net801 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_150_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4790_ net1209 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3810_ _0481_ _0094_ _0483_ _0485_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0
+ sky130_fd_sc_hd__o22a_4
X_3741_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q _0418_ _0422_
+ _0397_ _0395_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ sky130_fd_sc_hd__o32a_4
XANTENNA_18 Tile_X0Y0_E6END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 Tile_X0Y0_EE4END[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _0357_ _0356_ _0358_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a22oi_4
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2623_ net632 VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__inv_2
X_5411_ net154 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__buf_1
X_2554_ _1132_ _1105_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__xor2_2
X_5273_ Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_4
X_2485_ net989 net1004 net864 net1008 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q VGND VGND VPWR VPWR
+ _1343_ sky130_fd_sc_hd__mux4_1
XFILLER_101_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4224_ _0869_ _0870_ _0871_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ _0138_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__a221o_1
X_4155_ _0617_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nand2_4
X_3106_ _1880_ _1879_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 sky130_fd_sc_hd__mux2_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4086_ _0733_ _0731_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q
+ _0738_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a32o_2
X_3037_ _1816_ _1822_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 sky130_fd_sc_hd__mux2_2
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4988_ net1198 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3939_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q _0606_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q
+ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput27 Tile_X0Y0_FrameData[0] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
Xinput16 Tile_X0Y0_E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_30_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput49 Tile_X0Y0_FrameData[31] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
Xinput38 Tile_X0Y0_FrameData[1] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XFILLER_155_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2270_ _0998_ _1000_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__o21a_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4911_ net1187 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4842_ net1216 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_290 _0554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4773_ net154 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3724_ net973 net970 net997 net990 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0407_ sky130_fd_sc_hd__mux4_1
XFILLER_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3655_ _0332_ _0318_ net640 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a21oi_4
XFILLER_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2606_ net187 net132 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net223
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q
+ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__mux4_2
X_3586_ _0273_ _0272_ _0276_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__o22a_1
X_5325_ Tile_X0Y0_W6END[10] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_4
X_2537_ Tile_X0Y1_DSP_bot.C7 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\] net1063 VGND
+ VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux2_4
XFILLER_114_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5256_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net348
+ sky130_fd_sc_hd__buf_2
X_2468_ _1324_ _1325_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__nor2_1
X_4207_ net811 net869 net997 net988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0856_ sky130_fd_sc_hd__mux4_2
X_5187_ Tile_X0Y0_EE4END[15] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
X_2399_ net176 net1224 net184 net129 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q VGND VGND VPWR VPWR
+ _1264_ sky130_fd_sc_hd__mux4_1
X_4138_ net104 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4069_ _0708_ _0709_ _0725_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__and3_1
XFILLER_83_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1103 net1104 VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__buf_2
Xfanout1114 net1115 VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__buf_2
Xfanout1147 net1150 VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1125 net1126 VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1136 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout1158 net1159 VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__buf_1
Xfanout1169 net1170 VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__buf_2
XFILLER_93_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ net202 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_1
X_3371_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR
+ VPWR _0066_ sky130_fd_sc_hd__inv_2
X_2322_ net26 net77 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q VGND
+ VGND VPWR VPWR _1192_ sky130_fd_sc_hd__mux2_1
XFILLER_111_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5110_ net1209 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5041_ net1189 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2253_ _1123_ _1120_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__and2b_1
X_2184_ net618 net832 VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4825_ net1194 net1132 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4756_ net167 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4687_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0015_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3707_ net177 net185 net122 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q VGND VGND VPWR VPWR
+ _0392_ sky130_fd_sc_hd__mux4_1
X_3638_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0327_ VGND VGND
+ VPWR VPWR _0328_ sky130_fd_sc_hd__or2_1
X_3569_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q _0260_ VGND VGND
+ VPWR VPWR _0261_ sky130_fd_sc_hd__and2b_1
X_5308_ net104 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_2
XFILLER_108_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput217 Tile_X0Y1_W2END[3] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_4
Xinput206 Tile_X0Y1_NN4END[4] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
X_5239_ Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
Xinput228 Tile_X0Y1_W2MID[6] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_2
XFILLER_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone1 net1060 _0529_ _0574_ _0575_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_67_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_Tile_X0Y1_UserCLK_regs clknet_0_Tile_X0Y1_UserCLK_regs VGND VGND VPWR
+ VPWR clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_104_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_113_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2940_ net187 net113 net198 net1028 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2871_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q _1694_ VGND VGND
+ VPWR VPWR _1695_ sky130_fd_sc_hd__or2_1
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4610_ net1229 net1174 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4541_ net1257 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4472_ net1252 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3423_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q VGND VGND VPWR
+ VPWR _0118_ sky130_fd_sc_hd__inv_2
X_3354_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q VGND VGND VPWR
+ VPWR _0049_ sky130_fd_sc_hd__inv_1
X_2305_ net1044 net1030 net1048 net1058 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q VGND VGND VPWR VPWR
+ _1176_ sky130_fd_sc_hd__mux4_1
X_3285_ net978 net990 net998 net994 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _2018_ sky130_fd_sc_hd__mux4_1
X_5024_ net1203 net1076 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2236_ _1091_ _1098_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_127_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _1034_ _1035_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__xor2_1
X_2098_ _0969_ _0144_ _0971_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_64_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4808_ net1214 net1134 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_154_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4739_ net1208 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q net626 VGND VGND
+ VPWR VPWR _1849_ sky130_fd_sc_hd__or2_1
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3972_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q _0637_ _0636_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q VGND VGND VPWR VPWR
+ _0638_ sky130_fd_sc_hd__o211a_1
XFILLER_50_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2923_ _1736_ _1737_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q
+ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__mux2_1
X_2854_ _1677_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__a21o_1
XFILLER_148_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2785_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q _1614_ VGND VGND
+ VPWR VPWR _1615_ sky130_fd_sc_hd__nand2_1
X_4524_ net46 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4455_ net1236 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_133_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3406_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR
+ VPWR _0101_ sky130_fd_sc_hd__inv_1
X_4386_ net1229 net1129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3337_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q VGND VGND VPWR
+ VPWR _0032_ sky130_fd_sc_hd__inv_2
X_3268_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q _1998_ _2002_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o21a_1
X_2219_ _1080_ _1070_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__xnor2_2
X_3199_ _1939_ _1942_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q
+ _1943_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3
+ sky130_fd_sc_hd__o22a_4
X_5007_ net1187 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_38_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_119 Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 net513 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer310 net946 VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__clkbuf_2
Xrebuffer332 net950 VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__clkbuf_2
XFILLER_154_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer365 net1282 VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__clkbuf_2
XFILLER_107_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_150_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput307 net307 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[30] sky130_fd_sc_hd__buf_2
X_2570_ _1422_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q VGND VGND
+ VPWR VPWR _1423_ sky130_fd_sc_hd__nand2b_1
Xoutput329 net329 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput318 net318 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4240_ _0884_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nand2b_1
XFILLER_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4171_ net189 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 net225
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__mux4_2
X_3122_ net993 net1022 net1003 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _1887_ sky130_fd_sc_hd__mux4_1
X_3053_ _1834_ _1835_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3955_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net223 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux2_1
X_2906_ _1375_ _1529_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__xor2_1
X_3886_ _0448_ _0446_ _0452_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a211o_4
X_2837_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__nand2_4
XFILLER_136_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2768_ net1068 Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\] _1597_ _1598_ VGND VGND VPWR
+ VPWR _1599_ sky130_fd_sc_hd__a22o_1
XFILLER_144_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2699_ _1544_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] net1068 VGND VGND VPWR VPWR
+ _1545_ sky130_fd_sc_hd__mux2_2
X_4507_ net1255 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5487_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net579
+ sky130_fd_sc_hd__buf_6
X_4438_ net1250 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4369_ net1243 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer50 net826 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_6
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer173 net791 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer162 net780 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer151 net769 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer184 net802 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_110_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3740_ _0112_ _0421_ _0420_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o211a_1
XANTENNA_19 Tile_X0Y0_EE4END[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3671_ net74 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q VGND
+ VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux2_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2622_ _1471_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q _1470_
+ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__a21oi_4
X_5410_ net153 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_1
X_5341_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net424
+ sky130_fd_sc_hd__clkbuf_2
X_2553_ _1405_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] net1066 VGND VGND VPWR VPWR
+ _1406_ sky130_fd_sc_hd__mux2_1
XFILLER_114_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_4
X_2484_ net974 net969 net978 net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q VGND VGND VPWR VPWR
+ _1342_ sky130_fd_sc_hd__mux4_1
X_4223_ net211 net1072 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__mux2_1
X_4154_ _0615_ _0616_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or2_1
X_4085_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q _0742_ VGND VGND
+ VPWR VPWR _0743_ sky130_fd_sc_hd__nor2_1
X_3105_ net866 net670 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__mux2_1
X_3036_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q _1821_ _1820_
+ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__o21ba_1
XFILLER_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4987_ net162 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3938_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__inv_2
X_3869_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q _0538_ _0540_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q VGND VGND VPWR VPWR
+ _0541_ sky130_fd_sc_hd__o211a_1
XFILLER_117_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 Tile_X0Y0_FrameData[10] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput17 Tile_X0Y0_E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
Xinput39 Tile_X0Y0_FrameData[20] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_6_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4910_ net173 net1111 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4841_ net1215 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_280 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _0554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4772_ net155 net1145 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3723_ net993 net1023 net1004 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q VGND VGND VPWR VPWR
+ _0406_ sky130_fd_sc_hd__mux4_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3654_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q _0341_ VGND VGND
+ VPWR VPWR _0342_ sky130_fd_sc_hd__and2b_1
XFILLER_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2605_ net131 net222 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux4_2
X_3585_ _0275_ _0274_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q
+ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
X_5324_ Tile_X0Y0_W6END[9] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_4
XFILLER_114_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2536_ _1385_ _0164_ _1390_ _1381_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C7 sky130_fd_sc_hd__a31o_1
X_5255_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 VGND VGND VPWR VPWR net347
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2467_ _1325_ _1324_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__nand2_4
X_4206_ _0852_ _0853_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__xnor2_1
X_5186_ Tile_X0Y0_EE4END[14] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
X_2398_ _0442_ _0344_ net75 net1073 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1263_ sky130_fd_sc_hd__mux4_2
X_4137_ _0789_ _0788_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux2_1
XFILLER_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4068_ net1059 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] _0724_ VGND VGND VPWR VPWR
+ _0726_ sky130_fd_sc_hd__a21oi_4
X_3019_ net1034 net984 net1043 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1806_ sky130_fd_sc_hd__mux4_1
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_154_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1104 net1105 VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__buf_1
Xfanout1115 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1126 net1132 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__clkbuf_2
Xoutput490 net490 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[14] sky130_fd_sc_hd__buf_2
Xfanout1137 net1138 VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__clkbuf_2
Xfanout1148 net1150 VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__buf_2
Xfanout1159 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__buf_2
XFILLER_59_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3370_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR
+ VPWR _0065_ sky130_fd_sc_hd__inv_1
X_2321_ net116 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__o211a_1
X_5040_ net1188 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2252_ _1110_ _1121_ _1122_ _1093_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__a22oi_2
X_2183_ _1044_ _1046_ _1005_ _1047_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__a22o_4
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4824_ net1193 net1127 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4755_ net1191 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3706_ _0388_ _0389_ _0390_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0087_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a221o_1
X_4686_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0014_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3637_ net21 net63 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q VGND
+ VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
X_3568_ net909 net970 net977 net987 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q VGND VGND VPWR VPWR
+ _0260_ sky130_fd_sc_hd__mux4_1
X_5307_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR net399
+ sky130_fd_sc_hd__buf_4
XFILLER_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2519_ _1371_ _1373_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__and2_4
XFILLER_124_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput218 Tile_X0Y1_W2END[4] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_4
Xinput207 Tile_X0Y1_NN4END[5] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_4
X_3499_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q VGND VGND VPWR
+ VPWR _0194_ sky130_fd_sc_hd__inv_1
X_5238_ Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
Xinput229 Tile_X0Y1_W2MID[7] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_4
X_5169_ Tile_X0Y0_E6END[7] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone2 net636 _0336_ _0339_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__o22a_4
XFILLER_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2870_ net57 net59 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q VGND
+ VGND VPWR VPWR _1694_ sky130_fd_sc_hd__mux2_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4540_ net1256 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4471_ net1251 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3422_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q VGND VGND VPWR
+ VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3353_ net189 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
X_2304_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q _1174_ VGND VGND
+ VPWR VPWR _1175_ sky130_fd_sc_hd__nand2b_1
X_3284_ net1224 net1073 net974 net969 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _2017_ sky130_fd_sc_hd__mux4_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5023_ net1201 net1077 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2235_ _1101_ _1100_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_127_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _1012_ _1031_ _1030_ _1013_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_88_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2097_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _0970_ VGND VGND
+ VPWR VPWR _0971_ sky130_fd_sc_hd__or2_1
XFILLER_65_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4807_ net1213 net1136 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2999_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q net1030 VGND
+ VGND VPWR VPWR _1789_ sky130_fd_sc_hd__nor2_1
X_4738_ net1207 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4669_ net1257 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3971_ net178 net69 net123 net235 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q VGND VGND VPWR VPWR
+ _0637_ sky130_fd_sc_hd__mux4_2
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2922_ net1054 net1048 net1029 net1014 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _1737_ sky130_fd_sc_hd__mux4_1
X_2853_ net57 net61 net59 net93 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q VGND VGND VPWR VPWR
+ _1677_ sky130_fd_sc_hd__mux4_2
X_2784_ net74 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q
+ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__mux2_1
XFILLER_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4523_ net1235 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4454_ net1233 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_133_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3405_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR
+ VPWR _0100_ sky130_fd_sc_hd__inv_2
X_4385_ net1228 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3336_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q VGND VGND VPWR
+ VPWR _0031_ sky130_fd_sc_hd__inv_2
X_3267_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q _1999_ _2000_
+ _2001_ _0195_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__a221o_1
X_5006_ net1186 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2218_ _1083_ _1084_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__xnor2_2
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3198_ net175 net120 _0563_ net995 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1943_ sky130_fd_sc_hd__mux4_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_109 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2149_ _0569_ _0567_ _0146_ _0541_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a211o_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer333 net951 VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__clkbuf_2
Xrebuffer366 net1283 VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__clkbuf_2
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_141_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput308 net308 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput319 net319 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4170_ _0821_ _0617_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__xnor2_4
XFILLER_96_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3121_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q _1885_ VGND VGND
+ VPWR VPWR _1886_ sky130_fd_sc_hd__or2_1
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3052_ net968 _0659_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3954_ _0618_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q _0620_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q VGND VGND VPWR VPWR
+ _0621_ sky130_fd_sc_hd__a211o_1
XFILLER_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2905_ _1722_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 sky130_fd_sc_hd__mux2_4
XFILLER_50_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3885_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q
+ _0555_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q VGND VGND VPWR
+ VPWR _0556_ sky130_fd_sc_hd__o211a_4
X_2836_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q _0744_ _1660_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q VGND VGND VPWR VPWR
+ _1661_ sky130_fd_sc_hd__o211a_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2767_ net1064 _0172_ net1068 VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2698_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\] net1064 VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__mux2_1
X_4506_ net1254 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5486_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net578
+ sky130_fd_sc_hd__buf_6
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4437_ net1248 net1113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_92_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ net1241 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3319_ net967 _1553_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__and2b_1
X_4299_ net1235 net1149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer51 _0225_ VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer152 net770 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer163 net781 VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer174 net792 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer185 net803 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3670_ _0070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q
+ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a21oi_2
X_2621_ net226 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__mux2_4
X_5340_ Tile_X0Y0_WW4END[15] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_4
X_2552_ Tile_X0Y1_DSP_bot.C6 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\] net1063 VGND
+ VGND VPWR VPWR _1405_ sky130_fd_sc_hd__mux2_1
X_5271_ Tile_X0Y1_N4END[15] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_1
XFILLER_126_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2483_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q _1333_ _1335_
+ _1341_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 sky130_fd_sc_hd__a31o_4
X_4222_ _0071_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_130_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4153_ _0787_ _0803_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__xnor2_1
X_4084_ _0101_ _0741_ _0740_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q
+ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__o211a_1
X_3104_ _1878_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__inv_1
X_3035_ net1047 net1030 net1014 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q VGND VGND VPWR VPWR
+ _1821_ sky130_fd_sc_hd__mux4_1
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4986_ net163 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3937_ net194 net89 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux2_1
X_3868_ _0091_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or2_1
X_2819_ _1643_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q _1645_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR VPWR
+ _1646_ sky130_fd_sc_hd__a211o_1
X_3799_ _0098_ _0473_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__o21a_1
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5469_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net567
+ sky130_fd_sc_hd__buf_4
XFILLER_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 Tile_X0Y0_E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xinput29 Tile_X0Y0_FrameData[11] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_270 Tile_X0Y0_W6END[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4840_ net1214 net1124 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_281 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_292 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4771_ net1208 net1144 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3722_ net205 net232 net84 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q VGND VGND VPWR VPWR
+ _0405_ sky130_fd_sc_hd__mux4_2
X_3653_ net1046 net968 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
XFILLER_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2604_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q _1454_ VGND VGND
+ VPWR VPWR _1455_ sky130_fd_sc_hd__or2_1
X_5323_ Tile_X0Y0_W6END[8] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_4
X_3584_ net177 net179 net124 net140 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0275_ sky130_fd_sc_hd__mux4_1
X_2535_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q _1386_ _1389_
+ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5254_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 VGND VGND VPWR VPWR net346
+ sky130_fd_sc_hd__clkbuf_1
X_2466_ _1137_ _1041_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__xor2_4
X_5185_ Tile_X0Y0_EE4END[13] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_1
X_4205_ _0852_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__or2_1
X_4136_ net15 net107 net71 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q VGND VGND VPWR VPWR
+ _0789_ sky130_fd_sc_hd__mux4_1
X_2397_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q _1261_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q
+ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__a21bo_1
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4067_ net1059 Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] _0724_ VGND VGND VPWR VPWR
+ _0725_ sky130_fd_sc_hd__a21o_1
XFILLER_83_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3018_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q _1804_ VGND
+ VGND VPWR VPWR _1805_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4969_ net150 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_138_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput480 net480 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_154_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout1138 net1139 VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout1105 net1106 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__clkbuf_2
Xfanout1116 net1119 VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__clkbuf_2
Xoutput491 net491 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[15] sky130_fd_sc_hd__buf_2
Xfanout1127 net1132 VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__buf_2
Xfanout1149 net1150 VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2320_ _0494_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q VGND VGND
+ VPWR VPWR _1190_ sky130_fd_sc_hd__nand2_4
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2251_ _1110_ _1121_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__xor2_1
X_2182_ _0799_ _0981_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__or2_4
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4823_ net1220 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4754_ net1190 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3705_ net211 net1072 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
X_4685_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0013_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3636_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q _0323_ _0325_
+ _0067_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o211a_1
X_3567_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q
+ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5306_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net398
+ sky130_fd_sc_hd__clkbuf_2
X_2518_ _1136_ _1372_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__nor2_1
X_5237_ Tile_X0Y1_FrameStrobe[13] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
X_3498_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q VGND VGND VPWR
+ VPWR _0193_ sky130_fd_sc_hd__inv_1
Xinput208 Tile_X0Y1_NN4END[6] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__buf_2
XFILLER_124_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput219 Tile_X0Y1_W2END[5] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlymetal6s2s_1
X_2449_ _0153_ _1308_ _1310_ _1304_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__a31o_1
X_5168_ Tile_X0Y0_E6END[6] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4119_ _0772_ _0773_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__mux2_1
X_5099_ net148 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_67_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone3 Tile_X0Y1_DSP_bot.A0 net1059 _0927_ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__o21ai_4
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4470_ net1250 net1103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3421_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR
+ VPWR _0116_ sky130_fd_sc_hd__inv_1
XPHY_EDGE_ROW_36_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3352_ net90 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_1
X_2303_ net1019 net1039 net1035 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1174_ sky130_fd_sc_hd__mux4_1
XFILLER_97_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3283_ _2013_ _2014_ _2015_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__o22a_1
X_2234_ _1103_ _1089_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__xnor2_2
X_5022_ net1200 net1077 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2165_ _1034_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_88_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone250 net1041 VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__buf_6
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2096_ net655 net971 net981 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0970_ sky130_fd_sc_hd__mux4_1
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4806_ net1212 net1136 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2998_ _1787_ _1788_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4737_ net1205 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4668_ net1256 net1157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3619_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND
+ VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
X_4599_ net36 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3970_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q _0633_ _0634_
+ _0635_ _0122_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a221o_1
X_2921_ net1036 net1032 net983 net1044 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _1736_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_61_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2852_ net626 net186 net1 net5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1676_ sky130_fd_sc_hd__mux4_1
XFILLER_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2783_ _0070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q
+ _1612_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4522_ net49 net1088 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_44_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4453_ net1232 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3404_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q VGND VGND VPWR
+ VPWR _0099_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4384_ net1227 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3335_ net223 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3266_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ _1082_ _1085_ _1068_ _1064_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__o211a_1
X_5005_ net1219 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_53_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3197_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q _1941_ VGND
+ VGND VPWR VPWR _1942_ sky130_fd_sc_hd__nand2_1
XFILLER_66_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2148_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q _1019_ VGND VGND
+ VPWR VPWR _1020_ sky130_fd_sc_hd__or2_1
X_2079_ _0952_ _0951_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__xnor2_2
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer301 _0413_ VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_32_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer334 net952 VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__clkbuf_2
Xrebuffer367 net1284 VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput309 net309 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[3] sky130_fd_sc_hd__buf_2
X_3120_ net869 net664 net830 net988 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q VGND VGND VPWR VPWR
+ _1885_ sky130_fd_sc_hd__mux4_1
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3051_ net669 _1204_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3953_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q _0619_ VGND VGND
+ VPWR VPWR _0620_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_46_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2904_ _1521_ _1519_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__xnor2_2
X_3884_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q _0554_ VGND VGND
+ VPWR VPWR _0555_ sky130_fd_sc_hd__nand2_1
X_2835_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6
+ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__nand2_1
X_2766_ net1064 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__or2_4
XFILLER_117_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4505_ net1253 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2697_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q _1534_ _1536_
+ _1543_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X
+ sky130_fd_sc_hd__a31o_1
X_5485_ net218 VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__buf_1
X_4436_ net1247 net1113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4367_ net1240 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3318_ net967 _1720_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__and2b_1
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4298_ net1234 net1149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3249_ net177 net1072 _0387_ net830 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q VGND VGND VPWR VPWR
+ _1986_ sky130_fd_sc_hd__mux4_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer30 _1537_ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_6
XFILLER_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer164 net782 VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer153 net771 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer186 net804 VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer175 net793 VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer197 _0405_ VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__buf_6
XFILLER_123_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2620_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q _1469_ VGND VGND
+ VPWR VPWR _1470_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2551_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q _1399_ _1401_
+ _1404_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C6 sky130_fd_sc_hd__a22o_1
X_5270_ Tile_X0Y1_N4END[14] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_1
X_2482_ _1337_ _1339_ _1340_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q
+ _0158_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__o221a_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4221_ _0561_ _0562_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q
+ _0556_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__a211o_1
XFILLER_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4152_ _0803_ _0787_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nor2_1
X_4083_ net66 net94 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q VGND
+ VGND VPWR VPWR _0741_ sky130_fd_sc_hd__mux2_1
X_3103_ _0494_ _0428_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q
+ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__mux2_1
X_3034_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _1817_ _1819_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q VGND VGND VPWR VPWR
+ _1820_ sky130_fd_sc_hd__o211a_1
X_4985_ net165 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3936_ net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q
+ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux2_1
X_3867_ net995 net1025 net1005 net1012 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0539_ sky130_fd_sc_hd__mux4_1
X_2818_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q _1644_ VGND VGND
+ VPWR VPWR _1645_ sky130_fd_sc_hd__and2b_1
X_3798_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0474_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__o21ba_1
X_2749_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1581_ VGND VGND
+ VPWR VPWR _1582_ sky130_fd_sc_hd__or2_1
X_5468_ Tile_X0Y0_SS4END[15] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__buf_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4419_ net1230 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5399_ net170 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkbuf_2
XFILLER_98_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 Tile_X0Y0_E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_40_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_260 net231 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_271 Tile_X0Y0_W6END[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_282 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_293 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4770_ net1207 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3721_ _0399_ _0401_ _0404_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 sky130_fd_sc_hd__o22a_4
X_3652_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q VGND VGND VPWR VPWR
+ _0340_ sky130_fd_sc_hd__mux4_2
X_2603_ net204 net124 net70 net215 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q VGND VGND VPWR VPWR
+ _1454_ sky130_fd_sc_hd__mux4_2
X_3583_ net70 net82 net215 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0274_ sky130_fd_sc_hd__mux4_1
X_5322_ Tile_X0Y0_W6END[7] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_4
X_2534_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q _1388_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__o21ai_1
X_5253_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 VGND VGND VPWR VPWR net345
+ sky130_fd_sc_hd__clkbuf_2
X_2465_ _1323_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] net1067 VGND VGND VPWR VPWR
+ _1324_ sky130_fd_sc_hd__mux2_4
X_5184_ Tile_X0Y0_EE4END[12] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_1
XFILLER_114_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4204_ _0785_ _0786_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__xnor2_1
X_2396_ net991 net1025 net1006 net1012 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1261_ sky130_fd_sc_hd__mux4_1
X_4135_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 net16 net72 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q VGND VGND VPWR VPWR
+ _0788_ sky130_fd_sc_hd__mux4_2
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4066_ net1059 Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__and2b_1
X_3017_ net1263 net96 net1019 net1038 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1804_ sky130_fd_sc_hd__mux4_1
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ net151 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_11_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4899_ net1208 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3919_ _0581_ _0583_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__a21oi_4
XFILLER_137_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput470 net470 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[10] sky130_fd_sc_hd__buf_2
XFILLER_154_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1106 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__buf_1
Xoutput481 net481 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput492 net492 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[16] sky130_fd_sc_hd__buf_2
Xfanout1117 net1118 VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__clkbuf_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1128 net1129 VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__clkbuf_2
Xfanout1139 net1141 VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ _0848_ _0981_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_2
X_2181_ _1043_ _1050_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__xnor2_2
XFILLER_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4822_ net1209 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4753_ net1189 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3704_ _0053_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q
+ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__a21oi_1
X_4684_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0012_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3635_ _0066_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3566_ _0255_ net834 _0256_ _0044_ _0045_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a221o_1
X_2517_ _1087_ _1134_ _1067_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a21oi_1
X_5305_ net101 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3497_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q VGND VGND VPWR
+ VPWR _0192_ sky130_fd_sc_hd__inv_1
X_5236_ net1158 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__buf_1
Xinput209 Tile_X0Y1_NN4END[7] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_4
X_2448_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1309_ VGND VGND
+ VPWR VPWR _1310_ sky130_fd_sc_hd__or2_1
XFILLER_102_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2379_ net59 net67 net93 net1226 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ _1246_ sky130_fd_sc_hd__mux4_1
X_5167_ Tile_X0Y0_E6END[5] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
X_4118_ net1262 net65 net101 net113 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0773_ sky130_fd_sc_hd__mux4_1
X_5098_ net1216 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4049_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] net1062 VGND VGND VPWR VPWR _0709_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_67_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3420_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q VGND VGND VPWR
+ VPWR _0115_ sky130_fd_sc_hd__inv_2
XFILLER_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3351_ net195 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_1
X_2302_ _0459_ _1171_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__xnor2_4
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3282_ net1023 net1004 net1011 net1008 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q VGND VGND VPWR VPWR
+ _2015_ sky130_fd_sc_hd__mux4_1
X_2233_ _1089_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__and2b_1
X_5021_ net1199 net1074 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2164_ _0994_ _0995_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_88_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2095_ net995 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 net1005 net653 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0969_ sky130_fd_sc_hd__mux4_2
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4805_ net1211 net1136 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2997_ net1047 _0756_ _0788_ _0293_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _1788_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4736_ net1203 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4667_ net1255 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3618_ _0306_ _0305_ _0307_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q VGND VGND VPWR VPWR
+ _0308_ sky130_fd_sc_hd__a221oi_4
X_4598_ net37 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3549_ net1 net5 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q VGND
+ VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
XFILLER_88_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5219_ net1239 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2920_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q _1734_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2851_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 net876 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q
+ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__mux2_1
X_2782_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__nor2_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4521_ net1260 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4452_ net1231 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3403_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q VGND VGND VPWR
+ VPWR _0098_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4383_ net1259 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3334_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q VGND VGND VPWR
+ VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_85_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3265_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q _1472_ VGND VGND
+ VPWR VPWR _2000_ sky130_fd_sc_hd__nand2_2
X_2216_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__inv_2
X_5004_ net1218 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_0_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3196_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q net634 _1940_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1941_ sky130_fd_sc_hd__a211o_1
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2147_ net205 net129 net75 net220 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q VGND VGND VPWR VPWR
+ _1019_ sky130_fd_sc_hd__mux4_2
X_2078_ _0822_ _0889_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer302 _1566_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_32_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4719_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer335 net953 VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__clkbuf_2
XFILLER_146_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer368 net1285 VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__clkbuf_2
XFILLER_107_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3050_ _1830_ _1831_ _1832_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q VGND VGND VPWR VPWR
+ _1833_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3952_ net186 net131 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2903_ _1721_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 sky130_fd_sc_hd__mux2_4
X_3883_ _0058_ _0059_ _0023_ _0537_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q VGND VGND VPWR VPWR
+ _0554_ sky130_fd_sc_hd__mux4_2
X_2834_ _1658_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q VGND VGND
+ VPWR VPWR _1659_ sky130_fd_sc_hd__nor2_4
X_4504_ net1252 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2765_ _0116_ _1588_ _1589_ _1596_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X
+ sky130_fd_sc_hd__a31o_1
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2696_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q _1537_ _1542_
+ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__o21ba_1
X_5484_ net217 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkbuf_2
X_4435_ net1246 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_104_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4366_ net1239 net1130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3317_ net967 _1569_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__and2b_1
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4297_ net1260 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3248_ _1982_ _1980_ _1985_ _0192_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3179_ _1925_ _1926_ _0187_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__mux2_1
Xrebuffer31 _1537_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_6
Xrebuffer53 _0439_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer154 net772 VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer165 net783 VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer176 net794 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer187 net805 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_112_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2550_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q _1403_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q
+ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__a21oi_1
X_2481_ net177 net185 net1223 net130 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q VGND VGND VPWR VPWR
+ _1340_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_81_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4220_ _0138_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_130_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4151_ _0802_ _0800_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__xnor2_2
X_3102_ _1877_ _1874_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux2_2
X_4082_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0739_ VGND VGND
+ VPWR VPWR _0740_ sky130_fd_sc_hd__or2_1
X_3033_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q _1818_ VGND
+ VGND VPWR VPWR _1819_ sky130_fd_sc_hd__nand2_2
XFILLER_48_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4984_ net166 net1083 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3935_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q _0215_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q
+ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3866_ net922 net971 net980 net1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR VPWR
+ _0538_ sky130_fd_sc_hd__mux4_1
X_3797_ net19 net111 net75 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q VGND VGND VPWR VPWR
+ _0474_ sky130_fd_sc_hd__mux4_2
X_2817_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 net13 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__mux2_2
X_2748_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q VGND
+ VGND VPWR VPWR _1581_ sky130_fd_sc_hd__mux2_1
XFILLER_117_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5467_ Tile_X0Y0_SS4END[14] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__buf_4
XFILLER_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4418_ net54 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2679_ _1448_ _1525_ _1447_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__o21a_4
X_5398_ net1190 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_4
XFILLER_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4349_ net1257 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_129_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_250 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_261 net234 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_272 net422 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_283 net538 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_294 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3720_ _0402_ _0403_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3651_ _0336_ _0334_ _0339_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 sky130_fd_sc_hd__o22a_4
X_2602_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q _1449_ _1452_
+ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__a21o_1
X_3582_ _0270_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q
+ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a21bo_1
X_5321_ Tile_X0Y0_W6END[6] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_4
X_2533_ _1387_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__inv_1
X_5252_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 VGND VGND VPWR VPWR net344
+ sky130_fd_sc_hd__clkbuf_1
X_2464_ Tile_X0Y1_DSP_bot.C9 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\] net1063 VGND
+ VGND VPWR VPWR _1323_ sky130_fd_sc_hd__mux2_4
X_5183_ Tile_X0Y0_EE4END[11] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
X_4203_ _0727_ _0849_ _0850_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__o2bb2a_1
X_2395_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q _1259_ VGND VGND
+ VPWR VPWR _1260_ sky130_fd_sc_hd__and2b_1
XFILLER_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4134_ _0728_ _0729_ _0785_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ _0723_ _0722_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A2 sky130_fd_sc_hd__mux2_4
X_3016_ _1802_ _1800_ _1803_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 sky130_fd_sc_hd__o22a_1
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4967_ net1213 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4898_ net1207 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3918_ _0584_ _0133_ _0586_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__o211a_4
XFILLER_137_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3849_ _0478_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__or2_4
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5519_ Tile_X0Y1_WW4END[14] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_150_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput460 net460 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[1] sky130_fd_sc_hd__buf_2
Xoutput471 net471 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_154_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1107 net1110 VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__clkbuf_2
Xoutput482 net482 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput493 net493 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[17] sky130_fd_sc_hd__buf_2
Xfanout1118 net1119 VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__buf_2
Xfanout1129 net1132 VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_155_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2180_ _1043_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__nand2_4
XFILLER_77_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4821_ net1195 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_16_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4752_ net1188 net1178 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_21_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4683_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0011_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3703_ _0360_ _0361_ _0386_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q
+ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a211o_1
X_3634_ net200 net7 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q VGND
+ VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
X_3565_ net639 _0255_ _0256_ _0044_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a22oi_4
X_5304_ net100 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_2
X_3496_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q VGND VGND VPWR
+ VPWR _0191_ sky130_fd_sc_hd__inv_1
X_2516_ _1370_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] net1066 VGND VGND VPWR VPWR
+ _1371_ sky130_fd_sc_hd__mux2_4
X_5235_ net1166 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_1
X_2447_ net174 net178 net119 net123 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q VGND VGND VPWR VPWR
+ _1309_ sky130_fd_sc_hd__mux4_1
X_2378_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q _1244_ VGND VGND
+ VPWR VPWR _1245_ sky130_fd_sc_hd__and2b_1
X_5166_ Tile_X0Y0_E6END[4] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4117_ net190 net198 net1264 net9 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0772_ sky130_fd_sc_hd__mux4_1
X_5097_ net1215 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
Xclone5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X
+ net1061 _0761_ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__o21ai_4
X_4048_ _0702_ _0707_ net1062 _0684_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_67_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_149_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_152_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput290 net290 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[15] sky130_fd_sc_hd__buf_2
XFILLER_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3350_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q VGND VGND VPWR
+ VPWR _0045_ sky130_fd_sc_hd__inv_2
X_2301_ _1171_ _0459_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__and2b_1
XFILLER_151_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5020_ net1198 net1075 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2011_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q
+ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__a21bo_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2232_ _1090_ _1099_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2163_ _0990_ _1008_ _1009_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_88_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone252 net972 VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__buf_6
X_2094_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q _0967_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q
+ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_64_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4804_ net1210 net1136 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2996_ net637 net59 net1264 net1034 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q VGND VGND VPWR VPWR
+ _1787_ sky130_fd_sc_hd__mux4_1
X_4735_ net1202 net1181 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_138_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4666_ net1254 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4597_ net1248 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3617_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q VGND
+ VGND VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_1
X_3548_ _0040_ net617 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3479_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q VGND VGND VPWR
+ VPWR _0174_ sky130_fd_sc_hd__inv_2
XFILLER_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5218_ net1240 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_2
XFILLER_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5149_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net241
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2850_ _1653_ _1671_ _1672_ _1669_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_122_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q _1610_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__o21ai_1
X_4520_ net1249 net1094 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4451_ net1230 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_7_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3402_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q VGND VGND VPWR
+ VPWR _0097_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ net1258 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3333_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q VGND VGND VPWR
+ VPWR _0028_ sky130_fd_sc_hd__inv_1
XFILLER_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3264_ _1400_ _0721_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q
+ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ _1068_ _1064_ _1082_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__a211oi_4
X_5003_ net148 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3195_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q net653 VGND
+ VGND VPWR VPWR _1940_ sky130_fd_sc_hd__nor2_1
XFILLER_26_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2146_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q _1014_ _1017_
+ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_144_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2077_ _0949_ _0945_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_24_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2979_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q _0571_ _1772_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q VGND VGND VPWR VPWR
+ _1773_ sky130_fd_sc_hd__a211oi_1
Xrebuffer303 net813 VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_32_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4718_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_101_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer336 net954 VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__clkbuf_2
XFILLER_135_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4649_ net1260 net1165 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
Xrebuffer369 net1286 VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__clkbuf_2
XFILLER_146_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_110_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3951_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 net819 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q
+ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux2_2
X_2902_ _1673_ _1671_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_46_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3882_ _0090_ _0549_ _0553_ _0545_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0
+ sky130_fd_sc_hd__a31o_4
X_2833_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR VPWR
+ _1658_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_135_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2764_ _1591_ _1594_ _1595_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q VGND VGND VPWR VPWR
+ _1596_ sky130_fd_sc_hd__o221a_1
X_4503_ net36 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2695_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q _1539_ _1541_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q VGND VGND VPWR VPWR
+ _1542_ sky130_fd_sc_hd__a31o_1
X_5483_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net575
+ sky130_fd_sc_hd__buf_1
X_4434_ net1245 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4365_ net1238 net1131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3316_ net967 _1568_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__and2b_1
X_4296_ net1249 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3247_ _1983_ _1984_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q
+ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__mux2_1
Xrebuffer21 net912 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_6
Xrebuffer10 net667 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd1_1
X_3178_ net1025 _0823_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__mux2_1
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer32 net648 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_2
X_2129_ _0999_ _0983_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__xor2_4
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer43 _0268_ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_37_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer155 net773 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_153_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer199 _0413_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__buf_6
Xrebuffer177 net795 VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer166 net784 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer188 net806 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2480_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q _1338_ _0157_
+ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__a21o_1
XFILLER_141_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4150_ _0801_ _0668_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_91_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3101_ _1875_ _1876_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q
+ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__mux2_1
X_4081_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q VGND
+ VGND VPWR VPWR _0739_ sky130_fd_sc_hd__mux2_1
X_3032_ net648 _1616_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__mux2_1
Xinput190 Tile_X0Y1_N2MID[4] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_34_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4983_ net1220 net1093 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3934_ _0589_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q _0590_
+ _0601_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q VGND VGND VPWR
+ VPWR _0602_ sky130_fd_sc_hd__a311o_1
X_3865_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR _0537_
+ sky130_fd_sc_hd__inv_2
X_2816_ net105 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q
+ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__mux2_4
X_3796_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 net76 net20 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q VGND VGND VPWR VPWR
+ _0473_ sky130_fd_sc_hd__mux4_2
X_2747_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q _1577_ _1579_
+ _0115_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__o211a_1
X_5466_ Tile_X0Y0_SS4END[13] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_4
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2678_ _1463_ _1464_ _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__o21ba_4
X_4417_ net55 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5397_ net1191 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_4
X_4348_ net1256 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4279_ net36 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_251 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_240 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_273 net435 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_284 net614 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_295 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3650_ _0337_ _0338_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q
+ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux2_1
X_2601_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q _1451_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__o21ai_1
X_3581_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q _0271_ VGND VGND
+ VPWR VPWR _0272_ sky130_fd_sc_hd__and2b_1
X_5320_ Tile_X0Y0_W6END[5] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_4
X_2532_ net187 net132 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__mux2_1
X_5251_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR net343
+ sky130_fd_sc_hd__clkbuf_2
X_4202_ _0727_ _0849_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2463_ _0150_ _1279_ _1298_ _1322_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C9 sky130_fd_sc_hd__o31a_1
X_5182_ Tile_X0Y0_EE4END[10] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
X_2394_ net922 net971 net981 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1259_ sky130_fd_sc_hd__mux4_1
X_4133_ _0729_ _0728_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__xnor2_4
XFILLER_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4064_ _0712_ net816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__mux2_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3015_ _0279_ net58 net2 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q VGND VGND VPWR VPWR
+ _1803_ sky130_fd_sc_hd__mux4_1
XFILLER_113_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4966_ net1212 net1092 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_149_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4897_ net1206 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3917_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q _0585_ VGND VGND
+ VPWR VPWR _0586_ sky130_fd_sc_hd__or2_1
XFILLER_149_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ net1060 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__o21ai_4
X_3779_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q _0292_ _0294_
+ _0457_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X
+ sky130_fd_sc_hd__a31o_1
XFILLER_105_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5518_ Tile_X0Y1_WW4END[13] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_150_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5449_ Tile_X0Y0_S4END[12] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__buf_1
Xoutput450 net450 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput461 net461 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[2] sky130_fd_sc_hd__buf_2
Xfanout1108 net1110 VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__buf_1
Xoutput483 net483 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput472 net472 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput494 net494 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[18] sky130_fd_sc_hd__buf_2
Xfanout1119 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4820_ net1192 net1133 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ net172 net1181 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4682_ clknet_2_3__leaf_Tile_X0Y1_UserCLK_regs _0010_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3702_ _0360_ _0361_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a21o_4
X_3633_ _0239_ net188 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
X_3564_ net193 net138 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_142_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5303_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR net395
+ sky130_fd_sc_hd__buf_1
X_3495_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q VGND VGND VPWR
+ VPWR _0190_ sky130_fd_sc_hd__inv_1
X_2515_ Tile_X0Y1_DSP_bot.C8 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\] net1065 VGND
+ VGND VPWR VPWR _1370_ sky130_fd_sc_hd__mux2_4
X_5234_ net1176 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
X_2446_ _1305_ _1306_ _1307_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0152_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__a221o_1
X_5165_ Tile_X0Y0_E6END[3] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
X_2377_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net1264 net192 net11 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _1244_ sky130_fd_sc_hd__mux4_1
XFILLER_110_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4116_ _0079_ _0770_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q
+ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__o21a_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5096_ net1214 net1162 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4047_ _0702_ _0707_ _0684_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X
+ sky130_fd_sc_hd__a21o_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4949_ net1195 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_130_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput280 net280 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_58_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput291 net291 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[16] sky130_fd_sc_hd__buf_2
XFILLER_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2300_ _1169_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__nand2_4
XFILLER_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3280_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q _2012_ VGND VGND
+ VPWR VPWR _2013_ sky130_fd_sc_hd__and2b_1
X_2231_ _1101_ _1100_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nand2b_1
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2162_ _1032_ _1011_ _1010_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__and3_4
X_2093_ net175 net183 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q VGND VGND VPWR VPWR
+ _0967_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_64_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4803_ net1208 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2995_ _1785_ _1783_ _1786_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 sky130_fd_sc_hd__o22a_1
X_4734_ net159 net1181 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_138_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4665_ net1253 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4596_ net1247 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3616_ _0054_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q
+ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3547_ _0217_ _0216_ _0229_ _0238_ net617 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a221o_1
XFILLER_142_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3478_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q VGND VGND VPWR
+ VPWR _0173_ sky130_fd_sc_hd__inv_1
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5217_ net1242 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_1
XFILLER_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2429_ _0155_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__or2_1
XFILLER_76_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5148_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net240
+ sky130_fd_sc_hd__buf_4
X_5079_ net1220 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2780_ net207 net66 net10 net102 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q VGND VGND VPWR VPWR
+ _1610_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4450_ net1229 net1112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3401_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q VGND VGND VPWR
+ VPWR _0096_ sky130_fd_sc_hd__inv_2
X_4381_ net1257 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3332_ net1 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3263_ net175 net211 _0563_ net864 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q VGND VGND VPWR VPWR
+ _1998_ sky130_fd_sc_hd__mux4_2
X_2214_ _1083_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__nor2_1
X_3194_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q _1400_ _1938_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q VGND VGND VPWR VPWR
+ _1939_ sky130_fd_sc_hd__o211a_1
X_5002_ net1216 net1082 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2145_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q _1016_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q
+ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o21ai_1
X_2076_ _0887_ _0888_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2978_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q net1030 VGND
+ VGND VPWR VPWR _1772_ sky130_fd_sc_hd__nor2_1
Xrebuffer304 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 VGND VGND VPWR VPWR net921
+ sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_32_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer337 net955 VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__clkbuf_2
X_4717_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C9 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\] sky130_fd_sc_hd__dfxtp_1
X_4648_ net1249 net1165 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4579_ net1230 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3950_ _0615_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__nand2_4
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2901_ _1720_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 sky130_fd_sc_hd__mux2_4
X_3881_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q _0552_ _0551_
+ _0089_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__a211o_1
X_2832_ _1657_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 sky130_fd_sc_hd__mux2_4
XFILLER_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2763_ net189 net8 net85 net100 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q VGND VGND VPWR VPWR
+ _1595_ sky130_fd_sc_hd__mux4_2
XFILLER_144_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4502_ net37 net1096 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2694_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q _1540_ VGND VGND
+ VPWR VPWR _1541_ sky130_fd_sc_hd__nand2_1
X_5482_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net574
+ sky130_fd_sc_hd__clkbuf_1
X_4433_ net1243 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4364_ net1237 net1131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3315_ net967 _1567_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__and2b_1
X_4295_ net1236 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3246_ _0977_ _1398_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__mux2_1
XFILLER_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer11 _0216_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd1_1
X_3177_ _0977_ _1436_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__mux2_1
X_2128_ _0983_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__nor2_1
Xrebuffer33 _0238_ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_37_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer44 _0268_ VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_2
Xrebuffer22 net820 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_6
X_2059_ _0930_ _0931_ _0932_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nand3_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer156 net774 VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_153_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer189 net807 VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer167 net785 VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer178 net796 VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_112_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3100_ net1032 net983 net1042 net1053 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q VGND VGND VPWR VPWR
+ _1876_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_8_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4080_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q _0737_ _0735_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q VGND VGND VPWR VPWR
+ _0738_ sky130_fd_sc_hd__a211o_1
X_3031_ _0571_ _0701_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q
+ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__mux2_1
Xinput180 Tile_X0Y1_N2END[2] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
Xinput191 Tile_X0Y1_N2MID[5] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_141_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4982_ net1209 net1093 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3933_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q _0599_ _0600_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q VGND VGND VPWR VPWR
+ _0601_ sky130_fd_sc_hd__a211oi_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3864_ _0532_ _0061_ _0534_ _0536_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__o22a_4
X_2815_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q _1638_ _1642_
+ _1634_ _1632_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__o32a_4
X_3795_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q _0471_ VGND VGND
+ VPWR VPWR _0472_ sky130_fd_sc_hd__or2_1
X_2746_ _0114_ _1578_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__or2_1
X_5465_ Tile_X0Y0_SS4END[12] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_4
XFILLER_117_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput610 net610 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[3] sky130_fd_sc_hd__buf_2
X_2677_ _1483_ _1523_ _1465_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__a21oi_4
X_4416_ net56 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5396_ net167 VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_1
X_4347_ net1255 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4278_ net37 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3229_ net213 net1000 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__mux2_1
XFILLER_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_252 net199 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_230 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_263 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_274 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_285 _0344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_296 net1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2600_ _1450_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__inv_2
X_3580_ net969 net978 net998 net989 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q VGND VGND VPWR VPWR
+ _0271_ sky130_fd_sc_hd__mux4_1
X_2531_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 net223 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q
+ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__mux2_1
X_5250_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR net342
+ sky130_fd_sc_hd__buf_1
X_4201_ _0640_ _0762_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__or2_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2462_ _1299_ _1300_ _1321_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q VGND VGND VPWR VPWR
+ _1322_ sky130_fd_sc_hd__a221o_1
X_5181_ Tile_X0Y0_EE4END[9] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_1
X_2393_ _1256_ _1254_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__xnor2_4
X_4132_ net622 _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__or2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4063_ _0721_ _0720_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q
+ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_4
X_3014_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q _1801_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q
+ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__a21bo_1
X_4965_ net1211 net1093 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3916_ net655 net971 net980 net1001 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0585_ sky130_fd_sc_hd__mux4_1
X_4896_ net1204 net1107 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3847_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] net1060 VGND VGND VPWR VPWR _0520_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3778_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q _0423_ _0456_
+ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__o21a_1
XFILLER_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2729_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 _1378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__mux2_4
X_5517_ Tile_X0Y1_WW4END[12] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_150_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5448_ Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__buf_1
Xoutput440 net440 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput451 net451 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput462 net462 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[3] sky130_fd_sc_hd__buf_2
X_5379_ Tile_X0Y1_EE4END[6] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
Xfanout1109 net1110 VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__clkbuf_2
Xoutput484 net484 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[9] sky130_fd_sc_hd__buf_2
Xoutput473 net473 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[13] sky130_fd_sc_hd__buf_4
Xoutput495 net495 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4750_ net1186 net1181 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3701_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q
+ _0385_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q VGND VGND VPWR
+ VPWR _0386_ sky130_fd_sc_hd__o211a_4
X_4681_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0009_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_78_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3632_ _0321_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q
+ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a21bo_1
X_5302_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR net394
+ sky130_fd_sc_hd__buf_1
X_3563_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q _0043_ _0044_
+ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a21oi_2
XFILLER_154_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3494_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q VGND VGND VPWR
+ VPWR _0189_ sky130_fd_sc_hd__inv_1
X_2514_ _0159_ _1331_ _1355_ _1357_ _1369_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C8
+ sky130_fd_sc_hd__o32a_4
X_5233_ net1081 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_2
X_2445_ net210 net1073 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q
+ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5164_ Tile_X0Y0_E6END[2] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_1
XFILLER_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ _1241_ _1242_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q
+ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__mux2_1
X_4115_ net1051 net1045 net1027 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0770_ sky130_fd_sc_hd__mux4_1
X_5095_ net1213 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4046_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q _0704_ _0706_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q VGND VGND VPWR VPWR
+ _0707_ sky130_fd_sc_hd__a31oi_1
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_96_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4948_ net1192 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4879_ net1187 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput270 net270 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput292 net292 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[17] sky130_fd_sc_hd__buf_2
Xoutput281 net281 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_58_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2230_ _1099_ _1090_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__xnor2_2
X_2161_ _1012_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_127_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2092_ _0143_ _0962_ _0963_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a31o_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2994_ _0279_ net94 net2 net1055 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q VGND VGND VPWR VPWR
+ _1786_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4802_ net1207 net1135 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4733_ net1199 net1180 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_99_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4664_ net1252 net1159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4595_ net1246 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_134_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3615_ net652 _0259_ _0278_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a211o_4
XFILLER_115_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3546_ _0216_ _0217_ net667 _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a22o_4
X_5216_ net1244 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_1
X_3477_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\] VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__inv_1
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2428_ _0442_ _0344_ net69 net210 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q VGND VGND VPWR VPWR
+ _1290_ sky130_fd_sc_hd__mux4_1
XFILLER_130_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2359_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\] net1064 VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__mux2_4
X_5147_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 VGND VGND VPWR VPWR net239
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5078_ net1209 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4029_ _0104_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__or2_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4380_ net1256 net1128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3400_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q VGND VGND VPWR
+ VPWR _0095_ sky130_fd_sc_hd__inv_2
X_3331_ net187 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_1
XTAP_TAPCELL_ROW_133_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3262_ _1992_ _1994_ _1997_ _0194_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2
+ sky130_fd_sc_hd__o22a_1
X_2213_ _1069_ _1081_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__xnor2_2
X_3193_ _0906_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q VGND
+ VGND VPWR VPWR _1938_ sky130_fd_sc_hd__nand2b_1
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5001_ net150 net1085 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2144_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__inv_1
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2075_ _0948_ _0946_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_24_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2977_ _1768_ _1771_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 sky130_fd_sc_hd__mux2_1
Xrebuffer305 net976 VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_32_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer338 net956 VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__clkbuf_2
X_4716_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C8 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\] sky130_fd_sc_hd__dfxtp_1
X_4647_ net1236 net1165 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_146_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4578_ net54 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3529_ net1221 net72 net217 net231 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0223_ sky130_fd_sc_hd__mux4_1
XFILLER_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2900_ _1719_ _1203_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__xnor2_2
XFILLER_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3880_ net98 net114 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q VGND
+ VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux2_1
X_2831_ _1627_ _1656_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2762_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q _1593_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__o21ai_1
XFILLER_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4501_ net39 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5481_ net214 VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__buf_1
X_4432_ net1241 net1115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2693_ net74 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q
+ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__mux2_1
XFILLER_132_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4363_ net1235 net1131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4294_ net1233 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3314_ net966 _1564_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__and2b_1
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3245_ net1024 _0823_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__mux2_1
XFILLER_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3176_ _0187_ _1923_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q
+ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__a21o_1
XFILLER_39_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer12 _0343_ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_6
X_2127_ _0996_ _0997_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__xnor2_2
Xrebuffer34 _0211_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_37_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer45 _0268_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_2
Xrebuffer23 _0342_ VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_6
X_2058_ _0708_ _0709_ _0847_ _0929_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__a31o_1
XFILLER_26_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer157 net775 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer168 net786 VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer179 net797 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3030_ _1814_ _1815_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q
+ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__mux2_1
Xinput181 Tile_X0Y1_N2END[3] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__buf_2
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput170 Tile_X0Y1_FrameData[6] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_2
Xinput192 Tile_X0Y1_N2MID[6] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_141_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4981_ net1195 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3932_ net186 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q VGND VGND
+ VPWR VPWR _0600_ sky130_fd_sc_hd__nor2_1
X_3863_ _0060_ _0535_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__a21o_1
X_2814_ _0119_ _1641_ _1640_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q
+ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__o211a_1
X_3794_ net209 net67 net11 net103 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q VGND VGND VPWR VPWR
+ _0471_ sky130_fd_sc_hd__mux4_2
X_2745_ net1263 net12 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__mux2_1
XFILLER_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5464_ Tile_X0Y0_SS4END[11] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_4
Xoutput611 net611 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput600 net600 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[9] sky130_fd_sc_hd__buf_2
X_2676_ _1522_ _1484_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__or2_4
X_4415_ net1259 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5395_ net164 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkbuf_1
X_4346_ net1254 net1137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4277_ net1248 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3228_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q _1968_ VGND
+ VGND VPWR VPWR _1969_ sky130_fd_sc_hd__and2b_1
X_3159_ net176 net1224 net1073 net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q VGND VGND VPWR VPWR
+ _1911_ sky130_fd_sc_hd__mux4_1
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_220 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_242 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_231 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_253 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_286 _0344_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_297 net1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2530_ _1383_ _1382_ _1384_ _0163_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q
+ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__a221o_1
XFILLER_114_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2461_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ _0148_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__mux2_1
XFILLER_114_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4200_ _0667_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__nor2_1
X_2392_ _1254_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__nand2_1
X_5180_ Tile_X0Y0_EE4END[8] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4131_ _0782_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nand2_8
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4062_ net182 net73 net141 net218 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q VGND VGND VPWR VPWR
+ _0721_ sky130_fd_sc_hd__mux4_2
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3013_ _1616_ _0764_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__mux2_4
XPHY_EDGE_ROW_134_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4964_ net1210 net1093 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3915_ net995 net1025 net1005 net653 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0584_ sky130_fd_sc_hd__mux4_2
X_4895_ net1201 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3846_ _0517_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q _0519_
+ _0497_ _0500_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X
+ sky130_fd_sc_hd__a32o_2
X_3777_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q _0455_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a21oi_1
X_2728_ net987 net1013 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q
+ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__mux2_4
X_5516_ Tile_X0Y1_WW4END[11] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_150_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5447_ Tile_X0Y0_S4END[10] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__buf_1
Xoutput430 net430 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput441 net441 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput452 net452 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[3] sky130_fd_sc_hd__buf_2
X_2659_ _1506_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__inv_1
XFILLER_154_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5378_ Tile_X0Y1_EE4END[5] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_1
Xoutput496 net496 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput474 net474 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput485 net485 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput463 net463 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[4] sky130_fd_sc_hd__buf_2
X_4329_ net1260 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q _0384_ VGND VGND
+ VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
X_4680_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs _0008_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3631_ net1052 net828 net1027 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q VGND VGND VPWR VPWR
+ _0321_ sky130_fd_sc_hd__mux4_2
X_3562_ _0243_ _0249_ _0253_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q
+ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a211o_1
X_5301_ net97 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_1
X_2513_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q _1368_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q
+ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__a21o_1
X_3493_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q VGND VGND VPWR
+ VPWR _0188_ sky130_fd_sc_hd__inv_1
X_5232_ net1088 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_1
X_2444_ _0050_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q
+ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__a21oi_1
X_2375_ net1043 net1030 net1047 net1015 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q VGND VGND VPWR VPWR
+ _1242_ sky130_fd_sc_hd__mux4_1
X_5163_ net20 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4114_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q _0768_ VGND VGND
+ VPWR VPWR _0769_ sky130_fd_sc_hd__or2_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5094_ net1212 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4045_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q _0705_ VGND VGND
+ VPWR VPWR _0706_ sky130_fd_sc_hd__nand2_1
XFILLER_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ net168 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4878_ net1186 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3829_ _0501_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q _0503_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q VGND VGND VPWR VPWR
+ _0504_ sky130_fd_sc_hd__o211a_1
Xoutput260 net260 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_133_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput271 net271 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput293 net293 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput282 net282 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[8] sky130_fd_sc_hd__buf_2
XFILLER_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone211 net1049 VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__buf_6
X_2160_ _1013_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2091_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q _0964_ _0144_
+ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21o_1
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2993_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q _1784_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4801_ net1206 net1136 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4732_ net161 net1180 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4663_ net1251 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_99_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3614_ _0065_ _0302_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__o21ai_4
X_4594_ net1245 net1175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3545_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q _0237_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q
+ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__o21a_4
X_3476_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\] VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_1
X_5215_ net1245 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
X_2427_ _1285_ _1283_ _1288_ _1289_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_149_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2358_ _0111_ _1218_ _1222_ _1225_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X
+ sky130_fd_sc_hd__a31o_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2289_ _1159_ _1158_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__xnor2_4
X_5077_ net1195 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4028_ net2 net10 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q VGND
+ VGND VPWR VPWR _0690_ sky130_fd_sc_hd__mux2_1
XFILLER_37_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3330_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q VGND VGND VPWR
+ VPWR _0025_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _1995_ _1996_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q
+ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__mux2_1
X_5000_ net1214 net1084 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2212_ _1077_ _1078_ _1079_ _1071_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__a22oi_2
X_3192_ _0190_ _1937_ _1936_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2
+ sky130_fd_sc_hd__o21a_1
Xfanout1260 net27 VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__buf_4
X_2143_ net126 net92 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q VGND
+ VGND VPWR VPWR _1015_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2074_ _0945_ _0947_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__nand2_2
XFILLER_93_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2976_ _1769_ _1770_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q
+ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__mux2_1
X_4715_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C7 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer339 net957 VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__clkbuf_2
Xrebuffer306 net922 VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd1_1
X_4646_ net1233 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4577_ net1228 net1081 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3528_ net175 net181 net197 net126 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0222_ sky130_fd_sc_hd__mux4_1
X_3459_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q VGND VGND VPWR
+ VPWR _0154_ sky130_fd_sc_hd__inv_2
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5129_ net1215 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_153_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2830_ _1653_ _1655_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__nand2_4
XFILLER_31_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2761_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2692_ _0070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q
+ _1538_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__a211o_1
X_4500_ net40 net1095 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5480_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net572
+ sky130_fd_sc_hd__clkbuf_2
X_4431_ net1240 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4362_ net1234 net1131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4293_ net1232 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3313_ net966 _1723_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__and2b_1
XFILLER_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3244_ _1981_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q
+ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__a21oi_2
Xfanout1090 net1091 VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__clkbuf_2
X_3175_ net176 net121 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q
+ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__mux2_1
X_2126_ _0996_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer13 net629 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer46 _0446_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer35 _0258_ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd1_1
X_2057_ _0726_ _0762_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2959_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q _0384_ _1762_
+ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer169 net787 VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer158 net776 VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd1_1
X_4629_ net39 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_112_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput171 Tile_X0Y1_FrameData[7] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xinput160 Tile_X0Y1_FrameData[26] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
Xinput182 Tile_X0Y1_N2END[4] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xinput193 Tile_X0Y1_N2MID[7] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_4
XFILLER_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4980_ net1192 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3931_ _0599_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__inv_2
X_3862_ net190 net9 net1264 net1262 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0535_ sky130_fd_sc_hd__mux4_1
X_2813_ net68 net1225 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q
+ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__mux2_1
X_3793_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q _0467_ _0469_
+ _0098_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a211o_1
X_2744_ net920 net193 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q
+ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__mux2_4
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5463_ Tile_X0Y0_SS4END[10] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__buf_4
Xoutput601 net601 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[0] sky130_fd_sc_hd__buf_2
X_2675_ _1520_ _1521_ _1504_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__o21a_1
X_4414_ net1258 net1120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput612 net612 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[5] sky130_fd_sc_hd__buf_2
X_5394_ net1209 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4345_ net1253 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4276_ net1247 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3227_ net177 net1223 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__mux2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3158_ net975 net816 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 _0405_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_54_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2109_ Tile_X0Y1_DSP_bot.B1 net1061 _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__o21ai_4
X_3089_ _0788_ _1204_ _0756_ net968 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q VGND VGND VPWR VPWR
+ _1866_ sky130_fd_sc_hd__mux4_2
XFILLER_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_210 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_232 net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_243 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 net243 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_254 net203 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_276 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_298 net1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_287 _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer4 _0359_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q _1320_ _1318_
+ _1314_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ sky130_fd_sc_hd__o31ai_4
X_2391_ _1255_ _1144_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__nor2_8
X_4130_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] net1060 VGND VGND VPWR VPWR _0783_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4061_ net195 net231 net1221 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q
+ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux4_2
X_3012_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q _1799_ VGND
+ VGND VPWR VPWR _1800_ sky130_fd_sc_hd__and2b_1
XFILLER_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4963_ net1208 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3914_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q _0582_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o21ba_1
X_4894_ net159 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3845_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q _0518_ VGND VGND
+ VPWR VPWR _0519_ sky130_fd_sc_hd__or2_1
XFILLER_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3776_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__inv_2
X_5515_ Tile_X0Y1_WW4END[10] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__buf_4
X_2727_ _1564_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 sky130_fd_sc_hd__mux2_4
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput420 net420 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[9] sky130_fd_sc_hd__buf_2
X_5446_ Tile_X0Y0_S4END[9] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__buf_1
Xoutput431 net431 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput442 net442 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput453 net453 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[4] sky130_fd_sc_hd__buf_2
X_2658_ net197 net126 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__mux2_1
XFILLER_120_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5377_ Tile_X0Y1_EE4END[4] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_1
Xoutput475 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR
+ Tile_X0Y1_EE4BEG[15] sky130_fd_sc_hd__buf_8
Xoutput464 net464 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput486 net486 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[10] sky130_fd_sc_hd__buf_2
X_2589_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q _1440_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q
+ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__a21oi_1
X_4328_ net1249 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput497 net497 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[20] sky130_fd_sc_hd__buf_2
X_4259_ _0890_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nor2_1
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_155_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3630_ _0067_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__and2_1
X_3561_ net825 _0249_ _0253_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__a21o_4
X_5300_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net392
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2512_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q VGND VGND VPWR VPWR
+ _1368_ sky130_fd_sc_hd__mux2_1
XFILLER_142_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3492_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q VGND VGND VPWR
+ VPWR _0187_ sky130_fd_sc_hd__inv_2
X_5231_ net1097 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_2
X_2443_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q _0442_ VGND VGND
+ VPWR VPWR _1305_ sky130_fd_sc_hd__or2_1
X_2374_ net1020 net1038 net1035 net985 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q VGND VGND VPWR VPWR
+ _1241_ sky130_fd_sc_hd__mux4_1
X_5162_ net19 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_1
X_4113_ net1017 net1037 net1031 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q VGND VGND VPWR VPWR
+ _0768_ sky130_fd_sc_hd__mux4_1
X_5093_ net1211 net1163 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4044_ net74 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q
+ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__mux2_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone9 net628 net821 net627 net650 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__a22o_1
XFILLER_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4946_ net169 net1100 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4877_ net1219 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3828_ _0063_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or2_4
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3759_ net868 net70 net14 net106 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q VGND VGND VPWR VPWR
+ _0439_ sky130_fd_sc_hd__mux4_2
Xoutput261 net261 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[3] sky130_fd_sc_hd__buf_2
Xoutput250 net250 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[2] sky130_fd_sc_hd__buf_2
X_5429_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 VGND VGND VPWR VPWR net521
+ sky130_fd_sc_hd__clkbuf_2
Xoutput294 net294 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput272 net272 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[13] sky130_fd_sc_hd__buf_8
Xoutput283 net283 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2090_ net74 net211 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q
+ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__mux2_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ net1204 net1136 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2992_ _1616_ _0796_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__mux2_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4731_ net1197 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4662_ net1250 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3613_ _0301_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q
+ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__o21a_1
X_4593_ net1244 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3544_ _0233_ _0231_ _0236_ _0035_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a22o_4
XFILLER_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3475_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q VGND VGND VPWR
+ VPWR _0170_ sky130_fd_sc_hd__inv_1
X_5214_ net1246 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_2
X_2426_ _0154_ _1286_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q
+ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_149_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5145_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net237
+ sky130_fd_sc_hd__clkbuf_2
X_2357_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q _1217_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q
+ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__o211a_1
X_2288_ _0903_ _0900_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__nor2_8
XFILLER_96_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5076_ net1192 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4027_ _0279_ net191 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__mux2_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4929_ net1205 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_10_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_156_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3260_ net666 _0864_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q
+ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__mux2_1
Xfanout1250 net37 VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__clkbuf_4
X_2211_ _1069_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__and2_1
X_3191_ net812 net666 _1497_ _1019_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q VGND VGND VPWR VPWR
+ _1937_ sky130_fd_sc_hd__mux4_1
Xfanout1261 net22 VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2142_ net234 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q
+ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2073_ _0936_ _0943_ _0944_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__or3_1
XFILLER_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2975_ _0756_ _1595_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__mux2_4
X_4714_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C6 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer307 net976 VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer329 net947 VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__clkbuf_2
XFILLER_147_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4645_ net1232 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4576_ net1227 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3527_ _0037_ _0220_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q
+ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__o21a_1
XFILLER_115_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3458_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q VGND VGND VPWR
+ VPWR _0153_ sky130_fd_sc_hd__inv_1
X_3389_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q VGND VGND VPWR
+ VPWR _0084_ sky130_fd_sc_hd__inv_1
X_2409_ net991 net1023 net996 net812 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q VGND VGND VPWR VPWR
+ _1273_ sky130_fd_sc_hd__mux4_2
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5128_ net1214 net1154 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5059_ net1208 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2760_ net200 net87 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q
+ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__mux2_1
XFILLER_144_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2691_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__nor2_1
XFILLER_144_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4430_ net1239 net1114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
XANTENNA_2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4361_ net1260 net1138 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4292_ net1231 net1182 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3312_ net928 _1563_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__and2b_1
XFILLER_112_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3243_ net1073 net979 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q
+ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__mux2_2
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout1080 net1081 VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__clkbuf_4
X_3174_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q _0344_ _1921_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q VGND VGND VPWR VPWR
+ _1922_ sky130_fd_sc_hd__o211a_1
Xfanout1091 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer25 net911 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__buf_6
X_2125_ _0946_ _0948_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer14 net630 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2056_ net620 _0709_ _0708_ _0849_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nand4b_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q VGND VGND VPWR VPWR
+ _1762_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4628_ net1247 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2889_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q _1707_ _1711_
+ _1701_ _1703_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ sky130_fd_sc_hd__o32a_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer159 net777 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer148 net766 VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_112_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4559_ net43 net1079 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput172 Tile_X0Y1_FrameData[8] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xinput150 Tile_X0Y1_FrameData[14] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
Xinput161 Tile_X0Y1_FrameData[27] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
Xinput194 Tile_X0Y1_N4END[0] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_2
Xinput183 Tile_X0Y1_N2END[5] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_2
X_3930_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q _0596_ _0598_
+ _0594_ _0592_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__o32a_4
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3861_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q _0533_ VGND VGND
+ VPWR VPWR _0534_ sky130_fd_sc_hd__and2_1
X_2812_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1639_ VGND VGND
+ VPWR VPWR _1640_ sky130_fd_sc_hd__or2_1
X_3792_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q _0468_ VGND VGND
+ VPWR VPWR _0469_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_42_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2743_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q _1575_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q
+ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__a21bo_1
X_5462_ Tile_X0Y0_SS4END[9] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__buf_4
Xoutput602 net602 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[10] sky130_fd_sc_hd__buf_2
X_2674_ _1503_ _1501_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__xnor2_4
X_4413_ net1257 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
X_5393_ net145 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__buf_1
Xoutput613 net613 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[6] sky130_fd_sc_hd__buf_2
X_4344_ net35 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4275_ net1246 net1185 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3226_ _1965_ _1966_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q
+ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__mux2_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3157_ _1909_ _1910_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 sky130_fd_sc_hd__mux2_1
X_2108_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] net1061 VGND VGND VPWR VPWR _0980_
+ sky130_fd_sc_hd__nand2b_1
X_3088_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q _1864_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q
+ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__a21oi_1
X_2039_ net1044 net1029 net1054 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q VGND VGND VPWR VPWR
+ _0915_ sky130_fd_sc_hd__mux4_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_200 net1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_222 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_233 net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 net292 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_277 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_244 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_255 net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_288 _0494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_299 net1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2390_ _1138_ _1143_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__nor2_4
XFILLER_95_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4060_ _0716_ _0714_ _0719_ _0129_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__a22o_1
X_3011_ net1057 net648 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__mux2_4
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4962_ net1207 net1091 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4893_ net160 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3913_ net175 net183 net120 net128 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0582_ sky130_fd_sc_hd__mux4_1
X_3844_ net186 net5 net61 net118 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q VGND VGND VPWR VPWR
+ _0518_ sky130_fd_sc_hd__mux4_2
X_3775_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 net76 net20 net112 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q VGND VGND VPWR VPWR
+ _0454_ sky130_fd_sc_hd__mux4_2
XFILLER_145_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5514_ Tile_X0Y1_WW4END[9] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__buf_4
X_2726_ _1329_ _1530_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__xnor2_2
Xoutput410 net410 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[10] sky130_fd_sc_hd__buf_8
X_5445_ Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__buf_1
X_2657_ net217 net619 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q
+ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__mux2_4
XFILLER_154_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput432 net432 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput421 net421 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput443 net443 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5376_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 VGND VGND VPWR VPWR net459
+ sky130_fd_sc_hd__clkbuf_2
Xoutput476 net476 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput454 net454 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput465 net465 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput487 net487 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[11] sky130_fd_sc_hd__buf_2
X_2588_ _1439_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__inv_2
X_4327_ net47 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput498 net498 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[21] sky130_fd_sc_hd__buf_2
XFILLER_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4258_ _0901_ _0902_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__xnor2_2
X_3209_ net1224 net212 net924 net971 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q VGND VGND VPWR VPWR
+ _1952_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4189_ _0838_ _0839_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q
+ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__mux2_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3560_ _0042_ _0250_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q
+ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_47_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ _1365_ _0161_ _1367_ _1361_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__a31o_4
X_5230_ net1105 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_2
X_3491_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q VGND VGND VPWR
+ VPWR _0186_ sky130_fd_sc_hd__inv_1
XFILLER_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2442_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q _1301_ _1303_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q VGND VGND VPWR VPWR
+ _1304_ sky130_fd_sc_hd__o211a_1
X_2373_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 net19 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q
+ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux2_4
X_5161_ net18 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_1
X_5092_ net155 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4112_ _0068_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q
+ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__a21oi_1
X_4043_ _0070_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q
+ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__a211o_1
XFILLER_56_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4945_ net1189 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4876_ net1218 net1119 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3827_ net1051 net1046 net1027 net1056 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0502_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3758_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or2_1
X_2709_ _1484_ _1522_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__nand2_2
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3689_ _0365_ _0371_ _0375_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2
+ sky130_fd_sc_hd__a21o_1
Xoutput262 net262 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput251 net251 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput240 net240 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[0] sky130_fd_sc_hd__buf_2
X_5428_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net520
+ sky130_fd_sc_hd__buf_1
Xoutput284 net284 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput295 net295 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[1] sky130_fd_sc_hd__buf_2
Xoutput273 net273 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5359_ net133 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone213 net999 VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__clkbuf_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2991_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q _1782_ VGND VGND
+ VPWR VPWR _1783_ sky130_fd_sc_hd__and2b_1
X_4730_ net1196 net1179 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4661_ net1248 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3612_ net1051 net828 net1026 net1016 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0302_ sky130_fd_sc_hd__mux4_2
X_4592_ net1242 net1176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3543_ _0234_ _0235_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q
+ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
XFILLER_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3474_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q VGND VGND VPWR
+ VPWR _0169_ sky130_fd_sc_hd__inv_1
X_5213_ net40 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
X_2425_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q _1287_ VGND VGND
+ VPWR VPWR _1288_ sky130_fd_sc_hd__or2_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5144_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net236
+ sky130_fd_sc_hd__buf_2
X_2356_ _1205_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q _1223_
+ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a21o_1
XFILLER_56_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2287_ _1157_ _1156_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__and2_4
X_5075_ net1191 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4026_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q _0687_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a21bo_1
XFILLER_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4928_ net1203 net1099 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4859_ net1197 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ _1070_ _1080_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__and2b_1
Xfanout1240 net43 VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__buf_2
X_3190_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q _1933_ _1935_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q VGND VGND VPWR VPWR
+ _1936_ sky130_fd_sc_hd__a211o_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout1251 net36 VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__clkbuf_4
Xfanout1262 net21 VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__clkbuf_4
X_2141_ _0955_ _1005_ _1006_ _1004_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2072_ _0881_ _0939_ _0941_ _0938_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2974_ net1047 _0788_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__mux2_4
X_4713_ clknet_2_1__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C5 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer308 net975 VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd1_1
X_4644_ net1231 net1164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4575_ net1259 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3526_ net993 net1021 net1003 net1007 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q VGND VGND VPWR VPWR
+ _0220_ sky130_fd_sc_hd__mux4_1
XFILLER_115_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3457_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q VGND VGND VPWR
+ VPWR _0152_ sky130_fd_sc_hd__inv_2
X_3388_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q VGND VGND VPWR
+ VPWR _0083_ sky130_fd_sc_hd__inv_1
X_2408_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q _1271_ VGND VGND
+ VPWR VPWR _1272_ sky130_fd_sc_hd__nor2_1
X_2339_ net1019 net1038 net1034 net984 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q VGND VGND VPWR VPWR
+ _1208_ sky130_fd_sc_hd__mux4_1
X_5127_ net1213 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5058_ net1207 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4009_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q _0671_ VGND VGND
+ VPWR VPWR _0672_ sky130_fd_sc_hd__nand2_1
XFILLER_25_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 net109 net73 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q
+ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__mux4_2
XANTENNA_3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_4360_ net1249 net1138 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_20_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3311_ net928 _1562_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__and2b_1
X_4291_ net53 net1185 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_140_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3242_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q net631 _1979_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q VGND VGND VPWR VPWR
+ _1980_ sky130_fd_sc_hd__a211o_1
X_3173_ net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q VGND
+ VGND VPWR VPWR _1921_ sky130_fd_sc_hd__nand2b_1
X_2124_ _0994_ _0995_ _0993_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__o21ai_2
Xfanout1081 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__buf_2
Xfanout1092 net1093 VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__buf_2
Xfanout1070 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q VGND VGND
+ VPWR VPWR net1070 sky130_fd_sc_hd__clkbuf_4
Xrebuffer15 _1472_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__buf_6
Xrebuffer37 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 VGND VGND VPWR VPWR
+ net654 sky130_fd_sc_hd__dlygate4sd1_1
X_2055_ net620 _0667_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__nor2_1
XFILLER_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer48 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 VGND VGND VPWR VPWR
+ net665 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer59 net765 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_37_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2957_ net1053 net641 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 _0317_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 sky130_fd_sc_hd__mux4_2
X_2888_ _0174_ _1710_ _1709_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q
+ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__o211a_1
X_4627_ net1246 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer149 net767 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd1_1
X_4558_ net44 net1079 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3509_ net1018 net1033 net982 net1040 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q VGND VGND VPWR VPWR
+ _0204_ sky130_fd_sc_hd__mux4_2
X_4489_ net1260 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput140 Tile_X0Y1_E6END[1] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_1
Xinput151 Tile_X0Y1_FrameData[15] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xinput162 Tile_X0Y1_FrameData[28] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_4
Xinput195 Tile_X0Y1_N4END[1] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
Xinput184 Tile_X0Y1_N2END[6] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_2
XFILLER_36_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput173 Tile_X0Y1_FrameData[9] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3860_ net65 net101 net77 net117 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q VGND VGND VPWR VPWR
+ _0533_ sky130_fd_sc_hd__mux4_1
X_2811_ net58 net60 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q VGND
+ VGND VPWR VPWR _1639_ sky130_fd_sc_hd__mux2_1
X_3791_ net8 net88 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q VGND
+ VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ net1042 net1029 net1054 net669 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q VGND VGND VPWR VPWR
+ _1575_ sky130_fd_sc_hd__mux4_2
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5461_ Tile_X0Y0_SS4END[8] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__buf_4
X_4412_ net1256 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2673_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput614 net614 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput603 net603 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[11] sky130_fd_sc_hd__buf_2
X_4343_ net1251 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4274_ net42 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3225_ _0875_ _1454_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__mux2_1
X_3156_ net665 _1378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q
+ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__mux2_1
X_3087_ _1863_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__inv_1
XFILLER_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2107_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q _0961_ _0979_
+ _0976_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B1 sky130_fd_sc_hd__a22o_4
X_2038_ _0118_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__and2_1
XFILLER_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3989_ _0074_ _0649_ _0653_ _0645_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2
+ sky130_fd_sc_hd__a31o_1
XFILLER_148_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_212 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_201 net1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_223 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_234 net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 net330 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_256 net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_289 _0554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_278 net488 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3010_ _0180_ _1798_ _1797_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2
+ sky130_fd_sc_hd__o21a_1
XFILLER_67_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_103_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4961_ net1205 net1090 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4892_ net161 net1109 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3912_ _0578_ _0577_ _0132_ _0580_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a31o_4
X_3843_ _0513_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q _0516_
+ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK VGND VGND VPWR VPWR clknet_0_Tile_X0Y1_UserCLK
+ sky130_fd_sc_hd__clkbuf_16
X_3774_ _0453_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7
+ sky130_fd_sc_hd__inv_2
X_5513_ Tile_X0Y1_WW4END[8] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_4
X_2725_ _1563_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] net1070 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 sky130_fd_sc_hd__mux2_4
Xoutput411 net411 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[11] sky130_fd_sc_hd__buf_6
Xoutput400 net400 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[7] sky130_fd_sc_hd__buf_2
X_2656_ _1501_ _1503_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__or2_1
X_5444_ net876 VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_6
Xoutput422 net422 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput433 net433 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput444 net444 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput477 net477 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput455 net455 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput466 net466 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[7] sky130_fd_sc_hd__buf_2
X_5375_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net458
+ sky130_fd_sc_hd__clkbuf_1
X_2587_ net193 net138 net874 net229 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q VGND VGND VPWR VPWR
+ _1439_ sky130_fd_sc_hd__mux4_1
X_4326_ net50 net1148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q
+ sky130_fd_sc_hd__dlxtp_1
Xoutput488 net488 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput499 net499 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[22] sky130_fd_sc_hd__buf_2
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4257_ _0901_ _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nor2_2
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4188_ net1222 net73 net218 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q VGND VGND VPWR VPWR
+ _0839_ sky130_fd_sc_hd__mux4_1
X_3208_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q _1946_ _1948_
+ _1951_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3139_ net69 net84 net231 net980 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3490_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q VGND VGND VPWR
+ VPWR _0185_ sky130_fd_sc_hd__inv_2
X_2510_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q _1366_ VGND VGND
+ VPWR VPWR _1367_ sky130_fd_sc_hd__or2_1
XFILLER_154_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2441_ _0152_ _1302_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__or2_1
X_2372_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q _1238_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q
+ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__o21a_1
X_5160_ net17 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_1
X_5091_ net157 net1160 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4111_ _0391_ _0393_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q
+ _0298_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__a211o_1
X_4042_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5
+ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__nor2_1
XFILLER_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4944_ net1188 net1098 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_24_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4875_ net1217 net1116 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_50_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3826_ net1017 net866 net865 net1041 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q VGND VGND VPWR VPWR
+ _0501_ sky130_fd_sc_hd__mux4_2
X_3757_ _0433_ _0024_ _0435_ _0437_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3
+ sky130_fd_sc_hd__o22a_4
X_2708_ _1553_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] net1071 VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 sky130_fd_sc_hd__mux2_4
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3688_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q _0374_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q
+ _0373_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__o211a_1
XFILLER_145_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput252 net252 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput241 net241 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[1] sky130_fd_sc_hd__buf_2
X_5427_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net519
+ sky130_fd_sc_hd__buf_1
X_2639_ _0170_ _1485_ _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__o21ai_1
Xoutput285 net285 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput263 net263 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[15] sky130_fd_sc_hd__buf_8
X_5358_ net132 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput296 net296 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[20] sky130_fd_sc_hd__buf_2
XFILLER_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4309_ net39 net1149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5289_ Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_4
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_151_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone214 net1001 VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__buf_6
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone247 net996 VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2990_ net1057 net648 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q
+ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__mux2_4
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4660_ net1247 net1156 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3611_ net1017 net1037 net866 net865 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q VGND VGND VPWR VPWR
+ _0301_ sky130_fd_sc_hd__mux4_2
X_4591_ net43 net1177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_115_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3542_ net73 net81 net218 net230 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q VGND VGND VPWR VPWR
+ _0235_ sky130_fd_sc_hd__mux4_1
X_3473_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\] VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_1
XFILLER_142_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5212_ net1248 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_2
X_2424_ net974 net969 net978 net998 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q VGND VGND VPWR VPWR
+ _1287_ sky130_fd_sc_hd__mux4_1
X_2355_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q _1207_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q
+ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__o21ai_1
X_5143_ net145 net1155 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2286_ _0896_ _1155_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__or2_1
X_5074_ net1190 net1169 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4025_ net1053 net1048 net1028 net1058 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q VGND VGND VPWR VPWR
+ _0687_ sky130_fd_sc_hd__mux4_1
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4927_ net1201 net1101 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4858_ net1196 net1117 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_10_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3809_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q _0484_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21o_1
X_4789_ net1195 net1143 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_115_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1241 net1242 VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__buf_4
Xfanout1230 net53 VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__buf_4
Xfanout1263 net4 VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__clkbuf_4
Xfanout1252 net35 VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__buf_4
X_2140_ net618 _0981_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__or2_1
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2071_ _0936_ _0943_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__o21ai_4
XFILLER_38_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2973_ net637 net1264 net1226 net1034 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q VGND VGND VPWR VPWR
+ _1768_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_103_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4712_ clknet_2_0__leaf_Tile_X0Y1_UserCLK_regs Tile_X0Y1_DSP_bot.C4 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer309 net925 VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd1_1
X_4643_ net1230 net1168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4574_ net1258 net1080 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3525_ _0218_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q VGND VGND
+ VPWR VPWR _0219_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3456_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q VGND VGND VPWR
+ VPWR _0151_ sky130_fd_sc_hd__inv_1
X_3387_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q VGND VGND VPWR
+ VPWR _0082_ sky130_fd_sc_hd__inv_1
X_2407_ net174 net178 net119 net123 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q VGND VGND VPWR VPWR
+ _1271_ sky130_fd_sc_hd__mux4_1
X_2338_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__inv_2
X_5126_ net1212 net1151 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2269_ _0951_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__nor2_2
X_5057_ net1205 net1171 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4008_ net1052 net1046 net1027 net1057 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q
+ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q VGND VGND VPWR VPWR
+ _0671_ sky130_fd_sc_hd__mux4_1
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3310_ net928 _1561_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__and2b_1
XFILLER_152_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4290_ net1229 net1183 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_98_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3241_ net176 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q VGND VGND
+ VPWR VPWR _1979_ sky130_fd_sc_hd__nor2_1
X_3172_ _1919_ _1920_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A sky130_fd_sc_hd__mux2_1
X_2123_ _0959_ _0982_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__xnor2_1
Xfanout1071 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q VGND VGND
+ VPWR VPWR net1071 sky130_fd_sc_hd__clkbuf_4
Xfanout1060 Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q VGND VGND
+ VPWR VPWR net1060 sky130_fd_sc_hd__buf_2
Xfanout1082 net1085 VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__buf_2
Xrebuffer16 net632 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd1_1
Xfanout1093 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__clkbuf_2
X_2054_ Tile_X0Y1_DSP_bot.A0 net1059 _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__o21ai_4
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2956_ _1759_ _1761_ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__nand2_1
X_2887_ net93 net1226 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q
+ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__mux2_1
X_4626_ net1245 net1166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4557_ net1238 net1079 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3508_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q _0202_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q
+ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a21bo_1
XFILLER_89_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4488_ net1249 net1102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q
+ sky130_fd_sc_hd__dlxtp_1
X_3439_ net214 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5109_ net1195 net1161 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_123_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_149_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput130 Tile_X0Y1_E2END[7] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
Xinput141 Tile_X0Y1_EE4END[0] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xinput152 Tile_X0Y1_FrameData[16] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_2
Xinput163 Tile_X0Y1_FrameData[29] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_4
Xinput196 Tile_X0Y1_N4END[2] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
Xinput185 Tile_X0Y1_N2END[7] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_4
Xinput174 Tile_X0Y1_N1END[0] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2810_ Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q _1635_ _1637_
+ _0120_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__o211a_1
X_3790_ net117 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q
+ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _0115_ _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__and2_1
X_5460_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net543
+ sky130_fd_sc_hd__clkbuf_1
X_4411_ net1255 net1123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q
+ sky130_fd_sc_hd__dlxtp_1
X_2672_ net829 _1518_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_152_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput615 net615 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput604 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR
+ Tile_X0Y1_WW4BEG[12] sky130_fd_sc_hd__buf_6
X_5391_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net474
+ sky130_fd_sc_hd__clkbuf_2
X_4342_ net1250 net1140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q
+ sky130_fd_sc_hd__dlxtp_1
X_4273_ net1243 net1184 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_86_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3224_ net1005 _0712_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q
+ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__mux2_1
.ends

