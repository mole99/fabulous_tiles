VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IHP_SRAM
  CLASS BLOCK ;
  FOREIGN IHP_SRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 108.000 BY 483.840 ;
  PIN ADDR_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 102.700 108.000 103.100 ;
    END
  END ADDR_SRAM0
  PIN ADDR_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 105.220 108.000 105.620 ;
    END
  END ADDR_SRAM1
  PIN ADDR_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 107.740 108.000 108.140 ;
    END
  END ADDR_SRAM2
  PIN ADDR_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 110.260 108.000 110.660 ;
    END
  END ADDR_SRAM3
  PIN ADDR_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 112.780 108.000 113.180 ;
    END
  END ADDR_SRAM4
  PIN ADDR_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 115.300 108.000 115.700 ;
    END
  END ADDR_SRAM5
  PIN ADDR_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 117.820 108.000 118.220 ;
    END
  END ADDR_SRAM6
  PIN ADDR_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 120.340 108.000 120.740 ;
    END
  END ADDR_SRAM7
  PIN ADDR_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 122.860 108.000 123.260 ;
    END
  END ADDR_SRAM8
  PIN ADDR_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 125.380 108.000 125.780 ;
    END
  END ADDR_SRAM9
  PIN BM_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 127.900 108.000 128.300 ;
    END
  END BM_SRAM0
  PIN BM_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 130.420 108.000 130.820 ;
    END
  END BM_SRAM1
  PIN BM_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 153.100 108.000 153.500 ;
    END
  END BM_SRAM10
  PIN BM_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 155.620 108.000 156.020 ;
    END
  END BM_SRAM11
  PIN BM_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 158.140 108.000 158.540 ;
    END
  END BM_SRAM12
  PIN BM_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 160.660 108.000 161.060 ;
    END
  END BM_SRAM13
  PIN BM_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 163.180 108.000 163.580 ;
    END
  END BM_SRAM14
  PIN BM_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 165.700 108.000 166.100 ;
    END
  END BM_SRAM15
  PIN BM_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 168.220 108.000 168.620 ;
    END
  END BM_SRAM16
  PIN BM_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 170.740 108.000 171.140 ;
    END
  END BM_SRAM17
  PIN BM_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 173.260 108.000 173.660 ;
    END
  END BM_SRAM18
  PIN BM_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 175.780 108.000 176.180 ;
    END
  END BM_SRAM19
  PIN BM_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 132.940 108.000 133.340 ;
    END
  END BM_SRAM2
  PIN BM_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 178.300 108.000 178.700 ;
    END
  END BM_SRAM20
  PIN BM_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 180.820 108.000 181.220 ;
    END
  END BM_SRAM21
  PIN BM_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 183.340 108.000 183.740 ;
    END
  END BM_SRAM22
  PIN BM_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 185.860 108.000 186.260 ;
    END
  END BM_SRAM23
  PIN BM_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 188.380 108.000 188.780 ;
    END
  END BM_SRAM24
  PIN BM_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 190.900 108.000 191.300 ;
    END
  END BM_SRAM25
  PIN BM_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 193.420 108.000 193.820 ;
    END
  END BM_SRAM26
  PIN BM_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 195.940 108.000 196.340 ;
    END
  END BM_SRAM27
  PIN BM_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 198.460 108.000 198.860 ;
    END
  END BM_SRAM28
  PIN BM_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 200.980 108.000 201.380 ;
    END
  END BM_SRAM29
  PIN BM_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 135.460 108.000 135.860 ;
    END
  END BM_SRAM3
  PIN BM_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 203.500 108.000 203.900 ;
    END
  END BM_SRAM30
  PIN BM_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 206.020 108.000 206.420 ;
    END
  END BM_SRAM31
  PIN BM_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 137.980 108.000 138.380 ;
    END
  END BM_SRAM4
  PIN BM_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 140.500 108.000 140.900 ;
    END
  END BM_SRAM5
  PIN BM_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 143.020 108.000 143.420 ;
    END
  END BM_SRAM6
  PIN BM_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 145.540 108.000 145.940 ;
    END
  END BM_SRAM7
  PIN BM_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 148.060 108.000 148.460 ;
    END
  END BM_SRAM8
  PIN BM_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 150.580 108.000 150.980 ;
    END
  END BM_SRAM9
  PIN CLK_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 208.540 108.000 208.940 ;
    END
  END CLK_SRAM
  PIN CONFIGURED_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 19.540 108.000 19.940 ;
    END
  END CONFIGURED_top
  PIN DIN_SRAM0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 211.060 108.000 211.460 ;
    END
  END DIN_SRAM0
  PIN DIN_SRAM1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 213.580 108.000 213.980 ;
    END
  END DIN_SRAM1
  PIN DIN_SRAM10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 236.260 108.000 236.660 ;
    END
  END DIN_SRAM10
  PIN DIN_SRAM11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 238.780 108.000 239.180 ;
    END
  END DIN_SRAM11
  PIN DIN_SRAM12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 241.300 108.000 241.700 ;
    END
  END DIN_SRAM12
  PIN DIN_SRAM13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 243.820 108.000 244.220 ;
    END
  END DIN_SRAM13
  PIN DIN_SRAM14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 246.340 108.000 246.740 ;
    END
  END DIN_SRAM14
  PIN DIN_SRAM15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 248.860 108.000 249.260 ;
    END
  END DIN_SRAM15
  PIN DIN_SRAM16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 251.380 108.000 251.780 ;
    END
  END DIN_SRAM16
  PIN DIN_SRAM17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 253.900 108.000 254.300 ;
    END
  END DIN_SRAM17
  PIN DIN_SRAM18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 256.420 108.000 256.820 ;
    END
  END DIN_SRAM18
  PIN DIN_SRAM19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 258.940 108.000 259.340 ;
    END
  END DIN_SRAM19
  PIN DIN_SRAM2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 216.100 108.000 216.500 ;
    END
  END DIN_SRAM2
  PIN DIN_SRAM20
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 261.460 108.000 261.860 ;
    END
  END DIN_SRAM20
  PIN DIN_SRAM21
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 263.980 108.000 264.380 ;
    END
  END DIN_SRAM21
  PIN DIN_SRAM22
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 266.500 108.000 266.900 ;
    END
  END DIN_SRAM22
  PIN DIN_SRAM23
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 269.020 108.000 269.420 ;
    END
  END DIN_SRAM23
  PIN DIN_SRAM24
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 271.540 108.000 271.940 ;
    END
  END DIN_SRAM24
  PIN DIN_SRAM25
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 274.060 108.000 274.460 ;
    END
  END DIN_SRAM25
  PIN DIN_SRAM26
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 276.580 108.000 276.980 ;
    END
  END DIN_SRAM26
  PIN DIN_SRAM27
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 279.100 108.000 279.500 ;
    END
  END DIN_SRAM27
  PIN DIN_SRAM28
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 281.620 108.000 282.020 ;
    END
  END DIN_SRAM28
  PIN DIN_SRAM29
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 284.140 108.000 284.540 ;
    END
  END DIN_SRAM29
  PIN DIN_SRAM3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 218.620 108.000 219.020 ;
    END
  END DIN_SRAM3
  PIN DIN_SRAM30
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 286.660 108.000 287.060 ;
    END
  END DIN_SRAM30
  PIN DIN_SRAM31
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 289.180 108.000 289.580 ;
    END
  END DIN_SRAM31
  PIN DIN_SRAM4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 221.140 108.000 221.540 ;
    END
  END DIN_SRAM4
  PIN DIN_SRAM5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 223.660 108.000 224.060 ;
    END
  END DIN_SRAM5
  PIN DIN_SRAM6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 226.180 108.000 226.580 ;
    END
  END DIN_SRAM6
  PIN DIN_SRAM7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 228.700 108.000 229.100 ;
    END
  END DIN_SRAM7
  PIN DIN_SRAM8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 231.220 108.000 231.620 ;
    END
  END DIN_SRAM8
  PIN DIN_SRAM9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 233.740 108.000 234.140 ;
    END
  END DIN_SRAM9
  PIN DOUT_SRAM0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 22.060 108.000 22.460 ;
    END
  END DOUT_SRAM0
  PIN DOUT_SRAM1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 24.580 108.000 24.980 ;
    END
  END DOUT_SRAM1
  PIN DOUT_SRAM10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 47.260 108.000 47.660 ;
    END
  END DOUT_SRAM10
  PIN DOUT_SRAM11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 49.780 108.000 50.180 ;
    END
  END DOUT_SRAM11
  PIN DOUT_SRAM12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 52.300 108.000 52.700 ;
    END
  END DOUT_SRAM12
  PIN DOUT_SRAM13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 54.820 108.000 55.220 ;
    END
  END DOUT_SRAM13
  PIN DOUT_SRAM14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 57.340 108.000 57.740 ;
    END
  END DOUT_SRAM14
  PIN DOUT_SRAM15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 59.860 108.000 60.260 ;
    END
  END DOUT_SRAM15
  PIN DOUT_SRAM16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 62.380 108.000 62.780 ;
    END
  END DOUT_SRAM16
  PIN DOUT_SRAM17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 64.900 108.000 65.300 ;
    END
  END DOUT_SRAM17
  PIN DOUT_SRAM18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 67.420 108.000 67.820 ;
    END
  END DOUT_SRAM18
  PIN DOUT_SRAM19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 69.940 108.000 70.340 ;
    END
  END DOUT_SRAM19
  PIN DOUT_SRAM2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 27.100 108.000 27.500 ;
    END
  END DOUT_SRAM2
  PIN DOUT_SRAM20
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 72.460 108.000 72.860 ;
    END
  END DOUT_SRAM20
  PIN DOUT_SRAM21
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 74.980 108.000 75.380 ;
    END
  END DOUT_SRAM21
  PIN DOUT_SRAM22
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 77.500 108.000 77.900 ;
    END
  END DOUT_SRAM22
  PIN DOUT_SRAM23
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 80.020 108.000 80.420 ;
    END
  END DOUT_SRAM23
  PIN DOUT_SRAM24
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 82.540 108.000 82.940 ;
    END
  END DOUT_SRAM24
  PIN DOUT_SRAM25
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 85.060 108.000 85.460 ;
    END
  END DOUT_SRAM25
  PIN DOUT_SRAM26
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 87.580 108.000 87.980 ;
    END
  END DOUT_SRAM26
  PIN DOUT_SRAM27
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 90.100 108.000 90.500 ;
    END
  END DOUT_SRAM27
  PIN DOUT_SRAM28
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 92.620 108.000 93.020 ;
    END
  END DOUT_SRAM28
  PIN DOUT_SRAM29
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 95.140 108.000 95.540 ;
    END
  END DOUT_SRAM29
  PIN DOUT_SRAM3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 29.620 108.000 30.020 ;
    END
  END DOUT_SRAM3
  PIN DOUT_SRAM30
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 97.660 108.000 98.060 ;
    END
  END DOUT_SRAM30
  PIN DOUT_SRAM31
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 100.180 108.000 100.580 ;
    END
  END DOUT_SRAM31
  PIN DOUT_SRAM4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 32.140 108.000 32.540 ;
    END
  END DOUT_SRAM4
  PIN DOUT_SRAM5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 34.660 108.000 35.060 ;
    END
  END DOUT_SRAM5
  PIN DOUT_SRAM6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 37.180 108.000 37.580 ;
    END
  END DOUT_SRAM6
  PIN DOUT_SRAM7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 39.700 108.000 40.100 ;
    END
  END DOUT_SRAM7
  PIN DOUT_SRAM8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 42.220 108.000 42.620 ;
    END
  END DOUT_SRAM8
  PIN DOUT_SRAM9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 44.740 108.000 45.140 ;
    END
  END DOUT_SRAM9
  PIN MEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 291.700 108.000 292.100 ;
    END
  END MEN_SRAM
  PIN REN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 294.220 108.000 294.620 ;
    END
  END REN_SRAM
  PIN TIE_HIGH_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 296.740 108.000 297.140 ;
    END
  END TIE_HIGH_SRAM
  PIN TIE_LOW_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 299.260 108.000 299.660 ;
    END
  END TIE_LOW_SRAM
  PIN Tile_X0Y0_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 336.220 0.450 336.620 ;
    END
  END Tile_X0Y0_E1END[0]
  PIN Tile_X0Y0_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 337.900 0.450 338.300 ;
    END
  END Tile_X0Y0_E1END[1]
  PIN Tile_X0Y0_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 339.580 0.450 339.980 ;
    END
  END Tile_X0Y0_E1END[2]
  PIN Tile_X0Y0_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 341.260 0.450 341.660 ;
    END
  END Tile_X0Y0_E1END[3]
  PIN Tile_X0Y0_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 356.380 0.450 356.780 ;
    END
  END Tile_X0Y0_E2END[0]
  PIN Tile_X0Y0_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 358.060 0.450 358.460 ;
    END
  END Tile_X0Y0_E2END[1]
  PIN Tile_X0Y0_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 359.740 0.450 360.140 ;
    END
  END Tile_X0Y0_E2END[2]
  PIN Tile_X0Y0_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 361.420 0.450 361.820 ;
    END
  END Tile_X0Y0_E2END[3]
  PIN Tile_X0Y0_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 363.100 0.450 363.500 ;
    END
  END Tile_X0Y0_E2END[4]
  PIN Tile_X0Y0_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 364.780 0.450 365.180 ;
    END
  END Tile_X0Y0_E2END[5]
  PIN Tile_X0Y0_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 366.460 0.450 366.860 ;
    END
  END Tile_X0Y0_E2END[6]
  PIN Tile_X0Y0_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 368.140 0.450 368.540 ;
    END
  END Tile_X0Y0_E2END[7]
  PIN Tile_X0Y0_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 342.940 0.450 343.340 ;
    END
  END Tile_X0Y0_E2MID[0]
  PIN Tile_X0Y0_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 344.620 0.450 345.020 ;
    END
  END Tile_X0Y0_E2MID[1]
  PIN Tile_X0Y0_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 346.300 0.450 346.700 ;
    END
  END Tile_X0Y0_E2MID[2]
  PIN Tile_X0Y0_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 347.980 0.450 348.380 ;
    END
  END Tile_X0Y0_E2MID[3]
  PIN Tile_X0Y0_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 349.660 0.450 350.060 ;
    END
  END Tile_X0Y0_E2MID[4]
  PIN Tile_X0Y0_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 351.340 0.450 351.740 ;
    END
  END Tile_X0Y0_E2MID[5]
  PIN Tile_X0Y0_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 353.020 0.450 353.420 ;
    END
  END Tile_X0Y0_E2MID[6]
  PIN Tile_X0Y0_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 354.700 0.450 355.100 ;
    END
  END Tile_X0Y0_E2MID[7]
  PIN Tile_X0Y0_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 396.700 0.450 397.100 ;
    END
  END Tile_X0Y0_E6END[0]
  PIN Tile_X0Y0_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 413.500 0.450 413.900 ;
    END
  END Tile_X0Y0_E6END[10]
  PIN Tile_X0Y0_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 415.180 0.450 415.580 ;
    END
  END Tile_X0Y0_E6END[11]
  PIN Tile_X0Y0_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 398.380 0.450 398.780 ;
    END
  END Tile_X0Y0_E6END[1]
  PIN Tile_X0Y0_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 400.060 0.450 400.460 ;
    END
  END Tile_X0Y0_E6END[2]
  PIN Tile_X0Y0_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 401.740 0.450 402.140 ;
    END
  END Tile_X0Y0_E6END[3]
  PIN Tile_X0Y0_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 403.420 0.450 403.820 ;
    END
  END Tile_X0Y0_E6END[4]
  PIN Tile_X0Y0_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 405.100 0.450 405.500 ;
    END
  END Tile_X0Y0_E6END[5]
  PIN Tile_X0Y0_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 406.780 0.450 407.180 ;
    END
  END Tile_X0Y0_E6END[6]
  PIN Tile_X0Y0_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 408.460 0.450 408.860 ;
    END
  END Tile_X0Y0_E6END[7]
  PIN Tile_X0Y0_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 410.140 0.450 410.540 ;
    END
  END Tile_X0Y0_E6END[8]
  PIN Tile_X0Y0_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 411.820 0.450 412.220 ;
    END
  END Tile_X0Y0_E6END[9]
  PIN Tile_X0Y0_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 369.820 0.450 370.220 ;
    END
  END Tile_X0Y0_EE4END[0]
  PIN Tile_X0Y0_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 386.620 0.450 387.020 ;
    END
  END Tile_X0Y0_EE4END[10]
  PIN Tile_X0Y0_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 388.300 0.450 388.700 ;
    END
  END Tile_X0Y0_EE4END[11]
  PIN Tile_X0Y0_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 389.980 0.450 390.380 ;
    END
  END Tile_X0Y0_EE4END[12]
  PIN Tile_X0Y0_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 391.660 0.450 392.060 ;
    END
  END Tile_X0Y0_EE4END[13]
  PIN Tile_X0Y0_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 393.340 0.450 393.740 ;
    END
  END Tile_X0Y0_EE4END[14]
  PIN Tile_X0Y0_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 395.020 0.450 395.420 ;
    END
  END Tile_X0Y0_EE4END[15]
  PIN Tile_X0Y0_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 371.500 0.450 371.900 ;
    END
  END Tile_X0Y0_EE4END[1]
  PIN Tile_X0Y0_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 373.180 0.450 373.580 ;
    END
  END Tile_X0Y0_EE4END[2]
  PIN Tile_X0Y0_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 374.860 0.450 375.260 ;
    END
  END Tile_X0Y0_EE4END[3]
  PIN Tile_X0Y0_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 376.540 0.450 376.940 ;
    END
  END Tile_X0Y0_EE4END[4]
  PIN Tile_X0Y0_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 378.220 0.450 378.620 ;
    END
  END Tile_X0Y0_EE4END[5]
  PIN Tile_X0Y0_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 379.900 0.450 380.300 ;
    END
  END Tile_X0Y0_EE4END[6]
  PIN Tile_X0Y0_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 381.580 0.450 381.980 ;
    END
  END Tile_X0Y0_EE4END[7]
  PIN Tile_X0Y0_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 383.260 0.450 383.660 ;
    END
  END Tile_X0Y0_EE4END[8]
  PIN Tile_X0Y0_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 384.940 0.450 385.340 ;
    END
  END Tile_X0Y0_EE4END[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 416.860 0.450 417.260 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 433.660 0.450 434.060 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 435.340 0.450 435.740 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 437.020 0.450 437.420 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 438.700 0.450 439.100 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 440.380 0.450 440.780 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 442.060 0.450 442.460 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 443.740 0.450 444.140 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 445.420 0.450 445.820 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 447.100 0.450 447.500 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 448.780 0.450 449.180 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 418.540 0.450 418.940 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 450.460 0.450 450.860 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 452.140 0.450 452.540 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 453.820 0.450 454.220 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 455.500 0.450 455.900 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 457.180 0.450 457.580 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 458.860 0.450 459.260 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 460.540 0.450 460.940 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 462.220 0.450 462.620 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 463.900 0.450 464.300 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 465.580 0.450 465.980 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 420.220 0.450 420.620 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 467.260 0.450 467.660 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 468.940 0.450 469.340 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 421.900 0.450 422.300 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 423.580 0.450 423.980 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 425.260 0.450 425.660 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 426.940 0.450 427.340 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 428.620 0.450 429.020 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 430.300 0.450 430.700 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 431.980 0.450 432.380 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 304.300 108.000 304.700 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 329.500 108.000 329.900 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 332.020 108.000 332.420 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 334.540 108.000 334.940 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 337.060 108.000 337.460 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 339.580 108.000 339.980 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 342.100 108.000 342.500 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 344.620 108.000 345.020 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 347.140 108.000 347.540 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 349.660 108.000 350.060 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 352.180 108.000 352.580 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 306.820 108.000 307.220 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 354.700 108.000 355.100 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 357.220 108.000 357.620 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 359.740 108.000 360.140 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 362.260 108.000 362.660 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 364.780 108.000 365.180 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 367.300 108.000 367.700 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 369.820 108.000 370.220 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 372.340 108.000 372.740 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 374.860 108.000 375.260 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 377.380 108.000 377.780 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 309.340 108.000 309.740 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 379.900 108.000 380.300 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 382.420 108.000 382.820 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 311.860 108.000 312.260 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 314.380 108.000 314.780 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 316.900 108.000 317.300 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 319.420 108.000 319.820 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 321.940 108.000 322.340 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 324.460 108.000 324.860 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 326.980 108.000 327.380 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 483.440 79.400 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 483.440 89.000 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 89.560 483.440 89.960 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 483.440 90.920 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 91.480 483.440 91.880 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 483.440 92.840 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 93.400 483.440 93.800 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 483.440 94.760 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 95.320 483.440 95.720 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 483.440 96.680 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 97.240 483.440 97.640 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.960 483.440 80.360 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 483.440 81.320 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 81.880 483.440 82.280 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 483.440 83.240 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 83.800 483.440 84.200 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 483.440 85.160 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 85.720 483.440 86.120 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 483.440 87.080 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 87.640 483.440 88.040 483.840 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 8.920 483.440 9.320 483.840 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 9.880 483.440 10.280 483.840 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 10.840 483.440 11.240 483.840 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 11.800 483.440 12.200 483.840 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 12.760 483.440 13.160 483.840 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 483.440 14.120 483.840 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 14.680 483.440 15.080 483.840 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 483.440 16.040 483.840 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 16.600 483.440 17.000 483.840 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 483.440 17.960 483.840 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 18.520 483.440 18.920 483.840 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 483.440 19.880 483.840 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 20.440 483.440 20.840 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 483.440 21.800 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 22.360 483.440 22.760 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 483.440 23.720 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 24.280 483.440 24.680 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 483.440 25.640 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 26.200 483.440 26.600 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 483.440 27.560 483.840 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 28.120 483.440 28.520 483.840 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 37.720 483.440 38.120 483.840 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 483.440 39.080 483.840 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 39.640 483.440 40.040 483.840 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 483.440 41.000 483.840 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 41.560 483.440 41.960 483.840 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 483.440 42.920 483.840 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 483.440 29.480 483.840 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 30.040 483.440 30.440 483.840 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 483.440 31.400 483.840 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 31.960 483.440 32.360 483.840 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 483.440 33.320 483.840 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 33.880 483.440 34.280 483.840 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 483.440 35.240 483.840 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 35.800 483.440 36.200 483.840 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 483.440 37.160 483.840 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 43.480 483.440 43.880 483.840 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 483.440 44.840 483.840 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 483.440 45.800 483.840 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 483.440 46.760 483.840 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.000 483.440 55.400 483.840 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 483.440 56.360 483.840 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 483.440 57.320 483.840 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 483.440 58.280 483.840 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 58.840 483.440 59.240 483.840 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 483.440 60.200 483.840 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 60.760 483.440 61.160 483.840 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 483.440 62.120 483.840 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 47.320 483.440 47.720 483.840 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 483.440 48.680 483.840 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 49.240 483.440 49.640 483.840 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 483.440 50.600 483.840 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 51.160 483.440 51.560 483.840 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 483.440 52.520 483.840 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 53.080 483.440 53.480 483.840 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 483.440 54.440 483.840 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 483.440 63.080 483.840 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 72.280 483.440 72.680 483.840 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 483.440 73.640 483.840 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 74.200 483.440 74.600 483.840 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 483.440 75.560 483.840 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 76.120 483.440 76.520 483.840 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 483.440 77.480 483.840 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 483.440 64.040 483.840 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 64.600 483.440 65.000 483.840 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 483.440 65.960 483.840 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 66.520 483.440 66.920 483.840 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 483.440 67.880 483.840 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 68.440 483.440 68.840 483.840 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 483.440 69.800 483.840 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 70.360 483.440 70.760 483.840 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 483.440 71.720 483.840 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 78.040 483.440 78.440 483.840 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 255.580 0.450 255.980 ;
    END
  END Tile_X0Y0_W1BEG[0]
  PIN Tile_X0Y0_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 257.260 0.450 257.660 ;
    END
  END Tile_X0Y0_W1BEG[1]
  PIN Tile_X0Y0_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 258.940 0.450 259.340 ;
    END
  END Tile_X0Y0_W1BEG[2]
  PIN Tile_X0Y0_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 260.620 0.450 261.020 ;
    END
  END Tile_X0Y0_W1BEG[3]
  PIN Tile_X0Y0_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 262.300 0.450 262.700 ;
    END
  END Tile_X0Y0_W2BEG[0]
  PIN Tile_X0Y0_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 263.980 0.450 264.380 ;
    END
  END Tile_X0Y0_W2BEG[1]
  PIN Tile_X0Y0_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 265.660 0.450 266.060 ;
    END
  END Tile_X0Y0_W2BEG[2]
  PIN Tile_X0Y0_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 267.340 0.450 267.740 ;
    END
  END Tile_X0Y0_W2BEG[3]
  PIN Tile_X0Y0_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 269.020 0.450 269.420 ;
    END
  END Tile_X0Y0_W2BEG[4]
  PIN Tile_X0Y0_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 270.700 0.450 271.100 ;
    END
  END Tile_X0Y0_W2BEG[5]
  PIN Tile_X0Y0_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 272.380 0.450 272.780 ;
    END
  END Tile_X0Y0_W2BEG[6]
  PIN Tile_X0Y0_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 274.060 0.450 274.460 ;
    END
  END Tile_X0Y0_W2BEG[7]
  PIN Tile_X0Y0_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 275.740 0.450 276.140 ;
    END
  END Tile_X0Y0_W2BEGb[0]
  PIN Tile_X0Y0_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 277.420 0.450 277.820 ;
    END
  END Tile_X0Y0_W2BEGb[1]
  PIN Tile_X0Y0_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 279.100 0.450 279.500 ;
    END
  END Tile_X0Y0_W2BEGb[2]
  PIN Tile_X0Y0_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 280.780 0.450 281.180 ;
    END
  END Tile_X0Y0_W2BEGb[3]
  PIN Tile_X0Y0_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 282.460 0.450 282.860 ;
    END
  END Tile_X0Y0_W2BEGb[4]
  PIN Tile_X0Y0_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 284.140 0.450 284.540 ;
    END
  END Tile_X0Y0_W2BEGb[5]
  PIN Tile_X0Y0_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 285.820 0.450 286.220 ;
    END
  END Tile_X0Y0_W2BEGb[6]
  PIN Tile_X0Y0_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 287.500 0.450 287.900 ;
    END
  END Tile_X0Y0_W2BEGb[7]
  PIN Tile_X0Y0_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 316.060 0.450 316.460 ;
    END
  END Tile_X0Y0_W6BEG[0]
  PIN Tile_X0Y0_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 332.860 0.450 333.260 ;
    END
  END Tile_X0Y0_W6BEG[10]
  PIN Tile_X0Y0_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 334.540 0.450 334.940 ;
    END
  END Tile_X0Y0_W6BEG[11]
  PIN Tile_X0Y0_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 317.740 0.450 318.140 ;
    END
  END Tile_X0Y0_W6BEG[1]
  PIN Tile_X0Y0_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 319.420 0.450 319.820 ;
    END
  END Tile_X0Y0_W6BEG[2]
  PIN Tile_X0Y0_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 321.100 0.450 321.500 ;
    END
  END Tile_X0Y0_W6BEG[3]
  PIN Tile_X0Y0_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 322.780 0.450 323.180 ;
    END
  END Tile_X0Y0_W6BEG[4]
  PIN Tile_X0Y0_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 324.460 0.450 324.860 ;
    END
  END Tile_X0Y0_W6BEG[5]
  PIN Tile_X0Y0_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 326.140 0.450 326.540 ;
    END
  END Tile_X0Y0_W6BEG[6]
  PIN Tile_X0Y0_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 327.820 0.450 328.220 ;
    END
  END Tile_X0Y0_W6BEG[7]
  PIN Tile_X0Y0_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 329.500 0.450 329.900 ;
    END
  END Tile_X0Y0_W6BEG[8]
  PIN Tile_X0Y0_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 331.180 0.450 331.580 ;
    END
  END Tile_X0Y0_W6BEG[9]
  PIN Tile_X0Y0_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 289.180 0.450 289.580 ;
    END
  END Tile_X0Y0_WW4BEG[0]
  PIN Tile_X0Y0_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 305.980 0.450 306.380 ;
    END
  END Tile_X0Y0_WW4BEG[10]
  PIN Tile_X0Y0_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 307.660 0.450 308.060 ;
    END
  END Tile_X0Y0_WW4BEG[11]
  PIN Tile_X0Y0_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 309.340 0.450 309.740 ;
    END
  END Tile_X0Y0_WW4BEG[12]
  PIN Tile_X0Y0_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 311.020 0.450 311.420 ;
    END
  END Tile_X0Y0_WW4BEG[13]
  PIN Tile_X0Y0_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 312.700 0.450 313.100 ;
    END
  END Tile_X0Y0_WW4BEG[14]
  PIN Tile_X0Y0_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 314.380 0.450 314.780 ;
    END
  END Tile_X0Y0_WW4BEG[15]
  PIN Tile_X0Y0_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 290.860 0.450 291.260 ;
    END
  END Tile_X0Y0_WW4BEG[1]
  PIN Tile_X0Y0_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 292.540 0.450 292.940 ;
    END
  END Tile_X0Y0_WW4BEG[2]
  PIN Tile_X0Y0_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 294.220 0.450 294.620 ;
    END
  END Tile_X0Y0_WW4BEG[3]
  PIN Tile_X0Y0_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 295.900 0.450 296.300 ;
    END
  END Tile_X0Y0_WW4BEG[4]
  PIN Tile_X0Y0_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 297.580 0.450 297.980 ;
    END
  END Tile_X0Y0_WW4BEG[5]
  PIN Tile_X0Y0_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 299.260 0.450 299.660 ;
    END
  END Tile_X0Y0_WW4BEG[6]
  PIN Tile_X0Y0_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 300.940 0.450 301.340 ;
    END
  END Tile_X0Y0_WW4BEG[7]
  PIN Tile_X0Y0_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 302.620 0.450 303.020 ;
    END
  END Tile_X0Y0_WW4BEG[8]
  PIN Tile_X0Y0_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 304.300 0.450 304.700 ;
    END
  END Tile_X0Y0_WW4BEG[9]
  PIN Tile_X0Y1_E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 94.300 0.450 94.700 ;
    END
  END Tile_X0Y1_E1END[0]
  PIN Tile_X0Y1_E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 95.980 0.450 96.380 ;
    END
  END Tile_X0Y1_E1END[1]
  PIN Tile_X0Y1_E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 97.660 0.450 98.060 ;
    END
  END Tile_X0Y1_E1END[2]
  PIN Tile_X0Y1_E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 99.340 0.450 99.740 ;
    END
  END Tile_X0Y1_E1END[3]
  PIN Tile_X0Y1_E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 114.460 0.450 114.860 ;
    END
  END Tile_X0Y1_E2END[0]
  PIN Tile_X0Y1_E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 116.140 0.450 116.540 ;
    END
  END Tile_X0Y1_E2END[1]
  PIN Tile_X0Y1_E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 117.820 0.450 118.220 ;
    END
  END Tile_X0Y1_E2END[2]
  PIN Tile_X0Y1_E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 119.500 0.450 119.900 ;
    END
  END Tile_X0Y1_E2END[3]
  PIN Tile_X0Y1_E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 121.180 0.450 121.580 ;
    END
  END Tile_X0Y1_E2END[4]
  PIN Tile_X0Y1_E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 122.860 0.450 123.260 ;
    END
  END Tile_X0Y1_E2END[5]
  PIN Tile_X0Y1_E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 124.540 0.450 124.940 ;
    END
  END Tile_X0Y1_E2END[6]
  PIN Tile_X0Y1_E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 126.220 0.450 126.620 ;
    END
  END Tile_X0Y1_E2END[7]
  PIN Tile_X0Y1_E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 101.020 0.450 101.420 ;
    END
  END Tile_X0Y1_E2MID[0]
  PIN Tile_X0Y1_E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 102.700 0.450 103.100 ;
    END
  END Tile_X0Y1_E2MID[1]
  PIN Tile_X0Y1_E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 104.380 0.450 104.780 ;
    END
  END Tile_X0Y1_E2MID[2]
  PIN Tile_X0Y1_E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 106.060 0.450 106.460 ;
    END
  END Tile_X0Y1_E2MID[3]
  PIN Tile_X0Y1_E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 107.740 0.450 108.140 ;
    END
  END Tile_X0Y1_E2MID[4]
  PIN Tile_X0Y1_E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 109.420 0.450 109.820 ;
    END
  END Tile_X0Y1_E2MID[5]
  PIN Tile_X0Y1_E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 111.100 0.450 111.500 ;
    END
  END Tile_X0Y1_E2MID[6]
  PIN Tile_X0Y1_E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 112.780 0.450 113.180 ;
    END
  END Tile_X0Y1_E2MID[7]
  PIN Tile_X0Y1_E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 154.780 0.450 155.180 ;
    END
  END Tile_X0Y1_E6END[0]
  PIN Tile_X0Y1_E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 171.580 0.450 171.980 ;
    END
  END Tile_X0Y1_E6END[10]
  PIN Tile_X0Y1_E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 173.260 0.450 173.660 ;
    END
  END Tile_X0Y1_E6END[11]
  PIN Tile_X0Y1_E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 156.460 0.450 156.860 ;
    END
  END Tile_X0Y1_E6END[1]
  PIN Tile_X0Y1_E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 158.140 0.450 158.540 ;
    END
  END Tile_X0Y1_E6END[2]
  PIN Tile_X0Y1_E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 159.820 0.450 160.220 ;
    END
  END Tile_X0Y1_E6END[3]
  PIN Tile_X0Y1_E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 161.500 0.450 161.900 ;
    END
  END Tile_X0Y1_E6END[4]
  PIN Tile_X0Y1_E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 163.180 0.450 163.580 ;
    END
  END Tile_X0Y1_E6END[5]
  PIN Tile_X0Y1_E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 164.860 0.450 165.260 ;
    END
  END Tile_X0Y1_E6END[6]
  PIN Tile_X0Y1_E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 166.540 0.450 166.940 ;
    END
  END Tile_X0Y1_E6END[7]
  PIN Tile_X0Y1_E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 168.220 0.450 168.620 ;
    END
  END Tile_X0Y1_E6END[8]
  PIN Tile_X0Y1_E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 169.900 0.450 170.300 ;
    END
  END Tile_X0Y1_E6END[9]
  PIN Tile_X0Y1_EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 127.900 0.450 128.300 ;
    END
  END Tile_X0Y1_EE4END[0]
  PIN Tile_X0Y1_EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 144.700 0.450 145.100 ;
    END
  END Tile_X0Y1_EE4END[10]
  PIN Tile_X0Y1_EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 146.380 0.450 146.780 ;
    END
  END Tile_X0Y1_EE4END[11]
  PIN Tile_X0Y1_EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 148.060 0.450 148.460 ;
    END
  END Tile_X0Y1_EE4END[12]
  PIN Tile_X0Y1_EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 149.740 0.450 150.140 ;
    END
  END Tile_X0Y1_EE4END[13]
  PIN Tile_X0Y1_EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 151.420 0.450 151.820 ;
    END
  END Tile_X0Y1_EE4END[14]
  PIN Tile_X0Y1_EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 153.100 0.450 153.500 ;
    END
  END Tile_X0Y1_EE4END[15]
  PIN Tile_X0Y1_EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 129.580 0.450 129.980 ;
    END
  END Tile_X0Y1_EE4END[1]
  PIN Tile_X0Y1_EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 131.260 0.450 131.660 ;
    END
  END Tile_X0Y1_EE4END[2]
  PIN Tile_X0Y1_EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 132.940 0.450 133.340 ;
    END
  END Tile_X0Y1_EE4END[3]
  PIN Tile_X0Y1_EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 134.620 0.450 135.020 ;
    END
  END Tile_X0Y1_EE4END[4]
  PIN Tile_X0Y1_EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 136.300 0.450 136.700 ;
    END
  END Tile_X0Y1_EE4END[5]
  PIN Tile_X0Y1_EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 137.980 0.450 138.380 ;
    END
  END Tile_X0Y1_EE4END[6]
  PIN Tile_X0Y1_EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 139.660 0.450 140.060 ;
    END
  END Tile_X0Y1_EE4END[7]
  PIN Tile_X0Y1_EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 141.340 0.450 141.740 ;
    END
  END Tile_X0Y1_EE4END[8]
  PIN Tile_X0Y1_EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 143.020 0.450 143.420 ;
    END
  END Tile_X0Y1_EE4END[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 174.940 0.450 175.340 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 191.740 0.450 192.140 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 193.420 0.450 193.820 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 195.100 0.450 195.500 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 196.780 0.450 197.180 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 198.460 0.450 198.860 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 200.140 0.450 200.540 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 201.820 0.450 202.220 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 203.500 0.450 203.900 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 205.180 0.450 205.580 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 206.860 0.450 207.260 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 176.620 0.450 177.020 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 208.540 0.450 208.940 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 210.220 0.450 210.620 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 211.900 0.450 212.300 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 213.580 0.450 213.980 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 215.260 0.450 215.660 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 216.940 0.450 217.340 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 218.620 0.450 219.020 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 220.300 0.450 220.700 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 221.980 0.450 222.380 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 223.660 0.450 224.060 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 178.300 0.450 178.700 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 225.340 0.450 225.740 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 227.020 0.450 227.420 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 179.980 0.450 180.380 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 181.660 0.450 182.060 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 183.340 0.450 183.740 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 185.020 0.450 185.420 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 186.700 0.450 187.100 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 188.380 0.450 188.780 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 190.060 0.450 190.460 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 384.940 108.000 385.340 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 410.140 108.000 410.540 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 412.660 108.000 413.060 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 415.180 108.000 415.580 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 417.700 108.000 418.100 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 420.220 108.000 420.620 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 422.740 108.000 423.140 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 425.260 108.000 425.660 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 427.780 108.000 428.180 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 430.300 108.000 430.700 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 432.820 108.000 433.220 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 387.460 108.000 387.860 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 435.340 108.000 435.740 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 437.860 108.000 438.260 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 440.380 108.000 440.780 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 442.900 108.000 443.300 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 445.420 108.000 445.820 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 447.940 108.000 448.340 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 450.460 108.000 450.860 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 452.980 108.000 453.380 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 455.500 108.000 455.900 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 458.020 108.000 458.420 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 389.980 108.000 390.380 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 460.540 108.000 460.940 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 463.060 108.000 463.460 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 392.500 108.000 392.900 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 395.020 108.000 395.420 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 397.540 108.000 397.940 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 400.060 108.000 400.460 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 402.580 108.000 402.980 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 405.100 108.000 405.500 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 407.620 108.000 408.020 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 91.480 0.000 91.880 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 93.400 0.000 93.800 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 97.240 0.000 97.640 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 79.960 0.000 80.360 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 81.880 0.000 82.280 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.542100 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 85.720 0.000 86.120 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 87.640 0.000 88.040 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 8.920 0.000 9.320 0.400 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 9.880 0.000 10.280 0.400 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 10.840 0.000 11.240 0.400 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 11.800 0.000 12.200 0.400 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 20.440 0.000 20.840 0.400 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 0.000 21.800 0.400 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 22.360 0.000 22.760 0.400 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 0.000 23.720 0.400 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 24.280 0.000 24.680 0.400 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 26.200 0.000 26.600 0.400 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 0.000 27.560 0.400 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 12.760 0.000 13.160 0.400 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 14.680 0.000 15.080 0.400 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 0.000 16.040 0.400 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 16.600 0.000 17.000 0.400 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 0.000 17.960 0.400 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 18.520 0.000 18.920 0.400 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 28.120 0.000 28.520 0.400 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 37.720 0.000 38.120 0.400 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 41.560 0.000 41.960 0.400 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 0.000 29.480 0.400 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 30.040 0.000 30.440 0.400 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 31.960 0.000 32.360 0.400 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 33.880 0.000 34.280 0.400 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 35.800 0.000 36.200 0.400 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 43.480 0.000 43.880 0.400 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 47.320 0.000 47.720 0.400 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 49.240 0.000 49.640 0.400 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 0.000 50.600 0.400 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 51.160 0.000 51.560 0.400 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 0.000 52.520 0.400 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 53.080 0.000 53.480 0.400 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 58.840 0.000 59.240 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 74.200 0.000 74.600 0.400 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 76.120 0.000 76.520 0.400 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 64.600 0.000 65.000 0.400 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 68.440 0.000 68.840 0.400 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.361400 ;
    PORT
      LAYER Metal3 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 13.660 0.450 14.060 ;
    END
  END Tile_X0Y1_W1BEG[0]
  PIN Tile_X0Y1_W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.340 0.450 15.740 ;
    END
  END Tile_X0Y1_W1BEG[1]
  PIN Tile_X0Y1_W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.020 0.450 17.420 ;
    END
  END Tile_X0Y1_W1BEG[2]
  PIN Tile_X0Y1_W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.700 0.450 19.100 ;
    END
  END Tile_X0Y1_W1BEG[3]
  PIN Tile_X0Y1_W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 20.380 0.450 20.780 ;
    END
  END Tile_X0Y1_W2BEG[0]
  PIN Tile_X0Y1_W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.060 0.450 22.460 ;
    END
  END Tile_X0Y1_W2BEG[1]
  PIN Tile_X0Y1_W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.740 0.450 24.140 ;
    END
  END Tile_X0Y1_W2BEG[2]
  PIN Tile_X0Y1_W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 25.420 0.450 25.820 ;
    END
  END Tile_X0Y1_W2BEG[3]
  PIN Tile_X0Y1_W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.100 0.450 27.500 ;
    END
  END Tile_X0Y1_W2BEG[4]
  PIN Tile_X0Y1_W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 28.780 0.450 29.180 ;
    END
  END Tile_X0Y1_W2BEG[5]
  PIN Tile_X0Y1_W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.460 0.450 30.860 ;
    END
  END Tile_X0Y1_W2BEG[6]
  PIN Tile_X0Y1_W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.140 0.450 32.540 ;
    END
  END Tile_X0Y1_W2BEG[7]
  PIN Tile_X0Y1_W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 33.820 0.450 34.220 ;
    END
  END Tile_X0Y1_W2BEGb[0]
  PIN Tile_X0Y1_W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 35.500 0.450 35.900 ;
    END
  END Tile_X0Y1_W2BEGb[1]
  PIN Tile_X0Y1_W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 37.180 0.450 37.580 ;
    END
  END Tile_X0Y1_W2BEGb[2]
  PIN Tile_X0Y1_W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.860 0.450 39.260 ;
    END
  END Tile_X0Y1_W2BEGb[3]
  PIN Tile_X0Y1_W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 40.540 0.450 40.940 ;
    END
  END Tile_X0Y1_W2BEGb[4]
  PIN Tile_X0Y1_W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 42.220 0.450 42.620 ;
    END
  END Tile_X0Y1_W2BEGb[5]
  PIN Tile_X0Y1_W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.900 0.450 44.300 ;
    END
  END Tile_X0Y1_W2BEGb[6]
  PIN Tile_X0Y1_W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 45.580 0.450 45.980 ;
    END
  END Tile_X0Y1_W2BEGb[7]
  PIN Tile_X0Y1_W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 74.140 0.450 74.540 ;
    END
  END Tile_X0Y1_W6BEG[0]
  PIN Tile_X0Y1_W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 90.940 0.450 91.340 ;
    END
  END Tile_X0Y1_W6BEG[10]
  PIN Tile_X0Y1_W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 92.620 0.450 93.020 ;
    END
  END Tile_X0Y1_W6BEG[11]
  PIN Tile_X0Y1_W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 75.820 0.450 76.220 ;
    END
  END Tile_X0Y1_W6BEG[1]
  PIN Tile_X0Y1_W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 77.500 0.450 77.900 ;
    END
  END Tile_X0Y1_W6BEG[2]
  PIN Tile_X0Y1_W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 79.180 0.450 79.580 ;
    END
  END Tile_X0Y1_W6BEG[3]
  PIN Tile_X0Y1_W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 80.860 0.450 81.260 ;
    END
  END Tile_X0Y1_W6BEG[4]
  PIN Tile_X0Y1_W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 82.540 0.450 82.940 ;
    END
  END Tile_X0Y1_W6BEG[5]
  PIN Tile_X0Y1_W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 84.220 0.450 84.620 ;
    END
  END Tile_X0Y1_W6BEG[6]
  PIN Tile_X0Y1_W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 85.900 0.450 86.300 ;
    END
  END Tile_X0Y1_W6BEG[7]
  PIN Tile_X0Y1_W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 87.580 0.450 87.980 ;
    END
  END Tile_X0Y1_W6BEG[8]
  PIN Tile_X0Y1_W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 89.260 0.450 89.660 ;
    END
  END Tile_X0Y1_W6BEG[9]
  PIN Tile_X0Y1_WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 47.260 0.450 47.660 ;
    END
  END Tile_X0Y1_WW4BEG[0]
  PIN Tile_X0Y1_WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 64.060 0.450 64.460 ;
    END
  END Tile_X0Y1_WW4BEG[10]
  PIN Tile_X0Y1_WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 65.740 0.450 66.140 ;
    END
  END Tile_X0Y1_WW4BEG[11]
  PIN Tile_X0Y1_WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 67.420 0.450 67.820 ;
    END
  END Tile_X0Y1_WW4BEG[12]
  PIN Tile_X0Y1_WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 69.100 0.450 69.500 ;
    END
  END Tile_X0Y1_WW4BEG[13]
  PIN Tile_X0Y1_WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 70.780 0.450 71.180 ;
    END
  END Tile_X0Y1_WW4BEG[14]
  PIN Tile_X0Y1_WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 72.460 0.450 72.860 ;
    END
  END Tile_X0Y1_WW4BEG[15]
  PIN Tile_X0Y1_WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.940 0.450 49.340 ;
    END
  END Tile_X0Y1_WW4BEG[1]
  PIN Tile_X0Y1_WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 50.620 0.450 51.020 ;
    END
  END Tile_X0Y1_WW4BEG[2]
  PIN Tile_X0Y1_WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.300 0.450 52.700 ;
    END
  END Tile_X0Y1_WW4BEG[3]
  PIN Tile_X0Y1_WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.980 0.450 54.380 ;
    END
  END Tile_X0Y1_WW4BEG[4]
  PIN Tile_X0Y1_WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 55.660 0.450 56.060 ;
    END
  END Tile_X0Y1_WW4BEG[5]
  PIN Tile_X0Y1_WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 57.340 0.450 57.740 ;
    END
  END Tile_X0Y1_WW4BEG[6]
  PIN Tile_X0Y1_WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 59.020 0.450 59.420 ;
    END
  END Tile_X0Y1_WW4BEG[7]
  PIN Tile_X0Y1_WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 60.700 0.450 61.100 ;
    END
  END Tile_X0Y1_WW4BEG[8]
  PIN Tile_X0Y1_WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 62.380 0.450 62.780 ;
    END
  END Tile_X0Y1_WW4BEG[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 483.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 100.060 0.000 102.260 483.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 483.840 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.860 0.000 96.060 483.840 ;
    END
  END VPWR
  PIN WEN_SRAM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.550 301.780 108.000 302.180 ;
    END
  END WEN_SRAM
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 102.240 476.430 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 102.260 476.500 ;
      LAYER Metal2 ;
        RECT 0.335 469.550 107.875 476.380 ;
        RECT 0.660 468.730 107.875 469.550 ;
        RECT 0.335 467.870 107.875 468.730 ;
        RECT 0.660 467.050 107.875 467.870 ;
        RECT 0.335 466.190 107.875 467.050 ;
        RECT 0.660 465.370 107.875 466.190 ;
        RECT 0.335 464.510 107.875 465.370 ;
        RECT 0.660 463.690 107.875 464.510 ;
        RECT 0.335 463.670 107.875 463.690 ;
        RECT 0.335 462.850 107.340 463.670 ;
        RECT 0.335 462.830 107.875 462.850 ;
        RECT 0.660 462.010 107.875 462.830 ;
        RECT 0.335 461.150 107.875 462.010 ;
        RECT 0.660 460.330 107.340 461.150 ;
        RECT 0.335 459.470 107.875 460.330 ;
        RECT 0.660 458.650 107.875 459.470 ;
        RECT 0.335 458.630 107.875 458.650 ;
        RECT 0.335 457.810 107.340 458.630 ;
        RECT 0.335 457.790 107.875 457.810 ;
        RECT 0.660 456.970 107.875 457.790 ;
        RECT 0.335 456.110 107.875 456.970 ;
        RECT 0.660 455.290 107.340 456.110 ;
        RECT 0.335 454.430 107.875 455.290 ;
        RECT 0.660 453.610 107.875 454.430 ;
        RECT 0.335 453.590 107.875 453.610 ;
        RECT 0.335 452.770 107.340 453.590 ;
        RECT 0.335 452.750 107.875 452.770 ;
        RECT 0.660 451.930 107.875 452.750 ;
        RECT 0.335 451.070 107.875 451.930 ;
        RECT 0.660 450.250 107.340 451.070 ;
        RECT 0.335 449.390 107.875 450.250 ;
        RECT 0.660 448.570 107.875 449.390 ;
        RECT 0.335 448.550 107.875 448.570 ;
        RECT 0.335 447.730 107.340 448.550 ;
        RECT 0.335 447.710 107.875 447.730 ;
        RECT 0.660 446.890 107.875 447.710 ;
        RECT 0.335 446.030 107.875 446.890 ;
        RECT 0.660 445.210 107.340 446.030 ;
        RECT 0.335 444.350 107.875 445.210 ;
        RECT 0.660 443.530 107.875 444.350 ;
        RECT 0.335 443.510 107.875 443.530 ;
        RECT 0.335 442.690 107.340 443.510 ;
        RECT 0.335 442.670 107.875 442.690 ;
        RECT 0.660 441.850 107.875 442.670 ;
        RECT 0.335 440.990 107.875 441.850 ;
        RECT 0.660 440.170 107.340 440.990 ;
        RECT 0.335 439.310 107.875 440.170 ;
        RECT 0.660 438.490 107.875 439.310 ;
        RECT 0.335 438.470 107.875 438.490 ;
        RECT 0.335 437.650 107.340 438.470 ;
        RECT 0.335 437.630 107.875 437.650 ;
        RECT 0.660 436.810 107.875 437.630 ;
        RECT 0.335 435.950 107.875 436.810 ;
        RECT 0.660 435.130 107.340 435.950 ;
        RECT 0.335 434.270 107.875 435.130 ;
        RECT 0.660 433.450 107.875 434.270 ;
        RECT 0.335 433.430 107.875 433.450 ;
        RECT 0.335 432.610 107.340 433.430 ;
        RECT 0.335 432.590 107.875 432.610 ;
        RECT 0.660 431.770 107.875 432.590 ;
        RECT 0.335 430.910 107.875 431.770 ;
        RECT 0.660 430.090 107.340 430.910 ;
        RECT 0.335 429.230 107.875 430.090 ;
        RECT 0.660 428.410 107.875 429.230 ;
        RECT 0.335 428.390 107.875 428.410 ;
        RECT 0.335 427.570 107.340 428.390 ;
        RECT 0.335 427.550 107.875 427.570 ;
        RECT 0.660 426.730 107.875 427.550 ;
        RECT 0.335 425.870 107.875 426.730 ;
        RECT 0.660 425.050 107.340 425.870 ;
        RECT 0.335 424.190 107.875 425.050 ;
        RECT 0.660 423.370 107.875 424.190 ;
        RECT 0.335 423.350 107.875 423.370 ;
        RECT 0.335 422.530 107.340 423.350 ;
        RECT 0.335 422.510 107.875 422.530 ;
        RECT 0.660 421.690 107.875 422.510 ;
        RECT 0.335 420.830 107.875 421.690 ;
        RECT 0.660 420.010 107.340 420.830 ;
        RECT 0.335 419.150 107.875 420.010 ;
        RECT 0.660 418.330 107.875 419.150 ;
        RECT 0.335 418.310 107.875 418.330 ;
        RECT 0.335 417.490 107.340 418.310 ;
        RECT 0.335 417.470 107.875 417.490 ;
        RECT 0.660 416.650 107.875 417.470 ;
        RECT 0.335 415.790 107.875 416.650 ;
        RECT 0.660 414.970 107.340 415.790 ;
        RECT 0.335 414.110 107.875 414.970 ;
        RECT 0.660 413.290 107.875 414.110 ;
        RECT 0.335 413.270 107.875 413.290 ;
        RECT 0.335 412.450 107.340 413.270 ;
        RECT 0.335 412.430 107.875 412.450 ;
        RECT 0.660 411.610 107.875 412.430 ;
        RECT 0.335 410.750 107.875 411.610 ;
        RECT 0.660 409.930 107.340 410.750 ;
        RECT 0.335 409.070 107.875 409.930 ;
        RECT 0.660 408.250 107.875 409.070 ;
        RECT 0.335 408.230 107.875 408.250 ;
        RECT 0.335 407.410 107.340 408.230 ;
        RECT 0.335 407.390 107.875 407.410 ;
        RECT 0.660 406.570 107.875 407.390 ;
        RECT 0.335 405.710 107.875 406.570 ;
        RECT 0.660 404.890 107.340 405.710 ;
        RECT 0.335 404.030 107.875 404.890 ;
        RECT 0.660 403.210 107.875 404.030 ;
        RECT 0.335 403.190 107.875 403.210 ;
        RECT 0.335 402.370 107.340 403.190 ;
        RECT 0.335 402.350 107.875 402.370 ;
        RECT 0.660 401.530 107.875 402.350 ;
        RECT 0.335 400.670 107.875 401.530 ;
        RECT 0.660 399.850 107.340 400.670 ;
        RECT 0.335 398.990 107.875 399.850 ;
        RECT 0.660 398.170 107.875 398.990 ;
        RECT 0.335 398.150 107.875 398.170 ;
        RECT 0.335 397.330 107.340 398.150 ;
        RECT 0.335 397.310 107.875 397.330 ;
        RECT 0.660 396.490 107.875 397.310 ;
        RECT 0.335 395.630 107.875 396.490 ;
        RECT 0.660 394.810 107.340 395.630 ;
        RECT 0.335 393.950 107.875 394.810 ;
        RECT 0.660 393.130 107.875 393.950 ;
        RECT 0.335 393.110 107.875 393.130 ;
        RECT 0.335 392.290 107.340 393.110 ;
        RECT 0.335 392.270 107.875 392.290 ;
        RECT 0.660 391.450 107.875 392.270 ;
        RECT 0.335 390.590 107.875 391.450 ;
        RECT 0.660 389.770 107.340 390.590 ;
        RECT 0.335 388.910 107.875 389.770 ;
        RECT 0.660 388.090 107.875 388.910 ;
        RECT 0.335 388.070 107.875 388.090 ;
        RECT 0.335 387.250 107.340 388.070 ;
        RECT 0.335 387.230 107.875 387.250 ;
        RECT 0.660 386.410 107.875 387.230 ;
        RECT 0.335 385.550 107.875 386.410 ;
        RECT 0.660 384.730 107.340 385.550 ;
        RECT 0.335 383.870 107.875 384.730 ;
        RECT 0.660 383.050 107.875 383.870 ;
        RECT 0.335 383.030 107.875 383.050 ;
        RECT 0.335 382.210 107.340 383.030 ;
        RECT 0.335 382.190 107.875 382.210 ;
        RECT 0.660 381.370 107.875 382.190 ;
        RECT 0.335 380.510 107.875 381.370 ;
        RECT 0.660 379.690 107.340 380.510 ;
        RECT 0.335 378.830 107.875 379.690 ;
        RECT 0.660 378.010 107.875 378.830 ;
        RECT 0.335 377.990 107.875 378.010 ;
        RECT 0.335 377.170 107.340 377.990 ;
        RECT 0.335 377.150 107.875 377.170 ;
        RECT 0.660 376.330 107.875 377.150 ;
        RECT 0.335 375.470 107.875 376.330 ;
        RECT 0.660 374.650 107.340 375.470 ;
        RECT 0.335 373.790 107.875 374.650 ;
        RECT 0.660 372.970 107.875 373.790 ;
        RECT 0.335 372.950 107.875 372.970 ;
        RECT 0.335 372.130 107.340 372.950 ;
        RECT 0.335 372.110 107.875 372.130 ;
        RECT 0.660 371.290 107.875 372.110 ;
        RECT 0.335 370.430 107.875 371.290 ;
        RECT 0.660 369.610 107.340 370.430 ;
        RECT 0.335 368.750 107.875 369.610 ;
        RECT 0.660 367.930 107.875 368.750 ;
        RECT 0.335 367.910 107.875 367.930 ;
        RECT 0.335 367.090 107.340 367.910 ;
        RECT 0.335 367.070 107.875 367.090 ;
        RECT 0.660 366.250 107.875 367.070 ;
        RECT 0.335 365.390 107.875 366.250 ;
        RECT 0.660 364.570 107.340 365.390 ;
        RECT 0.335 363.710 107.875 364.570 ;
        RECT 0.660 362.890 107.875 363.710 ;
        RECT 0.335 362.870 107.875 362.890 ;
        RECT 0.335 362.050 107.340 362.870 ;
        RECT 0.335 362.030 107.875 362.050 ;
        RECT 0.660 361.210 107.875 362.030 ;
        RECT 0.335 360.350 107.875 361.210 ;
        RECT 0.660 359.530 107.340 360.350 ;
        RECT 0.335 358.670 107.875 359.530 ;
        RECT 0.660 357.850 107.875 358.670 ;
        RECT 0.335 357.830 107.875 357.850 ;
        RECT 0.335 357.010 107.340 357.830 ;
        RECT 0.335 356.990 107.875 357.010 ;
        RECT 0.660 356.170 107.875 356.990 ;
        RECT 0.335 355.310 107.875 356.170 ;
        RECT 0.660 354.490 107.340 355.310 ;
        RECT 0.335 353.630 107.875 354.490 ;
        RECT 0.660 352.810 107.875 353.630 ;
        RECT 0.335 352.790 107.875 352.810 ;
        RECT 0.335 351.970 107.340 352.790 ;
        RECT 0.335 351.950 107.875 351.970 ;
        RECT 0.660 351.130 107.875 351.950 ;
        RECT 0.335 350.270 107.875 351.130 ;
        RECT 0.660 349.450 107.340 350.270 ;
        RECT 0.335 348.590 107.875 349.450 ;
        RECT 0.660 347.770 107.875 348.590 ;
        RECT 0.335 347.750 107.875 347.770 ;
        RECT 0.335 346.930 107.340 347.750 ;
        RECT 0.335 346.910 107.875 346.930 ;
        RECT 0.660 346.090 107.875 346.910 ;
        RECT 0.335 345.230 107.875 346.090 ;
        RECT 0.660 344.410 107.340 345.230 ;
        RECT 0.335 343.550 107.875 344.410 ;
        RECT 0.660 342.730 107.875 343.550 ;
        RECT 0.335 342.710 107.875 342.730 ;
        RECT 0.335 341.890 107.340 342.710 ;
        RECT 0.335 341.870 107.875 341.890 ;
        RECT 0.660 341.050 107.875 341.870 ;
        RECT 0.335 340.190 107.875 341.050 ;
        RECT 0.660 339.370 107.340 340.190 ;
        RECT 0.335 338.510 107.875 339.370 ;
        RECT 0.660 337.690 107.875 338.510 ;
        RECT 0.335 337.670 107.875 337.690 ;
        RECT 0.335 336.850 107.340 337.670 ;
        RECT 0.335 336.830 107.875 336.850 ;
        RECT 0.660 336.010 107.875 336.830 ;
        RECT 0.335 335.150 107.875 336.010 ;
        RECT 0.660 334.330 107.340 335.150 ;
        RECT 0.335 333.470 107.875 334.330 ;
        RECT 0.660 332.650 107.875 333.470 ;
        RECT 0.335 332.630 107.875 332.650 ;
        RECT 0.335 331.810 107.340 332.630 ;
        RECT 0.335 331.790 107.875 331.810 ;
        RECT 0.660 330.970 107.875 331.790 ;
        RECT 0.335 330.110 107.875 330.970 ;
        RECT 0.660 329.290 107.340 330.110 ;
        RECT 0.335 328.430 107.875 329.290 ;
        RECT 0.660 327.610 107.875 328.430 ;
        RECT 0.335 327.590 107.875 327.610 ;
        RECT 0.335 326.770 107.340 327.590 ;
        RECT 0.335 326.750 107.875 326.770 ;
        RECT 0.660 325.930 107.875 326.750 ;
        RECT 0.335 325.070 107.875 325.930 ;
        RECT 0.660 324.250 107.340 325.070 ;
        RECT 0.335 323.390 107.875 324.250 ;
        RECT 0.660 322.570 107.875 323.390 ;
        RECT 0.335 322.550 107.875 322.570 ;
        RECT 0.335 321.730 107.340 322.550 ;
        RECT 0.335 321.710 107.875 321.730 ;
        RECT 0.660 320.890 107.875 321.710 ;
        RECT 0.335 320.030 107.875 320.890 ;
        RECT 0.660 319.210 107.340 320.030 ;
        RECT 0.335 318.350 107.875 319.210 ;
        RECT 0.660 317.530 107.875 318.350 ;
        RECT 0.335 317.510 107.875 317.530 ;
        RECT 0.335 316.690 107.340 317.510 ;
        RECT 0.335 316.670 107.875 316.690 ;
        RECT 0.660 315.850 107.875 316.670 ;
        RECT 0.335 314.990 107.875 315.850 ;
        RECT 0.660 314.170 107.340 314.990 ;
        RECT 0.335 313.310 107.875 314.170 ;
        RECT 0.660 312.490 107.875 313.310 ;
        RECT 0.335 312.470 107.875 312.490 ;
        RECT 0.335 311.650 107.340 312.470 ;
        RECT 0.335 311.630 107.875 311.650 ;
        RECT 0.660 310.810 107.875 311.630 ;
        RECT 0.335 309.950 107.875 310.810 ;
        RECT 0.660 309.130 107.340 309.950 ;
        RECT 0.335 308.270 107.875 309.130 ;
        RECT 0.660 307.450 107.875 308.270 ;
        RECT 0.335 307.430 107.875 307.450 ;
        RECT 0.335 306.610 107.340 307.430 ;
        RECT 0.335 306.590 107.875 306.610 ;
        RECT 0.660 305.770 107.875 306.590 ;
        RECT 0.335 304.910 107.875 305.770 ;
        RECT 0.660 304.090 107.340 304.910 ;
        RECT 0.335 303.230 107.875 304.090 ;
        RECT 0.660 302.410 107.875 303.230 ;
        RECT 0.335 302.390 107.875 302.410 ;
        RECT 0.335 301.570 107.340 302.390 ;
        RECT 0.335 301.550 107.875 301.570 ;
        RECT 0.660 300.730 107.875 301.550 ;
        RECT 0.335 299.870 107.875 300.730 ;
        RECT 0.660 299.050 107.340 299.870 ;
        RECT 0.335 298.190 107.875 299.050 ;
        RECT 0.660 297.370 107.875 298.190 ;
        RECT 0.335 297.350 107.875 297.370 ;
        RECT 0.335 296.530 107.340 297.350 ;
        RECT 0.335 296.510 107.875 296.530 ;
        RECT 0.660 295.690 107.875 296.510 ;
        RECT 0.335 294.830 107.875 295.690 ;
        RECT 0.660 294.010 107.340 294.830 ;
        RECT 0.335 293.150 107.875 294.010 ;
        RECT 0.660 292.330 107.875 293.150 ;
        RECT 0.335 292.310 107.875 292.330 ;
        RECT 0.335 291.490 107.340 292.310 ;
        RECT 0.335 291.470 107.875 291.490 ;
        RECT 0.660 290.650 107.875 291.470 ;
        RECT 0.335 289.790 107.875 290.650 ;
        RECT 0.660 288.970 107.340 289.790 ;
        RECT 0.335 288.110 107.875 288.970 ;
        RECT 0.660 287.290 107.875 288.110 ;
        RECT 0.335 287.270 107.875 287.290 ;
        RECT 0.335 286.450 107.340 287.270 ;
        RECT 0.335 286.430 107.875 286.450 ;
        RECT 0.660 285.610 107.875 286.430 ;
        RECT 0.335 284.750 107.875 285.610 ;
        RECT 0.660 283.930 107.340 284.750 ;
        RECT 0.335 283.070 107.875 283.930 ;
        RECT 0.660 282.250 107.875 283.070 ;
        RECT 0.335 282.230 107.875 282.250 ;
        RECT 0.335 281.410 107.340 282.230 ;
        RECT 0.335 281.390 107.875 281.410 ;
        RECT 0.660 280.570 107.875 281.390 ;
        RECT 0.335 279.710 107.875 280.570 ;
        RECT 0.660 278.890 107.340 279.710 ;
        RECT 0.335 278.030 107.875 278.890 ;
        RECT 0.660 277.210 107.875 278.030 ;
        RECT 0.335 277.190 107.875 277.210 ;
        RECT 0.335 276.370 107.340 277.190 ;
        RECT 0.335 276.350 107.875 276.370 ;
        RECT 0.660 275.530 107.875 276.350 ;
        RECT 0.335 274.670 107.875 275.530 ;
        RECT 0.660 273.850 107.340 274.670 ;
        RECT 0.335 272.990 107.875 273.850 ;
        RECT 0.660 272.170 107.875 272.990 ;
        RECT 0.335 272.150 107.875 272.170 ;
        RECT 0.335 271.330 107.340 272.150 ;
        RECT 0.335 271.310 107.875 271.330 ;
        RECT 0.660 270.490 107.875 271.310 ;
        RECT 0.335 269.630 107.875 270.490 ;
        RECT 0.660 268.810 107.340 269.630 ;
        RECT 0.335 267.950 107.875 268.810 ;
        RECT 0.660 267.130 107.875 267.950 ;
        RECT 0.335 267.110 107.875 267.130 ;
        RECT 0.335 266.290 107.340 267.110 ;
        RECT 0.335 266.270 107.875 266.290 ;
        RECT 0.660 265.450 107.875 266.270 ;
        RECT 0.335 264.590 107.875 265.450 ;
        RECT 0.660 263.770 107.340 264.590 ;
        RECT 0.335 262.910 107.875 263.770 ;
        RECT 0.660 262.090 107.875 262.910 ;
        RECT 0.335 262.070 107.875 262.090 ;
        RECT 0.335 261.250 107.340 262.070 ;
        RECT 0.335 261.230 107.875 261.250 ;
        RECT 0.660 260.410 107.875 261.230 ;
        RECT 0.335 259.550 107.875 260.410 ;
        RECT 0.660 258.730 107.340 259.550 ;
        RECT 0.335 257.870 107.875 258.730 ;
        RECT 0.660 257.050 107.875 257.870 ;
        RECT 0.335 257.030 107.875 257.050 ;
        RECT 0.335 256.210 107.340 257.030 ;
        RECT 0.335 256.190 107.875 256.210 ;
        RECT 0.660 255.370 107.875 256.190 ;
        RECT 0.335 254.510 107.875 255.370 ;
        RECT 0.335 253.690 107.340 254.510 ;
        RECT 0.335 251.990 107.875 253.690 ;
        RECT 0.335 251.170 107.340 251.990 ;
        RECT 0.335 249.470 107.875 251.170 ;
        RECT 0.335 248.650 107.340 249.470 ;
        RECT 0.335 246.950 107.875 248.650 ;
        RECT 0.335 246.130 107.340 246.950 ;
        RECT 0.335 244.430 107.875 246.130 ;
        RECT 0.335 243.610 107.340 244.430 ;
        RECT 0.335 241.910 107.875 243.610 ;
        RECT 0.335 241.090 107.340 241.910 ;
        RECT 0.335 239.390 107.875 241.090 ;
        RECT 0.335 238.570 107.340 239.390 ;
        RECT 0.335 236.870 107.875 238.570 ;
        RECT 0.335 236.050 107.340 236.870 ;
        RECT 0.335 234.350 107.875 236.050 ;
        RECT 0.335 233.530 107.340 234.350 ;
        RECT 0.335 231.830 107.875 233.530 ;
        RECT 0.335 231.010 107.340 231.830 ;
        RECT 0.335 229.310 107.875 231.010 ;
        RECT 0.335 228.490 107.340 229.310 ;
        RECT 0.335 227.630 107.875 228.490 ;
        RECT 0.660 226.810 107.875 227.630 ;
        RECT 0.335 226.790 107.875 226.810 ;
        RECT 0.335 225.970 107.340 226.790 ;
        RECT 0.335 225.950 107.875 225.970 ;
        RECT 0.660 225.130 107.875 225.950 ;
        RECT 0.335 224.270 107.875 225.130 ;
        RECT 0.660 223.450 107.340 224.270 ;
        RECT 0.335 222.590 107.875 223.450 ;
        RECT 0.660 221.770 107.875 222.590 ;
        RECT 0.335 221.750 107.875 221.770 ;
        RECT 0.335 220.930 107.340 221.750 ;
        RECT 0.335 220.910 107.875 220.930 ;
        RECT 0.660 220.090 107.875 220.910 ;
        RECT 0.335 219.230 107.875 220.090 ;
        RECT 0.660 218.410 107.340 219.230 ;
        RECT 0.335 217.550 107.875 218.410 ;
        RECT 0.660 216.730 107.875 217.550 ;
        RECT 0.335 216.710 107.875 216.730 ;
        RECT 0.335 215.890 107.340 216.710 ;
        RECT 0.335 215.870 107.875 215.890 ;
        RECT 0.660 215.050 107.875 215.870 ;
        RECT 0.335 214.190 107.875 215.050 ;
        RECT 0.660 213.370 107.340 214.190 ;
        RECT 0.335 212.510 107.875 213.370 ;
        RECT 0.660 211.690 107.875 212.510 ;
        RECT 0.335 211.670 107.875 211.690 ;
        RECT 0.335 210.850 107.340 211.670 ;
        RECT 0.335 210.830 107.875 210.850 ;
        RECT 0.660 210.010 107.875 210.830 ;
        RECT 0.335 209.150 107.875 210.010 ;
        RECT 0.660 208.330 107.340 209.150 ;
        RECT 0.335 207.470 107.875 208.330 ;
        RECT 0.660 206.650 107.875 207.470 ;
        RECT 0.335 206.630 107.875 206.650 ;
        RECT 0.335 205.810 107.340 206.630 ;
        RECT 0.335 205.790 107.875 205.810 ;
        RECT 0.660 204.970 107.875 205.790 ;
        RECT 0.335 204.110 107.875 204.970 ;
        RECT 0.660 203.290 107.340 204.110 ;
        RECT 0.335 202.430 107.875 203.290 ;
        RECT 0.660 201.610 107.875 202.430 ;
        RECT 0.335 201.590 107.875 201.610 ;
        RECT 0.335 200.770 107.340 201.590 ;
        RECT 0.335 200.750 107.875 200.770 ;
        RECT 0.660 199.930 107.875 200.750 ;
        RECT 0.335 199.070 107.875 199.930 ;
        RECT 0.660 198.250 107.340 199.070 ;
        RECT 0.335 197.390 107.875 198.250 ;
        RECT 0.660 196.570 107.875 197.390 ;
        RECT 0.335 196.550 107.875 196.570 ;
        RECT 0.335 195.730 107.340 196.550 ;
        RECT 0.335 195.710 107.875 195.730 ;
        RECT 0.660 194.890 107.875 195.710 ;
        RECT 0.335 194.030 107.875 194.890 ;
        RECT 0.660 193.210 107.340 194.030 ;
        RECT 0.335 192.350 107.875 193.210 ;
        RECT 0.660 191.530 107.875 192.350 ;
        RECT 0.335 191.510 107.875 191.530 ;
        RECT 0.335 190.690 107.340 191.510 ;
        RECT 0.335 190.670 107.875 190.690 ;
        RECT 0.660 189.850 107.875 190.670 ;
        RECT 0.335 188.990 107.875 189.850 ;
        RECT 0.660 188.170 107.340 188.990 ;
        RECT 0.335 187.310 107.875 188.170 ;
        RECT 0.660 186.490 107.875 187.310 ;
        RECT 0.335 186.470 107.875 186.490 ;
        RECT 0.335 185.650 107.340 186.470 ;
        RECT 0.335 185.630 107.875 185.650 ;
        RECT 0.660 184.810 107.875 185.630 ;
        RECT 0.335 183.950 107.875 184.810 ;
        RECT 0.660 183.130 107.340 183.950 ;
        RECT 0.335 182.270 107.875 183.130 ;
        RECT 0.660 181.450 107.875 182.270 ;
        RECT 0.335 181.430 107.875 181.450 ;
        RECT 0.335 180.610 107.340 181.430 ;
        RECT 0.335 180.590 107.875 180.610 ;
        RECT 0.660 179.770 107.875 180.590 ;
        RECT 0.335 178.910 107.875 179.770 ;
        RECT 0.660 178.090 107.340 178.910 ;
        RECT 0.335 177.230 107.875 178.090 ;
        RECT 0.660 176.410 107.875 177.230 ;
        RECT 0.335 176.390 107.875 176.410 ;
        RECT 0.335 175.570 107.340 176.390 ;
        RECT 0.335 175.550 107.875 175.570 ;
        RECT 0.660 174.730 107.875 175.550 ;
        RECT 0.335 173.870 107.875 174.730 ;
        RECT 0.660 173.050 107.340 173.870 ;
        RECT 0.335 172.190 107.875 173.050 ;
        RECT 0.660 171.370 107.875 172.190 ;
        RECT 0.335 171.350 107.875 171.370 ;
        RECT 0.335 170.530 107.340 171.350 ;
        RECT 0.335 170.510 107.875 170.530 ;
        RECT 0.660 169.690 107.875 170.510 ;
        RECT 0.335 168.830 107.875 169.690 ;
        RECT 0.660 168.010 107.340 168.830 ;
        RECT 0.335 167.150 107.875 168.010 ;
        RECT 0.660 166.330 107.875 167.150 ;
        RECT 0.335 166.310 107.875 166.330 ;
        RECT 0.335 165.490 107.340 166.310 ;
        RECT 0.335 165.470 107.875 165.490 ;
        RECT 0.660 164.650 107.875 165.470 ;
        RECT 0.335 163.790 107.875 164.650 ;
        RECT 0.660 162.970 107.340 163.790 ;
        RECT 0.335 162.110 107.875 162.970 ;
        RECT 0.660 161.290 107.875 162.110 ;
        RECT 0.335 161.270 107.875 161.290 ;
        RECT 0.335 160.450 107.340 161.270 ;
        RECT 0.335 160.430 107.875 160.450 ;
        RECT 0.660 159.610 107.875 160.430 ;
        RECT 0.335 158.750 107.875 159.610 ;
        RECT 0.660 157.930 107.340 158.750 ;
        RECT 0.335 157.070 107.875 157.930 ;
        RECT 0.660 156.250 107.875 157.070 ;
        RECT 0.335 156.230 107.875 156.250 ;
        RECT 0.335 155.410 107.340 156.230 ;
        RECT 0.335 155.390 107.875 155.410 ;
        RECT 0.660 154.570 107.875 155.390 ;
        RECT 0.335 153.710 107.875 154.570 ;
        RECT 0.660 152.890 107.340 153.710 ;
        RECT 0.335 152.030 107.875 152.890 ;
        RECT 0.660 151.210 107.875 152.030 ;
        RECT 0.335 151.190 107.875 151.210 ;
        RECT 0.335 150.370 107.340 151.190 ;
        RECT 0.335 150.350 107.875 150.370 ;
        RECT 0.660 149.530 107.875 150.350 ;
        RECT 0.335 148.670 107.875 149.530 ;
        RECT 0.660 147.850 107.340 148.670 ;
        RECT 0.335 146.990 107.875 147.850 ;
        RECT 0.660 146.170 107.875 146.990 ;
        RECT 0.335 146.150 107.875 146.170 ;
        RECT 0.335 145.330 107.340 146.150 ;
        RECT 0.335 145.310 107.875 145.330 ;
        RECT 0.660 144.490 107.875 145.310 ;
        RECT 0.335 143.630 107.875 144.490 ;
        RECT 0.660 142.810 107.340 143.630 ;
        RECT 0.335 141.950 107.875 142.810 ;
        RECT 0.660 141.130 107.875 141.950 ;
        RECT 0.335 141.110 107.875 141.130 ;
        RECT 0.335 140.290 107.340 141.110 ;
        RECT 0.335 140.270 107.875 140.290 ;
        RECT 0.660 139.450 107.875 140.270 ;
        RECT 0.335 138.590 107.875 139.450 ;
        RECT 0.660 137.770 107.340 138.590 ;
        RECT 0.335 136.910 107.875 137.770 ;
        RECT 0.660 136.090 107.875 136.910 ;
        RECT 0.335 136.070 107.875 136.090 ;
        RECT 0.335 135.250 107.340 136.070 ;
        RECT 0.335 135.230 107.875 135.250 ;
        RECT 0.660 134.410 107.875 135.230 ;
        RECT 0.335 133.550 107.875 134.410 ;
        RECT 0.660 132.730 107.340 133.550 ;
        RECT 0.335 131.870 107.875 132.730 ;
        RECT 0.660 131.050 107.875 131.870 ;
        RECT 0.335 131.030 107.875 131.050 ;
        RECT 0.335 130.210 107.340 131.030 ;
        RECT 0.335 130.190 107.875 130.210 ;
        RECT 0.660 129.370 107.875 130.190 ;
        RECT 0.335 128.510 107.875 129.370 ;
        RECT 0.660 127.690 107.340 128.510 ;
        RECT 0.335 126.830 107.875 127.690 ;
        RECT 0.660 126.010 107.875 126.830 ;
        RECT 0.335 125.990 107.875 126.010 ;
        RECT 0.335 125.170 107.340 125.990 ;
        RECT 0.335 125.150 107.875 125.170 ;
        RECT 0.660 124.330 107.875 125.150 ;
        RECT 0.335 123.470 107.875 124.330 ;
        RECT 0.660 122.650 107.340 123.470 ;
        RECT 0.335 121.790 107.875 122.650 ;
        RECT 0.660 120.970 107.875 121.790 ;
        RECT 0.335 120.950 107.875 120.970 ;
        RECT 0.335 120.130 107.340 120.950 ;
        RECT 0.335 120.110 107.875 120.130 ;
        RECT 0.660 119.290 107.875 120.110 ;
        RECT 0.335 118.430 107.875 119.290 ;
        RECT 0.660 117.610 107.340 118.430 ;
        RECT 0.335 116.750 107.875 117.610 ;
        RECT 0.660 115.930 107.875 116.750 ;
        RECT 0.335 115.910 107.875 115.930 ;
        RECT 0.335 115.090 107.340 115.910 ;
        RECT 0.335 115.070 107.875 115.090 ;
        RECT 0.660 114.250 107.875 115.070 ;
        RECT 0.335 113.390 107.875 114.250 ;
        RECT 0.660 112.570 107.340 113.390 ;
        RECT 0.335 111.710 107.875 112.570 ;
        RECT 0.660 110.890 107.875 111.710 ;
        RECT 0.335 110.870 107.875 110.890 ;
        RECT 0.335 110.050 107.340 110.870 ;
        RECT 0.335 110.030 107.875 110.050 ;
        RECT 0.660 109.210 107.875 110.030 ;
        RECT 0.335 108.350 107.875 109.210 ;
        RECT 0.660 107.530 107.340 108.350 ;
        RECT 0.335 106.670 107.875 107.530 ;
        RECT 0.660 105.850 107.875 106.670 ;
        RECT 0.335 105.830 107.875 105.850 ;
        RECT 0.335 105.010 107.340 105.830 ;
        RECT 0.335 104.990 107.875 105.010 ;
        RECT 0.660 104.170 107.875 104.990 ;
        RECT 0.335 103.310 107.875 104.170 ;
        RECT 0.660 102.490 107.340 103.310 ;
        RECT 0.335 101.630 107.875 102.490 ;
        RECT 0.660 100.810 107.875 101.630 ;
        RECT 0.335 100.790 107.875 100.810 ;
        RECT 0.335 99.970 107.340 100.790 ;
        RECT 0.335 99.950 107.875 99.970 ;
        RECT 0.660 99.130 107.875 99.950 ;
        RECT 0.335 98.270 107.875 99.130 ;
        RECT 0.660 97.450 107.340 98.270 ;
        RECT 0.335 96.590 107.875 97.450 ;
        RECT 0.660 95.770 107.875 96.590 ;
        RECT 0.335 95.750 107.875 95.770 ;
        RECT 0.335 94.930 107.340 95.750 ;
        RECT 0.335 94.910 107.875 94.930 ;
        RECT 0.660 94.090 107.875 94.910 ;
        RECT 0.335 93.230 107.875 94.090 ;
        RECT 0.660 92.410 107.340 93.230 ;
        RECT 0.335 91.550 107.875 92.410 ;
        RECT 0.660 90.730 107.875 91.550 ;
        RECT 0.335 90.710 107.875 90.730 ;
        RECT 0.335 89.890 107.340 90.710 ;
        RECT 0.335 89.870 107.875 89.890 ;
        RECT 0.660 89.050 107.875 89.870 ;
        RECT 0.335 88.190 107.875 89.050 ;
        RECT 0.660 87.370 107.340 88.190 ;
        RECT 0.335 86.510 107.875 87.370 ;
        RECT 0.660 85.690 107.875 86.510 ;
        RECT 0.335 85.670 107.875 85.690 ;
        RECT 0.335 84.850 107.340 85.670 ;
        RECT 0.335 84.830 107.875 84.850 ;
        RECT 0.660 84.010 107.875 84.830 ;
        RECT 0.335 83.150 107.875 84.010 ;
        RECT 0.660 82.330 107.340 83.150 ;
        RECT 0.335 81.470 107.875 82.330 ;
        RECT 0.660 80.650 107.875 81.470 ;
        RECT 0.335 80.630 107.875 80.650 ;
        RECT 0.335 79.810 107.340 80.630 ;
        RECT 0.335 79.790 107.875 79.810 ;
        RECT 0.660 78.970 107.875 79.790 ;
        RECT 0.335 78.110 107.875 78.970 ;
        RECT 0.660 77.290 107.340 78.110 ;
        RECT 0.335 76.430 107.875 77.290 ;
        RECT 0.660 75.610 107.875 76.430 ;
        RECT 0.335 75.590 107.875 75.610 ;
        RECT 0.335 74.770 107.340 75.590 ;
        RECT 0.335 74.750 107.875 74.770 ;
        RECT 0.660 73.930 107.875 74.750 ;
        RECT 0.335 73.070 107.875 73.930 ;
        RECT 0.660 72.250 107.340 73.070 ;
        RECT 0.335 71.390 107.875 72.250 ;
        RECT 0.660 70.570 107.875 71.390 ;
        RECT 0.335 70.550 107.875 70.570 ;
        RECT 0.335 69.730 107.340 70.550 ;
        RECT 0.335 69.710 107.875 69.730 ;
        RECT 0.660 68.890 107.875 69.710 ;
        RECT 0.335 68.030 107.875 68.890 ;
        RECT 0.660 67.210 107.340 68.030 ;
        RECT 0.335 66.350 107.875 67.210 ;
        RECT 0.660 65.530 107.875 66.350 ;
        RECT 0.335 65.510 107.875 65.530 ;
        RECT 0.335 64.690 107.340 65.510 ;
        RECT 0.335 64.670 107.875 64.690 ;
        RECT 0.660 63.850 107.875 64.670 ;
        RECT 0.335 62.990 107.875 63.850 ;
        RECT 0.660 62.170 107.340 62.990 ;
        RECT 0.335 61.310 107.875 62.170 ;
        RECT 0.660 60.490 107.875 61.310 ;
        RECT 0.335 60.470 107.875 60.490 ;
        RECT 0.335 59.650 107.340 60.470 ;
        RECT 0.335 59.630 107.875 59.650 ;
        RECT 0.660 58.810 107.875 59.630 ;
        RECT 0.335 57.950 107.875 58.810 ;
        RECT 0.660 57.130 107.340 57.950 ;
        RECT 0.335 56.270 107.875 57.130 ;
        RECT 0.660 55.450 107.875 56.270 ;
        RECT 0.335 55.430 107.875 55.450 ;
        RECT 0.335 54.610 107.340 55.430 ;
        RECT 0.335 54.590 107.875 54.610 ;
        RECT 0.660 53.770 107.875 54.590 ;
        RECT 0.335 52.910 107.875 53.770 ;
        RECT 0.660 52.090 107.340 52.910 ;
        RECT 0.335 51.230 107.875 52.090 ;
        RECT 0.660 50.410 107.875 51.230 ;
        RECT 0.335 50.390 107.875 50.410 ;
        RECT 0.335 49.570 107.340 50.390 ;
        RECT 0.335 49.550 107.875 49.570 ;
        RECT 0.660 48.730 107.875 49.550 ;
        RECT 0.335 47.870 107.875 48.730 ;
        RECT 0.660 47.050 107.340 47.870 ;
        RECT 0.335 46.190 107.875 47.050 ;
        RECT 0.660 45.370 107.875 46.190 ;
        RECT 0.335 45.350 107.875 45.370 ;
        RECT 0.335 44.530 107.340 45.350 ;
        RECT 0.335 44.510 107.875 44.530 ;
        RECT 0.660 43.690 107.875 44.510 ;
        RECT 0.335 42.830 107.875 43.690 ;
        RECT 0.660 42.010 107.340 42.830 ;
        RECT 0.335 41.150 107.875 42.010 ;
        RECT 0.660 40.330 107.875 41.150 ;
        RECT 0.335 40.310 107.875 40.330 ;
        RECT 0.335 39.490 107.340 40.310 ;
        RECT 0.335 39.470 107.875 39.490 ;
        RECT 0.660 38.650 107.875 39.470 ;
        RECT 0.335 37.790 107.875 38.650 ;
        RECT 0.660 36.970 107.340 37.790 ;
        RECT 0.335 36.110 107.875 36.970 ;
        RECT 0.660 35.290 107.875 36.110 ;
        RECT 0.335 35.270 107.875 35.290 ;
        RECT 0.335 34.450 107.340 35.270 ;
        RECT 0.335 34.430 107.875 34.450 ;
        RECT 0.660 33.610 107.875 34.430 ;
        RECT 0.335 32.750 107.875 33.610 ;
        RECT 0.660 31.930 107.340 32.750 ;
        RECT 0.335 31.070 107.875 31.930 ;
        RECT 0.660 30.250 107.875 31.070 ;
        RECT 0.335 30.230 107.875 30.250 ;
        RECT 0.335 29.410 107.340 30.230 ;
        RECT 0.335 29.390 107.875 29.410 ;
        RECT 0.660 28.570 107.875 29.390 ;
        RECT 0.335 27.710 107.875 28.570 ;
        RECT 0.660 26.890 107.340 27.710 ;
        RECT 0.335 26.030 107.875 26.890 ;
        RECT 0.660 25.210 107.875 26.030 ;
        RECT 0.335 25.190 107.875 25.210 ;
        RECT 0.335 24.370 107.340 25.190 ;
        RECT 0.335 24.350 107.875 24.370 ;
        RECT 0.660 23.530 107.875 24.350 ;
        RECT 0.335 22.670 107.875 23.530 ;
        RECT 0.660 21.850 107.340 22.670 ;
        RECT 0.335 20.990 107.875 21.850 ;
        RECT 0.660 20.170 107.875 20.990 ;
        RECT 0.335 20.150 107.875 20.170 ;
        RECT 0.335 19.330 107.340 20.150 ;
        RECT 0.335 19.310 107.875 19.330 ;
        RECT 0.660 18.490 107.875 19.310 ;
        RECT 0.335 17.630 107.875 18.490 ;
        RECT 0.660 16.810 107.875 17.630 ;
        RECT 0.335 15.950 107.875 16.810 ;
        RECT 0.660 15.130 107.875 15.950 ;
        RECT 0.335 14.270 107.875 15.130 ;
        RECT 0.660 13.450 107.875 14.270 ;
        RECT 0.335 7.460 107.875 13.450 ;
      LAYER Metal3 ;
        RECT 0.380 483.230 8.710 483.440 ;
        RECT 9.530 483.230 9.670 483.440 ;
        RECT 10.490 483.230 10.630 483.440 ;
        RECT 11.450 483.230 11.590 483.440 ;
        RECT 12.410 483.230 12.550 483.440 ;
        RECT 13.370 483.230 13.510 483.440 ;
        RECT 14.330 483.230 14.470 483.440 ;
        RECT 15.290 483.230 15.430 483.440 ;
        RECT 16.250 483.230 16.390 483.440 ;
        RECT 17.210 483.230 17.350 483.440 ;
        RECT 18.170 483.230 18.310 483.440 ;
        RECT 19.130 483.230 19.270 483.440 ;
        RECT 20.090 483.230 20.230 483.440 ;
        RECT 21.050 483.230 21.190 483.440 ;
        RECT 22.010 483.230 22.150 483.440 ;
        RECT 22.970 483.230 23.110 483.440 ;
        RECT 23.930 483.230 24.070 483.440 ;
        RECT 24.890 483.230 25.030 483.440 ;
        RECT 25.850 483.230 25.990 483.440 ;
        RECT 26.810 483.230 26.950 483.440 ;
        RECT 27.770 483.230 27.910 483.440 ;
        RECT 28.730 483.230 28.870 483.440 ;
        RECT 29.690 483.230 29.830 483.440 ;
        RECT 30.650 483.230 30.790 483.440 ;
        RECT 31.610 483.230 31.750 483.440 ;
        RECT 32.570 483.230 32.710 483.440 ;
        RECT 33.530 483.230 33.670 483.440 ;
        RECT 34.490 483.230 34.630 483.440 ;
        RECT 35.450 483.230 35.590 483.440 ;
        RECT 36.410 483.230 36.550 483.440 ;
        RECT 37.370 483.230 37.510 483.440 ;
        RECT 38.330 483.230 38.470 483.440 ;
        RECT 39.290 483.230 39.430 483.440 ;
        RECT 40.250 483.230 40.390 483.440 ;
        RECT 41.210 483.230 41.350 483.440 ;
        RECT 42.170 483.230 42.310 483.440 ;
        RECT 43.130 483.230 43.270 483.440 ;
        RECT 44.090 483.230 44.230 483.440 ;
        RECT 45.050 483.230 45.190 483.440 ;
        RECT 46.010 483.230 46.150 483.440 ;
        RECT 46.970 483.230 47.110 483.440 ;
        RECT 47.930 483.230 48.070 483.440 ;
        RECT 48.890 483.230 49.030 483.440 ;
        RECT 49.850 483.230 49.990 483.440 ;
        RECT 50.810 483.230 50.950 483.440 ;
        RECT 51.770 483.230 51.910 483.440 ;
        RECT 52.730 483.230 52.870 483.440 ;
        RECT 53.690 483.230 53.830 483.440 ;
        RECT 54.650 483.230 54.790 483.440 ;
        RECT 55.610 483.230 55.750 483.440 ;
        RECT 56.570 483.230 56.710 483.440 ;
        RECT 57.530 483.230 57.670 483.440 ;
        RECT 58.490 483.230 58.630 483.440 ;
        RECT 59.450 483.230 59.590 483.440 ;
        RECT 60.410 483.230 60.550 483.440 ;
        RECT 61.370 483.230 61.510 483.440 ;
        RECT 62.330 483.230 62.470 483.440 ;
        RECT 63.290 483.230 63.430 483.440 ;
        RECT 64.250 483.230 64.390 483.440 ;
        RECT 65.210 483.230 65.350 483.440 ;
        RECT 66.170 483.230 66.310 483.440 ;
        RECT 67.130 483.230 67.270 483.440 ;
        RECT 68.090 483.230 68.230 483.440 ;
        RECT 69.050 483.230 69.190 483.440 ;
        RECT 70.010 483.230 70.150 483.440 ;
        RECT 70.970 483.230 71.110 483.440 ;
        RECT 71.930 483.230 72.070 483.440 ;
        RECT 72.890 483.230 73.030 483.440 ;
        RECT 73.850 483.230 73.990 483.440 ;
        RECT 74.810 483.230 74.950 483.440 ;
        RECT 75.770 483.230 75.910 483.440 ;
        RECT 76.730 483.230 76.870 483.440 ;
        RECT 77.690 483.230 77.830 483.440 ;
        RECT 78.650 483.230 78.790 483.440 ;
        RECT 79.610 483.230 79.750 483.440 ;
        RECT 80.570 483.230 80.710 483.440 ;
        RECT 81.530 483.230 81.670 483.440 ;
        RECT 82.490 483.230 82.630 483.440 ;
        RECT 83.450 483.230 83.590 483.440 ;
        RECT 84.410 483.230 84.550 483.440 ;
        RECT 85.370 483.230 85.510 483.440 ;
        RECT 86.330 483.230 86.470 483.440 ;
        RECT 87.290 483.230 87.430 483.440 ;
        RECT 88.250 483.230 88.390 483.440 ;
        RECT 89.210 483.230 89.350 483.440 ;
        RECT 90.170 483.230 90.310 483.440 ;
        RECT 91.130 483.230 91.270 483.440 ;
        RECT 92.090 483.230 92.230 483.440 ;
        RECT 93.050 483.230 93.190 483.440 ;
        RECT 94.010 483.230 94.150 483.440 ;
        RECT 94.970 483.230 95.110 483.440 ;
        RECT 95.930 483.230 96.070 483.440 ;
        RECT 96.890 483.230 97.030 483.440 ;
        RECT 97.850 483.230 107.620 483.440 ;
        RECT 0.380 0.610 107.620 483.230 ;
        RECT 0.380 0.400 8.710 0.610 ;
        RECT 9.530 0.400 9.670 0.610 ;
        RECT 10.490 0.400 10.630 0.610 ;
        RECT 11.450 0.400 11.590 0.610 ;
        RECT 12.410 0.400 12.550 0.610 ;
        RECT 13.370 0.400 13.510 0.610 ;
        RECT 14.330 0.400 14.470 0.610 ;
        RECT 15.290 0.400 15.430 0.610 ;
        RECT 16.250 0.400 16.390 0.610 ;
        RECT 17.210 0.400 17.350 0.610 ;
        RECT 18.170 0.400 18.310 0.610 ;
        RECT 19.130 0.400 19.270 0.610 ;
        RECT 20.090 0.400 20.230 0.610 ;
        RECT 21.050 0.400 21.190 0.610 ;
        RECT 22.010 0.400 22.150 0.610 ;
        RECT 22.970 0.400 23.110 0.610 ;
        RECT 23.930 0.400 24.070 0.610 ;
        RECT 24.890 0.400 25.030 0.610 ;
        RECT 25.850 0.400 25.990 0.610 ;
        RECT 26.810 0.400 26.950 0.610 ;
        RECT 27.770 0.400 27.910 0.610 ;
        RECT 28.730 0.400 28.870 0.610 ;
        RECT 29.690 0.400 29.830 0.610 ;
        RECT 30.650 0.400 30.790 0.610 ;
        RECT 31.610 0.400 31.750 0.610 ;
        RECT 32.570 0.400 32.710 0.610 ;
        RECT 33.530 0.400 33.670 0.610 ;
        RECT 34.490 0.400 34.630 0.610 ;
        RECT 35.450 0.400 35.590 0.610 ;
        RECT 36.410 0.400 36.550 0.610 ;
        RECT 37.370 0.400 37.510 0.610 ;
        RECT 38.330 0.400 38.470 0.610 ;
        RECT 39.290 0.400 39.430 0.610 ;
        RECT 40.250 0.400 40.390 0.610 ;
        RECT 41.210 0.400 41.350 0.610 ;
        RECT 42.170 0.400 42.310 0.610 ;
        RECT 43.130 0.400 43.270 0.610 ;
        RECT 44.090 0.400 44.230 0.610 ;
        RECT 45.050 0.400 45.190 0.610 ;
        RECT 46.010 0.400 46.150 0.610 ;
        RECT 46.970 0.400 47.110 0.610 ;
        RECT 47.930 0.400 48.070 0.610 ;
        RECT 48.890 0.400 49.030 0.610 ;
        RECT 49.850 0.400 49.990 0.610 ;
        RECT 50.810 0.400 50.950 0.610 ;
        RECT 51.770 0.400 51.910 0.610 ;
        RECT 52.730 0.400 52.870 0.610 ;
        RECT 53.690 0.400 53.830 0.610 ;
        RECT 54.650 0.400 54.790 0.610 ;
        RECT 55.610 0.400 55.750 0.610 ;
        RECT 56.570 0.400 56.710 0.610 ;
        RECT 57.530 0.400 57.670 0.610 ;
        RECT 58.490 0.400 58.630 0.610 ;
        RECT 59.450 0.400 59.590 0.610 ;
        RECT 60.410 0.400 60.550 0.610 ;
        RECT 61.370 0.400 61.510 0.610 ;
        RECT 62.330 0.400 62.470 0.610 ;
        RECT 63.290 0.400 63.430 0.610 ;
        RECT 64.250 0.400 64.390 0.610 ;
        RECT 65.210 0.400 65.350 0.610 ;
        RECT 66.170 0.400 66.310 0.610 ;
        RECT 67.130 0.400 67.270 0.610 ;
        RECT 68.090 0.400 68.230 0.610 ;
        RECT 69.050 0.400 69.190 0.610 ;
        RECT 70.010 0.400 70.150 0.610 ;
        RECT 70.970 0.400 71.110 0.610 ;
        RECT 71.930 0.400 72.070 0.610 ;
        RECT 72.890 0.400 73.030 0.610 ;
        RECT 73.850 0.400 73.990 0.610 ;
        RECT 74.810 0.400 74.950 0.610 ;
        RECT 75.770 0.400 75.910 0.610 ;
        RECT 76.730 0.400 76.870 0.610 ;
        RECT 77.690 0.400 77.830 0.610 ;
        RECT 78.650 0.400 78.790 0.610 ;
        RECT 79.610 0.400 79.750 0.610 ;
        RECT 80.570 0.400 80.710 0.610 ;
        RECT 81.530 0.400 81.670 0.610 ;
        RECT 82.490 0.400 82.630 0.610 ;
        RECT 83.450 0.400 83.590 0.610 ;
        RECT 84.410 0.400 84.550 0.610 ;
        RECT 85.370 0.400 85.510 0.610 ;
        RECT 86.330 0.400 86.470 0.610 ;
        RECT 87.290 0.400 87.430 0.610 ;
        RECT 88.250 0.400 88.390 0.610 ;
        RECT 89.210 0.400 89.350 0.610 ;
        RECT 90.170 0.400 90.310 0.610 ;
        RECT 91.130 0.400 91.270 0.610 ;
        RECT 92.090 0.400 92.230 0.610 ;
        RECT 93.050 0.400 93.190 0.610 ;
        RECT 94.010 0.400 94.150 0.610 ;
        RECT 94.970 0.400 95.110 0.610 ;
        RECT 95.930 0.400 96.070 0.610 ;
        RECT 96.890 0.400 97.030 0.610 ;
        RECT 97.850 0.400 107.620 0.610 ;
      LAYER Metal4 ;
        RECT 0.335 0.740 107.665 483.100 ;
      LAYER Metal5 ;
        RECT 1.820 0.695 18.050 483.145 ;
        RECT 20.670 0.695 24.250 483.145 ;
        RECT 26.870 0.695 93.650 483.145 ;
        RECT 96.270 0.695 99.850 483.145 ;
        RECT 102.470 0.695 107.620 483.145 ;
  END
END IHP_SRAM
END LIBRARY

