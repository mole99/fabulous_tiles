VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 205.000 BY 56.250 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 0.280 ;
    END
  END Ci
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 0.600 7.440 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 0.600 21.040 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 0.600 22.400 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 0.600 23.760 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 0.600 25.120 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 0.600 26.480 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 0.600 27.840 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.600 29.200 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 0.600 30.560 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 0.600 31.920 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 0.600 33.280 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 0.600 8.800 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 0.600 34.640 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.600 36.000 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 0.600 37.360 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 0.600 38.720 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 0.600 40.080 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 0.600 41.440 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.600 42.800 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 0.600 44.160 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 0.600 45.520 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 0.600 46.880 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 0.600 10.160 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.600 48.240 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.600 49.600 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 0.600 11.520 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 0.600 12.880 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 0.600 14.240 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 0.600 15.600 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 0.600 16.960 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 0.600 18.320 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 0.600 19.680 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 6.840 205.000 7.440 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 20.440 205.000 21.040 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 21.800 205.000 22.400 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 23.160 205.000 23.760 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 24.520 205.000 25.120 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 25.880 205.000 26.480 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 27.240 205.000 27.840 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 28.600 205.000 29.200 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 29.960 205.000 30.560 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 31.320 205.000 31.920 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 32.680 205.000 33.280 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 8.200 205.000 8.800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 34.040 205.000 34.640 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 35.400 205.000 36.000 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 36.760 205.000 37.360 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 38.120 205.000 38.720 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 39.480 205.000 40.080 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 40.840 205.000 41.440 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 42.200 205.000 42.800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 43.560 205.000 44.160 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 44.920 205.000 45.520 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 46.280 205.000 46.880 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 9.560 205.000 10.160 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 47.640 205.000 48.240 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 49.000 205.000 49.600 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 10.920 205.000 11.520 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 12.280 205.000 12.880 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 13.640 205.000 14.240 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 15.000 205.000 15.600 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 16.360 205.000 16.960 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 17.720 205.000 18.320 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 204.400 19.080 205.000 19.680 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 0.280 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 0.280 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 0.280 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 0.280 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 0.280 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 0.280 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 0.280 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 0.280 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 0.280 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 0.280 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 0.280 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 0.280 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 0.280 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 0.280 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 0.280 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 0.280 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 0.280 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 0.280 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 0.280 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 0.280 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 15.270 55.970 15.550 56.250 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.870 55.970 112.150 56.250 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.530 55.970 121.810 56.250 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 131.190 55.970 131.470 56.250 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.850 55.970 141.130 56.250 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.510 55.970 150.790 56.250 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.170 55.970 160.450 56.250 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 169.830 55.970 170.110 56.250 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 179.490 55.970 179.770 56.250 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 189.150 55.970 189.430 56.250 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 198.810 55.970 199.090 56.250 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.930 55.970 25.210 56.250 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 34.590 55.970 34.870 56.250 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 55.970 44.530 56.250 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.910 55.970 54.190 56.250 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 63.570 55.970 63.850 56.250 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.230 55.970 73.510 56.250 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.890 55.970 83.170 56.250 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.550 55.970 92.830 56.250 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.210 55.970 102.490 56.250 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 0.280 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 0.280 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 0.280 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 0.280 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 0.280 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 0.280 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.280 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 0.280 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.280 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.280 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 0.280 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 0.280 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 0.280 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 0.280 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 0.280 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 0.280 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 0.280 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 0.280 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 0.280 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 0.280 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.280 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 0.280 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.280 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 0.280 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 0.280 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 0.280 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 0.280 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 0.280 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 0.280 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 0.280 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 0.280 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 0.280 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 0.280 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 0.280 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 0.280 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 0.280 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 0.280 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 0.280 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 0.280 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 0.280 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 0.280 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 0.280 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 0.280 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 0.280 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 0.280 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 0.280 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 0.280 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 0.280 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 0.280 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 0.280 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 0.280 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 0.280 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 0.280 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 0.280 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 0.280 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 0.280 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 0.280 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 0.280 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 0.280 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 0.280 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 0.280 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 0.280 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 0.280 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 0.280 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 0.280 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 0.280 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 0.280 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 0.280 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 0.280 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 0.280 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 0.280 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 0.280 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 0.280 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 0.280 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 0.280 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 0.280 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.870 0.000 135.150 0.280 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 0.280 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 0.280 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 0.280 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 0.280 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 0.280 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 0.280 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 0.280 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 0.280 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 0.280 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 0.280 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 0.280 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 0.280 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 0.280 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 0.280 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 0.280 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 0.280 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 0.280 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 0.280 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 0.280 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 0.280 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 0.280 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 0.280 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 0.280 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 0.280 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 0.280 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 0.280 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 0.280 ;
    END
  END SS4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 0.280 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 5.610 55.970 5.890 56.250 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 0.000 16.620 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.020 0.000 46.620 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.020 0.000 76.620 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 105.020 0.000 106.620 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.020 0.000 136.620 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 165.020 0.000 166.620 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 195.020 0.000 196.620 56.250 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 0.000 11.320 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.720 0.000 41.320 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.720 0.000 71.320 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.720 0.000 101.320 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.720 0.000 131.320 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 0.000 161.320 56.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 0.000 191.320 56.250 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 199.370 43.605 ;
      LAYER li1 ;
        RECT 5.520 10.795 199.180 43.605 ;
      LAYER met1 ;
        RECT 2.830 0.040 202.330 46.880 ;
      LAYER met2 ;
        RECT 2.850 55.690 5.330 55.970 ;
        RECT 6.170 55.690 14.990 55.970 ;
        RECT 15.830 55.690 24.650 55.970 ;
        RECT 25.490 55.690 34.310 55.970 ;
        RECT 35.150 55.690 43.970 55.970 ;
        RECT 44.810 55.690 53.630 55.970 ;
        RECT 54.470 55.690 63.290 55.970 ;
        RECT 64.130 55.690 72.950 55.970 ;
        RECT 73.790 55.690 82.610 55.970 ;
        RECT 83.450 55.690 92.270 55.970 ;
        RECT 93.110 55.690 101.930 55.970 ;
        RECT 102.770 55.690 111.590 55.970 ;
        RECT 112.430 55.690 121.250 55.970 ;
        RECT 122.090 55.690 130.910 55.970 ;
        RECT 131.750 55.690 140.570 55.970 ;
        RECT 141.410 55.690 150.230 55.970 ;
        RECT 151.070 55.690 159.890 55.970 ;
        RECT 160.730 55.690 169.550 55.970 ;
        RECT 170.390 55.690 179.210 55.970 ;
        RECT 180.050 55.690 188.870 55.970 ;
        RECT 189.710 55.690 198.530 55.970 ;
        RECT 199.370 55.690 202.310 55.970 ;
        RECT 2.850 0.560 202.310 55.690 ;
        RECT 2.850 0.010 15.910 0.560 ;
        RECT 16.750 0.010 17.290 0.560 ;
        RECT 18.130 0.010 18.670 0.560 ;
        RECT 19.510 0.010 20.050 0.560 ;
        RECT 20.890 0.010 21.430 0.560 ;
        RECT 22.270 0.010 22.810 0.560 ;
        RECT 23.650 0.010 24.190 0.560 ;
        RECT 25.030 0.010 25.570 0.560 ;
        RECT 26.410 0.010 26.950 0.560 ;
        RECT 27.790 0.010 28.330 0.560 ;
        RECT 29.170 0.010 29.710 0.560 ;
        RECT 30.550 0.010 31.090 0.560 ;
        RECT 31.930 0.010 32.470 0.560 ;
        RECT 33.310 0.010 33.850 0.560 ;
        RECT 34.690 0.010 35.230 0.560 ;
        RECT 36.070 0.010 36.610 0.560 ;
        RECT 37.450 0.010 37.990 0.560 ;
        RECT 38.830 0.010 39.370 0.560 ;
        RECT 40.210 0.010 40.750 0.560 ;
        RECT 41.590 0.010 42.130 0.560 ;
        RECT 42.970 0.010 43.510 0.560 ;
        RECT 44.350 0.010 44.890 0.560 ;
        RECT 45.730 0.010 46.270 0.560 ;
        RECT 47.110 0.010 47.650 0.560 ;
        RECT 48.490 0.010 49.030 0.560 ;
        RECT 49.870 0.010 50.410 0.560 ;
        RECT 51.250 0.010 51.790 0.560 ;
        RECT 52.630 0.010 53.170 0.560 ;
        RECT 54.010 0.010 54.550 0.560 ;
        RECT 55.390 0.010 55.930 0.560 ;
        RECT 56.770 0.010 57.310 0.560 ;
        RECT 58.150 0.010 58.690 0.560 ;
        RECT 59.530 0.010 60.070 0.560 ;
        RECT 60.910 0.010 61.450 0.560 ;
        RECT 62.290 0.010 62.830 0.560 ;
        RECT 63.670 0.010 64.210 0.560 ;
        RECT 65.050 0.010 65.590 0.560 ;
        RECT 66.430 0.010 66.970 0.560 ;
        RECT 67.810 0.010 68.350 0.560 ;
        RECT 69.190 0.010 69.730 0.560 ;
        RECT 70.570 0.010 71.110 0.560 ;
        RECT 71.950 0.010 72.490 0.560 ;
        RECT 73.330 0.010 73.870 0.560 ;
        RECT 74.710 0.010 75.250 0.560 ;
        RECT 76.090 0.010 76.630 0.560 ;
        RECT 77.470 0.010 78.010 0.560 ;
        RECT 78.850 0.010 79.390 0.560 ;
        RECT 80.230 0.010 80.770 0.560 ;
        RECT 81.610 0.010 82.150 0.560 ;
        RECT 82.990 0.010 83.530 0.560 ;
        RECT 84.370 0.010 84.910 0.560 ;
        RECT 85.750 0.010 86.290 0.560 ;
        RECT 87.130 0.010 87.670 0.560 ;
        RECT 88.510 0.010 89.050 0.560 ;
        RECT 89.890 0.010 90.430 0.560 ;
        RECT 91.270 0.010 91.810 0.560 ;
        RECT 92.650 0.010 93.190 0.560 ;
        RECT 94.030 0.010 94.570 0.560 ;
        RECT 95.410 0.010 95.950 0.560 ;
        RECT 96.790 0.010 97.330 0.560 ;
        RECT 98.170 0.010 98.710 0.560 ;
        RECT 99.550 0.010 100.090 0.560 ;
        RECT 100.930 0.010 101.470 0.560 ;
        RECT 102.310 0.010 102.850 0.560 ;
        RECT 103.690 0.010 104.230 0.560 ;
        RECT 105.070 0.010 105.610 0.560 ;
        RECT 106.450 0.010 106.990 0.560 ;
        RECT 107.830 0.010 108.370 0.560 ;
        RECT 109.210 0.010 109.750 0.560 ;
        RECT 110.590 0.010 111.130 0.560 ;
        RECT 111.970 0.010 112.510 0.560 ;
        RECT 113.350 0.010 113.890 0.560 ;
        RECT 114.730 0.010 115.270 0.560 ;
        RECT 116.110 0.010 116.650 0.560 ;
        RECT 117.490 0.010 118.030 0.560 ;
        RECT 118.870 0.010 119.410 0.560 ;
        RECT 120.250 0.010 120.790 0.560 ;
        RECT 121.630 0.010 122.170 0.560 ;
        RECT 123.010 0.010 123.550 0.560 ;
        RECT 124.390 0.010 124.930 0.560 ;
        RECT 125.770 0.010 126.310 0.560 ;
        RECT 127.150 0.010 127.690 0.560 ;
        RECT 128.530 0.010 129.070 0.560 ;
        RECT 129.910 0.010 130.450 0.560 ;
        RECT 131.290 0.010 131.830 0.560 ;
        RECT 132.670 0.010 133.210 0.560 ;
        RECT 134.050 0.010 134.590 0.560 ;
        RECT 135.430 0.010 135.970 0.560 ;
        RECT 136.810 0.010 137.350 0.560 ;
        RECT 138.190 0.010 138.730 0.560 ;
        RECT 139.570 0.010 140.110 0.560 ;
        RECT 140.950 0.010 141.490 0.560 ;
        RECT 142.330 0.010 142.870 0.560 ;
        RECT 143.710 0.010 144.250 0.560 ;
        RECT 145.090 0.010 145.630 0.560 ;
        RECT 146.470 0.010 147.010 0.560 ;
        RECT 147.850 0.010 148.390 0.560 ;
        RECT 149.230 0.010 149.770 0.560 ;
        RECT 150.610 0.010 151.150 0.560 ;
        RECT 151.990 0.010 152.530 0.560 ;
        RECT 153.370 0.010 153.910 0.560 ;
        RECT 154.750 0.010 155.290 0.560 ;
        RECT 156.130 0.010 156.670 0.560 ;
        RECT 157.510 0.010 158.050 0.560 ;
        RECT 158.890 0.010 159.430 0.560 ;
        RECT 160.270 0.010 160.810 0.560 ;
        RECT 161.650 0.010 162.190 0.560 ;
        RECT 163.030 0.010 163.570 0.560 ;
        RECT 164.410 0.010 164.950 0.560 ;
        RECT 165.790 0.010 166.330 0.560 ;
        RECT 167.170 0.010 167.710 0.560 ;
        RECT 168.550 0.010 169.090 0.560 ;
        RECT 169.930 0.010 170.470 0.560 ;
        RECT 171.310 0.010 171.850 0.560 ;
        RECT 172.690 0.010 173.230 0.560 ;
        RECT 174.070 0.010 174.610 0.560 ;
        RECT 175.450 0.010 175.990 0.560 ;
        RECT 176.830 0.010 177.370 0.560 ;
        RECT 178.210 0.010 178.750 0.560 ;
        RECT 179.590 0.010 180.130 0.560 ;
        RECT 180.970 0.010 181.510 0.560 ;
        RECT 182.350 0.010 182.890 0.560 ;
        RECT 183.730 0.010 184.270 0.560 ;
        RECT 185.110 0.010 185.650 0.560 ;
        RECT 186.490 0.010 187.030 0.560 ;
        RECT 187.870 0.010 188.410 0.560 ;
        RECT 189.250 0.010 202.310 0.560 ;
      LAYER met3 ;
        RECT 1.000 6.440 204.000 49.465 ;
        RECT 0.600 0.175 204.400 6.440 ;
  END
END N_term_single
END LIBRARY

