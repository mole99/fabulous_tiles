magic
tech sky130A
magscale 1 2
timestamp 1740383690
<< viali >>
rect 2513 8585 2547 8619
rect 2789 8585 2823 8619
rect 3433 8585 3467 8619
rect 4169 8585 4203 8619
rect 4537 8585 4571 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7113 8585 7147 8619
rect 7849 8585 7883 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 9321 8585 9355 8619
rect 10057 8585 10091 8619
rect 10517 8585 10551 8619
rect 10885 8585 10919 8619
rect 11161 8585 11195 8619
rect 11989 8585 12023 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 13369 8585 13403 8619
rect 13737 8585 13771 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15301 8585 15335 8619
rect 15577 8585 15611 8619
rect 15945 8585 15979 8619
rect 16405 8585 16439 8619
rect 16957 8585 16991 8619
rect 22017 8585 22051 8619
rect 23121 8585 23155 8619
rect 25513 8585 25547 8619
rect 25789 8585 25823 8619
rect 27905 8585 27939 8619
rect 28733 8585 28767 8619
rect 30573 8585 30607 8619
rect 32321 8585 32355 8619
rect 32781 8585 32815 8619
rect 33425 8585 33459 8619
rect 33885 8585 33919 8619
rect 34805 8585 34839 8619
rect 35173 8585 35207 8619
rect 36737 8585 36771 8619
rect 37841 8585 37875 8619
rect 38577 8585 38611 8619
rect 30665 8517 30699 8551
rect 2329 8449 2363 8483
rect 2605 8449 2639 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10333 8449 10367 8483
rect 10701 8449 10735 8483
rect 11345 8449 11379 8483
rect 11805 8449 11839 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13553 8449 13587 8483
rect 13921 8449 13955 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15117 8449 15151 8483
rect 15761 8449 15795 8483
rect 16129 8449 16163 8483
rect 16221 8449 16255 8483
rect 17141 8449 17175 8483
rect 17693 8449 17727 8483
rect 18061 8449 18095 8483
rect 18337 8449 18371 8483
rect 18797 8449 18831 8483
rect 18889 8449 18923 8483
rect 19349 8449 19383 8483
rect 19625 8449 19659 8483
rect 20085 8449 20119 8483
rect 21281 8449 21315 8483
rect 21833 8449 21867 8483
rect 22109 8449 22143 8483
rect 22569 8449 22603 8483
rect 22661 8449 22695 8483
rect 22937 8449 22971 8483
rect 23213 8449 23247 8483
rect 23673 8449 23707 8483
rect 23949 8449 23983 8483
rect 24041 8449 24075 8483
rect 24593 8449 24627 8483
rect 24869 8449 24903 8483
rect 25145 8449 25179 8483
rect 25237 8449 25271 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 28089 8449 28123 8483
rect 28181 8449 28215 8483
rect 28641 8449 28675 8483
rect 28917 8449 28951 8483
rect 29193 8449 29227 8483
rect 32505 8449 32539 8483
rect 32597 8449 32631 8483
rect 32965 8449 32999 8483
rect 33609 8449 33643 8483
rect 33701 8449 33735 8483
rect 34345 8449 34379 8483
rect 34989 8449 35023 8483
rect 35357 8449 35391 8483
rect 35449 8449 35483 8483
rect 35817 8449 35851 8483
rect 36185 8449 36219 8483
rect 36553 8449 36587 8483
rect 37289 8449 37323 8483
rect 37657 8449 37691 8483
rect 38025 8449 38059 8483
rect 38393 8449 38427 8483
rect 38853 8449 38887 8483
rect 39221 8449 39255 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 29561 8381 29595 8415
rect 29837 8381 29871 8415
rect 3065 8313 3099 8347
rect 4905 8313 4939 8347
rect 5273 8313 5307 8347
rect 7481 8313 7515 8347
rect 9689 8313 9723 8347
rect 17509 8313 17543 8347
rect 17877 8313 17911 8347
rect 19809 8313 19843 8347
rect 21465 8313 21499 8347
rect 22845 8313 22879 8347
rect 23765 8313 23799 8347
rect 24409 8313 24443 8347
rect 24685 8313 24719 8347
rect 28365 8313 28399 8347
rect 33149 8313 33183 8347
rect 34161 8313 34195 8347
rect 35633 8313 35667 8347
rect 36001 8313 36035 8347
rect 38209 8313 38243 8347
rect 39037 8313 39071 8347
rect 39405 8313 39439 8347
rect 18521 8245 18555 8279
rect 18613 8245 18647 8279
rect 19073 8245 19107 8279
rect 19533 8245 19567 8279
rect 19901 8245 19935 8279
rect 22293 8245 22327 8279
rect 22385 8245 22419 8279
rect 23397 8245 23431 8279
rect 23489 8245 23523 8279
rect 24225 8245 24259 8279
rect 24961 8245 24995 8279
rect 25421 8245 25455 8279
rect 28457 8245 28491 8279
rect 29009 8245 29043 8279
rect 36369 8245 36403 8279
rect 37473 8245 37507 8279
rect 2145 8041 2179 8075
rect 3433 8041 3467 8075
rect 4261 8041 4295 8075
rect 4813 8041 4847 8075
rect 5365 8041 5399 8075
rect 6745 8041 6779 8075
rect 7297 8041 7331 8075
rect 7849 8041 7883 8075
rect 8401 8041 8435 8075
rect 9045 8041 9079 8075
rect 9505 8041 9539 8075
rect 10057 8041 10091 8075
rect 11437 8041 11471 8075
rect 11989 8041 12023 8075
rect 12817 8041 12851 8075
rect 14105 8041 14139 8075
rect 14473 8041 14507 8075
rect 15025 8041 15059 8075
rect 15301 8041 15335 8075
rect 16129 8041 16163 8075
rect 17509 8041 17543 8075
rect 23029 8041 23063 8075
rect 24409 8041 24443 8075
rect 34805 8041 34839 8075
rect 35725 8041 35759 8075
rect 36277 8041 36311 8075
rect 36921 8041 36955 8075
rect 38669 8041 38703 8075
rect 8585 7973 8619 8007
rect 10333 7973 10367 8007
rect 10793 7973 10827 8007
rect 21557 7973 21591 8007
rect 22201 7973 22235 8007
rect 29561 7973 29595 8007
rect 33057 7973 33091 8007
rect 38393 7973 38427 8007
rect 19901 7905 19935 7939
rect 23581 7905 23615 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 2789 7837 2823 7871
rect 3617 7837 3651 7871
rect 4445 7837 4479 7871
rect 4997 7837 5031 7871
rect 5549 7837 5583 7871
rect 6929 7837 6963 7871
rect 7481 7837 7515 7871
rect 8033 7837 8067 7871
rect 8309 7837 8343 7871
rect 8769 7837 8803 7871
rect 9229 7837 9263 7871
rect 9689 7837 9723 7871
rect 10241 7837 10275 7871
rect 11621 7837 11655 7871
rect 12173 7837 12207 7871
rect 13001 7837 13035 7871
rect 13829 7837 13863 7871
rect 14289 7837 14323 7871
rect 14657 7837 14691 7871
rect 15209 7837 15243 7871
rect 15485 7837 15519 7871
rect 16313 7837 16347 7871
rect 17601 7837 17635 7871
rect 17877 7837 17911 7871
rect 18153 7837 18187 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 19717 7837 19751 7871
rect 20453 7837 20487 7871
rect 20546 7837 20580 7871
rect 20918 7837 20952 7871
rect 21373 7837 21407 7871
rect 21649 7837 21683 7871
rect 21985 7837 22019 7871
rect 22109 7837 22143 7871
rect 22385 7837 22419 7871
rect 23489 7837 23523 7871
rect 24041 7837 24075 7871
rect 24593 7837 24627 7871
rect 25697 7837 25731 7871
rect 27077 7837 27111 7871
rect 28733 7837 28767 7871
rect 29009 7837 29043 7871
rect 29101 7837 29135 7871
rect 29745 7837 29779 7871
rect 32137 7837 32171 7871
rect 32781 7837 32815 7871
rect 32873 7837 32907 7871
rect 33149 7837 33183 7871
rect 33425 7837 33459 7871
rect 34989 7837 35023 7871
rect 35265 7837 35299 7871
rect 35909 7837 35943 7871
rect 36461 7837 36495 7871
rect 36737 7837 36771 7871
rect 38117 7837 38151 7871
rect 38209 7837 38243 7871
rect 38485 7837 38519 7871
rect 39221 7837 39255 7871
rect 5917 7769 5951 7803
rect 6285 7769 6319 7803
rect 6469 7769 6503 7803
rect 10425 7769 10459 7803
rect 10609 7769 10643 7803
rect 20729 7769 20763 7803
rect 20821 7769 20855 7803
rect 21741 7769 21775 7803
rect 39129 7769 39163 7803
rect 1593 7701 1627 7735
rect 1869 7701 1903 7735
rect 2421 7701 2455 7735
rect 2697 7701 2731 7735
rect 2973 7701 3007 7735
rect 6009 7701 6043 7735
rect 13645 7701 13679 7735
rect 17785 7701 17819 7735
rect 18889 7701 18923 7735
rect 21097 7701 21131 7735
rect 21189 7701 21223 7735
rect 23397 7701 23431 7735
rect 23857 7701 23891 7735
rect 25513 7701 25547 7735
rect 27261 7701 27295 7735
rect 28549 7701 28583 7735
rect 29009 7701 29043 7735
rect 29285 7701 29319 7735
rect 31953 7701 31987 7735
rect 32781 7701 32815 7735
rect 33333 7701 33367 7735
rect 33517 7701 33551 7735
rect 35081 7701 35115 7735
rect 38025 7701 38059 7735
rect 39405 7701 39439 7735
rect 1593 7497 1627 7531
rect 14933 7497 14967 7531
rect 20913 7497 20947 7531
rect 38301 7497 38335 7531
rect 38669 7497 38703 7531
rect 39037 7497 39071 7531
rect 39405 7497 39439 7531
rect 30021 7429 30055 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 7757 7361 7791 7395
rect 8769 7361 8803 7395
rect 10241 7361 10275 7395
rect 10701 7361 10735 7395
rect 13461 7361 13495 7395
rect 14013 7361 14047 7395
rect 15301 7361 15335 7395
rect 16313 7361 16347 7395
rect 16957 7361 16991 7395
rect 17969 7361 18003 7395
rect 18245 7361 18279 7395
rect 20821 7361 20855 7395
rect 25513 7361 25547 7395
rect 30113 7361 30147 7395
rect 30205 7361 30239 7395
rect 37749 7361 37783 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 10517 7293 10551 7327
rect 13737 7293 13771 7327
rect 15393 7293 15427 7327
rect 15485 7293 15519 7327
rect 16681 7293 16715 7327
rect 1869 7225 1903 7259
rect 8585 7225 8619 7259
rect 10885 7225 10919 7259
rect 14749 7225 14783 7259
rect 17693 7225 17727 7259
rect 37933 7225 37967 7259
rect 2145 7157 2179 7191
rect 7849 7157 7883 7191
rect 9505 7157 9539 7191
rect 13645 7157 13679 7191
rect 16497 7157 16531 7191
rect 18153 7157 18187 7191
rect 18429 7157 18463 7191
rect 25697 7157 25731 7191
rect 30389 7157 30423 7191
rect 1869 6885 1903 6919
rect 28273 6885 28307 6919
rect 28549 6885 28583 6919
rect 12449 6817 12483 6851
rect 27905 6817 27939 6851
rect 28043 6817 28077 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 12173 6749 12207 6783
rect 12541 6749 12575 6783
rect 25237 6749 25271 6783
rect 25513 6749 25547 6783
rect 28448 6745 28482 6779
rect 28733 6749 28767 6783
rect 37473 6749 37507 6783
rect 38209 6749 38243 6783
rect 38485 6749 38519 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 38117 6681 38151 6715
rect 1593 6613 1627 6647
rect 2145 6613 2179 6647
rect 8401 6613 8435 6647
rect 11437 6613 11471 6647
rect 12725 6613 12759 6647
rect 26249 6613 26283 6647
rect 27445 6613 27479 6647
rect 27813 6613 27847 6647
rect 37289 6613 37323 6647
rect 38025 6613 38059 6647
rect 38393 6613 38427 6647
rect 38669 6613 38703 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 1593 6409 1627 6443
rect 14749 6409 14783 6443
rect 16957 6409 16991 6443
rect 18981 6409 19015 6443
rect 21833 6409 21867 6443
rect 22109 6409 22143 6443
rect 37657 6409 37691 6443
rect 39405 6409 39439 6443
rect 2605 6341 2639 6375
rect 19809 6341 19843 6375
rect 1409 6273 1443 6307
rect 1685 6273 1719 6307
rect 3157 6273 3191 6307
rect 6009 6273 6043 6307
rect 6561 6273 6595 6307
rect 9535 6273 9569 6307
rect 10114 6272 10148 6306
rect 14565 6273 14599 6307
rect 15117 6273 15151 6307
rect 17141 6273 17175 6307
rect 17969 6273 18003 6307
rect 18245 6273 18279 6307
rect 19073 6273 19107 6307
rect 19717 6273 19751 6307
rect 20453 6273 20487 6307
rect 20612 6273 20646 6307
rect 21465 6273 21499 6307
rect 21649 6273 21683 6307
rect 22017 6273 22051 6307
rect 22293 6273 22327 6307
rect 30481 6273 30515 6307
rect 30665 6273 30699 6307
rect 33885 6273 33919 6307
rect 37473 6273 37507 6307
rect 37841 6273 37875 6307
rect 38485 6273 38519 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 2881 6205 2915 6239
rect 9781 6205 9815 6239
rect 10011 6205 10045 6239
rect 14841 6205 14875 6239
rect 20729 6205 20763 6239
rect 1869 6137 1903 6171
rect 2789 6137 2823 6171
rect 19533 6137 19567 6171
rect 21005 6137 21039 6171
rect 30297 6137 30331 6171
rect 34069 6137 34103 6171
rect 39037 6137 39071 6171
rect 3893 6069 3927 6103
rect 6193 6069 6227 6103
rect 6745 6069 6779 6103
rect 9321 6069 9355 6103
rect 9689 6069 9723 6103
rect 15853 6069 15887 6103
rect 19257 6069 19291 6103
rect 30849 6069 30883 6103
rect 37381 6069 37415 6103
rect 38669 6069 38703 6103
rect 1593 5865 1627 5899
rect 16957 5865 16991 5899
rect 38301 5865 38335 5899
rect 38577 5865 38611 5899
rect 39405 5865 39439 5899
rect 1869 5797 1903 5831
rect 10701 5797 10735 5831
rect 12357 5797 12391 5831
rect 25421 5797 25455 5831
rect 27813 5797 27847 5831
rect 39037 5797 39071 5831
rect 5089 5729 5123 5763
rect 5273 5729 5307 5763
rect 5733 5729 5767 5763
rect 13369 5729 13403 5763
rect 17509 5729 17543 5763
rect 27077 5729 27111 5763
rect 29193 5729 29227 5763
rect 29653 5729 29687 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 3157 5661 3191 5695
rect 6009 5661 6043 5695
rect 6126 5661 6160 5695
rect 6285 5661 6319 5695
rect 6929 5661 6963 5695
rect 10057 5661 10091 5695
rect 10150 5661 10184 5695
rect 10563 5661 10597 5695
rect 10885 5661 10919 5695
rect 11069 5661 11103 5695
rect 11345 5661 11379 5695
rect 11529 5661 11563 5695
rect 13093 5661 13127 5695
rect 20269 5661 20303 5695
rect 23581 5661 23615 5695
rect 23857 5661 23891 5695
rect 24409 5661 24443 5695
rect 24685 5661 24719 5695
rect 25973 5661 26007 5695
rect 26127 5661 26161 5695
rect 26433 5661 26467 5695
rect 26617 5661 26651 5695
rect 26893 5661 26927 5695
rect 27169 5661 27203 5695
rect 27317 5661 27351 5695
rect 27445 5661 27479 5695
rect 27634 5661 27668 5695
rect 28917 5661 28951 5695
rect 29101 5661 29135 5695
rect 29561 5661 29595 5695
rect 38485 5661 38519 5695
rect 38761 5661 38795 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 10333 5593 10367 5627
rect 10425 5593 10459 5627
rect 13553 5593 13587 5627
rect 13737 5593 13771 5627
rect 17417 5593 17451 5627
rect 26341 5593 26375 5627
rect 27537 5593 27571 5627
rect 3341 5525 3375 5559
rect 4997 5525 5031 5559
rect 17325 5525 17359 5559
rect 20085 5525 20119 5559
rect 23765 5525 23799 5559
rect 24041 5525 24075 5559
rect 28733 5525 28767 5559
rect 4445 5321 4479 5355
rect 26341 5321 26375 5355
rect 33425 5321 33459 5355
rect 39405 5321 39439 5355
rect 1409 5185 1443 5219
rect 4261 5185 4295 5219
rect 7906 5185 7940 5219
rect 8493 5185 8527 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 10639 5185 10673 5219
rect 10793 5185 10827 5219
rect 26525 5185 26559 5219
rect 32505 5185 32539 5219
rect 33241 5185 33275 5219
rect 33517 5185 33551 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 32689 5049 32723 5083
rect 1593 4981 1627 5015
rect 7803 4981 7837 5015
rect 8309 4981 8343 5015
rect 10609 4981 10643 5015
rect 33701 4981 33735 5015
rect 39037 4981 39071 5015
rect 10149 4777 10183 4811
rect 16129 4777 16163 4811
rect 19073 4777 19107 4811
rect 20637 4777 20671 4811
rect 20913 4777 20947 4811
rect 23121 4777 23155 4811
rect 23397 4777 23431 4811
rect 24869 4777 24903 4811
rect 29377 4777 29411 4811
rect 29929 4777 29963 4811
rect 33793 4777 33827 4811
rect 34989 4777 35023 4811
rect 35725 4777 35759 4811
rect 37105 4777 37139 4811
rect 38117 4777 38151 4811
rect 39405 4777 39439 4811
rect 13645 4709 13679 4743
rect 17233 4709 17267 4743
rect 22385 4709 22419 4743
rect 26065 4709 26099 4743
rect 28181 4709 28215 4743
rect 5089 4641 5123 4675
rect 5273 4641 5307 4675
rect 5733 4641 5767 4675
rect 6285 4641 6319 4675
rect 6929 4641 6963 4675
rect 7389 4641 7423 4675
rect 7481 4641 7515 4675
rect 9781 4641 9815 4675
rect 10701 4641 10735 4675
rect 14105 4641 14139 4675
rect 18061 4641 18095 4675
rect 21971 4641 22005 4675
rect 22109 4641 22143 4675
rect 22845 4641 22879 4675
rect 25053 4641 25087 4675
rect 28733 4641 28767 4675
rect 6009 4573 6043 4607
rect 6126 4573 6160 4607
rect 7205 4573 7239 4607
rect 8120 4573 8154 4607
rect 8492 4573 8526 4607
rect 8585 4573 8619 4607
rect 9689 4573 9723 4607
rect 12265 4573 12299 4607
rect 13461 4573 13495 4607
rect 14381 4573 14415 4607
rect 15393 4573 15427 4607
rect 15945 4573 15979 4607
rect 16221 4573 16255 4607
rect 16497 4573 16531 4607
rect 17877 4573 17911 4607
rect 18889 4573 18923 4607
rect 19257 4573 19291 4607
rect 19533 4573 19567 4607
rect 20821 4573 20855 4607
rect 21097 4573 21131 4607
rect 21833 4573 21867 4607
rect 23029 4573 23063 4607
rect 23305 4573 23339 4607
rect 23581 4573 23615 4607
rect 24961 4573 24995 4607
rect 25329 4573 25363 4607
rect 27537 4573 27571 4607
rect 27721 4573 27755 4607
rect 28457 4573 28491 4607
rect 28595 4573 28629 4607
rect 29745 4573 29779 4607
rect 30113 4573 30147 4607
rect 33609 4573 33643 4607
rect 34897 4573 34931 4607
rect 35173 4573 35207 4607
rect 35909 4573 35943 4607
rect 36921 4573 36955 4607
rect 38301 4573 38335 4607
rect 38577 4573 38611 4607
rect 39221 4573 39255 4607
rect 3341 4505 3375 4539
rect 3525 4505 3559 4539
rect 8217 4505 8251 4539
rect 8309 4505 8343 4539
rect 9597 4505 9631 4539
rect 10609 4505 10643 4539
rect 17969 4505 18003 4539
rect 38669 4505 38703 4539
rect 38853 4505 38887 4539
rect 7021 4437 7055 4471
rect 7941 4437 7975 4471
rect 9229 4437 9263 4471
rect 10517 4437 10551 4471
rect 12081 4437 12115 4471
rect 15117 4437 15151 4471
rect 15209 4437 15243 4471
rect 17509 4437 17543 4471
rect 20269 4437 20303 4471
rect 21189 4437 21223 4471
rect 29561 4437 29595 4471
rect 34805 4437 34839 4471
rect 38393 4437 38427 4471
rect 6193 4233 6227 4267
rect 8125 4233 8159 4267
rect 14657 4233 14691 4267
rect 27169 4233 27203 4267
rect 3617 4165 3651 4199
rect 37473 4165 37507 4199
rect 5457 4097 5491 4131
rect 8355 4097 8389 4131
rect 8493 4097 8527 4131
rect 10425 4097 10459 4131
rect 10701 4097 10735 4131
rect 14565 4097 14599 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 17877 4097 17911 4131
rect 25237 4097 25271 4131
rect 27353 4097 27387 4131
rect 27905 4097 27939 4131
rect 32479 4097 32513 4131
rect 38485 4097 38519 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 5181 4029 5215 4063
rect 14473 4029 14507 4063
rect 37289 4029 37323 4063
rect 3801 3961 3835 3995
rect 10517 3961 10551 3995
rect 15025 3961 15059 3995
rect 25421 3961 25455 3995
rect 27721 3961 27755 3995
rect 39037 3961 39071 3995
rect 39405 3961 39439 3995
rect 10241 3893 10275 3927
rect 17693 3893 17727 3927
rect 32321 3893 32355 3927
rect 38669 3893 38703 3927
rect 39405 3689 39439 3723
rect 39037 3621 39071 3655
rect 5641 3485 5675 3519
rect 11989 3485 12023 3519
rect 19625 3485 19659 3519
rect 19809 3485 19843 3519
rect 20085 3485 20119 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 5825 3417 5859 3451
rect 12173 3349 12207 3383
rect 20269 3349 20303 3383
rect 16865 3145 16899 3179
rect 18245 3145 18279 3179
rect 19349 3145 19383 3179
rect 24133 3145 24167 3179
rect 24593 3145 24627 3179
rect 25237 3145 25271 3179
rect 26617 3145 26651 3179
rect 27905 3145 27939 3179
rect 29193 3145 29227 3179
rect 29469 3145 29503 3179
rect 29745 3145 29779 3179
rect 30389 3145 30423 3179
rect 32413 3145 32447 3179
rect 34621 3145 34655 3179
rect 36369 3145 36403 3179
rect 38209 3145 38243 3179
rect 39405 3145 39439 3179
rect 22109 3077 22143 3111
rect 22221 3077 22255 3111
rect 23121 3077 23155 3111
rect 16681 3009 16715 3043
rect 16957 3009 16991 3043
rect 17509 3009 17543 3043
rect 19165 3009 19199 3043
rect 19717 3009 19751 3043
rect 21465 3009 21499 3043
rect 21833 3009 21867 3043
rect 21926 3009 21960 3043
rect 22298 3009 22332 3043
rect 22753 3009 22787 3043
rect 22937 3009 22971 3043
rect 23335 3009 23369 3043
rect 23489 3009 23523 3043
rect 23765 3009 23799 3043
rect 24501 3009 24535 3043
rect 25145 3009 25179 3043
rect 25421 3009 25455 3043
rect 26341 3009 26375 3043
rect 26433 3009 26467 3043
rect 28089 3009 28123 3043
rect 29009 3009 29043 3043
rect 29285 3009 29319 3043
rect 29561 3009 29595 3043
rect 30573 3009 30607 3043
rect 32229 3009 32263 3043
rect 34069 3009 34103 3043
rect 34805 3009 34839 3043
rect 36277 3009 36311 3043
rect 36553 3009 36587 3043
rect 38393 3009 38427 3043
rect 38485 3009 38519 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 17233 2941 17267 2975
rect 19441 2941 19475 2975
rect 23029 2941 23063 2975
rect 24593 2941 24627 2975
rect 24685 2941 24719 2975
rect 20453 2873 20487 2907
rect 21557 2873 21591 2907
rect 22477 2873 22511 2907
rect 24961 2873 24995 2907
rect 33885 2873 33919 2907
rect 36185 2873 36219 2907
rect 17141 2805 17175 2839
rect 22569 2805 22603 2839
rect 23581 2805 23615 2839
rect 38669 2805 38703 2839
rect 39037 2805 39071 2839
rect 39405 2601 39439 2635
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3157 2397 3191 2431
rect 4629 2397 4663 2431
rect 6101 2397 6135 2431
rect 7573 2397 7607 2431
rect 9229 2397 9263 2431
rect 11713 2397 11747 2431
rect 37749 2397 37783 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 2973 2261 3007 2295
rect 4445 2261 4479 2295
rect 5917 2261 5951 2295
rect 7389 2261 7423 2295
rect 9045 2261 9079 2295
rect 11897 2261 11931 2295
rect 37933 2261 37967 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
rect 39037 2261 39071 2295
<< metal1 >>
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 25590 11200 25596 11212
rect 1912 11172 25596 11200
rect 1912 11160 1918 11172
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 26418 10140 26424 10192
rect 26476 10180 26482 10192
rect 32582 10180 32588 10192
rect 26476 10152 32588 10180
rect 26476 10140 26482 10152
rect 32582 10140 32588 10152
rect 32640 10140 32646 10192
rect 24486 10004 24492 10056
rect 24544 10044 24550 10056
rect 25130 10044 25136 10056
rect 24544 10016 25136 10044
rect 24544 10004 24550 10016
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 17494 9868 17500 9920
rect 17552 9908 17558 9920
rect 20622 9908 20628 9920
rect 17552 9880 20628 9908
rect 17552 9868 17558 9880
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 2498 9800 2504 9852
rect 2556 9840 2562 9852
rect 24578 9840 24584 9852
rect 2556 9812 24584 9840
rect 2556 9800 2562 9812
rect 24578 9800 24584 9812
rect 24636 9800 24642 9852
rect 10042 9732 10048 9784
rect 10100 9772 10106 9784
rect 37274 9772 37280 9784
rect 10100 9744 37280 9772
rect 10100 9732 10106 9744
rect 37274 9732 37280 9744
rect 37332 9732 37338 9784
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 37642 9704 37648 9716
rect 9548 9676 37648 9704
rect 9548 9664 9554 9676
rect 37642 9664 37648 9676
rect 37700 9664 37706 9716
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 16390 9636 16396 9648
rect 5684 9608 16396 9636
rect 5684 9596 5690 9608
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 23106 9596 23112 9648
rect 23164 9636 23170 9648
rect 23474 9636 23480 9648
rect 23164 9608 23480 9636
rect 23164 9596 23170 9608
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 18046 9528 18052 9580
rect 18104 9568 18110 9580
rect 24486 9568 24492 9580
rect 18104 9540 24492 9568
rect 18104 9528 18110 9540
rect 24486 9528 24492 9540
rect 24544 9528 24550 9580
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 11974 9500 11980 9512
rect 5132 9472 11980 9500
rect 5132 9460 5138 9472
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 4798 9392 4804 9444
rect 4856 9432 4862 9444
rect 15470 9432 15476 9444
rect 4856 9404 15476 9432
rect 4856 9392 4862 9404
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 22646 9392 22652 9444
rect 22704 9432 22710 9444
rect 29178 9432 29184 9444
rect 22704 9404 29184 9432
rect 22704 9392 22710 9404
rect 29178 9392 29184 9404
rect 29236 9392 29242 9444
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4212 9336 12434 9364
rect 4212 9324 4218 9336
rect 6178 9256 6184 9308
rect 6236 9296 6242 9308
rect 10502 9296 10508 9308
rect 6236 9268 10508 9296
rect 6236 9256 6242 9268
rect 10502 9256 10508 9268
rect 10560 9256 10566 9308
rect 12158 9296 12164 9308
rect 10612 9268 12164 9296
rect 6086 9188 6092 9240
rect 6144 9228 6150 9240
rect 10612 9228 10640 9268
rect 12158 9256 12164 9268
rect 12216 9256 12222 9308
rect 12406 9296 12434 9336
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 21174 9364 21180 9376
rect 13688 9336 21180 9364
rect 13688 9324 13694 9336
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 38838 9364 38844 9376
rect 31726 9336 38844 9364
rect 13814 9296 13820 9308
rect 12406 9268 13820 9296
rect 13814 9256 13820 9268
rect 13872 9256 13878 9308
rect 17034 9256 17040 9308
rect 17092 9296 17098 9308
rect 17678 9296 17684 9308
rect 17092 9268 17684 9296
rect 17092 9256 17098 9268
rect 17678 9256 17684 9268
rect 17736 9256 17742 9308
rect 24394 9256 24400 9308
rect 24452 9296 24458 9308
rect 31726 9296 31754 9336
rect 38838 9324 38844 9336
rect 38896 9324 38902 9376
rect 24452 9268 31754 9296
rect 24452 9256 24458 9268
rect 6144 9200 10640 9228
rect 6144 9188 6150 9200
rect 13262 9188 13268 9240
rect 13320 9228 13326 9240
rect 17770 9228 17776 9240
rect 13320 9200 17776 9228
rect 13320 9188 13326 9200
rect 17770 9188 17776 9200
rect 17828 9188 17834 9240
rect 19306 9200 21404 9228
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 8570 9160 8576 9172
rect 4764 9132 8576 9160
rect 4764 9120 4770 9132
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 13354 9120 13360 9172
rect 13412 9160 13418 9172
rect 19306 9160 19334 9200
rect 13412 9132 19334 9160
rect 21376 9160 21404 9200
rect 28994 9188 29000 9240
rect 29052 9228 29058 9240
rect 29052 9200 31754 9228
rect 29052 9188 29058 9200
rect 28258 9160 28264 9172
rect 21376 9132 28264 9160
rect 13412 9120 13418 9132
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 29822 9120 29828 9172
rect 29880 9160 29886 9172
rect 31726 9160 31754 9200
rect 38746 9160 38752 9172
rect 29880 9132 30604 9160
rect 31726 9132 38752 9160
rect 29880 9120 29886 9132
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 10594 9092 10600 9104
rect 3660 9064 10600 9092
rect 3660 9052 3666 9064
rect 10594 9052 10600 9064
rect 10652 9052 10658 9104
rect 30374 9092 30380 9104
rect 17052 9064 30380 9092
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 17052 9024 17080 9064
rect 30374 9052 30380 9064
rect 30432 9052 30438 9104
rect 30576 9092 30604 9132
rect 38746 9120 38752 9132
rect 38804 9120 38810 9172
rect 35434 9092 35440 9104
rect 30576 9064 35440 9092
rect 35434 9052 35440 9064
rect 35492 9052 35498 9104
rect 37550 9024 37556 9036
rect 12216 8996 17080 9024
rect 19306 8996 37556 9024
rect 12216 8984 12222 8996
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 7282 8956 7288 8968
rect 4580 8928 7288 8956
rect 4580 8916 4586 8928
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 13630 8956 13636 8968
rect 7576 8928 13636 8956
rect 7576 8832 7604 8928
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 19306 8956 19334 8996
rect 37550 8984 37556 8996
rect 37608 8984 37614 9036
rect 13964 8928 19334 8956
rect 13964 8916 13970 8928
rect 24946 8916 24952 8968
rect 25004 8956 25010 8968
rect 25958 8956 25964 8968
rect 25004 8928 25964 8956
rect 25004 8916 25010 8928
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 34238 8916 34244 8968
rect 34296 8956 34302 8968
rect 37826 8956 37832 8968
rect 34296 8928 37832 8956
rect 34296 8916 34302 8928
rect 37826 8916 37832 8928
rect 37884 8916 37890 8968
rect 10226 8848 10232 8900
rect 10284 8888 10290 8900
rect 14642 8888 14648 8900
rect 10284 8860 14648 8888
rect 10284 8848 10290 8860
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 16114 8848 16120 8900
rect 16172 8888 16178 8900
rect 20714 8888 20720 8900
rect 16172 8860 20720 8888
rect 16172 8848 16178 8860
rect 20714 8848 20720 8860
rect 20772 8848 20778 8900
rect 27706 8848 27712 8900
rect 27764 8888 27770 8900
rect 32674 8888 32680 8900
rect 27764 8860 32680 8888
rect 27764 8848 27770 8860
rect 32674 8848 32680 8860
rect 32732 8848 32738 8900
rect 33778 8848 33784 8900
rect 33836 8888 33842 8900
rect 35618 8888 35624 8900
rect 33836 8860 35624 8888
rect 33836 8848 33842 8860
rect 35618 8848 35624 8860
rect 35676 8848 35682 8900
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 6730 8820 6736 8832
rect 2924 8792 6736 8820
rect 2924 8780 2930 8792
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7558 8780 7564 8832
rect 7616 8780 7622 8832
rect 8294 8780 8300 8832
rect 8352 8820 8358 8832
rect 11146 8820 11152 8832
rect 8352 8792 11152 8820
rect 8352 8780 8358 8792
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 15746 8780 15752 8832
rect 15804 8820 15810 8832
rect 19426 8820 19432 8832
rect 15804 8792 19432 8820
rect 15804 8780 15810 8792
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 24026 8820 24032 8832
rect 22152 8792 24032 8820
rect 22152 8780 22158 8792
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 24302 8780 24308 8832
rect 24360 8820 24366 8832
rect 26786 8820 26792 8832
rect 24360 8792 26792 8820
rect 24360 8780 24366 8792
rect 26786 8780 26792 8792
rect 26844 8780 26850 8832
rect 34054 8780 34060 8832
rect 34112 8820 34118 8832
rect 36170 8820 36176 8832
rect 34112 8792 36176 8820
rect 34112 8780 34118 8792
rect 36170 8780 36176 8792
rect 36228 8780 36234 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 2498 8576 2504 8628
rect 2556 8576 2562 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 2866 8616 2872 8628
rect 2823 8588 2872 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3786 8616 3792 8628
rect 3467 8588 3792 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4338 8616 4344 8628
rect 4203 8588 4344 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4890 8616 4896 8628
rect 4571 8588 4896 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5902 8616 5908 8628
rect 5675 8588 5908 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6270 8616 6276 8628
rect 6043 8588 6276 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6822 8616 6828 8628
rect 6779 8588 6828 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7374 8616 7380 8628
rect 7147 8588 7380 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 7558 8576 7564 8628
rect 7616 8576 7622 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8110 8616 8116 8628
rect 7883 8588 8116 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8478 8616 8484 8628
rect 8251 8588 8484 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8616 8631 8619
rect 8846 8616 8852 8628
rect 8619 8588 8852 8616
rect 8619 8585 8631 8588
rect 8573 8579 8631 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9582 8616 9588 8628
rect 9355 8588 9588 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10410 8616 10416 8628
rect 10091 8588 10416 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 10686 8616 10692 8628
rect 10551 8588 10692 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10873 8619 10931 8625
rect 10873 8585 10885 8619
rect 10919 8616 10931 8619
rect 10962 8616 10968 8628
rect 10919 8588 10968 8616
rect 10919 8585 10931 8588
rect 10873 8579 10931 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 11514 8616 11520 8628
rect 11195 8588 11520 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11977 8619 12035 8625
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12066 8616 12072 8628
rect 12023 8588 12072 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 12894 8616 12900 8628
rect 12667 8588 12900 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13170 8616 13176 8628
rect 13035 8588 13176 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13630 8616 13636 8628
rect 13403 8588 13636 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13998 8616 14004 8628
rect 13771 8588 14004 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14550 8616 14556 8628
rect 14507 8588 14556 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 15289 8619 15347 8625
rect 15068 8588 15240 8616
rect 15068 8576 15074 8588
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 7576 8548 7604 8576
rect 8294 8548 8300 8560
rect 1360 8520 2636 8548
rect 1360 8508 1366 8520
rect 1210 8440 1216 8492
rect 1268 8480 1274 8492
rect 2608 8489 2636 8520
rect 6196 8520 7604 8548
rect 7944 8520 8300 8548
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1268 8452 2329 8480
rect 1268 8440 1274 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 382 8372 388 8424
rect 440 8412 446 8424
rect 1397 8415 1455 8421
rect 1397 8412 1409 8415
rect 440 8384 1409 8412
rect 440 8372 446 8384
rect 1397 8381 1409 8384
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 3252 8412 3280 8443
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4522 8480 4528 8492
rect 4387 8452 4528 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5626 8480 5632 8492
rect 5491 8452 5632 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 6196 8489 6224 8520
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 6181 8443 6239 8449
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8480 7343 8483
rect 7558 8480 7564 8492
rect 7331 8452 7564 8480
rect 7331 8449 7343 8452
rect 7285 8443 7343 8449
rect 4798 8412 4804 8424
rect 3252 8384 4804 8412
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 5368 8412 5396 8440
rect 4908 8384 5396 8412
rect 566 8304 572 8356
rect 624 8344 630 8356
rect 1486 8344 1492 8356
rect 624 8316 1492 8344
rect 624 8304 630 8316
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3510 8344 3516 8356
rect 3099 8316 3516 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 4908 8353 4936 8384
rect 4893 8347 4951 8353
rect 4893 8313 4905 8347
rect 4939 8313 4951 8347
rect 4893 8307 4951 8313
rect 5261 8347 5319 8353
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 5718 8344 5724 8356
rect 5307 8316 5724 8344
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 5718 8304 5724 8316
rect 5776 8304 5782 8356
rect 6932 8344 6960 8443
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7944 8480 7972 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 13262 8548 13268 8560
rect 8404 8520 13268 8548
rect 7699 8452 7972 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8404 8489 8432 8520
rect 13262 8508 13268 8520
rect 13320 8508 13326 8560
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 15212 8548 15240 8588
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15654 8616 15660 8628
rect 15611 8588 15660 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 16206 8616 16212 8628
rect 15979 8588 16212 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16482 8616 16488 8628
rect 16439 8588 16488 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16816 8588 16957 8616
rect 16816 8576 16822 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 19610 8616 19616 8628
rect 16945 8579 17003 8585
rect 17512 8588 19616 8616
rect 17512 8548 17540 8588
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 22005 8619 22063 8625
rect 22005 8585 22017 8619
rect 22051 8616 22063 8619
rect 22462 8616 22468 8628
rect 22051 8588 22468 8616
rect 22051 8585 22063 8588
rect 22005 8579 22063 8585
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 22554 8576 22560 8628
rect 22612 8616 22618 8628
rect 23109 8619 23167 8625
rect 22612 8588 22784 8616
rect 22612 8576 22618 8588
rect 13872 8520 15148 8548
rect 15212 8520 16252 8548
rect 13872 8508 13878 8520
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 8846 8480 8852 8492
rect 8803 8452 8852 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 10042 8480 10048 8492
rect 9907 8452 10048 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10560 8452 10701 8480
rect 10560 8440 10566 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12710 8480 12716 8492
rect 12483 8452 12716 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 11054 8412 11060 8424
rect 8036 8384 11060 8412
rect 7469 8347 7527 8353
rect 6932 8316 7420 8344
rect 7392 8276 7420 8316
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7926 8344 7932 8356
rect 7515 8316 7932 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8036 8276 8064 8384
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 9677 8347 9735 8353
rect 8352 8316 9628 8344
rect 8352 8304 8358 8316
rect 7392 8248 8064 8276
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9030 8276 9036 8288
rect 8812 8248 9036 8276
rect 8812 8236 8818 8248
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 9600 8276 9628 8316
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 10134 8344 10140 8356
rect 9723 8316 10140 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 11808 8344 11836 8443
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13354 8480 13360 8492
rect 13219 8452 13360 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 14458 8440 14464 8492
rect 14516 8480 14522 8492
rect 15120 8489 15148 8520
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14516 8452 14657 8480
rect 14516 8440 14522 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15028 8412 15056 8443
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 16114 8440 16120 8492
rect 16172 8440 16178 8492
rect 16224 8489 16252 8520
rect 17144 8520 17540 8548
rect 17144 8489 17172 8520
rect 17770 8508 17776 8560
rect 17828 8548 17834 8560
rect 21634 8548 21640 8560
rect 17828 8520 21640 8548
rect 17828 8508 17834 8520
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21784 8520 22140 8548
rect 21784 8508 21790 8520
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17681 8483 17739 8489
rect 17368 8452 17540 8480
rect 17368 8440 17374 8452
rect 16022 8412 16028 8424
rect 15028 8384 16028 8412
rect 16022 8372 16028 8384
rect 16080 8372 16086 8424
rect 10566 8316 11836 8344
rect 10566 8276 10594 8316
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 13630 8344 13636 8356
rect 12768 8316 13636 8344
rect 12768 8304 12774 8316
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 17512 8353 17540 8452
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 17954 8480 17960 8492
rect 17727 8452 17960 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18046 8440 18052 8492
rect 18104 8440 18110 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18414 8480 18420 8492
rect 18371 8452 18420 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18785 8483 18843 8489
rect 18785 8480 18797 8483
rect 18748 8452 18797 8480
rect 18748 8440 18754 8452
rect 18785 8449 18797 8452
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18966 8480 18972 8492
rect 18923 8452 18972 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19242 8440 19248 8492
rect 19300 8480 19306 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19300 8452 19349 8480
rect 19300 8440 19306 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 19576 8452 19625 8480
rect 19576 8440 19582 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19852 8452 20085 8480
rect 19852 8440 19858 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21358 8480 21364 8492
rect 21315 8452 21364 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 21450 8440 21456 8492
rect 21508 8480 21514 8492
rect 22112 8489 22140 8520
rect 22278 8508 22284 8560
rect 22336 8548 22342 8560
rect 22336 8520 22692 8548
rect 22336 8508 22342 8520
rect 22664 8489 22692 8520
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21508 8452 21833 8480
rect 21508 8440 21514 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22557 8483 22615 8489
rect 22557 8449 22569 8483
rect 22603 8449 22615 8483
rect 22557 8443 22615 8449
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22756 8480 22784 8588
rect 23109 8585 23121 8619
rect 23155 8616 23167 8619
rect 23155 8588 23336 8616
rect 23155 8585 23167 8588
rect 23109 8579 23167 8585
rect 22830 8508 22836 8560
rect 22888 8548 22894 8560
rect 22888 8520 23244 8548
rect 22888 8508 22894 8520
rect 23216 8489 23244 8520
rect 22925 8483 22983 8489
rect 22925 8480 22937 8483
rect 22756 8452 22937 8480
rect 22649 8443 22707 8449
rect 22925 8449 22937 8452
rect 22971 8449 22983 8483
rect 22925 8443 22983 8449
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 20622 8412 20628 8424
rect 17828 8384 20628 8412
rect 17828 8372 17834 8384
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 20772 8384 21404 8412
rect 20772 8372 20778 8384
rect 21376 8356 21404 8384
rect 22002 8372 22008 8424
rect 22060 8412 22066 8424
rect 22572 8412 22600 8443
rect 22060 8384 22600 8412
rect 23308 8412 23336 8588
rect 23658 8576 23664 8628
rect 23716 8616 23722 8628
rect 23716 8588 24072 8616
rect 23716 8576 23722 8588
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 23440 8520 23980 8548
rect 23440 8508 23446 8520
rect 23474 8440 23480 8492
rect 23532 8480 23538 8492
rect 23952 8489 23980 8520
rect 24044 8489 24072 8588
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 24912 8588 25268 8616
rect 24912 8576 24918 8588
rect 24210 8508 24216 8560
rect 24268 8548 24274 8560
rect 24268 8520 24900 8548
rect 24268 8508 24274 8520
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23532 8452 23673 8480
rect 23532 8440 23538 8452
rect 23661 8449 23673 8452
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 24118 8440 24124 8492
rect 24176 8480 24182 8492
rect 24872 8489 24900 8520
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24176 8452 24593 8480
rect 24176 8440 24182 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 25130 8440 25136 8492
rect 25188 8440 25194 8492
rect 25240 8489 25268 8588
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 25464 8588 25513 8616
rect 25464 8576 25470 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 25501 8579 25559 8585
rect 25590 8576 25596 8628
rect 25648 8616 25654 8628
rect 25777 8619 25835 8625
rect 25777 8616 25789 8619
rect 25648 8588 25789 8616
rect 25648 8576 25654 8588
rect 25777 8585 25789 8588
rect 25823 8585 25835 8619
rect 25777 8579 25835 8585
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 27893 8619 27951 8625
rect 27893 8616 27905 8619
rect 26016 8588 27905 8616
rect 26016 8576 26022 8588
rect 27893 8585 27905 8588
rect 27939 8585 27951 8619
rect 27893 8579 27951 8585
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 28721 8619 28779 8625
rect 28721 8616 28733 8619
rect 28592 8588 28733 8616
rect 28592 8576 28598 8588
rect 28721 8585 28733 8588
rect 28767 8585 28779 8619
rect 28721 8579 28779 8585
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 28960 8588 29224 8616
rect 28960 8576 28966 8588
rect 25314 8508 25320 8560
rect 25372 8548 25378 8560
rect 25372 8520 26004 8548
rect 25372 8508 25378 8520
rect 25976 8489 26004 8520
rect 26418 8508 26424 8560
rect 26476 8548 26482 8560
rect 26476 8520 28304 8548
rect 26476 8508 26482 8520
rect 25225 8483 25283 8489
rect 25225 8449 25237 8483
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 23308 8384 24992 8412
rect 22060 8372 22066 8384
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8313 17555 8347
rect 17497 8307 17555 8313
rect 17678 8304 17684 8356
rect 17736 8344 17742 8356
rect 17865 8347 17923 8353
rect 17865 8344 17877 8347
rect 17736 8316 17877 8344
rect 17736 8304 17742 8316
rect 17865 8313 17877 8316
rect 17911 8313 17923 8347
rect 17865 8307 17923 8313
rect 17954 8304 17960 8356
rect 18012 8344 18018 8356
rect 19334 8344 19340 8356
rect 18012 8316 19340 8344
rect 18012 8304 18018 8316
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 19797 8347 19855 8353
rect 19797 8313 19809 8347
rect 19843 8344 19855 8347
rect 20990 8344 20996 8356
rect 19843 8316 20996 8344
rect 19843 8313 19855 8316
rect 19797 8307 19855 8313
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 21358 8304 21364 8356
rect 21416 8304 21422 8356
rect 21453 8347 21511 8353
rect 21453 8313 21465 8347
rect 21499 8344 21511 8347
rect 22094 8344 22100 8356
rect 21499 8316 22100 8344
rect 21499 8313 21511 8316
rect 21453 8307 21511 8313
rect 22094 8304 22100 8316
rect 22152 8304 22158 8356
rect 22833 8347 22891 8353
rect 22204 8316 22508 8344
rect 9600 8248 10594 8276
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 14550 8276 14556 8288
rect 11388 8248 14556 8276
rect 11388 8236 11394 8248
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 14642 8236 14648 8288
rect 14700 8276 14706 8288
rect 18414 8276 18420 8288
rect 14700 8248 18420 8276
rect 14700 8236 14706 8248
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 18506 8236 18512 8288
rect 18564 8236 18570 8288
rect 18598 8236 18604 8288
rect 18656 8236 18662 8288
rect 19061 8279 19119 8285
rect 19061 8245 19073 8279
rect 19107 8276 19119 8279
rect 19150 8276 19156 8288
rect 19107 8248 19156 8276
rect 19107 8245 19119 8248
rect 19061 8239 19119 8245
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 19518 8236 19524 8288
rect 19576 8236 19582 8288
rect 19889 8279 19947 8285
rect 19889 8245 19901 8279
rect 19935 8276 19947 8279
rect 20530 8276 20536 8288
rect 19935 8248 20536 8276
rect 19935 8245 19947 8248
rect 19889 8239 19947 8245
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 20898 8236 20904 8288
rect 20956 8276 20962 8288
rect 22204 8276 22232 8316
rect 22480 8288 22508 8316
rect 22833 8313 22845 8347
rect 22879 8344 22891 8347
rect 23290 8344 23296 8356
rect 22879 8316 23296 8344
rect 22879 8313 22891 8316
rect 22833 8307 22891 8313
rect 23290 8304 23296 8316
rect 23348 8304 23354 8356
rect 23566 8304 23572 8356
rect 23624 8344 23630 8356
rect 23753 8347 23811 8353
rect 23753 8344 23765 8347
rect 23624 8316 23765 8344
rect 23624 8304 23630 8316
rect 23753 8313 23765 8316
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 23934 8304 23940 8356
rect 23992 8344 23998 8356
rect 24397 8347 24455 8353
rect 24397 8344 24409 8347
rect 23992 8316 24409 8344
rect 23992 8304 23998 8316
rect 24397 8313 24409 8316
rect 24443 8313 24455 8347
rect 24397 8307 24455 8313
rect 24670 8304 24676 8356
rect 24728 8304 24734 8356
rect 24964 8344 24992 8384
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25700 8412 25728 8443
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 28077 8483 28135 8489
rect 28077 8480 28089 8483
rect 27856 8452 28089 8480
rect 27856 8440 27862 8452
rect 28077 8449 28089 8452
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 28166 8440 28172 8492
rect 28224 8440 28230 8492
rect 25096 8384 25728 8412
rect 25096 8372 25102 8384
rect 25866 8372 25872 8424
rect 25924 8412 25930 8424
rect 26510 8412 26516 8424
rect 25924 8384 26516 8412
rect 25924 8372 25930 8384
rect 26510 8372 26516 8384
rect 26568 8372 26574 8424
rect 28276 8412 28304 8520
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 28629 8483 28687 8489
rect 28629 8480 28641 8483
rect 28408 8452 28641 8480
rect 28408 8440 28414 8452
rect 28629 8449 28641 8452
rect 28675 8449 28687 8483
rect 28629 8443 28687 8449
rect 28905 8483 28963 8489
rect 28905 8449 28917 8483
rect 28951 8480 28963 8483
rect 29086 8480 29092 8492
rect 28951 8452 29092 8480
rect 28951 8449 28963 8452
rect 28905 8443 28963 8449
rect 29086 8440 29092 8452
rect 29144 8440 29150 8492
rect 29196 8489 29224 8588
rect 30374 8576 30380 8628
rect 30432 8616 30438 8628
rect 30561 8619 30619 8625
rect 30561 8616 30573 8619
rect 30432 8588 30573 8616
rect 30432 8576 30438 8588
rect 30561 8585 30573 8588
rect 30607 8585 30619 8619
rect 30561 8579 30619 8585
rect 32214 8576 32220 8628
rect 32272 8616 32278 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 32272 8588 32321 8616
rect 32272 8576 32278 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32548 8588 32781 8616
rect 32548 8576 32554 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33413 8619 33471 8625
rect 33413 8616 33425 8619
rect 32916 8588 33425 8616
rect 32916 8576 32922 8588
rect 33413 8585 33425 8588
rect 33459 8585 33471 8619
rect 33413 8579 33471 8585
rect 33502 8576 33508 8628
rect 33560 8616 33566 8628
rect 33873 8619 33931 8625
rect 33873 8616 33885 8619
rect 33560 8588 33885 8616
rect 33560 8576 33566 8588
rect 33873 8585 33885 8588
rect 33919 8585 33931 8619
rect 33873 8579 33931 8585
rect 33962 8576 33968 8628
rect 34020 8616 34026 8628
rect 34793 8619 34851 8625
rect 34793 8616 34805 8619
rect 34020 8588 34805 8616
rect 34020 8576 34026 8588
rect 34793 8585 34805 8588
rect 34839 8585 34851 8619
rect 34793 8579 34851 8585
rect 35161 8619 35219 8625
rect 35161 8585 35173 8619
rect 35207 8585 35219 8619
rect 35161 8579 35219 8585
rect 29730 8508 29736 8560
rect 29788 8548 29794 8560
rect 30653 8551 30711 8557
rect 30653 8548 30665 8551
rect 29788 8520 30665 8548
rect 29788 8508 29794 8520
rect 30653 8517 30665 8520
rect 30699 8517 30711 8551
rect 30653 8511 30711 8517
rect 34146 8508 34152 8560
rect 34204 8548 34210 8560
rect 35176 8548 35204 8579
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36725 8619 36783 8625
rect 36725 8616 36737 8619
rect 35860 8588 36737 8616
rect 35860 8576 35866 8588
rect 36725 8585 36737 8588
rect 36771 8585 36783 8619
rect 36725 8579 36783 8585
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 37829 8619 37887 8625
rect 37829 8616 37841 8619
rect 36964 8588 37841 8616
rect 36964 8576 36970 8588
rect 37829 8585 37841 8588
rect 37875 8585 37887 8619
rect 37829 8579 37887 8585
rect 38565 8619 38623 8625
rect 38565 8585 38577 8619
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 34204 8520 35204 8548
rect 34204 8508 34210 8520
rect 35250 8508 35256 8560
rect 35308 8548 35314 8560
rect 35308 8520 36124 8548
rect 35308 8508 35314 8520
rect 29181 8483 29239 8489
rect 29181 8449 29193 8483
rect 29227 8449 29239 8483
rect 29181 8443 29239 8449
rect 32490 8440 32496 8492
rect 32548 8440 32554 8492
rect 32585 8483 32643 8489
rect 32585 8449 32597 8483
rect 32631 8449 32643 8483
rect 32585 8443 32643 8449
rect 28276 8384 28488 8412
rect 27430 8344 27436 8356
rect 24964 8316 27436 8344
rect 27430 8304 27436 8316
rect 27488 8304 27494 8356
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 28353 8347 28411 8353
rect 28353 8344 28365 8347
rect 27672 8316 28365 8344
rect 27672 8304 27678 8316
rect 28353 8313 28365 8316
rect 28399 8313 28411 8347
rect 28460 8344 28488 8384
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 29549 8415 29607 8421
rect 29549 8412 29561 8415
rect 28776 8384 29561 8412
rect 28776 8372 28782 8384
rect 29549 8381 29561 8384
rect 29595 8381 29607 8415
rect 29549 8375 29607 8381
rect 29825 8415 29883 8421
rect 29825 8381 29837 8415
rect 29871 8381 29883 8415
rect 29825 8375 29883 8381
rect 29840 8344 29868 8375
rect 32398 8372 32404 8424
rect 32456 8412 32462 8424
rect 32600 8412 32628 8443
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 32953 8483 33011 8489
rect 32953 8480 32965 8483
rect 32732 8452 32965 8480
rect 32732 8440 32738 8452
rect 32953 8449 32965 8452
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 33597 8483 33655 8489
rect 33597 8449 33609 8483
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 32456 8384 32628 8412
rect 33612 8412 33640 8443
rect 33686 8440 33692 8492
rect 33744 8440 33750 8492
rect 34333 8483 34391 8489
rect 34333 8449 34345 8483
rect 34379 8449 34391 8483
rect 34333 8443 34391 8449
rect 34238 8412 34244 8424
rect 33612 8384 34244 8412
rect 32456 8372 32462 8384
rect 34238 8372 34244 8384
rect 34296 8372 34302 8424
rect 34348 8412 34376 8443
rect 34974 8440 34980 8492
rect 35032 8440 35038 8492
rect 35342 8440 35348 8492
rect 35400 8440 35406 8492
rect 35434 8440 35440 8492
rect 35492 8440 35498 8492
rect 35618 8440 35624 8492
rect 35676 8480 35682 8492
rect 35805 8483 35863 8489
rect 35805 8480 35817 8483
rect 35676 8452 35817 8480
rect 35676 8440 35682 8452
rect 35805 8449 35817 8452
rect 35851 8449 35863 8483
rect 35805 8443 35863 8449
rect 34348 8384 34652 8412
rect 28460 8316 29868 8344
rect 28353 8307 28411 8313
rect 32766 8304 32772 8356
rect 32824 8344 32830 8356
rect 33137 8347 33195 8353
rect 33137 8344 33149 8347
rect 32824 8316 33149 8344
rect 32824 8304 32830 8316
rect 33137 8313 33149 8316
rect 33183 8313 33195 8347
rect 33137 8307 33195 8313
rect 33594 8304 33600 8356
rect 33652 8344 33658 8356
rect 34149 8347 34207 8353
rect 34149 8344 34161 8347
rect 33652 8316 34161 8344
rect 33652 8304 33658 8316
rect 34149 8313 34161 8316
rect 34195 8313 34207 8347
rect 34149 8307 34207 8313
rect 20956 8248 22232 8276
rect 20956 8236 20962 8248
rect 22278 8236 22284 8288
rect 22336 8236 22342 8288
rect 22370 8236 22376 8288
rect 22428 8236 22434 8288
rect 22462 8236 22468 8288
rect 22520 8236 22526 8288
rect 23382 8236 23388 8288
rect 23440 8236 23446 8288
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23658 8276 23664 8288
rect 23523 8248 23664 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 24210 8236 24216 8288
rect 24268 8236 24274 8288
rect 24946 8236 24952 8288
rect 25004 8236 25010 8288
rect 25409 8279 25467 8285
rect 25409 8245 25421 8279
rect 25455 8276 25467 8279
rect 26326 8276 26332 8288
rect 25455 8248 26332 8276
rect 25455 8245 25467 8248
rect 25409 8239 25467 8245
rect 26326 8236 26332 8248
rect 26384 8236 26390 8288
rect 26602 8236 26608 8288
rect 26660 8276 26666 8288
rect 28445 8279 28503 8285
rect 28445 8276 28457 8279
rect 26660 8248 28457 8276
rect 26660 8236 26666 8248
rect 28445 8245 28457 8248
rect 28491 8245 28503 8279
rect 28445 8239 28503 8245
rect 28997 8279 29055 8285
rect 28997 8245 29009 8279
rect 29043 8276 29055 8279
rect 29178 8276 29184 8288
rect 29043 8248 29184 8276
rect 29043 8245 29055 8248
rect 28997 8239 29055 8245
rect 29178 8236 29184 8248
rect 29236 8236 29242 8288
rect 30190 8236 30196 8288
rect 30248 8276 30254 8288
rect 31938 8276 31944 8288
rect 30248 8248 31944 8276
rect 30248 8236 30254 8248
rect 31938 8236 31944 8248
rect 31996 8236 32002 8288
rect 34624 8276 34652 8384
rect 35066 8372 35072 8424
rect 35124 8412 35130 8424
rect 35124 8384 36032 8412
rect 35124 8372 35130 8384
rect 34698 8304 34704 8356
rect 34756 8344 34762 8356
rect 36004 8353 36032 8384
rect 35621 8347 35679 8353
rect 35621 8344 35633 8347
rect 34756 8316 35633 8344
rect 34756 8304 34762 8316
rect 35621 8313 35633 8316
rect 35667 8313 35679 8347
rect 35621 8307 35679 8313
rect 35989 8347 36047 8353
rect 35989 8313 36001 8347
rect 36035 8313 36047 8347
rect 36096 8344 36124 8520
rect 36814 8508 36820 8560
rect 36872 8548 36878 8560
rect 36872 8520 37412 8548
rect 36872 8508 36878 8520
rect 36170 8440 36176 8492
rect 36228 8440 36234 8492
rect 36538 8440 36544 8492
rect 36596 8440 36602 8492
rect 37090 8440 37096 8492
rect 37148 8480 37154 8492
rect 37277 8483 37335 8489
rect 37277 8480 37289 8483
rect 37148 8452 37289 8480
rect 37148 8440 37154 8452
rect 37277 8449 37289 8452
rect 37323 8449 37335 8483
rect 37384 8480 37412 8520
rect 37458 8508 37464 8560
rect 37516 8548 37522 8560
rect 38580 8548 38608 8579
rect 37516 8520 38608 8548
rect 37516 8508 37522 8520
rect 38746 8508 38752 8560
rect 38804 8548 38810 8560
rect 38804 8520 39252 8548
rect 38804 8508 38810 8520
rect 37645 8483 37703 8489
rect 37645 8480 37657 8483
rect 37384 8452 37657 8480
rect 37277 8443 37335 8449
rect 37645 8449 37657 8452
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 38013 8483 38071 8489
rect 38013 8449 38025 8483
rect 38059 8449 38071 8483
rect 38013 8443 38071 8449
rect 38381 8483 38439 8489
rect 38381 8449 38393 8483
rect 38427 8480 38439 8483
rect 38470 8480 38476 8492
rect 38427 8452 38476 8480
rect 38427 8449 38439 8452
rect 38381 8443 38439 8449
rect 36354 8372 36360 8424
rect 36412 8412 36418 8424
rect 36412 8384 37136 8412
rect 36412 8372 36418 8384
rect 36096 8316 36400 8344
rect 35989 8307 36047 8313
rect 35894 8276 35900 8288
rect 34624 8248 35900 8276
rect 35894 8236 35900 8248
rect 35952 8236 35958 8288
rect 36372 8285 36400 8316
rect 36357 8279 36415 8285
rect 36357 8245 36369 8279
rect 36403 8245 36415 8279
rect 37108 8276 37136 8384
rect 37458 8372 37464 8424
rect 37516 8412 37522 8424
rect 38028 8412 38056 8443
rect 38470 8440 38476 8452
rect 38528 8440 38534 8492
rect 38838 8440 38844 8492
rect 38896 8440 38902 8492
rect 39224 8489 39252 8520
rect 39209 8483 39267 8489
rect 39209 8449 39221 8483
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 37516 8384 38056 8412
rect 37516 8372 37522 8384
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 37240 8316 38209 8344
rect 37240 8304 37246 8316
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 39022 8304 39028 8356
rect 39080 8304 39086 8356
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37108 8248 37473 8276
rect 36357 8239 36415 8245
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 3326 8072 3332 8084
rect 2179 8044 3332 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4120 8044 4261 8072
rect 4120 8032 4126 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4672 8044 4813 8072
rect 4672 8032 4678 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 5224 8044 5365 8072
rect 5224 8032 5230 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6604 8044 6745 8072
rect 6604 8032 6610 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7285 8075 7343 8081
rect 7285 8072 7297 8075
rect 7156 8044 7297 8072
rect 7156 8032 7162 8044
rect 7285 8041 7297 8044
rect 7331 8041 7343 8075
rect 7285 8035 7343 8041
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7708 8044 7849 8072
rect 7708 8032 7714 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 8389 8075 8447 8081
rect 8389 8041 8401 8075
rect 8435 8072 8447 8075
rect 8754 8072 8760 8084
rect 8435 8044 8760 8072
rect 8435 8041 8447 8044
rect 8389 8035 8447 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9030 8032 9036 8084
rect 9088 8032 9094 8084
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 9456 8044 9505 8072
rect 9456 8032 9462 8044
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 9916 8044 10057 8072
rect 9916 8032 9922 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 10045 8035 10103 8041
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11296 8044 11437 8072
rect 11296 8032 11302 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11848 8044 11989 8072
rect 11848 8032 11854 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12676 8044 12817 8072
rect 12676 8032 12682 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 12805 8035 12863 8041
rect 13648 8044 14105 8072
rect 1026 7964 1032 8016
rect 1084 8004 1090 8016
rect 8573 8007 8631 8013
rect 1084 7976 2544 8004
rect 1084 7964 1090 7976
rect 1118 7896 1124 7948
rect 1176 7936 1182 7948
rect 1176 7908 2268 7936
rect 1176 7896 1182 7908
rect 750 7828 756 7880
rect 808 7868 814 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 808 7840 1409 7868
rect 808 7828 814 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 842 7760 848 7812
rect 900 7800 906 7812
rect 1688 7800 1716 7831
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2240 7877 2268 7908
rect 2516 7877 2544 7976
rect 8573 7973 8585 8007
rect 8619 7973 8631 8007
rect 8573 7967 8631 7973
rect 8588 7936 8616 7967
rect 9122 7964 9128 8016
rect 9180 8004 9186 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9180 7976 10333 8004
rect 9180 7964 9186 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 10778 7964 10784 8016
rect 10836 7964 10842 8016
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 13648 8004 13676 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14461 8075 14519 8081
rect 14461 8072 14473 8075
rect 14332 8044 14473 8072
rect 14332 8032 14338 8044
rect 14461 8041 14473 8044
rect 14507 8041 14519 8075
rect 14461 8035 14519 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14884 8044 15025 8072
rect 14884 8032 14890 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15289 8075 15347 8081
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 15470 8072 15476 8084
rect 15335 8044 15476 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 15988 8044 16129 8072
rect 15988 8032 15994 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 17586 8072 17592 8084
rect 17543 8044 17592 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 20622 8072 20628 8084
rect 19576 8044 20628 8072
rect 19576 8032 19582 8044
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 23017 8075 23075 8081
rect 23017 8072 23029 8075
rect 20772 8044 23029 8072
rect 20772 8032 20778 8044
rect 23017 8041 23029 8044
rect 23063 8041 23075 8075
rect 23017 8035 23075 8041
rect 24394 8032 24400 8084
rect 24452 8032 24458 8084
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 26568 8044 31754 8072
rect 26568 8032 26574 8044
rect 12952 7976 13676 8004
rect 12952 7964 12958 7976
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 16298 8004 16304 8016
rect 13780 7976 16304 8004
rect 13780 7964 13786 7976
rect 16298 7964 16304 7976
rect 16356 7964 16362 8016
rect 19794 7964 19800 8016
rect 19852 8004 19858 8016
rect 21545 8007 21603 8013
rect 21545 8004 21557 8007
rect 19852 7976 21557 8004
rect 19852 7964 19858 7976
rect 21545 7973 21557 7976
rect 21591 7973 21603 8007
rect 21545 7967 21603 7973
rect 22186 7964 22192 8016
rect 22244 7964 22250 8016
rect 22462 7964 22468 8016
rect 22520 8004 22526 8016
rect 22520 7976 25728 8004
rect 22520 7964 22526 7976
rect 5552 7908 8616 7936
rect 8864 7908 10732 7936
rect 1949 7871 2007 7877
rect 1949 7868 1961 7871
rect 1912 7840 1961 7868
rect 1912 7828 1918 7840
rect 1949 7837 1961 7840
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 4430 7828 4436 7880
rect 4488 7828 4494 7880
rect 5552 7877 5580 7908
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 5828 7840 6868 7868
rect 2866 7800 2872 7812
rect 900 7772 1716 7800
rect 1872 7772 2872 7800
rect 900 7760 906 7772
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 1872 7741 1900 7772
rect 2866 7760 2872 7772
rect 2924 7760 2930 7812
rect 5000 7800 5028 7831
rect 5828 7800 5856 7840
rect 5000 7772 5856 7800
rect 5902 7760 5908 7812
rect 5960 7760 5966 7812
rect 6270 7760 6276 7812
rect 6328 7760 6334 7812
rect 6454 7760 6460 7812
rect 6512 7760 6518 7812
rect 6840 7800 6868 7840
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 8018 7828 8024 7880
rect 8076 7828 8082 7880
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7868 8355 7871
rect 8478 7868 8484 7880
rect 8343 7840 8484 7868
rect 8343 7837 8355 7840
rect 8297 7831 8355 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 8757 7871 8815 7877
rect 8757 7868 8769 7871
rect 8720 7840 8769 7868
rect 8720 7828 8726 7840
rect 8757 7837 8769 7840
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 8864 7800 8892 7908
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9398 7868 9404 7880
rect 9263 7840 9404 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9674 7828 9680 7880
rect 9732 7828 9738 7880
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 6840 7772 8892 7800
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 10318 7800 10324 7812
rect 8996 7772 10324 7800
rect 8996 7760 9002 7772
rect 10318 7760 10324 7772
rect 10376 7760 10382 7812
rect 10413 7803 10471 7809
rect 10413 7769 10425 7803
rect 10459 7800 10471 7803
rect 10597 7803 10655 7809
rect 10597 7800 10609 7803
rect 10459 7772 10609 7800
rect 10459 7769 10471 7772
rect 10413 7763 10471 7769
rect 10597 7769 10609 7772
rect 10643 7769 10655 7803
rect 10597 7763 10655 7769
rect 1857 7735 1915 7741
rect 1857 7701 1869 7735
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 2961 7735 3019 7741
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 5810 7732 5816 7744
rect 3007 7704 5816 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 5997 7735 6055 7741
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 6362 7732 6368 7744
rect 6043 7704 6368 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 10042 7732 10048 7744
rect 8076 7704 10048 7732
rect 8076 7692 8082 7704
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10704 7732 10732 7908
rect 10870 7896 10876 7948
rect 10928 7936 10934 7948
rect 19889 7939 19947 7945
rect 10928 7908 17632 7936
rect 10928 7896 10934 7908
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11624 7800 11652 7831
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 13817 7871 13875 7877
rect 13035 7840 13768 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 12618 7800 12624 7812
rect 11624 7772 12624 7800
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 13446 7760 13452 7812
rect 13504 7800 13510 7812
rect 13504 7772 13676 7800
rect 13504 7760 13510 7772
rect 12894 7732 12900 7744
rect 10704 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13648 7741 13676 7772
rect 13633 7735 13691 7741
rect 13633 7701 13645 7735
rect 13679 7701 13691 7735
rect 13740 7732 13768 7840
rect 13817 7837 13829 7871
rect 13863 7868 13875 7871
rect 14182 7868 14188 7880
rect 13863 7840 14188 7868
rect 13863 7837 13875 7840
rect 13817 7831 13875 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14292 7800 14320 7831
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 15197 7871 15255 7877
rect 15197 7837 15209 7871
rect 15243 7868 15255 7871
rect 15378 7868 15384 7880
rect 15243 7840 15384 7868
rect 15243 7837 15255 7840
rect 15197 7831 15255 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 16301 7871 16359 7877
rect 16301 7837 16313 7871
rect 16347 7868 16359 7871
rect 16390 7868 16396 7880
rect 16347 7840 16396 7868
rect 16347 7837 16359 7840
rect 16301 7831 16359 7837
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 17604 7877 17632 7908
rect 19889 7905 19901 7939
rect 19935 7936 19947 7939
rect 19935 7908 20760 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 17494 7800 17500 7812
rect 14292 7772 17500 7800
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 17604 7800 17632 7831
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 17865 7871 17923 7877
rect 17865 7868 17877 7871
rect 17736 7840 17877 7868
rect 17736 7828 17742 7840
rect 17865 7837 17877 7840
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18141 7831 18199 7837
rect 18340 7840 19257 7868
rect 18156 7800 18184 7831
rect 18340 7812 18368 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 19518 7868 19524 7880
rect 19475 7840 19524 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 19518 7828 19524 7840
rect 19576 7828 19582 7880
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 20438 7868 20444 7880
rect 20180 7840 20444 7868
rect 17604 7772 18184 7800
rect 18322 7760 18328 7812
rect 18380 7760 18386 7812
rect 20180 7800 20208 7840
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20534 7871 20592 7877
rect 20534 7837 20546 7871
rect 20580 7837 20592 7871
rect 20732 7868 20760 7908
rect 20990 7896 20996 7948
rect 21048 7936 21054 7948
rect 23569 7939 23627 7945
rect 23569 7936 23581 7939
rect 21048 7908 22140 7936
rect 21048 7896 21054 7908
rect 20906 7871 20964 7877
rect 20906 7868 20918 7871
rect 20732 7840 20918 7868
rect 20534 7831 20592 7837
rect 20906 7837 20918 7840
rect 20952 7837 20964 7871
rect 20906 7831 20964 7837
rect 18892 7772 20208 7800
rect 15562 7732 15568 7744
rect 13740 7704 15568 7732
rect 13633 7695 13691 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 17678 7732 17684 7744
rect 16724 7704 17684 7732
rect 16724 7692 16730 7704
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17770 7692 17776 7744
rect 17828 7692 17834 7744
rect 18892 7741 18920 7772
rect 18877 7735 18935 7741
rect 18877 7701 18889 7735
rect 18923 7701 18935 7735
rect 18877 7695 18935 7701
rect 19702 7692 19708 7744
rect 19760 7732 19766 7744
rect 20548 7732 20576 7831
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21140 7840 21373 7868
rect 21140 7828 21146 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21634 7828 21640 7880
rect 21692 7828 21698 7880
rect 22112 7877 22140 7908
rect 22480 7908 23581 7936
rect 21973 7871 22031 7877
rect 21973 7837 21985 7871
rect 22019 7868 22031 7871
rect 22097 7871 22155 7877
rect 22019 7837 22047 7868
rect 21973 7831 22047 7837
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22143 7840 22385 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 20714 7760 20720 7812
rect 20772 7760 20778 7812
rect 20809 7803 20867 7809
rect 20809 7769 20821 7803
rect 20855 7800 20867 7803
rect 21729 7803 21787 7809
rect 21729 7800 21741 7803
rect 20855 7772 21741 7800
rect 20855 7769 20867 7772
rect 20809 7763 20867 7769
rect 21729 7769 21741 7772
rect 21775 7769 21787 7803
rect 21729 7763 21787 7769
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 22019 7800 22047 7831
rect 22480 7800 22508 7908
rect 23569 7905 23581 7908
rect 23615 7905 23627 7939
rect 23569 7899 23627 7905
rect 23676 7908 24624 7936
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 23440 7840 23489 7868
rect 23440 7828 23446 7840
rect 23477 7837 23489 7840
rect 23523 7868 23535 7871
rect 23676 7868 23704 7908
rect 24596 7877 24624 7908
rect 25700 7877 25728 7976
rect 25774 7964 25780 8016
rect 25832 8004 25838 8016
rect 29549 8007 29607 8013
rect 29549 8004 29561 8007
rect 25832 7976 29561 8004
rect 25832 7964 25838 7976
rect 29549 7973 29561 7976
rect 29595 7973 29607 8007
rect 29549 7967 29607 7973
rect 30190 7936 30196 7948
rect 27080 7908 28672 7936
rect 27080 7877 27108 7908
rect 24029 7871 24087 7877
rect 24029 7868 24041 7871
rect 23523 7840 23704 7868
rect 23768 7840 24041 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 21876 7772 22508 7800
rect 21876 7760 21882 7772
rect 19760 7704 20576 7732
rect 19760 7692 19766 7704
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 21177 7735 21235 7741
rect 21177 7701 21189 7735
rect 21223 7732 21235 7735
rect 21450 7732 21456 7744
rect 21223 7704 21456 7732
rect 21223 7701 21235 7704
rect 21177 7695 21235 7701
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 23385 7735 23443 7741
rect 23385 7732 23397 7735
rect 22336 7704 23397 7732
rect 22336 7692 22342 7704
rect 23385 7701 23397 7704
rect 23431 7732 23443 7735
rect 23768 7732 23796 7840
rect 24029 7837 24041 7840
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 25685 7871 25743 7877
rect 25685 7837 25697 7871
rect 25731 7837 25743 7871
rect 25685 7831 25743 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 28258 7760 28264 7812
rect 28316 7800 28322 7812
rect 28644 7800 28672 7908
rect 28828 7908 30196 7936
rect 28721 7871 28779 7877
rect 28721 7837 28733 7871
rect 28767 7868 28779 7871
rect 28828 7868 28856 7908
rect 30190 7896 30196 7908
rect 30248 7896 30254 7948
rect 28767 7840 28856 7868
rect 28997 7871 29055 7877
rect 28767 7837 28779 7840
rect 28721 7831 28779 7837
rect 28997 7837 29009 7871
rect 29043 7868 29055 7871
rect 29089 7871 29147 7877
rect 29089 7868 29101 7871
rect 29043 7840 29101 7868
rect 29043 7837 29055 7840
rect 28997 7831 29055 7837
rect 29089 7837 29101 7840
rect 29135 7837 29147 7871
rect 29089 7831 29147 7837
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29512 7840 29745 7868
rect 29512 7828 29518 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 31726 7868 31754 8044
rect 34422 8032 34428 8084
rect 34480 8072 34486 8084
rect 34793 8075 34851 8081
rect 34793 8072 34805 8075
rect 34480 8044 34805 8072
rect 34480 8032 34486 8044
rect 34793 8041 34805 8044
rect 34839 8041 34851 8075
rect 34793 8035 34851 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35713 8075 35771 8081
rect 35713 8072 35725 8075
rect 35584 8044 35725 8072
rect 35584 8032 35590 8044
rect 35713 8041 35725 8044
rect 35759 8041 35771 8075
rect 35713 8035 35771 8041
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36265 8075 36323 8081
rect 36265 8072 36277 8075
rect 36136 8044 36277 8072
rect 36136 8032 36142 8044
rect 36265 8041 36277 8044
rect 36311 8041 36323 8075
rect 36265 8035 36323 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36909 8075 36967 8081
rect 36909 8072 36921 8075
rect 36688 8044 36921 8072
rect 36688 8032 36694 8044
rect 36909 8041 36921 8044
rect 36955 8041 36967 8075
rect 36909 8035 36967 8041
rect 37734 8032 37740 8084
rect 37792 8072 37798 8084
rect 38657 8075 38715 8081
rect 38657 8072 38669 8075
rect 37792 8044 38669 8072
rect 37792 8032 37798 8044
rect 38657 8041 38669 8044
rect 38703 8041 38715 8075
rect 38657 8035 38715 8041
rect 33045 8007 33103 8013
rect 33045 7973 33057 8007
rect 33091 8004 33103 8007
rect 36998 8004 37004 8016
rect 33091 7976 37004 8004
rect 33091 7973 33103 7976
rect 33045 7967 33103 7973
rect 36998 7964 37004 7976
rect 37056 7964 37062 8016
rect 38381 8007 38439 8013
rect 38381 7973 38393 8007
rect 38427 8004 38439 8007
rect 39758 8004 39764 8016
rect 38427 7976 39764 8004
rect 38427 7973 38439 7976
rect 38381 7967 38439 7973
rect 39758 7964 39764 7976
rect 39816 7964 39822 8016
rect 32582 7896 32588 7948
rect 32640 7936 32646 7948
rect 32640 7908 35296 7936
rect 32640 7896 32646 7908
rect 32125 7871 32183 7877
rect 32125 7868 32137 7871
rect 31726 7840 32137 7868
rect 29733 7831 29791 7837
rect 32125 7837 32137 7840
rect 32171 7837 32183 7871
rect 32125 7831 32183 7837
rect 32769 7871 32827 7877
rect 32769 7837 32781 7871
rect 32815 7868 32827 7871
rect 32861 7871 32919 7877
rect 32861 7868 32873 7871
rect 32815 7840 32873 7868
rect 32815 7837 32827 7840
rect 32769 7831 32827 7837
rect 32861 7837 32873 7840
rect 32907 7837 32919 7871
rect 32861 7831 32919 7837
rect 33137 7871 33195 7877
rect 33137 7837 33149 7871
rect 33183 7868 33195 7871
rect 33413 7871 33471 7877
rect 33413 7868 33425 7871
rect 33183 7840 33425 7868
rect 33183 7837 33195 7840
rect 33137 7831 33195 7837
rect 33413 7837 33425 7840
rect 33459 7837 33471 7871
rect 33413 7831 33471 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7868 35035 7871
rect 35158 7868 35164 7880
rect 35023 7840 35164 7868
rect 35023 7837 35035 7840
rect 34977 7831 35035 7837
rect 35158 7828 35164 7840
rect 35216 7828 35222 7880
rect 35268 7877 35296 7908
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7837 35311 7871
rect 35253 7831 35311 7837
rect 35897 7871 35955 7877
rect 35897 7837 35909 7871
rect 35943 7837 35955 7871
rect 35897 7831 35955 7837
rect 28810 7800 28816 7812
rect 28316 7772 28580 7800
rect 28644 7772 28816 7800
rect 28316 7760 28322 7772
rect 23431 7704 23796 7732
rect 23431 7701 23443 7704
rect 23385 7695 23443 7701
rect 23842 7692 23848 7744
rect 23900 7692 23906 7744
rect 25498 7692 25504 7744
rect 25556 7692 25562 7744
rect 27249 7735 27307 7741
rect 27249 7701 27261 7735
rect 27295 7732 27307 7735
rect 28442 7732 28448 7744
rect 27295 7704 28448 7732
rect 27295 7701 27307 7704
rect 27249 7695 27307 7701
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 28552 7741 28580 7772
rect 28810 7760 28816 7772
rect 28868 7760 28874 7812
rect 29178 7760 29184 7812
rect 29236 7800 29242 7812
rect 35912 7800 35940 7831
rect 36446 7828 36452 7880
rect 36504 7828 36510 7880
rect 36722 7828 36728 7880
rect 36780 7828 36786 7880
rect 38105 7871 38163 7877
rect 38105 7837 38117 7871
rect 38151 7868 38163 7871
rect 38197 7871 38255 7877
rect 38197 7868 38209 7871
rect 38151 7840 38209 7868
rect 38151 7837 38163 7840
rect 38105 7831 38163 7837
rect 38197 7837 38209 7840
rect 38243 7837 38255 7871
rect 38197 7831 38255 7837
rect 38286 7828 38292 7880
rect 38344 7868 38350 7880
rect 38473 7871 38531 7877
rect 38473 7868 38485 7871
rect 38344 7840 38485 7868
rect 38344 7828 38350 7840
rect 38473 7837 38485 7840
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7868 39267 7871
rect 39255 7840 39289 7868
rect 39255 7837 39267 7840
rect 39209 7831 39267 7837
rect 37642 7800 37648 7812
rect 29236 7772 35848 7800
rect 35912 7772 37648 7800
rect 29236 7760 29242 7772
rect 28537 7735 28595 7741
rect 28537 7701 28549 7735
rect 28583 7701 28595 7735
rect 28537 7695 28595 7701
rect 28997 7735 29055 7741
rect 28997 7701 29009 7735
rect 29043 7732 29055 7735
rect 29086 7732 29092 7744
rect 29043 7704 29092 7732
rect 29043 7701 29055 7704
rect 28997 7695 29055 7701
rect 29086 7692 29092 7704
rect 29144 7692 29150 7744
rect 29273 7735 29331 7741
rect 29273 7701 29285 7735
rect 29319 7732 29331 7735
rect 30466 7732 30472 7744
rect 29319 7704 30472 7732
rect 29319 7701 29331 7704
rect 29273 7695 29331 7701
rect 30466 7692 30472 7704
rect 30524 7692 30530 7744
rect 31938 7692 31944 7744
rect 31996 7692 32002 7744
rect 32766 7692 32772 7744
rect 32824 7692 32830 7744
rect 33321 7735 33379 7741
rect 33321 7701 33333 7735
rect 33367 7732 33379 7735
rect 33410 7732 33416 7744
rect 33367 7704 33416 7732
rect 33367 7701 33379 7704
rect 33321 7695 33379 7701
rect 33410 7692 33416 7704
rect 33468 7692 33474 7744
rect 33502 7692 33508 7744
rect 33560 7692 33566 7744
rect 35066 7692 35072 7744
rect 35124 7692 35130 7744
rect 35820 7732 35848 7772
rect 37642 7760 37648 7772
rect 37700 7760 37706 7812
rect 39117 7803 39175 7809
rect 39117 7769 39129 7803
rect 39163 7800 39175 7803
rect 39224 7800 39252 7831
rect 40126 7800 40132 7812
rect 39163 7772 40132 7800
rect 39163 7769 39175 7772
rect 39117 7763 39175 7769
rect 40126 7760 40132 7772
rect 40184 7760 40190 7812
rect 38013 7735 38071 7741
rect 38013 7732 38025 7735
rect 35820 7704 38025 7732
rect 38013 7701 38025 7704
rect 38059 7701 38071 7735
rect 38013 7695 38071 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 5534 7528 5540 7540
rect 1627 7500 5540 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 14921 7531 14979 7537
rect 7892 7500 14780 7528
rect 7892 7488 7898 7500
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 992 7432 1716 7460
rect 992 7420 998 7432
rect 750 7352 756 7404
rect 808 7392 814 7404
rect 1688 7401 1716 7432
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 10870 7460 10876 7472
rect 2464 7432 10876 7460
rect 2464 7420 2470 7432
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 14752 7460 14780 7500
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15470 7528 15476 7540
rect 14967 7500 15476 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 20901 7531 20959 7537
rect 20901 7497 20913 7531
rect 20947 7528 20959 7531
rect 21634 7528 21640 7540
rect 20947 7500 21640 7528
rect 20947 7497 20959 7500
rect 20901 7491 20959 7497
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 25682 7488 25688 7540
rect 25740 7528 25746 7540
rect 29178 7528 29184 7540
rect 25740 7500 29184 7528
rect 25740 7488 25746 7500
rect 29178 7488 29184 7500
rect 29236 7488 29242 7540
rect 29270 7488 29276 7540
rect 29328 7528 29334 7540
rect 38289 7531 38347 7537
rect 29328 7500 31754 7528
rect 29328 7488 29334 7500
rect 12216 7432 14688 7460
rect 14752 7432 15424 7460
rect 12216 7420 12222 7432
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 808 7364 1409 7392
rect 808 7352 814 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 658 7284 664 7336
rect 716 7324 722 7336
rect 1964 7324 1992 7355
rect 7742 7352 7748 7404
rect 7800 7352 7806 7404
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8444 7364 8769 7392
rect 8444 7352 8450 7364
rect 8757 7361 8769 7364
rect 8803 7361 8815 7395
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 8757 7355 8815 7361
rect 8864 7364 10241 7392
rect 716 7296 1992 7324
rect 716 7284 722 7296
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 2924 7296 4108 7324
rect 2924 7284 2930 7296
rect 1857 7259 1915 7265
rect 1857 7225 1869 7259
rect 1903 7256 1915 7259
rect 3878 7256 3884 7268
rect 1903 7228 3884 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 3878 7216 3884 7228
rect 3936 7216 3942 7268
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 3970 7188 3976 7200
rect 2179 7160 3976 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4080 7188 4108 7296
rect 5810 7284 5816 7336
rect 5868 7324 5874 7336
rect 8864 7324 8892 7364
rect 10229 7361 10241 7364
rect 10275 7392 10287 7395
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 10275 7364 10701 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13504 7364 14013 7392
rect 13504 7352 13510 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 5868 7296 8892 7324
rect 10505 7327 10563 7333
rect 5868 7284 5874 7296
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 10551 7296 12434 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 12406 7268 12434 7296
rect 13722 7284 13728 7336
rect 13780 7284 13786 7336
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 6972 7228 8524 7256
rect 6972 7216 6978 7228
rect 7282 7188 7288 7200
rect 4080 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 7834 7148 7840 7200
rect 7892 7148 7898 7200
rect 8496 7188 8524 7228
rect 8570 7216 8576 7268
rect 8628 7216 8634 7268
rect 9766 7256 9772 7268
rect 9324 7228 9772 7256
rect 9324 7188 9352 7228
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 10870 7216 10876 7268
rect 10928 7216 10934 7268
rect 12406 7228 12440 7268
rect 12434 7216 12440 7228
rect 12492 7216 12498 7268
rect 8496 7160 9352 7188
rect 9493 7191 9551 7197
rect 9493 7157 9505 7191
rect 9539 7188 9551 7191
rect 10134 7188 10140 7200
rect 9539 7160 10140 7188
rect 9539 7157 9551 7160
rect 9493 7151 9551 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 13630 7148 13636 7200
rect 13688 7148 13694 7200
rect 14660 7188 14688 7432
rect 15286 7352 15292 7404
rect 15344 7352 15350 7404
rect 15396 7392 15424 7432
rect 16132 7432 22094 7460
rect 16132 7392 16160 7432
rect 15396 7364 16160 7392
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16356 7364 16957 7392
rect 16356 7352 16362 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17920 7364 17969 7392
rect 17920 7352 17926 7364
rect 17957 7361 17969 7364
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 18138 7352 18144 7404
rect 18196 7392 18202 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 18196 7364 18245 7392
rect 18196 7352 18202 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 20438 7352 20444 7404
rect 20496 7392 20502 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20496 7364 20821 7392
rect 20496 7352 20502 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 22066 7392 22094 7432
rect 24762 7420 24768 7472
rect 24820 7460 24826 7472
rect 29086 7460 29092 7472
rect 24820 7432 29092 7460
rect 24820 7420 24826 7432
rect 29086 7420 29092 7432
rect 29144 7420 29150 7472
rect 29914 7420 29920 7472
rect 29972 7460 29978 7472
rect 30009 7463 30067 7469
rect 30009 7460 30021 7463
rect 29972 7432 30021 7460
rect 29972 7420 29978 7432
rect 30009 7429 30021 7432
rect 30055 7429 30067 7463
rect 30009 7423 30067 7429
rect 25498 7392 25504 7404
rect 22066 7364 25504 7392
rect 20809 7355 20867 7361
rect 25498 7352 25504 7364
rect 25556 7352 25562 7404
rect 25682 7352 25688 7404
rect 25740 7392 25746 7404
rect 25866 7392 25872 7404
rect 25740 7364 25872 7392
rect 25740 7352 25746 7364
rect 25866 7352 25872 7364
rect 25924 7352 25930 7404
rect 30101 7395 30159 7401
rect 30101 7361 30113 7395
rect 30147 7392 30159 7395
rect 30193 7395 30251 7401
rect 30193 7392 30205 7395
rect 30147 7364 30205 7392
rect 30147 7361 30159 7364
rect 30101 7355 30159 7361
rect 30193 7361 30205 7364
rect 30239 7361 30251 7395
rect 31726 7392 31754 7500
rect 38289 7497 38301 7531
rect 38335 7528 38347 7531
rect 38378 7528 38384 7540
rect 38335 7500 38384 7528
rect 38335 7497 38347 7500
rect 38289 7491 38347 7497
rect 38378 7488 38384 7500
rect 38436 7488 38442 7540
rect 38654 7488 38660 7540
rect 38712 7488 38718 7540
rect 38930 7488 38936 7540
rect 38988 7528 38994 7540
rect 39025 7531 39083 7537
rect 39025 7528 39037 7531
rect 38988 7500 39037 7528
rect 38988 7488 38994 7500
rect 39025 7497 39037 7500
rect 39071 7497 39083 7531
rect 39025 7491 39083 7497
rect 39393 7531 39451 7537
rect 39393 7497 39405 7531
rect 39439 7528 39451 7531
rect 39574 7528 39580 7540
rect 39439 7500 39580 7528
rect 39439 7497 39451 7500
rect 39393 7491 39451 7497
rect 39574 7488 39580 7500
rect 39632 7488 39638 7540
rect 37366 7420 37372 7472
rect 37424 7460 37430 7472
rect 37424 7432 39252 7460
rect 37424 7420 37430 7432
rect 37737 7395 37795 7401
rect 37737 7392 37749 7395
rect 31726 7364 37749 7392
rect 30193 7355 30251 7361
rect 37737 7361 37749 7364
rect 37783 7361 37795 7395
rect 37737 7355 37795 7361
rect 38102 7352 38108 7404
rect 38160 7352 38166 7404
rect 38473 7395 38531 7401
rect 38473 7361 38485 7395
rect 38519 7392 38531 7395
rect 38562 7392 38568 7404
rect 38519 7364 38568 7392
rect 38519 7361 38531 7364
rect 38473 7355 38531 7361
rect 38562 7352 38568 7364
rect 38620 7352 38626 7404
rect 38838 7352 38844 7404
rect 38896 7352 38902 7404
rect 39224 7401 39252 7432
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 15378 7284 15384 7336
rect 15436 7284 15442 7336
rect 15473 7327 15531 7333
rect 15473 7293 15485 7327
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 14737 7259 14795 7265
rect 14737 7225 14749 7259
rect 14783 7256 14795 7259
rect 15488 7256 15516 7287
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 23106 7324 23112 7336
rect 17328 7296 23112 7324
rect 14783 7228 15516 7256
rect 15580 7228 16620 7256
rect 14783 7225 14795 7228
rect 14737 7219 14795 7225
rect 15580 7188 15608 7228
rect 14660 7160 15608 7188
rect 16482 7148 16488 7200
rect 16540 7148 16546 7200
rect 16592 7188 16620 7228
rect 17328 7188 17356 7296
rect 23106 7284 23112 7296
rect 23164 7284 23170 7336
rect 23198 7284 23204 7336
rect 23256 7324 23262 7336
rect 26510 7324 26516 7336
rect 23256 7296 26516 7324
rect 23256 7284 23262 7296
rect 26510 7284 26516 7296
rect 26568 7284 26574 7336
rect 27430 7284 27436 7336
rect 27488 7324 27494 7336
rect 28166 7324 28172 7336
rect 27488 7296 28172 7324
rect 27488 7284 27494 7296
rect 28166 7284 28172 7296
rect 28224 7284 28230 7336
rect 28442 7284 28448 7336
rect 28500 7324 28506 7336
rect 38286 7324 38292 7336
rect 28500 7296 38292 7324
rect 28500 7284 28506 7296
rect 38286 7284 38292 7296
rect 38344 7284 38350 7336
rect 17681 7259 17739 7265
rect 17681 7225 17693 7259
rect 17727 7256 17739 7259
rect 19518 7256 19524 7268
rect 17727 7228 19524 7256
rect 17727 7225 17739 7228
rect 17681 7219 17739 7225
rect 19518 7216 19524 7228
rect 19576 7256 19582 7268
rect 20898 7256 20904 7268
rect 19576 7228 20904 7256
rect 19576 7216 19582 7228
rect 20898 7216 20904 7228
rect 20956 7256 20962 7268
rect 21818 7256 21824 7268
rect 20956 7228 21824 7256
rect 20956 7216 20962 7228
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 31938 7256 31944 7268
rect 25608 7228 31944 7256
rect 16592 7160 17356 7188
rect 18138 7148 18144 7200
rect 18196 7148 18202 7200
rect 18414 7148 18420 7200
rect 18472 7148 18478 7200
rect 18506 7148 18512 7200
rect 18564 7188 18570 7200
rect 25608 7188 25636 7228
rect 31938 7216 31944 7228
rect 31996 7216 32002 7268
rect 37921 7259 37979 7265
rect 37921 7225 37933 7259
rect 37967 7256 37979 7259
rect 39298 7256 39304 7268
rect 37967 7228 39304 7256
rect 37967 7225 37979 7228
rect 37921 7219 37979 7225
rect 39298 7216 39304 7228
rect 39356 7216 39362 7268
rect 18564 7160 25636 7188
rect 25685 7191 25743 7197
rect 18564 7148 18570 7160
rect 25685 7157 25697 7191
rect 25731 7188 25743 7191
rect 28350 7188 28356 7200
rect 25731 7160 28356 7188
rect 25731 7157 25743 7160
rect 25685 7151 25743 7157
rect 28350 7148 28356 7160
rect 28408 7148 28414 7200
rect 28442 7148 28448 7200
rect 28500 7188 28506 7200
rect 28718 7188 28724 7200
rect 28500 7160 28724 7188
rect 28500 7148 28506 7160
rect 28718 7148 28724 7160
rect 28776 7148 28782 7200
rect 30374 7148 30380 7200
rect 30432 7148 30438 7200
rect 33410 7148 33416 7200
rect 33468 7188 33474 7200
rect 39850 7188 39856 7200
rect 33468 7160 39856 7188
rect 33468 7148 33474 7160
rect 39850 7148 39856 7160
rect 39908 7148 39914 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 1118 6944 1124 6996
rect 1176 6984 1182 6996
rect 1176 6956 1992 6984
rect 1176 6944 1182 6956
rect 1857 6919 1915 6925
rect 1857 6885 1869 6919
rect 1903 6885 1915 6919
rect 1964 6916 1992 6956
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 2740 6956 8248 6984
rect 2740 6944 2746 6956
rect 5902 6916 5908 6928
rect 1964 6888 5908 6916
rect 1857 6879 1915 6885
rect 1026 6808 1032 6860
rect 1084 6848 1090 6860
rect 1872 6848 1900 6879
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 1084 6820 1808 6848
rect 1872 6820 6132 6848
rect 1084 6808 1090 6820
rect 750 6740 756 6792
rect 808 6780 814 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 808 6752 1409 6780
rect 808 6740 814 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1780 6780 1808 6820
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1780 6752 1961 6780
rect 1673 6743 1731 6749
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 5350 6780 5356 6792
rect 1949 6743 2007 6749
rect 2056 6752 5356 6780
rect 842 6672 848 6724
rect 900 6712 906 6724
rect 1688 6712 1716 6743
rect 900 6684 1716 6712
rect 900 6672 906 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2056 6644 2084 6752
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 6104 6712 6132 6820
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 6880 6752 7389 6780
rect 6880 6740 6886 6752
rect 7377 6749 7389 6752
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7742 6780 7748 6792
rect 7699 6752 7748 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 7668 6712 7696 6743
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8220 6780 8248 6956
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 9732 6956 10181 6984
rect 9732 6944 9738 6956
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9950 6916 9956 6928
rect 9824 6888 9956 6916
rect 9824 6876 9830 6888
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 10153 6916 10181 6956
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10284 6956 12434 6984
rect 10284 6944 10290 6956
rect 11422 6916 11428 6928
rect 10153 6888 11428 6916
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 11514 6876 11520 6928
rect 11572 6916 11578 6928
rect 12406 6916 12434 6956
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 38838 6984 38844 6996
rect 16540 6956 38844 6984
rect 16540 6944 16546 6956
rect 38838 6944 38844 6956
rect 38896 6944 38902 6996
rect 11572 6888 11836 6916
rect 12406 6888 24808 6916
rect 11572 6876 11578 6888
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 11698 6848 11704 6860
rect 8536 6820 11704 6848
rect 8536 6808 8542 6820
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11514 6780 11520 6792
rect 8220 6752 11520 6780
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 11808 6780 11836 6888
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13722 6848 13728 6860
rect 12492 6820 13728 6848
rect 12492 6808 12498 6820
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 22094 6848 22100 6860
rect 13872 6820 22100 6848
rect 13872 6808 13878 6820
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 12161 6783 12219 6789
rect 12161 6780 12173 6783
rect 11808 6752 12173 6780
rect 12161 6749 12173 6752
rect 12207 6780 12219 6783
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12207 6752 12541 6780
rect 12207 6749 12219 6752
rect 12161 6743 12219 6749
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 21818 6780 21824 6792
rect 12676 6752 21824 6780
rect 12676 6740 12682 6752
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 23842 6740 23848 6792
rect 23900 6780 23906 6792
rect 24302 6780 24308 6792
rect 23900 6752 24308 6780
rect 23900 6740 23906 6752
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 11606 6712 11612 6724
rect 6104 6684 7696 6712
rect 7760 6684 11612 6712
rect 1627 6616 2084 6644
rect 2133 6647 2191 6653
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2590 6644 2596 6656
rect 2179 6616 2596 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2590 6604 2596 6616
rect 2648 6604 2654 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 7760 6644 7788 6684
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 24670 6712 24676 6724
rect 11756 6684 24676 6712
rect 11756 6672 11762 6684
rect 24670 6672 24676 6684
rect 24728 6672 24734 6724
rect 24780 6712 24808 6888
rect 25958 6876 25964 6928
rect 26016 6916 26022 6928
rect 28261 6919 28319 6925
rect 28261 6916 28273 6919
rect 26016 6888 28273 6916
rect 26016 6876 26022 6888
rect 28261 6885 28273 6888
rect 28307 6885 28319 6919
rect 28261 6879 28319 6885
rect 28442 6876 28448 6928
rect 28500 6916 28506 6928
rect 28537 6919 28595 6925
rect 28537 6916 28549 6919
rect 28500 6888 28549 6916
rect 28500 6876 28506 6888
rect 28537 6885 28549 6888
rect 28583 6885 28595 6919
rect 28537 6879 28595 6885
rect 28626 6876 28632 6928
rect 28684 6916 28690 6928
rect 35066 6916 35072 6928
rect 28684 6888 35072 6916
rect 28684 6876 28690 6888
rect 35066 6876 35072 6888
rect 35124 6876 35130 6928
rect 27430 6808 27436 6860
rect 27488 6848 27494 6860
rect 27893 6851 27951 6857
rect 27893 6848 27905 6851
rect 27488 6820 27905 6848
rect 27488 6808 27494 6820
rect 27893 6817 27905 6820
rect 27939 6817 27951 6851
rect 27893 6811 27951 6817
rect 27982 6808 27988 6860
rect 28040 6857 28046 6860
rect 28040 6851 28089 6857
rect 28040 6817 28043 6851
rect 28077 6817 28089 6851
rect 28040 6811 28089 6817
rect 28040 6808 28046 6811
rect 28902 6808 28908 6860
rect 28960 6848 28966 6860
rect 28960 6820 39252 6848
rect 28960 6808 28966 6820
rect 25222 6740 25228 6792
rect 25280 6740 25286 6792
rect 25498 6740 25504 6792
rect 25556 6740 25562 6792
rect 27798 6780 27804 6792
rect 25608 6752 27804 6780
rect 25608 6712 25636 6752
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 28166 6740 28172 6792
rect 28224 6780 28230 6792
rect 28224 6776 28396 6780
rect 28436 6779 28494 6785
rect 28436 6776 28448 6779
rect 28224 6752 28448 6776
rect 28224 6740 28230 6752
rect 28368 6748 28448 6752
rect 28436 6745 28448 6748
rect 28482 6745 28494 6779
rect 28436 6739 28494 6745
rect 28718 6740 28724 6792
rect 28776 6740 28782 6792
rect 30834 6740 30840 6792
rect 30892 6780 30898 6792
rect 37461 6783 37519 6789
rect 37461 6780 37473 6783
rect 30892 6752 37473 6780
rect 30892 6740 30898 6752
rect 37461 6749 37473 6752
rect 37507 6749 37519 6783
rect 37461 6743 37519 6749
rect 37550 6740 37556 6792
rect 37608 6780 37614 6792
rect 38010 6780 38016 6792
rect 37608 6752 38016 6780
rect 37608 6740 37614 6752
rect 38010 6740 38016 6752
rect 38068 6740 38074 6792
rect 38194 6740 38200 6792
rect 38252 6740 38258 6792
rect 38470 6740 38476 6792
rect 38528 6740 38534 6792
rect 39224 6789 39252 6820
rect 38841 6783 38899 6789
rect 38841 6749 38853 6783
rect 38887 6749 38899 6783
rect 38841 6743 38899 6749
rect 39209 6783 39267 6789
rect 39209 6749 39221 6783
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 27982 6712 27988 6724
rect 24780 6684 25636 6712
rect 26620 6684 27988 6712
rect 26620 6656 26648 6684
rect 27982 6672 27988 6684
rect 28040 6672 28046 6724
rect 38105 6715 38163 6721
rect 38105 6681 38117 6715
rect 38151 6712 38163 6715
rect 38856 6712 38884 6743
rect 40034 6712 40040 6724
rect 38151 6684 38884 6712
rect 39040 6684 40040 6712
rect 38151 6681 38163 6684
rect 38105 6675 38163 6681
rect 4028 6616 7788 6644
rect 4028 6604 4034 6616
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11020 6616 11437 6644
rect 11020 6604 11026 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 12710 6604 12716 6656
rect 12768 6604 12774 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 14826 6644 14832 6656
rect 13780 6616 14832 6644
rect 13780 6604 13786 6616
rect 14826 6604 14832 6616
rect 14884 6644 14890 6656
rect 16666 6644 16672 6656
rect 14884 6616 16672 6644
rect 14884 6604 14890 6616
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 21910 6644 21916 6656
rect 17828 6616 21916 6644
rect 17828 6604 17834 6616
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 24578 6644 24584 6656
rect 23348 6616 24584 6644
rect 23348 6604 23354 6616
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 25038 6604 25044 6656
rect 25096 6644 25102 6656
rect 25222 6644 25228 6656
rect 25096 6616 25228 6644
rect 25096 6604 25102 6616
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 25314 6604 25320 6656
rect 25372 6644 25378 6656
rect 25958 6644 25964 6656
rect 25372 6616 25964 6644
rect 25372 6604 25378 6616
rect 25958 6604 25964 6616
rect 26016 6604 26022 6656
rect 26237 6647 26295 6653
rect 26237 6613 26249 6647
rect 26283 6644 26295 6647
rect 26602 6644 26608 6656
rect 26283 6616 26608 6644
rect 26283 6613 26295 6616
rect 26237 6607 26295 6613
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 27430 6604 27436 6656
rect 27488 6604 27494 6656
rect 27801 6647 27859 6653
rect 27801 6613 27813 6647
rect 27847 6644 27859 6647
rect 27890 6644 27896 6656
rect 27847 6616 27896 6644
rect 27847 6613 27859 6616
rect 27801 6607 27859 6613
rect 27890 6604 27896 6616
rect 27948 6604 27954 6656
rect 37274 6604 37280 6656
rect 37332 6604 37338 6656
rect 37550 6604 37556 6656
rect 37608 6644 37614 6656
rect 38013 6647 38071 6653
rect 38013 6644 38025 6647
rect 37608 6616 38025 6644
rect 37608 6604 37614 6616
rect 38013 6613 38025 6616
rect 38059 6613 38071 6647
rect 38013 6607 38071 6613
rect 38378 6604 38384 6656
rect 38436 6604 38442 6656
rect 38654 6604 38660 6656
rect 38712 6604 38718 6656
rect 39040 6653 39068 6684
rect 40034 6672 40040 6684
rect 40092 6672 40098 6724
rect 39025 6647 39083 6653
rect 39025 6613 39037 6647
rect 39071 6613 39083 6647
rect 39025 6607 39083 6613
rect 39393 6647 39451 6653
rect 39393 6613 39405 6647
rect 39439 6644 39451 6647
rect 39482 6644 39488 6656
rect 39439 6616 39488 6644
rect 39439 6613 39451 6616
rect 39393 6607 39451 6613
rect 39482 6604 39488 6616
rect 39540 6604 39546 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 5442 6440 5448 6452
rect 1627 6412 5448 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 13446 6440 13452 6452
rect 5684 6412 13452 6440
rect 5684 6400 5690 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 15102 6440 15108 6452
rect 14783 6412 15108 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 16206 6400 16212 6452
rect 16264 6440 16270 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16264 6412 16957 6440
rect 16264 6400 16270 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 16945 6403 17003 6409
rect 18969 6443 19027 6449
rect 18969 6409 18981 6443
rect 19015 6440 19027 6443
rect 19702 6440 19708 6452
rect 19015 6412 19708 6440
rect 19015 6409 19027 6412
rect 18969 6403 19027 6409
rect 19702 6400 19708 6412
rect 19760 6440 19766 6452
rect 20438 6440 20444 6452
rect 19760 6412 20444 6440
rect 19760 6400 19766 6412
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 21542 6440 21548 6452
rect 20680 6412 21548 6440
rect 20680 6400 20686 6412
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 21818 6400 21824 6452
rect 21876 6400 21882 6452
rect 22094 6400 22100 6452
rect 22152 6400 22158 6452
rect 24302 6400 24308 6452
rect 24360 6440 24366 6452
rect 37550 6440 37556 6452
rect 24360 6412 37556 6440
rect 24360 6400 24366 6412
rect 37550 6400 37556 6412
rect 37608 6400 37614 6452
rect 37642 6400 37648 6452
rect 37700 6400 37706 6452
rect 39393 6443 39451 6449
rect 39393 6409 39405 6443
rect 39439 6440 39451 6443
rect 39574 6440 39580 6452
rect 39439 6412 39580 6440
rect 39439 6409 39451 6412
rect 39393 6403 39451 6409
rect 39574 6400 39580 6412
rect 39632 6400 39638 6452
rect 2590 6332 2596 6384
rect 2648 6372 2654 6384
rect 2648 6344 2774 6372
rect 2648 6332 2654 6344
rect 198 6264 204 6316
rect 256 6304 262 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 256 6276 1409 6304
rect 256 6264 262 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 2746 6304 2774 6344
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 9398 6372 9404 6384
rect 5592 6344 9404 6372
rect 5592 6332 5598 6344
rect 9398 6332 9404 6344
rect 9456 6332 9462 6384
rect 10686 6372 10692 6384
rect 9568 6344 10692 6372
rect 3145 6307 3203 6313
rect 3145 6304 3157 6307
rect 2746 6276 3157 6304
rect 1673 6267 1731 6273
rect 3145 6273 3157 6276
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6304 6055 6307
rect 6043 6276 6500 6304
rect 6043 6273 6055 6276
rect 5997 6267 6055 6273
rect 842 6196 848 6248
rect 900 6236 906 6248
rect 1688 6236 1716 6267
rect 900 6208 1716 6236
rect 900 6196 906 6208
rect 2498 6196 2504 6248
rect 2556 6236 2562 6248
rect 2869 6239 2927 6245
rect 2869 6236 2881 6239
rect 2556 6208 2881 6236
rect 2556 6196 2562 6208
rect 2869 6205 2881 6208
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 6129 6236 6157 6276
rect 5132 6208 6157 6236
rect 6472 6236 6500 6276
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 8478 6304 8484 6316
rect 6604 6276 8484 6304
rect 6604 6264 6610 6276
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9568 6313 9596 6344
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15068 6344 18276 6372
rect 15068 6332 15074 6344
rect 9523 6307 9596 6313
rect 10134 6312 10140 6316
rect 9523 6273 9535 6307
rect 9569 6276 9596 6307
rect 10102 6306 10140 6312
rect 9569 6273 9581 6276
rect 9523 6267 9581 6273
rect 10102 6272 10114 6306
rect 10102 6266 10140 6272
rect 10134 6264 10140 6266
rect 10192 6264 10198 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 13872 6276 14565 6304
rect 13872 6264 13878 6276
rect 14553 6273 14565 6276
rect 14599 6304 14611 6307
rect 15105 6307 15163 6313
rect 15105 6304 15117 6307
rect 14599 6276 15117 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 15105 6273 15117 6276
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 16942 6264 16948 6316
rect 17000 6304 17006 6316
rect 17129 6307 17187 6313
rect 17129 6304 17141 6307
rect 17000 6276 17141 6304
rect 17000 6264 17006 6276
rect 17129 6273 17141 6276
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 18248 6313 18276 6344
rect 19794 6332 19800 6384
rect 19852 6332 19858 6384
rect 21468 6344 22324 6372
rect 17957 6307 18015 6313
rect 17957 6304 17969 6307
rect 17736 6276 17969 6304
rect 17736 6264 17742 6276
rect 17957 6273 17969 6276
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 18279 6276 19073 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 19061 6273 19073 6276
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 19751 6276 19932 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 9769 6239 9827 6245
rect 6472 6208 9444 6236
rect 5132 6196 5138 6208
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6168 1915 6171
rect 2682 6168 2688 6180
rect 1903 6140 2688 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 2682 6128 2688 6140
rect 2740 6128 2746 6180
rect 2774 6128 2780 6180
rect 2832 6128 2838 6180
rect 9214 6168 9220 6180
rect 3528 6140 9220 6168
rect 1578 6060 1584 6112
rect 1636 6100 1642 6112
rect 3528 6100 3556 6140
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 9416 6168 9444 6208
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 9999 6239 10057 6245
rect 9999 6236 10011 6239
rect 9815 6208 10011 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 9999 6205 10011 6208
rect 10045 6205 10057 6239
rect 9999 6199 10057 6205
rect 14826 6196 14832 6248
rect 14884 6196 14890 6248
rect 13446 6168 13452 6180
rect 9416 6140 13452 6168
rect 13446 6128 13452 6140
rect 13504 6128 13510 6180
rect 19426 6128 19432 6180
rect 19484 6168 19490 6180
rect 19521 6171 19579 6177
rect 19521 6168 19533 6171
rect 19484 6140 19533 6168
rect 19484 6128 19490 6140
rect 19521 6137 19533 6140
rect 19567 6137 19579 6171
rect 19521 6131 19579 6137
rect 1636 6072 3556 6100
rect 3881 6103 3939 6109
rect 1636 6060 1642 6072
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 5810 6100 5816 6112
rect 3927 6072 5816 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 5810 6060 5816 6072
rect 5868 6060 5874 6112
rect 6178 6060 6184 6112
rect 6236 6060 6242 6112
rect 6733 6103 6791 6109
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 8294 6100 8300 6112
rect 6779 6072 8300 6100
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 9309 6103 9367 6109
rect 9309 6100 9321 6103
rect 9180 6072 9321 6100
rect 9180 6060 9186 6072
rect 9309 6069 9321 6072
rect 9355 6069 9367 6103
rect 9309 6063 9367 6069
rect 9674 6060 9680 6112
rect 9732 6060 9738 6112
rect 15838 6060 15844 6112
rect 15896 6060 15902 6112
rect 19242 6060 19248 6112
rect 19300 6060 19306 6112
rect 19904 6100 19932 6276
rect 20438 6264 20444 6316
rect 20496 6264 20502 6316
rect 20622 6313 20628 6316
rect 20600 6307 20628 6313
rect 20600 6273 20612 6307
rect 20600 6267 20628 6273
rect 20622 6264 20628 6267
rect 20680 6264 20686 6316
rect 21468 6313 21496 6344
rect 22296 6313 22324 6344
rect 23382 6332 23388 6384
rect 23440 6372 23446 6384
rect 25590 6372 25596 6384
rect 23440 6344 25596 6372
rect 23440 6332 23446 6344
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 25866 6332 25872 6384
rect 25924 6372 25930 6384
rect 27706 6372 27712 6384
rect 25924 6344 27712 6372
rect 25924 6332 25930 6344
rect 27706 6332 27712 6344
rect 27764 6332 27770 6384
rect 27982 6332 27988 6384
rect 28040 6372 28046 6384
rect 28040 6344 37872 6372
rect 28040 6332 28046 6344
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 21637 6307 21695 6313
rect 21637 6273 21649 6307
rect 21683 6304 21695 6307
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21683 6276 22017 6304
rect 21683 6273 21695 6276
rect 21637 6267 21695 6273
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6304 22339 6307
rect 23934 6304 23940 6316
rect 22327 6276 23940 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 20717 6239 20775 6245
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 22020 6236 22048 6267
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 24210 6264 24216 6316
rect 24268 6304 24274 6316
rect 26418 6304 26424 6316
rect 24268 6276 26424 6304
rect 24268 6264 24274 6276
rect 26418 6264 26424 6276
rect 26476 6264 26482 6316
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 30469 6307 30527 6313
rect 30469 6304 30481 6307
rect 27580 6276 30481 6304
rect 27580 6264 27586 6276
rect 30469 6273 30481 6276
rect 30515 6273 30527 6307
rect 30469 6267 30527 6273
rect 30650 6264 30656 6316
rect 30708 6264 30714 6316
rect 30742 6264 30748 6316
rect 30800 6304 30806 6316
rect 37844 6313 37872 6344
rect 38378 6332 38384 6384
rect 38436 6372 38442 6384
rect 39482 6372 39488 6384
rect 38436 6344 39488 6372
rect 38436 6332 38442 6344
rect 39482 6332 39488 6344
rect 39540 6332 39546 6384
rect 33873 6307 33931 6313
rect 33873 6304 33885 6307
rect 30800 6276 33885 6304
rect 30800 6264 30806 6276
rect 33873 6273 33885 6276
rect 33919 6273 33931 6307
rect 33873 6267 33931 6273
rect 37461 6307 37519 6313
rect 37461 6273 37473 6307
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 37829 6307 37887 6313
rect 37829 6273 37841 6307
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 38473 6307 38531 6313
rect 38473 6273 38485 6307
rect 38519 6273 38531 6307
rect 38473 6267 38531 6273
rect 25406 6236 25412 6248
rect 20763 6208 21128 6236
rect 22020 6208 25412 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 20898 6128 20904 6180
rect 20956 6168 20962 6180
rect 20993 6171 21051 6177
rect 20993 6168 21005 6171
rect 20956 6140 21005 6168
rect 20956 6128 20962 6140
rect 20993 6137 21005 6140
rect 21039 6137 21051 6171
rect 20993 6131 21051 6137
rect 21100 6168 21128 6208
rect 25406 6196 25412 6208
rect 25464 6196 25470 6248
rect 26694 6196 26700 6248
rect 26752 6236 26758 6248
rect 37476 6236 37504 6267
rect 26752 6208 37504 6236
rect 26752 6196 26758 6208
rect 37550 6196 37556 6248
rect 37608 6236 37614 6248
rect 38488 6236 38516 6267
rect 38838 6264 38844 6316
rect 38896 6264 38902 6316
rect 38930 6264 38936 6316
rect 38988 6304 38994 6316
rect 39209 6307 39267 6313
rect 39209 6304 39221 6307
rect 38988 6276 39221 6304
rect 38988 6264 38994 6276
rect 39209 6273 39221 6276
rect 39255 6273 39267 6307
rect 39209 6267 39267 6273
rect 37608 6208 38516 6236
rect 37608 6196 37614 6208
rect 25774 6168 25780 6180
rect 21100 6140 25780 6168
rect 21100 6100 21128 6140
rect 25774 6128 25780 6140
rect 25832 6128 25838 6180
rect 27338 6128 27344 6180
rect 27396 6168 27402 6180
rect 27522 6168 27528 6180
rect 27396 6140 27528 6168
rect 27396 6128 27402 6140
rect 27522 6128 27528 6140
rect 27580 6128 27586 6180
rect 27798 6128 27804 6180
rect 27856 6168 27862 6180
rect 30285 6171 30343 6177
rect 30285 6168 30297 6171
rect 27856 6140 30297 6168
rect 27856 6128 27862 6140
rect 30285 6137 30297 6140
rect 30331 6137 30343 6171
rect 30285 6131 30343 6137
rect 34054 6128 34060 6180
rect 34112 6128 34118 6180
rect 39025 6171 39083 6177
rect 39025 6137 39037 6171
rect 39071 6168 39083 6171
rect 39666 6168 39672 6180
rect 39071 6140 39672 6168
rect 39071 6137 39083 6140
rect 39025 6131 39083 6137
rect 39666 6128 39672 6140
rect 39724 6128 39730 6180
rect 19904 6072 21128 6100
rect 21910 6060 21916 6112
rect 21968 6100 21974 6112
rect 24210 6100 24216 6112
rect 21968 6072 24216 6100
rect 21968 6060 21974 6072
rect 24210 6060 24216 6072
rect 24268 6060 24274 6112
rect 24394 6060 24400 6112
rect 24452 6100 24458 6112
rect 29730 6100 29736 6112
rect 24452 6072 29736 6100
rect 24452 6060 24458 6072
rect 29730 6060 29736 6072
rect 29788 6060 29794 6112
rect 30834 6060 30840 6112
rect 30892 6060 30898 6112
rect 37369 6103 37427 6109
rect 37369 6069 37381 6103
rect 37415 6100 37427 6103
rect 37734 6100 37740 6112
rect 37415 6072 37740 6100
rect 37415 6069 37427 6072
rect 37369 6063 37427 6069
rect 37734 6060 37740 6072
rect 37792 6060 37798 6112
rect 38010 6060 38016 6112
rect 38068 6100 38074 6112
rect 38470 6100 38476 6112
rect 38068 6072 38476 6100
rect 38068 6060 38074 6072
rect 38470 6060 38476 6072
rect 38528 6060 38534 6112
rect 38654 6060 38660 6112
rect 38712 6060 38718 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 6822 5896 6828 5908
rect 2556 5868 6828 5896
rect 2556 5856 2562 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 14550 5896 14556 5908
rect 8956 5868 14556 5896
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 5626 5828 5632 5840
rect 1903 5800 5632 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 5626 5788 5632 5800
rect 5684 5788 5690 5840
rect 6730 5788 6736 5840
rect 6788 5828 6794 5840
rect 8956 5828 8984 5868
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 16942 5856 16948 5908
rect 17000 5856 17006 5908
rect 23382 5896 23388 5908
rect 17926 5868 23388 5896
rect 6788 5800 8984 5828
rect 6788 5788 6794 5800
rect 10134 5788 10140 5840
rect 10192 5788 10198 5840
rect 10686 5788 10692 5840
rect 10744 5788 10750 5840
rect 12345 5831 12403 5837
rect 12345 5797 12357 5831
rect 12391 5797 12403 5831
rect 12345 5791 12403 5797
rect 5074 5720 5080 5772
rect 5132 5720 5138 5772
rect 5258 5720 5264 5772
rect 5316 5720 5322 5772
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 10152 5760 10180 5788
rect 10962 5760 10968 5772
rect 5767 5732 9904 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 750 5652 756 5704
rect 808 5692 814 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 808 5664 1409 5692
rect 808 5652 814 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 842 5584 848 5636
rect 900 5624 906 5636
rect 1688 5624 1716 5655
rect 3142 5652 3148 5704
rect 3200 5652 3206 5704
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 6086 5652 6092 5704
rect 6144 5701 6150 5704
rect 6144 5695 6172 5701
rect 6160 5661 6172 5695
rect 6144 5655 6172 5661
rect 6144 5652 6150 5655
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 9674 5692 9680 5704
rect 6963 5664 9680 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 900 5596 1716 5624
rect 900 5584 906 5596
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 4154 5556 4160 5568
rect 3375 5528 4160 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 6086 5556 6092 5568
rect 5031 5528 6092 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 6086 5516 6092 5528
rect 6144 5556 6150 5568
rect 6730 5556 6736 5568
rect 6144 5528 6736 5556
rect 6144 5516 6150 5528
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 9876 5556 9904 5732
rect 10060 5732 10180 5760
rect 10428 5732 10968 5760
rect 10060 5701 10088 5732
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 10428 5692 10456 5732
rect 10962 5720 10968 5732
rect 11020 5760 11026 5772
rect 12360 5760 12388 5791
rect 13446 5788 13452 5840
rect 13504 5828 13510 5840
rect 17926 5828 17954 5868
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 37826 5856 37832 5908
rect 37884 5896 37890 5908
rect 38289 5899 38347 5905
rect 38289 5896 38301 5899
rect 37884 5868 38301 5896
rect 37884 5856 37890 5868
rect 38289 5865 38301 5868
rect 38335 5865 38347 5899
rect 38289 5859 38347 5865
rect 38470 5856 38476 5908
rect 38528 5896 38534 5908
rect 38565 5899 38623 5905
rect 38565 5896 38577 5899
rect 38528 5868 38577 5896
rect 38528 5856 38534 5868
rect 38565 5865 38577 5868
rect 38611 5865 38623 5899
rect 38565 5859 38623 5865
rect 39390 5856 39396 5908
rect 39448 5856 39454 5908
rect 13504 5800 17954 5828
rect 13504 5788 13510 5800
rect 19242 5788 19248 5840
rect 19300 5828 19306 5840
rect 24394 5828 24400 5840
rect 19300 5800 24400 5828
rect 19300 5788 19306 5800
rect 24394 5788 24400 5800
rect 24452 5788 24458 5840
rect 25409 5831 25467 5837
rect 25409 5797 25421 5831
rect 25455 5828 25467 5831
rect 27801 5831 27859 5837
rect 25455 5800 27752 5828
rect 25455 5797 25467 5800
rect 25409 5791 25467 5797
rect 11020 5732 11100 5760
rect 11020 5720 11026 5732
rect 11072 5701 11100 5732
rect 11348 5732 12388 5760
rect 13357 5763 13415 5769
rect 11348 5701 11376 5732
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13722 5760 13728 5772
rect 13403 5732 13728 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 15896 5732 17509 5760
rect 15896 5720 15902 5732
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 21910 5760 21916 5772
rect 17497 5723 17555 5729
rect 19306 5732 21916 5760
rect 10192 5664 10456 5692
rect 10551 5695 10609 5701
rect 10192 5652 10198 5664
rect 10551 5661 10563 5695
rect 10597 5692 10609 5695
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10597 5664 10885 5692
rect 10597 5661 10609 5664
rect 10551 5655 10609 5661
rect 10873 5661 10885 5664
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 10318 5584 10324 5636
rect 10376 5584 10382 5636
rect 10410 5584 10416 5636
rect 10468 5584 10474 5636
rect 10594 5556 10600 5568
rect 9876 5528 10600 5556
rect 10594 5516 10600 5528
rect 10652 5556 10658 5568
rect 11348 5556 11376 5655
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 11664 5664 13093 5692
rect 11664 5652 11670 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13096 5624 13124 5655
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 19306 5692 19334 5732
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 22002 5720 22008 5772
rect 22060 5760 22066 5772
rect 24302 5760 24308 5772
rect 22060 5732 24308 5760
rect 22060 5720 22066 5732
rect 24302 5720 24308 5732
rect 24360 5720 24366 5772
rect 26528 5732 26832 5760
rect 14608 5664 19334 5692
rect 20257 5695 20315 5701
rect 14608 5652 14614 5664
rect 20257 5661 20269 5695
rect 20303 5692 20315 5695
rect 20622 5692 20628 5704
rect 20303 5664 20628 5692
rect 20303 5661 20315 5664
rect 20257 5655 20315 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 23290 5652 23296 5704
rect 23348 5692 23354 5704
rect 23569 5695 23627 5701
rect 23569 5692 23581 5695
rect 23348 5664 23581 5692
rect 23348 5652 23354 5664
rect 23569 5661 23581 5664
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 23845 5695 23903 5701
rect 23845 5661 23857 5695
rect 23891 5694 23903 5695
rect 23934 5694 23940 5704
rect 23891 5666 23940 5694
rect 23891 5661 23903 5666
rect 23845 5655 23903 5661
rect 23934 5652 23940 5666
rect 23992 5692 23998 5704
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 23992 5664 24409 5692
rect 23992 5652 23998 5664
rect 24397 5661 24409 5664
rect 24443 5661 24455 5695
rect 24397 5655 24455 5661
rect 24578 5652 24584 5704
rect 24636 5692 24642 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 24636 5664 24685 5692
rect 24636 5652 24642 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25958 5692 25964 5704
rect 24820 5664 25964 5692
rect 24820 5652 24826 5664
rect 25958 5652 25964 5664
rect 26016 5652 26022 5704
rect 26142 5701 26148 5704
rect 26115 5695 26148 5701
rect 26115 5661 26127 5695
rect 26115 5655 26148 5661
rect 26142 5652 26148 5655
rect 26200 5652 26206 5704
rect 26421 5695 26479 5701
rect 26421 5692 26433 5695
rect 26252 5664 26433 5692
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13096 5596 13553 5624
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 13722 5584 13728 5636
rect 13780 5584 13786 5636
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 15378 5624 15384 5636
rect 14424 5596 15384 5624
rect 14424 5584 14430 5596
rect 15378 5584 15384 5596
rect 15436 5624 15442 5636
rect 17402 5624 17408 5636
rect 15436 5596 17408 5624
rect 15436 5584 15442 5596
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 26252 5624 26280 5664
rect 26421 5661 26433 5664
rect 26467 5661 26479 5695
rect 26421 5655 26479 5661
rect 19260 5596 20208 5624
rect 10652 5528 11376 5556
rect 17313 5559 17371 5565
rect 10652 5516 10658 5528
rect 17313 5525 17325 5559
rect 17359 5556 17371 5559
rect 18414 5556 18420 5568
rect 17359 5528 18420 5556
rect 17359 5525 17371 5528
rect 17313 5519 17371 5525
rect 18414 5516 18420 5528
rect 18472 5556 18478 5568
rect 19260 5556 19288 5596
rect 18472 5528 19288 5556
rect 18472 5516 18478 5528
rect 19610 5516 19616 5568
rect 19668 5556 19674 5568
rect 20073 5559 20131 5565
rect 20073 5556 20085 5559
rect 19668 5528 20085 5556
rect 19668 5516 19674 5528
rect 20073 5525 20085 5528
rect 20119 5525 20131 5559
rect 20180 5556 20208 5596
rect 20456 5596 26280 5624
rect 26329 5627 26387 5633
rect 20456 5556 20484 5596
rect 26329 5593 26341 5627
rect 26375 5624 26387 5627
rect 26528 5624 26556 5732
rect 26602 5652 26608 5704
rect 26660 5652 26666 5704
rect 26375 5596 26556 5624
rect 26804 5624 26832 5732
rect 26878 5652 26884 5704
rect 26936 5652 26942 5704
rect 26988 5692 27016 5800
rect 27065 5763 27123 5769
rect 27065 5729 27077 5763
rect 27111 5760 27123 5763
rect 27111 5732 27568 5760
rect 27111 5729 27123 5732
rect 27065 5723 27123 5729
rect 27338 5701 27344 5704
rect 27157 5695 27215 5701
rect 27157 5692 27169 5695
rect 26988 5664 27169 5692
rect 27157 5661 27169 5664
rect 27203 5661 27215 5695
rect 27157 5655 27215 5661
rect 27305 5695 27344 5701
rect 27305 5661 27317 5695
rect 27305 5655 27344 5661
rect 27338 5652 27344 5655
rect 27396 5652 27402 5704
rect 27430 5652 27436 5704
rect 27488 5652 27494 5704
rect 27540 5692 27568 5732
rect 27622 5695 27680 5701
rect 27622 5692 27634 5695
rect 27540 5664 27634 5692
rect 27622 5661 27634 5664
rect 27668 5661 27680 5695
rect 27622 5655 27680 5661
rect 27525 5627 27583 5633
rect 27525 5624 27537 5627
rect 26804 5596 27537 5624
rect 26375 5593 26387 5596
rect 26329 5587 26387 5593
rect 27525 5593 27537 5596
rect 27571 5593 27583 5627
rect 27724 5624 27752 5800
rect 27801 5797 27813 5831
rect 27847 5797 27859 5831
rect 27801 5791 27859 5797
rect 27816 5692 27844 5791
rect 28074 5788 28080 5840
rect 28132 5828 28138 5840
rect 30742 5828 30748 5840
rect 28132 5800 30748 5828
rect 28132 5788 28138 5800
rect 30742 5788 30748 5800
rect 30800 5788 30806 5840
rect 30834 5788 30840 5840
rect 30892 5828 30898 5840
rect 38654 5828 38660 5840
rect 30892 5800 38660 5828
rect 30892 5788 30898 5800
rect 38654 5788 38660 5800
rect 38712 5788 38718 5840
rect 39025 5831 39083 5837
rect 39025 5797 39037 5831
rect 39071 5828 39083 5831
rect 39942 5828 39948 5840
rect 39071 5800 39948 5828
rect 39071 5797 39083 5800
rect 39025 5791 39083 5797
rect 39942 5788 39948 5800
rect 40000 5788 40006 5840
rect 29181 5763 29239 5769
rect 29181 5729 29193 5763
rect 29227 5760 29239 5763
rect 29641 5763 29699 5769
rect 29641 5760 29653 5763
rect 29227 5732 29653 5760
rect 29227 5729 29239 5732
rect 29181 5723 29239 5729
rect 29641 5729 29653 5732
rect 29687 5729 29699 5763
rect 29641 5723 29699 5729
rect 31110 5720 31116 5772
rect 31168 5760 31174 5772
rect 31168 5732 38792 5760
rect 31168 5720 31174 5732
rect 28905 5695 28963 5701
rect 28905 5692 28917 5695
rect 27816 5664 28917 5692
rect 28905 5661 28917 5664
rect 28951 5661 28963 5695
rect 28905 5655 28963 5661
rect 29089 5695 29147 5701
rect 29089 5661 29101 5695
rect 29135 5692 29147 5695
rect 29362 5692 29368 5704
rect 29135 5664 29368 5692
rect 29135 5661 29147 5664
rect 29089 5655 29147 5661
rect 29362 5652 29368 5664
rect 29420 5652 29426 5704
rect 29549 5695 29607 5701
rect 29549 5661 29561 5695
rect 29595 5661 29607 5695
rect 29549 5655 29607 5661
rect 29564 5624 29592 5655
rect 29730 5652 29736 5704
rect 29788 5692 29794 5704
rect 37274 5692 37280 5704
rect 29788 5664 37280 5692
rect 29788 5652 29794 5664
rect 37274 5652 37280 5664
rect 37332 5652 37338 5704
rect 37366 5652 37372 5704
rect 37424 5692 37430 5704
rect 38764 5701 38792 5732
rect 38473 5695 38531 5701
rect 38473 5692 38485 5695
rect 37424 5664 38485 5692
rect 37424 5652 37430 5664
rect 38473 5661 38485 5664
rect 38519 5661 38531 5695
rect 38473 5655 38531 5661
rect 38749 5695 38807 5701
rect 38749 5661 38761 5695
rect 38795 5661 38807 5695
rect 38749 5655 38807 5661
rect 38838 5652 38844 5704
rect 38896 5652 38902 5704
rect 39206 5652 39212 5704
rect 39264 5652 39270 5704
rect 27724 5596 29592 5624
rect 27525 5587 27583 5593
rect 20180 5528 20484 5556
rect 23753 5559 23811 5565
rect 20073 5519 20131 5525
rect 23753 5525 23765 5559
rect 23799 5556 23811 5559
rect 23842 5556 23848 5568
rect 23799 5528 23848 5556
rect 23799 5525 23811 5528
rect 23753 5519 23811 5525
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 24029 5559 24087 5565
rect 24029 5525 24041 5559
rect 24075 5556 24087 5559
rect 24118 5556 24124 5568
rect 24075 5528 24124 5556
rect 24075 5525 24087 5528
rect 24029 5519 24087 5525
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 26142 5516 26148 5568
rect 26200 5556 26206 5568
rect 26602 5556 26608 5568
rect 26200 5528 26608 5556
rect 26200 5516 26206 5528
rect 26602 5516 26608 5528
rect 26660 5516 26666 5568
rect 27890 5516 27896 5568
rect 27948 5556 27954 5568
rect 28721 5559 28779 5565
rect 28721 5556 28733 5559
rect 27948 5528 28733 5556
rect 27948 5516 27954 5528
rect 28721 5525 28733 5528
rect 28767 5525 28779 5559
rect 28721 5519 28779 5525
rect 30006 5516 30012 5568
rect 30064 5556 30070 5568
rect 34146 5556 34152 5568
rect 30064 5528 34152 5556
rect 30064 5516 30070 5528
rect 34146 5516 34152 5528
rect 34204 5516 34210 5568
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 14918 5352 14924 5364
rect 4479 5324 14924 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 24854 5352 24860 5364
rect 17236 5324 24860 5352
rect 1670 5244 1676 5296
rect 1728 5284 1734 5296
rect 17236 5284 17264 5324
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 26329 5355 26387 5361
rect 26329 5321 26341 5355
rect 26375 5352 26387 5355
rect 26418 5352 26424 5364
rect 26375 5324 26424 5352
rect 26375 5321 26387 5324
rect 26329 5315 26387 5321
rect 26418 5312 26424 5324
rect 26476 5312 26482 5364
rect 26878 5312 26884 5364
rect 26936 5352 26942 5364
rect 28074 5352 28080 5364
rect 26936 5324 28080 5352
rect 26936 5312 26942 5324
rect 28074 5312 28080 5324
rect 28132 5312 28138 5364
rect 33413 5355 33471 5361
rect 33413 5321 33425 5355
rect 33459 5352 33471 5355
rect 33686 5352 33692 5364
rect 33459 5324 33692 5352
rect 33459 5321 33471 5324
rect 33413 5315 33471 5321
rect 33686 5312 33692 5324
rect 33744 5312 33750 5364
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 1728 5256 17264 5284
rect 1728 5244 1734 5256
rect 19426 5244 19432 5296
rect 19484 5284 19490 5296
rect 24118 5284 24124 5296
rect 19484 5256 24124 5284
rect 19484 5244 19490 5256
rect 24118 5244 24124 5256
rect 24176 5284 24182 5296
rect 25038 5284 25044 5296
rect 24176 5256 25044 5284
rect 24176 5244 24182 5256
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 25130 5244 25136 5296
rect 25188 5284 25194 5296
rect 25188 5256 26648 5284
rect 25188 5244 25194 5256
rect 750 5176 756 5228
rect 808 5216 814 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 808 5188 1409 5216
rect 808 5176 814 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 6086 5216 6092 5228
rect 4295 5188 6092 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 7894 5219 7952 5225
rect 7894 5185 7906 5219
rect 7940 5216 7952 5219
rect 8386 5216 8392 5228
rect 7940 5188 8392 5216
rect 7940 5185 7952 5188
rect 7894 5179 7952 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8754 5176 8760 5228
rect 8812 5176 8818 5228
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5216 8999 5219
rect 8987 5188 10088 5216
rect 8987 5185 8999 5188
rect 8941 5179 8999 5185
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 8495 5148 8523 5176
rect 5868 5120 8523 5148
rect 5868 5108 5874 5120
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 10060 5080 10088 5188
rect 10594 5176 10600 5228
rect 10652 5225 10658 5228
rect 10652 5219 10685 5225
rect 10673 5185 10685 5219
rect 10652 5179 10685 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10652 5176 10658 5179
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10796 5148 10824 5179
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 23750 5216 23756 5228
rect 11020 5188 23756 5216
rect 11020 5176 11026 5188
rect 23750 5176 23756 5188
rect 23808 5176 23814 5228
rect 25958 5176 25964 5228
rect 26016 5216 26022 5228
rect 26513 5219 26571 5225
rect 26513 5216 26525 5219
rect 26016 5188 26525 5216
rect 26016 5176 26022 5188
rect 26513 5185 26525 5188
rect 26559 5185 26571 5219
rect 26620 5216 26648 5256
rect 27522 5244 27528 5296
rect 27580 5284 27586 5296
rect 38930 5284 38936 5296
rect 27580 5256 38936 5284
rect 27580 5244 27586 5256
rect 38930 5244 38936 5256
rect 38988 5244 38994 5296
rect 28718 5216 28724 5228
rect 26620 5188 28724 5216
rect 26513 5179 26571 5185
rect 28718 5176 28724 5188
rect 28776 5176 28782 5228
rect 32493 5219 32551 5225
rect 32493 5216 32505 5219
rect 31726 5188 32505 5216
rect 12250 5148 12256 5160
rect 10284 5120 12256 5148
rect 10284 5108 10290 5120
rect 12250 5108 12256 5120
rect 12308 5148 12314 5160
rect 20530 5148 20536 5160
rect 12308 5120 20536 5148
rect 12308 5108 12314 5120
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 21542 5148 21548 5160
rect 20864 5120 21548 5148
rect 20864 5108 20870 5120
rect 21542 5108 21548 5120
rect 21600 5108 21606 5160
rect 22002 5108 22008 5160
rect 22060 5148 22066 5160
rect 24762 5148 24768 5160
rect 22060 5120 24768 5148
rect 22060 5108 22066 5120
rect 24762 5108 24768 5120
rect 24820 5108 24826 5160
rect 25130 5108 25136 5160
rect 25188 5148 25194 5160
rect 31726 5148 31754 5188
rect 32493 5185 32505 5188
rect 32539 5185 32551 5219
rect 32493 5179 32551 5185
rect 33229 5219 33287 5225
rect 33229 5185 33241 5219
rect 33275 5216 33287 5219
rect 33410 5216 33416 5228
rect 33275 5188 33416 5216
rect 33275 5185 33287 5188
rect 33229 5179 33287 5185
rect 33410 5176 33416 5188
rect 33468 5176 33474 5228
rect 33505 5219 33563 5225
rect 33505 5185 33517 5219
rect 33551 5216 33563 5219
rect 37734 5216 37740 5228
rect 33551 5188 37740 5216
rect 33551 5185 33563 5188
rect 33505 5179 33563 5185
rect 37734 5176 37740 5188
rect 37792 5176 37798 5228
rect 38838 5176 38844 5228
rect 38896 5176 38902 5228
rect 39206 5176 39212 5228
rect 39264 5176 39270 5228
rect 38746 5148 38752 5160
rect 25188 5120 31754 5148
rect 32600 5120 38752 5148
rect 25188 5108 25194 5120
rect 11514 5080 11520 5092
rect 2832 5052 8432 5080
rect 10060 5052 11520 5080
rect 2832 5040 2838 5052
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 7190 5012 7196 5024
rect 1627 4984 7196 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7791 5015 7849 5021
rect 7791 5012 7803 5015
rect 7524 4984 7803 5012
rect 7524 4972 7530 4984
rect 7791 4981 7803 4984
rect 7837 4981 7849 5015
rect 7791 4975 7849 4981
rect 8294 4972 8300 5024
rect 8352 4972 8358 5024
rect 8404 5012 8432 5052
rect 11514 5040 11520 5052
rect 11572 5040 11578 5092
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 12860 5052 18736 5080
rect 12860 5040 12866 5052
rect 10410 5012 10416 5024
rect 8404 4984 10416 5012
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 10560 4984 10609 5012
rect 10560 4972 10566 4984
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 10597 4975 10655 4981
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 18598 5012 18604 5024
rect 14700 4984 18604 5012
rect 14700 4972 14706 4984
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 18708 5012 18736 5052
rect 19058 5040 19064 5092
rect 19116 5080 19122 5092
rect 32600 5080 32628 5120
rect 38746 5108 38752 5120
rect 38804 5108 38810 5160
rect 19116 5052 32628 5080
rect 32677 5083 32735 5089
rect 19116 5040 19122 5052
rect 32677 5049 32689 5083
rect 32723 5080 32735 5083
rect 33778 5080 33784 5092
rect 32723 5052 33784 5080
rect 32723 5049 32735 5052
rect 32677 5043 32735 5049
rect 33778 5040 33784 5052
rect 33836 5040 33842 5092
rect 38286 5080 38292 5092
rect 33888 5052 38292 5080
rect 20806 5012 20812 5024
rect 18708 4984 20812 5012
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21358 5012 21364 5024
rect 20956 4984 21364 5012
rect 20956 4972 20962 4984
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 21542 4972 21548 5024
rect 21600 5012 21606 5024
rect 23382 5012 23388 5024
rect 21600 4984 23388 5012
rect 21600 4972 21606 4984
rect 23382 4972 23388 4984
rect 23440 4972 23446 5024
rect 25498 4972 25504 5024
rect 25556 5012 25562 5024
rect 27706 5012 27712 5024
rect 25556 4984 27712 5012
rect 25556 4972 25562 4984
rect 27706 4972 27712 4984
rect 27764 4972 27770 5024
rect 33689 5015 33747 5021
rect 33689 4981 33701 5015
rect 33735 5012 33747 5015
rect 33888 5012 33916 5052
rect 38286 5040 38292 5052
rect 38344 5040 38350 5092
rect 33735 4984 33916 5012
rect 33735 4981 33747 4984
rect 33689 4975 33747 4981
rect 33962 4972 33968 5024
rect 34020 5012 34026 5024
rect 37458 5012 37464 5024
rect 34020 4984 37464 5012
rect 34020 4972 34026 4984
rect 37458 4972 37464 4984
rect 37516 4972 37522 5024
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 10137 4811 10195 4817
rect 7248 4780 8524 4808
rect 7248 4768 7254 4780
rect 8386 4700 8392 4752
rect 8444 4700 8450 4752
rect 8496 4740 8524 4780
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10318 4808 10324 4820
rect 10183 4780 10324 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 16117 4811 16175 4817
rect 10468 4780 15976 4808
rect 10468 4768 10474 4780
rect 8496 4712 13492 4740
rect 5074 4632 5080 4684
rect 5132 4632 5138 4684
rect 5258 4632 5264 4684
rect 5316 4632 5322 4684
rect 5718 4632 5724 4684
rect 5776 4632 5782 4684
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6273 4675 6331 4681
rect 6273 4672 6285 4675
rect 5868 4644 6285 4672
rect 5868 4632 5874 4644
rect 6273 4641 6285 4644
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6963 4644 7389 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 7466 4632 7472 4684
rect 7524 4632 7530 4684
rect 8294 4632 8300 4684
rect 8352 4632 8358 4684
rect 8404 4672 8432 4700
rect 8404 4644 8616 4672
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6086 4564 6092 4616
rect 6144 4613 6150 4616
rect 6144 4607 6172 4613
rect 6160 4573 6172 4607
rect 6144 4567 6172 4573
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 8108 4607 8166 4613
rect 8108 4573 8120 4607
rect 8154 4604 8166 4607
rect 8312 4604 8340 4632
rect 8478 4604 8484 4616
rect 8154 4576 8340 4604
rect 8439 4576 8484 4604
rect 8154 4573 8166 4576
rect 8108 4567 8166 4573
rect 6144 4564 6150 4567
rect 382 4496 388 4548
rect 440 4536 446 4548
rect 3329 4539 3387 4545
rect 3329 4536 3341 4539
rect 440 4508 3341 4536
rect 440 4496 446 4508
rect 3329 4505 3341 4508
rect 3375 4505 3387 4539
rect 3329 4499 3387 4505
rect 3510 4496 3516 4548
rect 3568 4496 3574 4548
rect 4522 4428 4528 4480
rect 4580 4468 4586 4480
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 4580 4440 7021 4468
rect 4580 4428 4586 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7208 4468 7236 4567
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 8588 4613 8616 4644
rect 8754 4632 8760 4684
rect 8812 4672 8818 4684
rect 9769 4675 9827 4681
rect 9769 4672 9781 4675
rect 8812 4644 9781 4672
rect 8812 4632 8818 4644
rect 9769 4641 9781 4644
rect 9815 4641 9827 4675
rect 9769 4635 9827 4641
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 10689 4675 10747 4681
rect 10689 4672 10701 4675
rect 10652 4644 10701 4672
rect 10652 4632 10658 4644
rect 10689 4641 10701 4644
rect 10735 4641 10747 4675
rect 10689 4635 10747 4641
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 9677 4607 9735 4613
rect 9677 4573 9689 4607
rect 9723 4604 9735 4607
rect 9723 4576 10640 4604
rect 9723 4573 9735 4576
rect 9677 4567 9735 4573
rect 10612 4548 10640 4576
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 10928 4576 12204 4604
rect 10928 4564 10934 4576
rect 8202 4496 8208 4548
rect 8260 4496 8266 4548
rect 8297 4539 8355 4545
rect 8297 4505 8309 4539
rect 8343 4505 8355 4539
rect 8297 4499 8355 4505
rect 9585 4539 9643 4545
rect 9585 4505 9597 4539
rect 9631 4536 9643 4539
rect 9631 4508 10548 4536
rect 9631 4505 9643 4508
rect 9585 4499 9643 4505
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 7208 4440 7941 4468
rect 7009 4431 7067 4437
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 8312 4468 8340 4499
rect 10520 4480 10548 4508
rect 10594 4496 10600 4548
rect 10652 4536 10658 4548
rect 10962 4536 10968 4548
rect 10652 4508 10968 4536
rect 10652 4496 10658 4508
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 8312 4440 9229 4468
rect 7929 4431 7987 4437
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 9217 4431 9275 4437
rect 10502 4428 10508 4480
rect 10560 4428 10566 4480
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 12069 4471 12127 4477
rect 12069 4468 12081 4471
rect 12032 4440 12081 4468
rect 12032 4428 12038 4440
rect 12069 4437 12081 4440
rect 12115 4437 12127 4471
rect 12176 4468 12204 4576
rect 12250 4564 12256 4616
rect 12308 4564 12314 4616
rect 13464 4613 13492 4712
rect 13630 4700 13636 4752
rect 13688 4700 13694 4752
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13872 4644 14105 4672
rect 13872 4632 13878 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 13449 4607 13507 4613
rect 13449 4573 13461 4607
rect 13495 4604 13507 4607
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 13495 4576 14381 4604
rect 13495 4573 13507 4576
rect 13449 4567 13507 4573
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 14734 4604 14740 4616
rect 14516 4576 14740 4604
rect 14516 4564 14522 4576
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15378 4564 15384 4616
rect 15436 4564 15442 4616
rect 15948 4613 15976 4780
rect 16117 4777 16129 4811
rect 16163 4808 16175 4811
rect 17954 4808 17960 4820
rect 16163 4780 17960 4808
rect 16163 4777 16175 4780
rect 16117 4771 16175 4777
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 19058 4768 19064 4820
rect 19116 4768 19122 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 19392 4780 20637 4808
rect 19392 4768 19398 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 20898 4768 20904 4820
rect 20956 4768 20962 4820
rect 21100 4780 22324 4808
rect 17221 4743 17279 4749
rect 17221 4709 17233 4743
rect 17267 4709 17279 4743
rect 17221 4703 17279 4709
rect 17236 4672 17264 4703
rect 18049 4675 18107 4681
rect 18049 4672 18061 4675
rect 17236 4644 18061 4672
rect 18049 4641 18061 4644
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 16390 4604 16396 4616
rect 16255 4576 16396 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 15948 4536 15976 4567
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4604 17923 4607
rect 18138 4604 18144 4616
rect 17911 4576 18144 4604
rect 17911 4573 17923 4576
rect 17865 4567 17923 4573
rect 16500 4536 16528 4567
rect 18138 4564 18144 4576
rect 18196 4604 18202 4616
rect 18782 4604 18788 4616
rect 18196 4576 18788 4604
rect 18196 4564 18202 4576
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 18874 4564 18880 4616
rect 18932 4564 18938 4616
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4604 19303 4607
rect 19426 4604 19432 4616
rect 19291 4576 19432 4604
rect 19291 4573 19303 4576
rect 19245 4567 19303 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 21100 4613 21128 4780
rect 22002 4681 22008 4684
rect 21959 4675 22008 4681
rect 21959 4672 21971 4675
rect 21284 4644 21971 4672
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 20809 4607 20867 4613
rect 20809 4573 20821 4607
rect 20855 4573 20867 4607
rect 20809 4567 20867 4573
rect 21085 4607 21143 4613
rect 21085 4573 21097 4607
rect 21131 4573 21143 4607
rect 21085 4567 21143 4573
rect 13556 4508 15240 4536
rect 15948 4508 16528 4536
rect 13556 4468 13584 4508
rect 12176 4440 13584 4468
rect 12069 4431 12127 4437
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 15212 4477 15240 4508
rect 17402 4496 17408 4548
rect 17460 4536 17466 4548
rect 17957 4539 18015 4545
rect 17957 4536 17969 4539
rect 17460 4508 17969 4536
rect 17460 4496 17466 4508
rect 17957 4505 17969 4508
rect 18003 4505 18015 4539
rect 18892 4536 18920 4564
rect 19536 4536 19564 4567
rect 18892 4508 19564 4536
rect 20824 4536 20852 4567
rect 21284 4536 21312 4644
rect 21959 4641 21971 4644
rect 22005 4641 22008 4675
rect 21959 4635 22008 4641
rect 22002 4632 22008 4635
rect 22060 4632 22066 4684
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4672 22155 4675
rect 22296 4672 22324 4780
rect 23106 4768 23112 4820
rect 23164 4768 23170 4820
rect 23382 4768 23388 4820
rect 23440 4768 23446 4820
rect 24854 4768 24860 4820
rect 24912 4768 24918 4820
rect 27522 4768 27528 4820
rect 27580 4808 27586 4820
rect 27580 4780 29132 4808
rect 27580 4768 27586 4780
rect 22373 4743 22431 4749
rect 22373 4709 22385 4743
rect 22419 4740 22431 4743
rect 23290 4740 23296 4752
rect 22419 4712 23296 4740
rect 22419 4709 22431 4712
rect 22373 4703 22431 4709
rect 23290 4700 23296 4712
rect 23348 4700 23354 4752
rect 26053 4743 26111 4749
rect 26053 4709 26065 4743
rect 26099 4709 26111 4743
rect 26053 4703 26111 4709
rect 22646 4672 22652 4684
rect 22143 4644 22652 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 22646 4632 22652 4644
rect 22704 4632 22710 4684
rect 22833 4675 22891 4681
rect 22833 4641 22845 4675
rect 22879 4672 22891 4675
rect 22879 4644 23612 4672
rect 22879 4641 22891 4644
rect 22833 4635 22891 4641
rect 23584 4616 23612 4644
rect 25038 4632 25044 4684
rect 25096 4632 25102 4684
rect 26068 4672 26096 4703
rect 26602 4700 26608 4752
rect 26660 4740 26666 4752
rect 28169 4743 28227 4749
rect 28169 4740 28181 4743
rect 26660 4712 28181 4740
rect 26660 4700 26666 4712
rect 28169 4709 28181 4712
rect 28215 4709 28227 4743
rect 28169 4703 28227 4709
rect 27338 4672 27344 4684
rect 26068 4644 27344 4672
rect 27338 4632 27344 4644
rect 27396 4672 27402 4684
rect 28721 4675 28779 4681
rect 28721 4672 28733 4675
rect 27396 4644 28733 4672
rect 27396 4632 27402 4644
rect 28721 4641 28733 4644
rect 28767 4641 28779 4675
rect 29104 4672 29132 4780
rect 29362 4768 29368 4820
rect 29420 4768 29426 4820
rect 29914 4768 29920 4820
rect 29972 4768 29978 4820
rect 33781 4811 33839 4817
rect 33781 4777 33793 4811
rect 33827 4808 33839 4811
rect 33962 4808 33968 4820
rect 33827 4780 33968 4808
rect 33827 4777 33839 4780
rect 33781 4771 33839 4777
rect 33962 4768 33968 4780
rect 34020 4768 34026 4820
rect 34974 4768 34980 4820
rect 35032 4768 35038 4820
rect 35158 4768 35164 4820
rect 35216 4808 35222 4820
rect 35713 4811 35771 4817
rect 35713 4808 35725 4811
rect 35216 4780 35725 4808
rect 35216 4768 35222 4780
rect 35713 4777 35725 4780
rect 35759 4777 35771 4811
rect 35713 4771 35771 4777
rect 37090 4768 37096 4820
rect 37148 4768 37154 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 38105 4811 38163 4817
rect 38105 4808 38117 4811
rect 37884 4780 38117 4808
rect 37884 4768 37890 4780
rect 38105 4777 38117 4780
rect 38151 4777 38163 4811
rect 38105 4771 38163 4777
rect 39390 4768 39396 4820
rect 39448 4768 39454 4820
rect 31386 4700 31392 4752
rect 31444 4740 31450 4752
rect 31444 4712 38332 4740
rect 31444 4700 31450 4712
rect 29104 4644 29776 4672
rect 28721 4635 28779 4641
rect 21818 4564 21824 4616
rect 21876 4564 21882 4616
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4604 23075 4607
rect 23293 4607 23351 4613
rect 23293 4604 23305 4607
rect 23063 4576 23305 4604
rect 23063 4573 23075 4576
rect 23017 4567 23075 4573
rect 23293 4573 23305 4576
rect 23339 4573 23351 4607
rect 23293 4567 23351 4573
rect 20824 4508 21312 4536
rect 23308 4536 23336 4567
rect 23566 4564 23572 4616
rect 23624 4564 23630 4616
rect 24949 4607 25007 4613
rect 24949 4573 24961 4607
rect 24995 4604 25007 4607
rect 25222 4604 25228 4616
rect 24995 4576 25228 4604
rect 24995 4573 25007 4576
rect 24949 4567 25007 4573
rect 25222 4564 25228 4576
rect 25280 4604 25286 4616
rect 25317 4607 25375 4613
rect 25317 4604 25329 4607
rect 25280 4576 25329 4604
rect 25280 4564 25286 4576
rect 25317 4573 25329 4576
rect 25363 4573 25375 4607
rect 25317 4567 25375 4573
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 27522 4604 27528 4616
rect 26384 4576 27528 4604
rect 26384 4564 26390 4576
rect 27522 4564 27528 4576
rect 27580 4564 27586 4616
rect 27709 4607 27767 4613
rect 27709 4573 27721 4607
rect 27755 4573 27767 4607
rect 27709 4567 27767 4573
rect 24854 4536 24860 4548
rect 23308 4508 24860 4536
rect 17957 4499 18015 4505
rect 24854 4496 24860 4508
rect 24912 4496 24918 4548
rect 26786 4496 26792 4548
rect 26844 4536 26850 4548
rect 27430 4536 27436 4548
rect 26844 4508 27436 4536
rect 26844 4496 26850 4508
rect 27430 4496 27436 4508
rect 27488 4536 27494 4548
rect 27724 4536 27752 4567
rect 28442 4564 28448 4616
rect 28500 4564 28506 4616
rect 28626 4613 28632 4616
rect 28583 4607 28632 4613
rect 28583 4573 28595 4607
rect 28629 4573 28632 4607
rect 28583 4567 28632 4573
rect 28626 4564 28632 4567
rect 28684 4564 28690 4616
rect 29748 4613 29776 4644
rect 32582 4632 32588 4684
rect 32640 4672 32646 4684
rect 32640 4644 36952 4672
rect 32640 4632 32646 4644
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 30098 4564 30104 4616
rect 30156 4564 30162 4616
rect 33597 4607 33655 4613
rect 33597 4573 33609 4607
rect 33643 4573 33655 4607
rect 33597 4567 33655 4573
rect 34885 4607 34943 4613
rect 34885 4573 34897 4607
rect 34931 4604 34943 4607
rect 35161 4607 35219 4613
rect 35161 4604 35173 4607
rect 34931 4576 35173 4604
rect 34931 4573 34943 4576
rect 34885 4567 34943 4573
rect 35161 4573 35173 4576
rect 35207 4573 35219 4607
rect 35161 4567 35219 4573
rect 35897 4607 35955 4613
rect 35897 4573 35909 4607
rect 35943 4604 35955 4607
rect 35986 4604 35992 4616
rect 35943 4576 35992 4604
rect 35943 4573 35955 4576
rect 35897 4567 35955 4573
rect 27488 4508 27752 4536
rect 33612 4536 33640 4567
rect 35986 4564 35992 4576
rect 36044 4564 36050 4616
rect 36924 4613 36952 4644
rect 38304 4613 38332 4712
rect 36909 4607 36967 4613
rect 36909 4573 36921 4607
rect 36955 4573 36967 4607
rect 36909 4567 36967 4573
rect 38289 4607 38347 4613
rect 38289 4573 38301 4607
rect 38335 4573 38347 4607
rect 38289 4567 38347 4573
rect 38562 4564 38568 4616
rect 38620 4564 38626 4616
rect 38746 4564 38752 4616
rect 38804 4604 38810 4616
rect 39209 4607 39267 4613
rect 39209 4604 39221 4607
rect 38804 4576 39221 4604
rect 38804 4564 38810 4576
rect 39209 4573 39221 4576
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 36262 4536 36268 4548
rect 33612 4508 36268 4536
rect 27488 4496 27494 4508
rect 36262 4496 36268 4508
rect 36320 4496 36326 4548
rect 38470 4496 38476 4548
rect 38528 4536 38534 4548
rect 38657 4539 38715 4545
rect 38657 4536 38669 4539
rect 38528 4508 38669 4536
rect 38528 4496 38534 4508
rect 38657 4505 38669 4508
rect 38703 4505 38715 4539
rect 38657 4499 38715 4505
rect 38841 4539 38899 4545
rect 38841 4505 38853 4539
rect 38887 4536 38899 4539
rect 38930 4536 38936 4548
rect 38887 4508 38936 4536
rect 38887 4505 38899 4508
rect 38841 4499 38899 4505
rect 38930 4496 38936 4508
rect 38988 4496 38994 4548
rect 15105 4471 15163 4477
rect 15105 4468 15117 4471
rect 14516 4440 15117 4468
rect 14516 4428 14522 4440
rect 15105 4437 15117 4440
rect 15151 4437 15163 4471
rect 15105 4431 15163 4437
rect 15197 4471 15255 4477
rect 15197 4437 15209 4471
rect 15243 4437 15255 4471
rect 15197 4431 15255 4437
rect 17494 4428 17500 4480
rect 17552 4428 17558 4480
rect 20254 4428 20260 4480
rect 20312 4428 20318 4480
rect 21177 4471 21235 4477
rect 21177 4437 21189 4471
rect 21223 4468 21235 4471
rect 21542 4468 21548 4480
rect 21223 4440 21548 4468
rect 21223 4437 21235 4440
rect 21177 4431 21235 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 21726 4428 21732 4480
rect 21784 4468 21790 4480
rect 25314 4468 25320 4480
rect 21784 4440 25320 4468
rect 21784 4428 21790 4440
rect 25314 4428 25320 4440
rect 25372 4428 25378 4480
rect 27614 4428 27620 4480
rect 27672 4468 27678 4480
rect 28626 4468 28632 4480
rect 27672 4440 28632 4468
rect 27672 4428 27678 4440
rect 28626 4428 28632 4440
rect 28684 4428 28690 4480
rect 28718 4428 28724 4480
rect 28776 4468 28782 4480
rect 29549 4471 29607 4477
rect 29549 4468 29561 4471
rect 28776 4440 29561 4468
rect 28776 4428 28782 4440
rect 29549 4437 29561 4440
rect 29595 4437 29607 4471
rect 29549 4431 29607 4437
rect 34790 4428 34796 4480
rect 34848 4428 34854 4480
rect 36446 4428 36452 4480
rect 36504 4468 36510 4480
rect 38381 4471 38439 4477
rect 38381 4468 38393 4471
rect 36504 4440 38393 4468
rect 36504 4428 36510 4440
rect 38381 4437 38393 4440
rect 38427 4437 38439 4471
rect 38381 4431 38439 4437
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 5776 4236 6193 4264
rect 5776 4224 5782 4236
rect 6181 4233 6193 4236
rect 6227 4233 6239 4267
rect 6181 4227 6239 4233
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8202 4264 8208 4276
rect 8159 4236 8208 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 1210 4156 1216 4208
rect 1268 4196 1274 4208
rect 3605 4199 3663 4205
rect 3605 4196 3617 4199
rect 1268 4168 3617 4196
rect 1268 4156 1274 4168
rect 3605 4165 3617 4168
rect 3651 4165 3663 4199
rect 3605 4159 3663 4165
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 6196 4128 6224 4227
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 10870 4264 10876 4276
rect 8352 4236 10876 4264
rect 8352 4224 8358 4236
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11514 4224 11520 4276
rect 11572 4264 11578 4276
rect 14642 4264 14648 4276
rect 11572 4236 14648 4264
rect 11572 4224 11578 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 19426 4264 19432 4276
rect 17276 4236 19432 4264
rect 17276 4224 17282 4236
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 20254 4224 20260 4276
rect 20312 4264 20318 4276
rect 21910 4264 21916 4276
rect 20312 4236 21916 4264
rect 20312 4224 20318 4236
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 24486 4224 24492 4276
rect 24544 4264 24550 4276
rect 27157 4267 27215 4273
rect 27157 4264 27169 4267
rect 24544 4236 27169 4264
rect 24544 4224 24550 4236
rect 27157 4233 27169 4236
rect 27203 4233 27215 4267
rect 27157 4227 27215 4233
rect 27430 4224 27436 4276
rect 27488 4264 27494 4276
rect 30098 4264 30104 4276
rect 27488 4236 30104 4264
rect 27488 4224 27494 4236
rect 30098 4224 30104 4236
rect 30156 4224 30162 4276
rect 8754 4196 8760 4208
rect 8404 4168 8760 4196
rect 8404 4158 8432 4168
rect 8342 4131 8432 4158
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 10502 4156 10508 4208
rect 10560 4196 10566 4208
rect 22370 4196 22376 4208
rect 10560 4168 22376 4196
rect 10560 4156 10566 4168
rect 8342 4128 8355 4131
rect 6196 4100 8355 4128
rect 8343 4097 8355 4100
rect 8389 4130 8432 4131
rect 8481 4131 8539 4137
rect 8389 4097 8401 4130
rect 8343 4091 8401 4097
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 10226 4128 10232 4140
rect 8527 4100 10232 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10594 4128 10600 4140
rect 10459 4100 10600 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10704 4137 10732 4168
rect 22370 4156 22376 4168
rect 22428 4156 22434 4208
rect 25682 4156 25688 4208
rect 25740 4196 25746 4208
rect 37461 4199 37519 4205
rect 37461 4196 37473 4199
rect 25740 4168 37473 4196
rect 25740 4156 25746 4168
rect 37461 4165 37473 4168
rect 37507 4165 37519 4199
rect 37461 4159 37519 4165
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14424 4100 14565 4128
rect 14424 4088 14430 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 17218 4128 17224 4140
rect 16899 4100 17224 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17552 4100 17877 4128
rect 17552 4088 17558 4100
rect 17865 4097 17877 4100
rect 17911 4097 17923 4131
rect 17865 4091 17923 4097
rect 25222 4088 25228 4140
rect 25280 4088 25286 4140
rect 27341 4131 27399 4137
rect 27341 4097 27353 4131
rect 27387 4128 27399 4131
rect 27614 4128 27620 4140
rect 27387 4100 27620 4128
rect 27387 4097 27399 4100
rect 27341 4091 27399 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 27893 4131 27951 4137
rect 27893 4097 27905 4131
rect 27939 4128 27951 4131
rect 28442 4128 28448 4140
rect 27939 4100 28448 4128
rect 27939 4097 27951 4100
rect 27893 4091 27951 4097
rect 28442 4088 28448 4100
rect 28500 4088 28506 4140
rect 29086 4088 29092 4140
rect 29144 4128 29150 4140
rect 30282 4128 30288 4140
rect 29144 4100 30288 4128
rect 29144 4088 29150 4100
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 32467 4131 32525 4137
rect 32467 4128 32479 4131
rect 31726 4100 32479 4128
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 3786 3952 3792 4004
rect 3844 3952 3850 4004
rect 5184 3924 5212 4023
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 7340 4032 12434 4060
rect 7340 4020 7346 4032
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10505 3995 10563 4001
rect 10505 3992 10517 3995
rect 10100 3964 10517 3992
rect 10100 3952 10106 3964
rect 10505 3961 10517 3964
rect 10551 3961 10563 3995
rect 10505 3955 10563 3961
rect 5902 3924 5908 3936
rect 5184 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 10008 3896 10241 3924
rect 10008 3884 10014 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 12406 3924 12434 4032
rect 14458 4020 14464 4072
rect 14516 4020 14522 4072
rect 14734 4020 14740 4072
rect 14792 4060 14798 4072
rect 14792 4032 16896 4060
rect 14792 4020 14798 4032
rect 15013 3995 15071 4001
rect 15013 3961 15025 3995
rect 15059 3992 15071 3995
rect 15378 3992 15384 4004
rect 15059 3964 15384 3992
rect 15059 3961 15071 3964
rect 15013 3955 15071 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 16868 3992 16896 4032
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 26878 4060 26884 4072
rect 17000 4032 26884 4060
rect 17000 4020 17006 4032
rect 26878 4020 26884 4032
rect 26936 4020 26942 4072
rect 28258 4020 28264 4072
rect 28316 4060 28322 4072
rect 31726 4060 31754 4100
rect 32467 4097 32479 4100
rect 32513 4097 32525 4131
rect 32467 4091 32525 4097
rect 38473 4131 38531 4137
rect 38473 4097 38485 4131
rect 38519 4097 38531 4131
rect 38473 4091 38531 4097
rect 28316 4032 31754 4060
rect 28316 4020 28322 4032
rect 37274 4020 37280 4072
rect 37332 4020 37338 4072
rect 21358 3992 21364 4004
rect 16868 3964 21364 3992
rect 21358 3952 21364 3964
rect 21416 3952 21422 4004
rect 21542 3952 21548 4004
rect 21600 3992 21606 4004
rect 22922 3992 22928 4004
rect 21600 3964 22928 3992
rect 21600 3952 21606 3964
rect 22922 3952 22928 3964
rect 22980 3952 22986 4004
rect 25409 3995 25467 4001
rect 25409 3961 25421 3995
rect 25455 3992 25467 3995
rect 25455 3964 27660 3992
rect 25455 3961 25467 3964
rect 25409 3955 25467 3961
rect 16574 3924 16580 3936
rect 12406 3896 16580 3924
rect 10229 3887 10287 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 17678 3884 17684 3936
rect 17736 3884 17742 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 23474 3924 23480 3936
rect 19208 3896 23480 3924
rect 19208 3884 19214 3896
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 27632 3924 27660 3964
rect 27706 3952 27712 4004
rect 27764 3952 27770 4004
rect 38488 3992 38516 4091
rect 38838 4088 38844 4140
rect 38896 4088 38902 4140
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4128 39267 4131
rect 39482 4128 39488 4140
rect 39255 4100 39488 4128
rect 39255 4097 39267 4100
rect 39209 4091 39267 4097
rect 39482 4088 39488 4100
rect 39540 4088 39546 4140
rect 31864 3964 38516 3992
rect 28994 3924 29000 3936
rect 27632 3896 29000 3924
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 30466 3884 30472 3936
rect 30524 3924 30530 3936
rect 31864 3924 31892 3964
rect 39022 3952 39028 4004
rect 39080 3952 39086 4004
rect 39390 3952 39396 4004
rect 39448 3952 39454 4004
rect 30524 3896 31892 3924
rect 30524 3884 30530 3896
rect 32306 3884 32312 3936
rect 32364 3884 32370 3936
rect 38654 3884 38660 3936
rect 38712 3884 38718 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 16080 3692 26740 3720
rect 16080 3680 16086 3692
rect 4430 3612 4436 3664
rect 4488 3652 4494 3664
rect 17678 3652 17684 3664
rect 4488 3624 17684 3652
rect 4488 3612 4494 3624
rect 17678 3612 17684 3624
rect 17736 3612 17742 3664
rect 26602 3652 26608 3664
rect 18800 3624 26608 3652
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5500 3488 5641 3516
rect 5500 3476 5506 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 11974 3476 11980 3528
rect 12032 3476 12038 3528
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 15528 3488 18092 3516
rect 15528 3476 15534 3488
rect 5810 3408 5816 3460
rect 5868 3408 5874 3460
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6822 3448 6828 3460
rect 5960 3420 6828 3448
rect 5960 3408 5966 3420
rect 6822 3408 6828 3420
rect 6880 3448 6886 3460
rect 16666 3448 16672 3460
rect 6880 3420 16672 3448
rect 6880 3408 6886 3420
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 18064 3448 18092 3488
rect 18800 3448 18828 3624
rect 26602 3612 26608 3624
rect 26660 3612 26666 3664
rect 26712 3652 26740 3692
rect 26970 3680 26976 3732
rect 27028 3720 27034 3732
rect 32398 3720 32404 3732
rect 27028 3692 32404 3720
rect 27028 3680 27034 3692
rect 32398 3680 32404 3692
rect 32456 3680 32462 3732
rect 39393 3723 39451 3729
rect 39393 3689 39405 3723
rect 39439 3720 39451 3723
rect 39574 3720 39580 3732
rect 39439 3692 39580 3720
rect 39439 3689 39451 3692
rect 39393 3683 39451 3689
rect 39574 3680 39580 3692
rect 39632 3680 39638 3732
rect 27062 3652 27068 3664
rect 26712 3624 27068 3652
rect 27062 3612 27068 3624
rect 27120 3612 27126 3664
rect 30374 3612 30380 3664
rect 30432 3652 30438 3664
rect 38930 3652 38936 3664
rect 30432 3624 38936 3652
rect 30432 3612 30438 3624
rect 38930 3612 38936 3624
rect 38988 3612 38994 3664
rect 39025 3655 39083 3661
rect 39025 3621 39037 3655
rect 39071 3652 39083 3655
rect 39942 3652 39948 3664
rect 39071 3624 39948 3652
rect 39071 3621 39083 3624
rect 39025 3615 39083 3621
rect 39942 3612 39948 3624
rect 40000 3612 40006 3664
rect 20438 3584 20444 3596
rect 19812 3556 20444 3584
rect 18874 3476 18880 3528
rect 18932 3516 18938 3528
rect 19812 3525 19840 3556
rect 20438 3544 20444 3556
rect 20496 3544 20502 3596
rect 21358 3544 21364 3596
rect 21416 3584 21422 3596
rect 30282 3584 30288 3596
rect 21416 3556 27016 3584
rect 21416 3544 21422 3556
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 18932 3488 19625 3516
rect 18932 3476 18938 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20346 3516 20352 3528
rect 20119 3488 20352 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 22370 3476 22376 3528
rect 22428 3516 22434 3528
rect 26510 3516 26516 3528
rect 22428 3488 26516 3516
rect 22428 3476 22434 3488
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 26988 3516 27016 3556
rect 29104 3556 30288 3584
rect 29104 3516 29132 3556
rect 30282 3544 30288 3556
rect 30340 3544 30346 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 36538 3584 36544 3596
rect 33928 3556 36544 3584
rect 33928 3544 33934 3556
rect 36538 3544 36544 3556
rect 36596 3544 36602 3596
rect 26988 3488 29132 3516
rect 29178 3476 29184 3528
rect 29236 3516 29242 3528
rect 36814 3516 36820 3528
rect 29236 3488 36820 3516
rect 29236 3476 29242 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 38746 3476 38752 3528
rect 38804 3516 38810 3528
rect 38841 3519 38899 3525
rect 38841 3516 38853 3519
rect 38804 3488 38853 3516
rect 38804 3476 38810 3488
rect 38841 3485 38853 3488
rect 38887 3485 38899 3519
rect 38841 3479 38899 3485
rect 39209 3519 39267 3525
rect 39209 3485 39221 3519
rect 39255 3516 39267 3519
rect 39758 3516 39764 3528
rect 39255 3488 39764 3516
rect 39255 3485 39267 3488
rect 39209 3479 39267 3485
rect 39758 3476 39764 3488
rect 39816 3476 39822 3528
rect 18064 3420 18828 3448
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 19392 3420 26740 3448
rect 19392 3408 19398 3420
rect 12158 3340 12164 3392
rect 12216 3340 12222 3392
rect 14274 3340 14280 3392
rect 14332 3380 14338 3392
rect 20162 3380 20168 3392
rect 14332 3352 20168 3380
rect 14332 3340 14338 3352
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 20257 3383 20315 3389
rect 20257 3349 20269 3383
rect 20303 3380 20315 3383
rect 22186 3380 22192 3392
rect 20303 3352 22192 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 22186 3340 22192 3352
rect 22244 3340 22250 3392
rect 23290 3340 23296 3392
rect 23348 3380 23354 3392
rect 24670 3380 24676 3392
rect 23348 3352 24676 3380
rect 23348 3340 23354 3352
rect 24670 3340 24676 3352
rect 24728 3340 24734 3392
rect 26712 3380 26740 3420
rect 27062 3408 27068 3460
rect 27120 3448 27126 3460
rect 34606 3448 34612 3460
rect 27120 3420 34612 3448
rect 27120 3408 27126 3420
rect 34606 3408 34612 3420
rect 34664 3408 34670 3460
rect 26878 3380 26884 3392
rect 26712 3352 26884 3380
rect 26878 3340 26884 3352
rect 26936 3340 26942 3392
rect 27338 3340 27344 3392
rect 27396 3380 27402 3392
rect 29270 3380 29276 3392
rect 27396 3352 29276 3380
rect 27396 3340 27402 3352
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 29454 3340 29460 3392
rect 29512 3380 29518 3392
rect 33870 3380 33876 3392
rect 29512 3352 33876 3380
rect 29512 3340 29518 3352
rect 33870 3340 33876 3352
rect 33928 3340 33934 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 16853 3179 16911 3185
rect 16853 3145 16865 3179
rect 16899 3176 16911 3179
rect 16942 3176 16948 3188
rect 16899 3148 16948 3176
rect 16899 3145 16911 3148
rect 16853 3139 16911 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18279 3148 19288 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 19260 3108 19288 3148
rect 19334 3136 19340 3188
rect 19392 3136 19398 3188
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 22002 3176 22008 3188
rect 20220 3148 22008 3176
rect 20220 3136 20226 3148
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 24121 3179 24179 3185
rect 24121 3176 24133 3179
rect 22112 3148 24133 3176
rect 20438 3108 20444 3120
rect 16632 3080 19196 3108
rect 19260 3080 20444 3108
rect 16632 3068 16638 3080
rect 16666 3000 16672 3052
rect 16724 3000 16730 3052
rect 19168 3049 19196 3080
rect 20438 3068 20444 3080
rect 20496 3068 20502 3120
rect 22112 3117 22140 3148
rect 24121 3145 24133 3148
rect 24167 3145 24179 3179
rect 24121 3139 24179 3145
rect 24581 3179 24639 3185
rect 24581 3145 24593 3179
rect 24627 3176 24639 3179
rect 25225 3179 25283 3185
rect 24627 3148 25176 3176
rect 24627 3145 24639 3148
rect 24581 3139 24639 3145
rect 22097 3111 22155 3117
rect 22097 3077 22109 3111
rect 22143 3077 22155 3111
rect 22097 3071 22155 3077
rect 22209 3111 22267 3117
rect 22209 3077 22221 3111
rect 22255 3108 22267 3111
rect 23109 3111 23167 3117
rect 23109 3108 23121 3111
rect 22255 3080 23121 3108
rect 22255 3077 22267 3080
rect 22209 3071 22267 3077
rect 23109 3077 23121 3080
rect 23155 3077 23167 3111
rect 23109 3071 23167 3077
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 16991 3012 17509 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3040 19211 3043
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19199 3012 19717 3040
rect 19199 3009 19211 3012
rect 19153 3003 19211 3009
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 21453 3043 21511 3049
rect 21453 3040 21465 3043
rect 19705 3003 19763 3009
rect 20456 3012 21465 3040
rect 5350 2932 5356 2984
rect 5408 2972 5414 2984
rect 16960 2972 16988 3003
rect 5408 2944 16988 2972
rect 5408 2932 5414 2944
rect 17218 2932 17224 2984
rect 17276 2932 17282 2984
rect 19426 2932 19432 2984
rect 19484 2932 19490 2984
rect 16666 2864 16672 2916
rect 16724 2904 16730 2916
rect 17236 2904 17264 2932
rect 20456 2913 20484 3012
rect 21453 3009 21465 3012
rect 21499 3040 21511 3043
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21499 3012 21833 3040
rect 21499 3009 21511 3012
rect 21453 3003 21511 3009
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 21910 3000 21916 3052
rect 21968 3000 21974 3052
rect 22286 3043 22344 3049
rect 22286 3009 22298 3043
rect 22332 3009 22344 3043
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22286 3003 22344 3009
rect 22480 3012 22753 3040
rect 22186 2932 22192 2984
rect 22244 2972 22250 2984
rect 22301 2972 22329 3003
rect 22480 2972 22508 3012
rect 22741 3009 22753 3012
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 22922 3000 22928 3052
rect 22980 3000 22986 3052
rect 23290 3000 23296 3052
rect 23348 3049 23354 3052
rect 23348 3043 23381 3049
rect 23369 3009 23381 3043
rect 23348 3003 23381 3009
rect 23348 3000 23354 3003
rect 23474 3000 23480 3052
rect 23532 3040 23538 3052
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23532 3012 23765 3040
rect 23532 3000 23538 3012
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 24026 3000 24032 3052
rect 24084 3040 24090 3052
rect 25148 3049 25176 3148
rect 25225 3145 25237 3179
rect 25271 3176 25283 3179
rect 25314 3176 25320 3188
rect 25271 3148 25320 3176
rect 25271 3145 25283 3148
rect 25225 3139 25283 3145
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 25866 3136 25872 3188
rect 25924 3176 25930 3188
rect 26605 3179 26663 3185
rect 26605 3176 26617 3179
rect 25924 3148 26617 3176
rect 25924 3136 25930 3148
rect 26605 3145 26617 3148
rect 26651 3145 26663 3179
rect 26605 3139 26663 3145
rect 26694 3136 26700 3188
rect 26752 3176 26758 3188
rect 27893 3179 27951 3185
rect 27893 3176 27905 3179
rect 26752 3148 27905 3176
rect 26752 3136 26758 3148
rect 27893 3145 27905 3148
rect 27939 3145 27951 3179
rect 29086 3176 29092 3188
rect 27893 3139 27951 3145
rect 28092 3148 29092 3176
rect 26510 3068 26516 3120
rect 26568 3108 26574 3120
rect 27338 3108 27344 3120
rect 26568 3080 27344 3108
rect 26568 3068 26574 3080
rect 27338 3068 27344 3080
rect 27396 3068 27402 3120
rect 24489 3043 24547 3049
rect 24489 3040 24501 3043
rect 24084 3012 24501 3040
rect 24084 3000 24090 3012
rect 24489 3009 24501 3012
rect 24535 3040 24547 3043
rect 25133 3043 25191 3049
rect 24535 3012 25084 3040
rect 24535 3009 24547 3012
rect 24489 3003 24547 3009
rect 22244 2944 22329 2972
rect 22388 2944 22508 2972
rect 22244 2932 22250 2944
rect 20441 2907 20499 2913
rect 16724 2876 17264 2904
rect 18156 2876 19564 2904
rect 16724 2864 16730 2876
rect 17129 2839 17187 2845
rect 17129 2805 17141 2839
rect 17175 2836 17187 2839
rect 18156 2836 18184 2876
rect 17175 2808 18184 2836
rect 19536 2836 19564 2876
rect 20441 2873 20453 2907
rect 20487 2873 20499 2907
rect 20441 2867 20499 2873
rect 21545 2907 21603 2913
rect 21545 2873 21557 2907
rect 21591 2904 21603 2907
rect 22278 2904 22284 2916
rect 21591 2876 22284 2904
rect 21591 2873 21603 2876
rect 21545 2867 21603 2873
rect 22278 2864 22284 2876
rect 22336 2864 22342 2916
rect 22388 2904 22416 2944
rect 22554 2932 22560 2984
rect 22612 2972 22618 2984
rect 23017 2975 23075 2981
rect 23017 2972 23029 2975
rect 22612 2944 23029 2972
rect 22612 2932 22618 2944
rect 23017 2941 23029 2944
rect 23063 2941 23075 2975
rect 23017 2935 23075 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 23624 2944 24593 2972
rect 23624 2932 23630 2944
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 24670 2932 24676 2984
rect 24728 2932 24734 2984
rect 25056 2972 25084 3012
rect 25133 3009 25145 3043
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 25409 3043 25467 3049
rect 25409 3009 25421 3043
rect 25455 3009 25467 3043
rect 25409 3003 25467 3009
rect 25424 2972 25452 3003
rect 26326 3000 26332 3052
rect 26384 3040 26390 3052
rect 28092 3049 28120 3148
rect 29086 3136 29092 3148
rect 29144 3136 29150 3188
rect 29178 3136 29184 3188
rect 29236 3136 29242 3188
rect 29454 3136 29460 3188
rect 29512 3136 29518 3188
rect 29733 3179 29791 3185
rect 29733 3145 29745 3179
rect 29779 3176 29791 3179
rect 29822 3176 29828 3188
rect 29779 3148 29828 3176
rect 29779 3145 29791 3148
rect 29733 3139 29791 3145
rect 29822 3136 29828 3148
rect 29880 3136 29886 3188
rect 30282 3136 30288 3188
rect 30340 3176 30346 3188
rect 30377 3179 30435 3185
rect 30377 3176 30389 3179
rect 30340 3148 30389 3176
rect 30340 3136 30346 3148
rect 30377 3145 30389 3148
rect 30423 3145 30435 3179
rect 30377 3139 30435 3145
rect 32401 3179 32459 3185
rect 32401 3145 32413 3179
rect 32447 3176 32459 3179
rect 32490 3176 32496 3188
rect 32447 3148 32496 3176
rect 32447 3145 32459 3148
rect 32401 3139 32459 3145
rect 32490 3136 32496 3148
rect 32548 3136 32554 3188
rect 34606 3136 34612 3188
rect 34664 3136 34670 3188
rect 35894 3136 35900 3188
rect 35952 3176 35958 3188
rect 36357 3179 36415 3185
rect 36357 3176 36369 3179
rect 35952 3148 36369 3176
rect 35952 3136 35958 3148
rect 36357 3145 36369 3148
rect 36403 3145 36415 3179
rect 36357 3139 36415 3145
rect 38197 3179 38255 3185
rect 38197 3145 38209 3179
rect 38243 3145 38255 3179
rect 38197 3139 38255 3145
rect 35158 3108 35164 3120
rect 29012 3080 35164 3108
rect 29012 3049 29040 3080
rect 35158 3068 35164 3080
rect 35216 3068 35222 3120
rect 35342 3068 35348 3120
rect 35400 3108 35406 3120
rect 38212 3108 38240 3139
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 35400 3080 38240 3108
rect 35400 3068 35406 3080
rect 26421 3043 26479 3049
rect 26421 3040 26433 3043
rect 26384 3012 26433 3040
rect 26384 3000 26390 3012
rect 26421 3009 26433 3012
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 28077 3043 28135 3049
rect 28077 3009 28089 3043
rect 28123 3009 28135 3043
rect 28077 3003 28135 3009
rect 28997 3043 29055 3049
rect 28997 3009 29009 3043
rect 29043 3009 29055 3043
rect 28997 3003 29055 3009
rect 29270 3000 29276 3052
rect 29328 3000 29334 3052
rect 29549 3043 29607 3049
rect 29549 3009 29561 3043
rect 29595 3009 29607 3043
rect 29549 3003 29607 3009
rect 25056 2944 25452 2972
rect 27706 2932 27712 2984
rect 27764 2972 27770 2984
rect 29564 2972 29592 3003
rect 30558 3000 30564 3052
rect 30616 3000 30622 3052
rect 31754 3000 31760 3052
rect 31812 3040 31818 3052
rect 32217 3043 32275 3049
rect 32217 3040 32229 3043
rect 31812 3012 32229 3040
rect 31812 3000 31818 3012
rect 32217 3009 32229 3012
rect 32263 3009 32275 3043
rect 32217 3003 32275 3009
rect 34057 3043 34115 3049
rect 34057 3009 34069 3043
rect 34103 3009 34115 3043
rect 34057 3003 34115 3009
rect 27764 2944 29592 2972
rect 27764 2932 27770 2944
rect 31846 2932 31852 2984
rect 31904 2972 31910 2984
rect 34072 2972 34100 3003
rect 34146 3000 34152 3052
rect 34204 3040 34210 3052
rect 34793 3043 34851 3049
rect 34793 3040 34805 3043
rect 34204 3012 34805 3040
rect 34204 3000 34210 3012
rect 34793 3009 34805 3012
rect 34839 3009 34851 3043
rect 34793 3003 34851 3009
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 36311 3012 36553 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 38381 3043 38439 3049
rect 38381 3009 38393 3043
rect 38427 3009 38439 3043
rect 38381 3003 38439 3009
rect 31904 2944 34100 2972
rect 31904 2932 31910 2944
rect 35250 2932 35256 2984
rect 35308 2972 35314 2984
rect 38396 2972 38424 3003
rect 38470 3000 38476 3052
rect 38528 3000 38534 3052
rect 38838 3000 38844 3052
rect 38896 3000 38902 3052
rect 38930 3000 38936 3052
rect 38988 3040 38994 3052
rect 39209 3043 39267 3049
rect 39209 3040 39221 3043
rect 38988 3012 39221 3040
rect 38988 3000 38994 3012
rect 39209 3009 39221 3012
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 35308 2944 38424 2972
rect 35308 2932 35314 2944
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 22388 2876 22477 2904
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 22465 2867 22523 2873
rect 23474 2864 23480 2916
rect 23532 2904 23538 2916
rect 24949 2907 25007 2913
rect 24949 2904 24961 2907
rect 23532 2876 24961 2904
rect 23532 2864 23538 2876
rect 24949 2873 24961 2876
rect 24995 2873 25007 2907
rect 24949 2867 25007 2873
rect 25038 2864 25044 2916
rect 25096 2904 25102 2916
rect 33873 2907 33931 2913
rect 33873 2904 33885 2907
rect 25096 2876 33885 2904
rect 25096 2864 25102 2876
rect 33873 2873 33885 2876
rect 33919 2873 33931 2907
rect 33873 2867 33931 2873
rect 34514 2864 34520 2916
rect 34572 2904 34578 2916
rect 36173 2907 36231 2913
rect 36173 2904 36185 2907
rect 34572 2876 36185 2904
rect 34572 2864 34578 2876
rect 36173 2873 36185 2876
rect 36219 2873 36231 2907
rect 40126 2904 40132 2916
rect 36173 2867 36231 2873
rect 38580 2876 40132 2904
rect 22370 2836 22376 2848
rect 19536 2808 22376 2836
rect 17175 2805 17187 2808
rect 17129 2799 17187 2805
rect 22370 2796 22376 2808
rect 22428 2796 22434 2848
rect 22554 2796 22560 2848
rect 22612 2796 22618 2848
rect 23014 2796 23020 2848
rect 23072 2836 23078 2848
rect 23569 2839 23627 2845
rect 23569 2836 23581 2839
rect 23072 2808 23581 2836
rect 23072 2796 23078 2808
rect 23569 2805 23581 2808
rect 23615 2805 23627 2839
rect 23569 2799 23627 2805
rect 26878 2796 26884 2848
rect 26936 2836 26942 2848
rect 38580 2836 38608 2876
rect 40126 2864 40132 2876
rect 40184 2864 40190 2916
rect 26936 2808 38608 2836
rect 26936 2796 26942 2808
rect 38654 2796 38660 2848
rect 38712 2796 38718 2848
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 22554 2632 22560 2644
rect 4632 2604 22560 2632
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 4522 2428 4528 2440
rect 3191 2400 4528 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 4522 2388 4528 2400
rect 4580 2388 4586 2440
rect 4632 2437 4660 2604
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 39390 2592 39396 2644
rect 39448 2592 39454 2644
rect 7558 2524 7564 2576
rect 7616 2564 7622 2576
rect 23474 2564 23480 2576
rect 7616 2536 23480 2564
rect 7616 2524 7622 2536
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 30742 2524 30748 2576
rect 30800 2564 30806 2576
rect 38562 2564 38568 2576
rect 30800 2536 38568 2564
rect 30800 2524 30806 2536
rect 38562 2524 38568 2536
rect 38620 2524 38626 2576
rect 6362 2456 6368 2508
rect 6420 2496 6426 2508
rect 6420 2468 22094 2496
rect 6420 2456 6426 2468
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9398 2428 9404 2440
rect 9263 2400 9404 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2832 2264 2973 2292
rect 2832 2252 2838 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 4246 2252 4252 2304
rect 4304 2292 4310 2304
rect 4433 2295 4491 2301
rect 4433 2292 4445 2295
rect 4304 2264 4445 2292
rect 4304 2252 4310 2264
rect 4433 2261 4445 2264
rect 4479 2261 4491 2295
rect 4433 2255 4491 2261
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5776 2264 5917 2292
rect 5776 2252 5782 2264
rect 5905 2261 5917 2264
rect 5951 2261 5963 2295
rect 6104 2292 6132 2391
rect 7576 2360 7604 2391
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 22066 2428 22094 2468
rect 36998 2456 37004 2508
rect 37056 2496 37062 2508
rect 39666 2496 39672 2508
rect 37056 2468 38148 2496
rect 37056 2456 37062 2468
rect 38120 2437 38148 2468
rect 38856 2468 39672 2496
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 22066 2400 37749 2428
rect 11701 2391 11759 2397
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38470 2388 38476 2440
rect 38528 2388 38534 2440
rect 38856 2437 38884 2468
rect 39666 2456 39672 2468
rect 39724 2456 39730 2508
rect 38841 2431 38899 2437
rect 38841 2397 38853 2431
rect 38887 2397 38899 2431
rect 38841 2391 38899 2397
rect 39206 2388 39212 2440
rect 39264 2388 39270 2440
rect 21450 2360 21456 2372
rect 7576 2332 21456 2360
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 6178 2292 6184 2304
rect 6104 2264 6184 2292
rect 5905 2255 5963 2261
rect 6178 2252 6184 2264
rect 6236 2252 6242 2304
rect 7190 2252 7196 2304
rect 7248 2292 7254 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7248 2264 7389 2292
rect 7248 2252 7254 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8720 2264 9045 2292
rect 8720 2252 8726 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 11885 2295 11943 2301
rect 11885 2261 11897 2295
rect 11931 2292 11943 2295
rect 23842 2292 23848 2304
rect 11931 2264 23848 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39025 2295 39083 2301
rect 39025 2261 39037 2295
rect 39071 2292 39083 2295
rect 39942 2292 39948 2304
rect 39071 2264 39948 2292
rect 39071 2261 39083 2264
rect 39025 2255 39083 2261
rect 39942 2252 39948 2264
rect 40000 2252 40006 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 2746 2060 6316 2088
rect 1026 1980 1032 2032
rect 1084 2020 1090 2032
rect 2746 2020 2774 2060
rect 1084 1992 2774 2020
rect 1084 1980 1090 1992
rect 6178 1980 6184 2032
rect 6236 1980 6242 2032
rect 6288 2020 6316 2060
rect 11422 2048 11428 2100
rect 11480 2088 11486 2100
rect 32306 2088 32312 2100
rect 11480 2060 32312 2088
rect 11480 2048 11486 2060
rect 32306 2048 32312 2060
rect 32364 2048 32370 2100
rect 30650 2020 30656 2032
rect 6288 1992 30656 2020
rect 30650 1980 30656 1992
rect 30708 1980 30714 2032
rect 6196 1952 6224 1980
rect 27890 1952 27896 1964
rect 6196 1924 27896 1952
rect 27890 1912 27896 1924
rect 27948 1912 27954 1964
rect 1670 1844 1676 1896
rect 1728 1884 1734 1896
rect 14366 1884 14372 1896
rect 1728 1856 14372 1884
rect 1728 1844 1734 1856
rect 14366 1844 14372 1856
rect 14424 1844 14430 1896
rect 3786 1776 3792 1828
rect 3844 1816 3850 1828
rect 38470 1816 38476 1828
rect 3844 1788 38476 1816
rect 3844 1776 3850 1788
rect 38470 1776 38476 1788
rect 38528 1776 38534 1828
rect 23382 824 23388 876
rect 23440 864 23446 876
rect 27706 864 27712 876
rect 23440 836 27712 864
rect 23440 824 23446 836
rect 27706 824 27712 836
rect 27764 824 27770 876
rect 20438 348 20444 400
rect 20496 388 20502 400
rect 35250 388 35256 400
rect 20496 360 35256 388
rect 20496 348 20502 360
rect 35250 348 35256 360
rect 35308 348 35314 400
rect 18966 280 18972 332
rect 19024 320 19030 332
rect 34790 320 34796 332
rect 19024 292 34796 320
rect 19024 280 19030 292
rect 34790 280 34796 292
rect 34848 280 34854 332
rect 16022 212 16028 264
rect 16080 252 16086 264
rect 33410 252 33416 264
rect 16080 224 33416 252
rect 16080 212 16086 224
rect 33410 212 33416 224
rect 33468 212 33474 264
rect 11974 144 11980 196
rect 12032 184 12038 196
rect 33686 184 33692 196
rect 12032 156 33692 184
rect 12032 144 12038 156
rect 33686 144 33692 156
rect 33744 144 33750 196
rect 14642 76 14648 128
rect 14700 116 14706 128
rect 37366 116 37372 128
rect 14700 88 37372 116
rect 14700 76 14706 88
rect 37366 76 37372 88
rect 37424 76 37430 128
rect 10226 8 10232 60
rect 10284 48 10290 60
rect 31754 48 31760 60
rect 10284 20 31760 48
rect 10284 8 10290 20
rect 31754 8 31760 20
rect 31812 8 31818 60
<< via1 >>
rect 1860 11160 1912 11212
rect 25596 11160 25648 11212
rect 26424 10140 26476 10192
rect 32588 10140 32640 10192
rect 24492 10004 24544 10056
rect 25136 10004 25188 10056
rect 17500 9868 17552 9920
rect 20628 9868 20680 9920
rect 2504 9800 2556 9852
rect 24584 9800 24636 9852
rect 10048 9732 10100 9784
rect 37280 9732 37332 9784
rect 9496 9664 9548 9716
rect 37648 9664 37700 9716
rect 5632 9596 5684 9648
rect 16396 9596 16448 9648
rect 23112 9596 23164 9648
rect 23480 9596 23532 9648
rect 18052 9528 18104 9580
rect 24492 9528 24544 9580
rect 5080 9460 5132 9512
rect 11980 9460 12032 9512
rect 4804 9392 4856 9444
rect 15476 9392 15528 9444
rect 22652 9392 22704 9444
rect 29184 9392 29236 9444
rect 4160 9324 4212 9376
rect 6184 9256 6236 9308
rect 10508 9256 10560 9308
rect 6092 9188 6144 9240
rect 12164 9256 12216 9308
rect 13636 9324 13688 9376
rect 21180 9324 21232 9376
rect 13820 9256 13872 9308
rect 17040 9256 17092 9308
rect 17684 9256 17736 9308
rect 24400 9256 24452 9308
rect 38844 9324 38896 9376
rect 13268 9188 13320 9240
rect 17776 9188 17828 9240
rect 4712 9120 4764 9172
rect 8576 9120 8628 9172
rect 13360 9120 13412 9172
rect 29000 9188 29052 9240
rect 28264 9120 28316 9172
rect 29828 9120 29880 9172
rect 3608 9052 3660 9104
rect 10600 9052 10652 9104
rect 12164 8984 12216 9036
rect 30380 9052 30432 9104
rect 38752 9120 38804 9172
rect 35440 9052 35492 9104
rect 4528 8916 4580 8968
rect 7288 8916 7340 8968
rect 13636 8916 13688 8968
rect 13912 8916 13964 8968
rect 37556 8984 37608 9036
rect 24952 8916 25004 8968
rect 25964 8916 26016 8968
rect 34244 8916 34296 8968
rect 37832 8916 37884 8968
rect 10232 8848 10284 8900
rect 14648 8848 14700 8900
rect 16120 8848 16172 8900
rect 20720 8848 20772 8900
rect 27712 8848 27764 8900
rect 32680 8848 32732 8900
rect 33784 8848 33836 8900
rect 35624 8848 35676 8900
rect 2872 8780 2924 8832
rect 6736 8780 6788 8832
rect 7564 8780 7616 8832
rect 8300 8780 8352 8832
rect 11152 8780 11204 8832
rect 15752 8780 15804 8832
rect 19432 8780 19484 8832
rect 22100 8780 22152 8832
rect 24032 8780 24084 8832
rect 24308 8780 24360 8832
rect 26792 8780 26844 8832
rect 34060 8780 34112 8832
rect 36176 8780 36228 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 2872 8576 2924 8628
rect 3792 8576 3844 8628
rect 4344 8576 4396 8628
rect 4896 8576 4948 8628
rect 5908 8576 5960 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7380 8576 7432 8628
rect 7564 8576 7616 8628
rect 8116 8576 8168 8628
rect 8484 8576 8536 8628
rect 8852 8576 8904 8628
rect 9588 8576 9640 8628
rect 10416 8576 10468 8628
rect 10692 8576 10744 8628
rect 10968 8576 11020 8628
rect 11520 8576 11572 8628
rect 12072 8576 12124 8628
rect 12348 8576 12400 8628
rect 12900 8576 12952 8628
rect 13176 8576 13228 8628
rect 13636 8576 13688 8628
rect 14004 8576 14056 8628
rect 14556 8576 14608 8628
rect 14924 8576 14976 8628
rect 15016 8576 15068 8628
rect 1308 8508 1360 8560
rect 1216 8440 1268 8492
rect 388 8372 440 8424
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 4528 8440 4580 8492
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5356 8440 5408 8492
rect 5632 8440 5684 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 4804 8372 4856 8424
rect 572 8304 624 8356
rect 1492 8304 1544 8356
rect 3516 8304 3568 8356
rect 5724 8304 5776 8356
rect 7564 8440 7616 8492
rect 8300 8508 8352 8560
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 13268 8508 13320 8560
rect 13820 8508 13872 8560
rect 15384 8576 15436 8628
rect 15660 8576 15712 8628
rect 16212 8576 16264 8628
rect 16488 8576 16540 8628
rect 16764 8576 16816 8628
rect 19616 8576 19668 8628
rect 22468 8576 22520 8628
rect 22560 8576 22612 8628
rect 8852 8440 8904 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 10048 8440 10100 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 10508 8440 10560 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 7932 8304 7984 8356
rect 11060 8372 11112 8424
rect 8300 8304 8352 8356
rect 8760 8236 8812 8288
rect 9036 8236 9088 8288
rect 10140 8304 10192 8356
rect 12716 8440 12768 8492
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13360 8440 13412 8492
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 14464 8440 14516 8492
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 17776 8508 17828 8560
rect 21640 8508 21692 8560
rect 21732 8508 21784 8560
rect 17316 8440 17368 8492
rect 16028 8372 16080 8424
rect 12716 8304 12768 8356
rect 13636 8304 13688 8356
rect 17960 8440 18012 8492
rect 18052 8483 18104 8492
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 18420 8440 18472 8492
rect 18696 8440 18748 8492
rect 18972 8440 19024 8492
rect 19248 8440 19300 8492
rect 19524 8440 19576 8492
rect 19800 8440 19852 8492
rect 21364 8440 21416 8492
rect 21456 8440 21508 8492
rect 22284 8508 22336 8560
rect 22836 8508 22888 8560
rect 17776 8372 17828 8424
rect 20628 8372 20680 8424
rect 20720 8372 20772 8424
rect 22008 8372 22060 8424
rect 23664 8576 23716 8628
rect 23388 8508 23440 8560
rect 23480 8440 23532 8492
rect 24860 8576 24912 8628
rect 24216 8508 24268 8560
rect 24124 8440 24176 8492
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 25412 8576 25464 8628
rect 25596 8576 25648 8628
rect 25964 8576 26016 8628
rect 28540 8576 28592 8628
rect 28908 8576 28960 8628
rect 25320 8508 25372 8560
rect 26424 8508 26476 8560
rect 17684 8304 17736 8356
rect 17960 8304 18012 8356
rect 19340 8304 19392 8356
rect 20996 8304 21048 8356
rect 21364 8304 21416 8356
rect 22100 8304 22152 8356
rect 11336 8236 11388 8288
rect 14556 8236 14608 8288
rect 14648 8236 14700 8288
rect 18420 8236 18472 8288
rect 18512 8279 18564 8288
rect 18512 8245 18521 8279
rect 18521 8245 18555 8279
rect 18555 8245 18564 8279
rect 18512 8236 18564 8245
rect 18604 8279 18656 8288
rect 18604 8245 18613 8279
rect 18613 8245 18647 8279
rect 18647 8245 18656 8279
rect 18604 8236 18656 8245
rect 19156 8236 19208 8288
rect 19524 8279 19576 8288
rect 19524 8245 19533 8279
rect 19533 8245 19567 8279
rect 19567 8245 19576 8279
rect 19524 8236 19576 8245
rect 20536 8236 20588 8288
rect 20904 8236 20956 8288
rect 23296 8304 23348 8356
rect 23572 8304 23624 8356
rect 23940 8304 23992 8356
rect 24676 8347 24728 8356
rect 24676 8313 24685 8347
rect 24685 8313 24719 8347
rect 24719 8313 24728 8347
rect 24676 8304 24728 8313
rect 25044 8372 25096 8424
rect 27804 8440 27856 8492
rect 28172 8483 28224 8492
rect 28172 8449 28181 8483
rect 28181 8449 28215 8483
rect 28215 8449 28224 8483
rect 28172 8440 28224 8449
rect 25872 8372 25924 8424
rect 26516 8372 26568 8424
rect 28356 8440 28408 8492
rect 29092 8440 29144 8492
rect 30380 8576 30432 8628
rect 32220 8576 32272 8628
rect 32496 8576 32548 8628
rect 32864 8576 32916 8628
rect 33508 8576 33560 8628
rect 33968 8576 34020 8628
rect 29736 8508 29788 8560
rect 34152 8508 34204 8560
rect 35808 8576 35860 8628
rect 36912 8576 36964 8628
rect 35256 8508 35308 8560
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 27436 8304 27488 8356
rect 27620 8304 27672 8356
rect 28724 8372 28776 8424
rect 32404 8372 32456 8424
rect 32680 8440 32732 8492
rect 33692 8483 33744 8492
rect 33692 8449 33701 8483
rect 33701 8449 33735 8483
rect 33735 8449 33744 8483
rect 33692 8440 33744 8449
rect 34244 8372 34296 8424
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35624 8440 35676 8492
rect 32772 8304 32824 8356
rect 33600 8304 33652 8356
rect 22284 8279 22336 8288
rect 22284 8245 22293 8279
rect 22293 8245 22327 8279
rect 22327 8245 22336 8279
rect 22284 8236 22336 8245
rect 22376 8279 22428 8288
rect 22376 8245 22385 8279
rect 22385 8245 22419 8279
rect 22419 8245 22428 8279
rect 22376 8236 22428 8245
rect 22468 8236 22520 8288
rect 23388 8279 23440 8288
rect 23388 8245 23397 8279
rect 23397 8245 23431 8279
rect 23431 8245 23440 8279
rect 23388 8236 23440 8245
rect 23664 8236 23716 8288
rect 24216 8279 24268 8288
rect 24216 8245 24225 8279
rect 24225 8245 24259 8279
rect 24259 8245 24268 8279
rect 24216 8236 24268 8245
rect 24952 8279 25004 8288
rect 24952 8245 24961 8279
rect 24961 8245 24995 8279
rect 24995 8245 25004 8279
rect 24952 8236 25004 8245
rect 26332 8236 26384 8288
rect 26608 8236 26660 8288
rect 29184 8236 29236 8288
rect 30196 8236 30248 8288
rect 31944 8236 31996 8288
rect 35072 8372 35124 8424
rect 34704 8304 34756 8356
rect 36820 8508 36872 8560
rect 36176 8483 36228 8492
rect 36176 8449 36185 8483
rect 36185 8449 36219 8483
rect 36219 8449 36228 8483
rect 36176 8440 36228 8449
rect 36544 8483 36596 8492
rect 36544 8449 36553 8483
rect 36553 8449 36587 8483
rect 36587 8449 36596 8483
rect 36544 8440 36596 8449
rect 37096 8440 37148 8492
rect 37464 8508 37516 8560
rect 38752 8508 38804 8560
rect 36360 8372 36412 8424
rect 35900 8236 35952 8288
rect 37464 8372 37516 8424
rect 38476 8440 38528 8492
rect 38844 8483 38896 8492
rect 38844 8449 38853 8483
rect 38853 8449 38887 8483
rect 38887 8449 38896 8483
rect 38844 8440 38896 8449
rect 37188 8304 37240 8356
rect 39028 8347 39080 8356
rect 39028 8313 39037 8347
rect 39037 8313 39071 8347
rect 39071 8313 39080 8347
rect 39028 8304 39080 8313
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 3332 8032 3384 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 4068 8032 4120 8084
rect 4620 8032 4672 8084
rect 5172 8032 5224 8084
rect 6552 8032 6604 8084
rect 7104 8032 7156 8084
rect 7656 8032 7708 8084
rect 8760 8032 8812 8084
rect 9036 8075 9088 8084
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 9404 8032 9456 8084
rect 9864 8032 9916 8084
rect 11244 8032 11296 8084
rect 11796 8032 11848 8084
rect 12624 8032 12676 8084
rect 1032 7964 1084 8016
rect 1124 7896 1176 7948
rect 756 7828 808 7880
rect 848 7760 900 7812
rect 1860 7828 1912 7880
rect 9128 7964 9180 8016
rect 10784 8007 10836 8016
rect 10784 7973 10793 8007
rect 10793 7973 10827 8007
rect 10827 7973 10836 8007
rect 10784 7964 10836 7973
rect 12900 7964 12952 8016
rect 14280 8032 14332 8084
rect 14832 8032 14884 8084
rect 15476 8032 15528 8084
rect 15936 8032 15988 8084
rect 17592 8032 17644 8084
rect 19524 8032 19576 8084
rect 20628 8032 20680 8084
rect 20720 8032 20772 8084
rect 24400 8075 24452 8084
rect 24400 8041 24409 8075
rect 24409 8041 24443 8075
rect 24443 8041 24452 8075
rect 24400 8032 24452 8041
rect 26516 8032 26568 8084
rect 13728 7964 13780 8016
rect 16304 7964 16356 8016
rect 19800 7964 19852 8016
rect 22192 8007 22244 8016
rect 22192 7973 22201 8007
rect 22201 7973 22235 8007
rect 22235 7973 22244 8007
rect 22192 7964 22244 7973
rect 22468 7964 22520 8016
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 2872 7760 2924 7812
rect 5908 7803 5960 7812
rect 5908 7769 5917 7803
rect 5917 7769 5951 7803
rect 5951 7769 5960 7803
rect 5908 7760 5960 7769
rect 6276 7803 6328 7812
rect 6276 7769 6285 7803
rect 6285 7769 6319 7803
rect 6319 7769 6328 7803
rect 6276 7760 6328 7769
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8484 7828 8536 7880
rect 8668 7828 8720 7880
rect 9404 7828 9456 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 8944 7760 8996 7812
rect 10324 7760 10376 7812
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 5816 7692 5868 7744
rect 6368 7692 6420 7744
rect 8024 7692 8076 7744
rect 10048 7692 10100 7744
rect 10876 7896 10928 7948
rect 12164 7871 12216 7880
rect 12164 7837 12173 7871
rect 12173 7837 12207 7871
rect 12207 7837 12216 7871
rect 12164 7828 12216 7837
rect 12624 7760 12676 7812
rect 13452 7760 13504 7812
rect 12900 7692 12952 7744
rect 14188 7828 14240 7880
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 15384 7828 15436 7880
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 16396 7828 16448 7880
rect 17500 7760 17552 7812
rect 17684 7828 17736 7880
rect 19524 7828 19576 7880
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 20444 7871 20496 7880
rect 18328 7760 18380 7812
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 20996 7896 21048 7948
rect 15568 7692 15620 7744
rect 16672 7692 16724 7744
rect 17684 7692 17736 7744
rect 17776 7735 17828 7744
rect 17776 7701 17785 7735
rect 17785 7701 17819 7735
rect 17819 7701 17828 7735
rect 17776 7692 17828 7701
rect 19708 7692 19760 7744
rect 21088 7828 21140 7880
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 20720 7803 20772 7812
rect 20720 7769 20729 7803
rect 20729 7769 20763 7803
rect 20763 7769 20772 7803
rect 20720 7760 20772 7769
rect 21824 7760 21876 7812
rect 23388 7828 23440 7880
rect 25780 7964 25832 8016
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 21456 7692 21508 7744
rect 22284 7692 22336 7744
rect 28264 7760 28316 7812
rect 30196 7896 30248 7948
rect 29460 7828 29512 7880
rect 34428 8032 34480 8084
rect 35532 8032 35584 8084
rect 36084 8032 36136 8084
rect 36636 8032 36688 8084
rect 37740 8032 37792 8084
rect 37004 7964 37056 8016
rect 39764 7964 39816 8016
rect 32588 7896 32640 7948
rect 35164 7828 35216 7880
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 25504 7735 25556 7744
rect 25504 7701 25513 7735
rect 25513 7701 25547 7735
rect 25547 7701 25556 7735
rect 25504 7692 25556 7701
rect 28448 7692 28500 7744
rect 28816 7760 28868 7812
rect 29184 7760 29236 7812
rect 36452 7871 36504 7880
rect 36452 7837 36461 7871
rect 36461 7837 36495 7871
rect 36495 7837 36504 7871
rect 36452 7828 36504 7837
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 38292 7828 38344 7880
rect 29092 7692 29144 7744
rect 30472 7692 30524 7744
rect 31944 7735 31996 7744
rect 31944 7701 31953 7735
rect 31953 7701 31987 7735
rect 31987 7701 31996 7735
rect 31944 7692 31996 7701
rect 32772 7735 32824 7744
rect 32772 7701 32781 7735
rect 32781 7701 32815 7735
rect 32815 7701 32824 7735
rect 32772 7692 32824 7701
rect 33416 7692 33468 7744
rect 33508 7735 33560 7744
rect 33508 7701 33517 7735
rect 33517 7701 33551 7735
rect 33551 7701 33560 7735
rect 33508 7692 33560 7701
rect 35072 7735 35124 7744
rect 35072 7701 35081 7735
rect 35081 7701 35115 7735
rect 35115 7701 35124 7735
rect 35072 7692 35124 7701
rect 37648 7760 37700 7812
rect 40132 7760 40184 7812
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 5540 7488 5592 7540
rect 7840 7488 7892 7540
rect 940 7420 992 7472
rect 756 7352 808 7404
rect 2412 7420 2464 7472
rect 10876 7420 10928 7472
rect 12164 7420 12216 7472
rect 15476 7488 15528 7540
rect 21640 7488 21692 7540
rect 25688 7488 25740 7540
rect 29184 7488 29236 7540
rect 29276 7488 29328 7540
rect 664 7284 716 7336
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 8392 7352 8444 7404
rect 2872 7284 2924 7336
rect 3884 7216 3936 7268
rect 3976 7148 4028 7200
rect 5816 7284 5868 7336
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 13728 7327 13780 7336
rect 13728 7293 13737 7327
rect 13737 7293 13771 7327
rect 13771 7293 13780 7327
rect 13728 7284 13780 7293
rect 6920 7216 6972 7268
rect 7288 7148 7340 7200
rect 7840 7191 7892 7200
rect 7840 7157 7849 7191
rect 7849 7157 7883 7191
rect 7883 7157 7892 7191
rect 7840 7148 7892 7157
rect 8576 7259 8628 7268
rect 8576 7225 8585 7259
rect 8585 7225 8619 7259
rect 8619 7225 8628 7259
rect 8576 7216 8628 7225
rect 9772 7216 9824 7268
rect 10876 7259 10928 7268
rect 10876 7225 10885 7259
rect 10885 7225 10919 7259
rect 10919 7225 10928 7259
rect 10876 7216 10928 7225
rect 12440 7216 12492 7268
rect 10140 7148 10192 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 17868 7352 17920 7404
rect 18144 7352 18196 7404
rect 20444 7352 20496 7404
rect 24768 7420 24820 7472
rect 29092 7420 29144 7472
rect 29920 7420 29972 7472
rect 25504 7395 25556 7404
rect 25504 7361 25513 7395
rect 25513 7361 25547 7395
rect 25547 7361 25556 7395
rect 25504 7352 25556 7361
rect 25688 7352 25740 7404
rect 25872 7352 25924 7404
rect 38384 7488 38436 7540
rect 38660 7531 38712 7540
rect 38660 7497 38669 7531
rect 38669 7497 38703 7531
rect 38703 7497 38712 7531
rect 38660 7488 38712 7497
rect 38936 7488 38988 7540
rect 39580 7488 39632 7540
rect 37372 7420 37424 7472
rect 38108 7395 38160 7404
rect 38108 7361 38117 7395
rect 38117 7361 38151 7395
rect 38151 7361 38160 7395
rect 38108 7352 38160 7361
rect 38568 7352 38620 7404
rect 38844 7395 38896 7404
rect 38844 7361 38853 7395
rect 38853 7361 38887 7395
rect 38887 7361 38896 7395
rect 38844 7352 38896 7361
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 16488 7191 16540 7200
rect 16488 7157 16497 7191
rect 16497 7157 16531 7191
rect 16531 7157 16540 7191
rect 16488 7148 16540 7157
rect 23112 7284 23164 7336
rect 23204 7284 23256 7336
rect 26516 7284 26568 7336
rect 27436 7284 27488 7336
rect 28172 7284 28224 7336
rect 28448 7284 28500 7336
rect 38292 7284 38344 7336
rect 19524 7216 19576 7268
rect 20904 7216 20956 7268
rect 21824 7216 21876 7268
rect 18144 7191 18196 7200
rect 18144 7157 18153 7191
rect 18153 7157 18187 7191
rect 18187 7157 18196 7191
rect 18144 7148 18196 7157
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 18512 7148 18564 7200
rect 31944 7216 31996 7268
rect 39304 7216 39356 7268
rect 28356 7148 28408 7200
rect 28448 7148 28500 7200
rect 28724 7148 28776 7200
rect 30380 7191 30432 7200
rect 30380 7157 30389 7191
rect 30389 7157 30423 7191
rect 30423 7157 30432 7191
rect 30380 7148 30432 7157
rect 33416 7148 33468 7200
rect 39856 7148 39908 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 1124 6944 1176 6996
rect 2688 6944 2740 6996
rect 1032 6808 1084 6860
rect 5908 6876 5960 6928
rect 756 6740 808 6792
rect 848 6672 900 6724
rect 5356 6740 5408 6792
rect 6828 6740 6880 6792
rect 7748 6740 7800 6792
rect 9680 6944 9732 6996
rect 9772 6876 9824 6928
rect 9956 6876 10008 6928
rect 10232 6944 10284 6996
rect 11428 6876 11480 6928
rect 11520 6876 11572 6928
rect 16488 6944 16540 6996
rect 38844 6944 38896 6996
rect 8484 6808 8536 6860
rect 11704 6808 11756 6860
rect 11520 6740 11572 6792
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12440 6808 12492 6817
rect 13728 6808 13780 6860
rect 13820 6808 13872 6860
rect 22100 6808 22152 6860
rect 12624 6740 12676 6792
rect 21824 6740 21876 6792
rect 23848 6740 23900 6792
rect 24308 6740 24360 6792
rect 2596 6604 2648 6656
rect 3976 6604 4028 6656
rect 11612 6672 11664 6724
rect 11704 6672 11756 6724
rect 24676 6672 24728 6724
rect 25964 6876 26016 6928
rect 28448 6876 28500 6928
rect 28632 6876 28684 6928
rect 35072 6876 35124 6928
rect 27436 6808 27488 6860
rect 27988 6808 28040 6860
rect 28908 6808 28960 6860
rect 25228 6783 25280 6792
rect 25228 6749 25237 6783
rect 25237 6749 25271 6783
rect 25271 6749 25280 6783
rect 25228 6740 25280 6749
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 27804 6740 27856 6792
rect 28172 6740 28224 6792
rect 28724 6783 28776 6792
rect 28724 6749 28733 6783
rect 28733 6749 28767 6783
rect 28767 6749 28776 6783
rect 28724 6740 28776 6749
rect 30840 6740 30892 6792
rect 37556 6740 37608 6792
rect 38016 6740 38068 6792
rect 38200 6783 38252 6792
rect 38200 6749 38209 6783
rect 38209 6749 38243 6783
rect 38243 6749 38252 6783
rect 38200 6740 38252 6749
rect 38476 6783 38528 6792
rect 38476 6749 38485 6783
rect 38485 6749 38519 6783
rect 38519 6749 38528 6783
rect 38476 6740 38528 6749
rect 27988 6672 28040 6724
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 10968 6604 11020 6656
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 13728 6604 13780 6656
rect 14832 6604 14884 6656
rect 16672 6604 16724 6656
rect 17776 6604 17828 6656
rect 21916 6604 21968 6656
rect 23296 6604 23348 6656
rect 24584 6604 24636 6656
rect 25044 6604 25096 6656
rect 25228 6604 25280 6656
rect 25320 6604 25372 6656
rect 25964 6604 26016 6656
rect 26608 6604 26660 6656
rect 27436 6647 27488 6656
rect 27436 6613 27445 6647
rect 27445 6613 27479 6647
rect 27479 6613 27488 6647
rect 27436 6604 27488 6613
rect 27896 6604 27948 6656
rect 37280 6647 37332 6656
rect 37280 6613 37289 6647
rect 37289 6613 37323 6647
rect 37323 6613 37332 6647
rect 37280 6604 37332 6613
rect 37556 6604 37608 6656
rect 38384 6647 38436 6656
rect 38384 6613 38393 6647
rect 38393 6613 38427 6647
rect 38427 6613 38436 6647
rect 38384 6604 38436 6613
rect 38660 6647 38712 6656
rect 38660 6613 38669 6647
rect 38669 6613 38703 6647
rect 38703 6613 38712 6647
rect 38660 6604 38712 6613
rect 40040 6672 40092 6724
rect 39488 6604 39540 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 5448 6400 5500 6452
rect 5632 6400 5684 6452
rect 13452 6400 13504 6452
rect 15108 6400 15160 6452
rect 16212 6400 16264 6452
rect 19708 6400 19760 6452
rect 20444 6400 20496 6452
rect 20628 6400 20680 6452
rect 21548 6400 21600 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 22100 6443 22152 6452
rect 22100 6409 22109 6443
rect 22109 6409 22143 6443
rect 22143 6409 22152 6443
rect 22100 6400 22152 6409
rect 24308 6400 24360 6452
rect 37556 6400 37608 6452
rect 37648 6443 37700 6452
rect 37648 6409 37657 6443
rect 37657 6409 37691 6443
rect 37691 6409 37700 6443
rect 37648 6400 37700 6409
rect 39580 6400 39632 6452
rect 2596 6375 2648 6384
rect 2596 6341 2605 6375
rect 2605 6341 2639 6375
rect 2639 6341 2648 6375
rect 2596 6332 2648 6341
rect 204 6264 256 6316
rect 5540 6332 5592 6384
rect 9404 6332 9456 6384
rect 848 6196 900 6248
rect 2504 6196 2556 6248
rect 5080 6196 5132 6248
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 8484 6264 8536 6316
rect 10692 6332 10744 6384
rect 15016 6332 15068 6384
rect 10140 6306 10192 6316
rect 10140 6272 10148 6306
rect 10148 6272 10192 6306
rect 10140 6264 10192 6272
rect 13820 6264 13872 6316
rect 16948 6264 17000 6316
rect 17684 6264 17736 6316
rect 19800 6375 19852 6384
rect 19800 6341 19809 6375
rect 19809 6341 19843 6375
rect 19843 6341 19852 6375
rect 19800 6332 19852 6341
rect 2688 6128 2740 6180
rect 2780 6171 2832 6180
rect 2780 6137 2789 6171
rect 2789 6137 2823 6171
rect 2823 6137 2832 6171
rect 2780 6128 2832 6137
rect 1584 6060 1636 6112
rect 9220 6128 9272 6180
rect 14832 6239 14884 6248
rect 14832 6205 14841 6239
rect 14841 6205 14875 6239
rect 14875 6205 14884 6239
rect 14832 6196 14884 6205
rect 13452 6128 13504 6180
rect 19432 6128 19484 6180
rect 5816 6060 5868 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 8300 6060 8352 6112
rect 9128 6060 9180 6112
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 19248 6103 19300 6112
rect 19248 6069 19257 6103
rect 19257 6069 19291 6103
rect 19291 6069 19300 6103
rect 19248 6060 19300 6069
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 20628 6307 20680 6316
rect 20628 6273 20646 6307
rect 20646 6273 20680 6307
rect 20628 6264 20680 6273
rect 23388 6332 23440 6384
rect 25596 6332 25648 6384
rect 25872 6332 25924 6384
rect 27712 6332 27764 6384
rect 27988 6332 28040 6384
rect 23940 6264 23992 6316
rect 24216 6264 24268 6316
rect 26424 6264 26476 6316
rect 27528 6264 27580 6316
rect 30656 6307 30708 6316
rect 30656 6273 30665 6307
rect 30665 6273 30699 6307
rect 30699 6273 30708 6307
rect 30656 6264 30708 6273
rect 30748 6264 30800 6316
rect 38384 6332 38436 6384
rect 39488 6332 39540 6384
rect 20904 6128 20956 6180
rect 25412 6196 25464 6248
rect 26700 6196 26752 6248
rect 37556 6196 37608 6248
rect 38844 6307 38896 6316
rect 38844 6273 38853 6307
rect 38853 6273 38887 6307
rect 38887 6273 38896 6307
rect 38844 6264 38896 6273
rect 38936 6264 38988 6316
rect 25780 6128 25832 6180
rect 27344 6128 27396 6180
rect 27528 6128 27580 6180
rect 27804 6128 27856 6180
rect 34060 6171 34112 6180
rect 34060 6137 34069 6171
rect 34069 6137 34103 6171
rect 34103 6137 34112 6171
rect 34060 6128 34112 6137
rect 39672 6128 39724 6180
rect 21916 6060 21968 6112
rect 24216 6060 24268 6112
rect 24400 6060 24452 6112
rect 29736 6060 29788 6112
rect 30840 6103 30892 6112
rect 30840 6069 30849 6103
rect 30849 6069 30883 6103
rect 30883 6069 30892 6103
rect 30840 6060 30892 6069
rect 37740 6060 37792 6112
rect 38016 6060 38068 6112
rect 38476 6060 38528 6112
rect 38660 6103 38712 6112
rect 38660 6069 38669 6103
rect 38669 6069 38703 6103
rect 38703 6069 38712 6103
rect 38660 6060 38712 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 2504 5856 2556 5908
rect 6828 5856 6880 5908
rect 5632 5788 5684 5840
rect 6736 5788 6788 5840
rect 14556 5856 14608 5908
rect 16948 5899 17000 5908
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 10140 5788 10192 5840
rect 10692 5831 10744 5840
rect 10692 5797 10701 5831
rect 10701 5797 10735 5831
rect 10735 5797 10744 5831
rect 10692 5788 10744 5797
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 5264 5763 5316 5772
rect 5264 5729 5273 5763
rect 5273 5729 5307 5763
rect 5307 5729 5316 5763
rect 5264 5720 5316 5729
rect 756 5652 808 5704
rect 848 5584 900 5636
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6092 5695 6144 5704
rect 6092 5661 6126 5695
rect 6126 5661 6144 5695
rect 6092 5652 6144 5661
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 9680 5652 9732 5704
rect 4160 5516 4212 5568
rect 6092 5516 6144 5568
rect 6736 5516 6788 5568
rect 10140 5695 10192 5704
rect 10140 5661 10150 5695
rect 10150 5661 10184 5695
rect 10184 5661 10192 5695
rect 10968 5720 11020 5772
rect 13452 5788 13504 5840
rect 23388 5856 23440 5908
rect 37832 5856 37884 5908
rect 38476 5856 38528 5908
rect 39396 5899 39448 5908
rect 39396 5865 39405 5899
rect 39405 5865 39439 5899
rect 39439 5865 39448 5899
rect 39396 5856 39448 5865
rect 19248 5788 19300 5840
rect 24400 5788 24452 5840
rect 13728 5720 13780 5772
rect 15844 5720 15896 5772
rect 10140 5652 10192 5661
rect 10324 5627 10376 5636
rect 10324 5593 10333 5627
rect 10333 5593 10367 5627
rect 10367 5593 10376 5627
rect 10324 5584 10376 5593
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 10600 5516 10652 5568
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11612 5652 11664 5704
rect 14556 5652 14608 5704
rect 21916 5720 21968 5772
rect 22008 5720 22060 5772
rect 24308 5720 24360 5772
rect 20628 5652 20680 5704
rect 23296 5652 23348 5704
rect 23940 5652 23992 5704
rect 24584 5652 24636 5704
rect 24768 5652 24820 5704
rect 25964 5695 26016 5704
rect 25964 5661 25973 5695
rect 25973 5661 26007 5695
rect 26007 5661 26016 5695
rect 25964 5652 26016 5661
rect 26148 5695 26200 5704
rect 26148 5661 26161 5695
rect 26161 5661 26200 5695
rect 26148 5652 26200 5661
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 14372 5584 14424 5636
rect 15384 5584 15436 5636
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 18420 5516 18472 5568
rect 19616 5516 19668 5568
rect 26608 5695 26660 5704
rect 26608 5661 26617 5695
rect 26617 5661 26651 5695
rect 26651 5661 26660 5695
rect 26608 5652 26660 5661
rect 26884 5695 26936 5704
rect 26884 5661 26893 5695
rect 26893 5661 26927 5695
rect 26927 5661 26936 5695
rect 26884 5652 26936 5661
rect 27344 5695 27396 5704
rect 27344 5661 27351 5695
rect 27351 5661 27396 5695
rect 27344 5652 27396 5661
rect 27436 5695 27488 5704
rect 27436 5661 27445 5695
rect 27445 5661 27479 5695
rect 27479 5661 27488 5695
rect 27436 5652 27488 5661
rect 28080 5788 28132 5840
rect 30748 5788 30800 5840
rect 30840 5788 30892 5840
rect 38660 5788 38712 5840
rect 39948 5788 40000 5840
rect 31116 5720 31168 5772
rect 29368 5652 29420 5704
rect 29736 5652 29788 5704
rect 37280 5652 37332 5704
rect 37372 5652 37424 5704
rect 38844 5695 38896 5704
rect 38844 5661 38853 5695
rect 38853 5661 38887 5695
rect 38887 5661 38896 5695
rect 38844 5652 38896 5661
rect 39212 5695 39264 5704
rect 39212 5661 39221 5695
rect 39221 5661 39255 5695
rect 39255 5661 39264 5695
rect 39212 5652 39264 5661
rect 23848 5516 23900 5568
rect 24124 5516 24176 5568
rect 26148 5516 26200 5568
rect 26608 5516 26660 5568
rect 27896 5516 27948 5568
rect 30012 5516 30064 5568
rect 34152 5516 34204 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 14924 5312 14976 5364
rect 1676 5244 1728 5296
rect 24860 5312 24912 5364
rect 26424 5312 26476 5364
rect 26884 5312 26936 5364
rect 28080 5312 28132 5364
rect 33692 5312 33744 5364
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 19432 5244 19484 5296
rect 24124 5244 24176 5296
rect 25044 5244 25096 5296
rect 25136 5244 25188 5296
rect 756 5176 808 5228
rect 6092 5176 6144 5228
rect 8392 5176 8444 5228
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 5816 5108 5868 5160
rect 2780 5040 2832 5092
rect 10600 5219 10652 5228
rect 10600 5185 10639 5219
rect 10639 5185 10652 5219
rect 10600 5176 10652 5185
rect 10232 5108 10284 5160
rect 10968 5176 11020 5228
rect 23756 5176 23808 5228
rect 25964 5176 26016 5228
rect 27528 5244 27580 5296
rect 38936 5244 38988 5296
rect 28724 5176 28776 5228
rect 12256 5108 12308 5160
rect 20536 5108 20588 5160
rect 20812 5108 20864 5160
rect 21548 5108 21600 5160
rect 22008 5108 22060 5160
rect 24768 5108 24820 5160
rect 25136 5108 25188 5160
rect 33416 5176 33468 5228
rect 37740 5176 37792 5228
rect 38844 5219 38896 5228
rect 38844 5185 38853 5219
rect 38853 5185 38887 5219
rect 38887 5185 38896 5219
rect 38844 5176 38896 5185
rect 39212 5219 39264 5228
rect 39212 5185 39221 5219
rect 39221 5185 39255 5219
rect 39255 5185 39264 5219
rect 39212 5176 39264 5185
rect 7196 4972 7248 5024
rect 7472 4972 7524 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 11520 5040 11572 5092
rect 12808 5040 12860 5092
rect 10416 4972 10468 5024
rect 10508 4972 10560 5024
rect 14648 4972 14700 5024
rect 18604 4972 18656 5024
rect 19064 5040 19116 5092
rect 38752 5108 38804 5160
rect 33784 5040 33836 5092
rect 20812 4972 20864 5024
rect 20904 4972 20956 5024
rect 21364 4972 21416 5024
rect 21548 4972 21600 5024
rect 23388 4972 23440 5024
rect 25504 4972 25556 5024
rect 27712 4972 27764 5024
rect 38292 5040 38344 5092
rect 33968 4972 34020 5024
rect 37464 4972 37516 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 7196 4768 7248 4820
rect 8392 4700 8444 4752
rect 10324 4768 10376 4820
rect 10416 4768 10468 4820
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 5264 4675 5316 4684
rect 5264 4641 5273 4675
rect 5273 4641 5307 4675
rect 5307 4641 5316 4675
rect 5264 4632 5316 4641
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 5816 4632 5868 4684
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 8300 4632 8352 4684
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6092 4607 6144 4616
rect 6092 4573 6126 4607
rect 6126 4573 6144 4607
rect 6092 4564 6144 4573
rect 8484 4607 8536 4616
rect 388 4496 440 4548
rect 3516 4539 3568 4548
rect 3516 4505 3525 4539
rect 3525 4505 3559 4539
rect 3559 4505 3568 4539
rect 3516 4496 3568 4505
rect 4528 4428 4580 4480
rect 8484 4573 8492 4607
rect 8492 4573 8526 4607
rect 8526 4573 8536 4607
rect 8484 4564 8536 4573
rect 8760 4632 8812 4684
rect 10600 4632 10652 4684
rect 10876 4564 10928 4616
rect 8208 4539 8260 4548
rect 8208 4505 8217 4539
rect 8217 4505 8251 4539
rect 8251 4505 8260 4539
rect 8208 4496 8260 4505
rect 10600 4539 10652 4548
rect 10600 4505 10609 4539
rect 10609 4505 10643 4539
rect 10643 4505 10652 4539
rect 10600 4496 10652 4505
rect 10968 4496 11020 4548
rect 10508 4471 10560 4480
rect 10508 4437 10517 4471
rect 10517 4437 10551 4471
rect 10551 4437 10560 4471
rect 10508 4428 10560 4437
rect 11980 4428 12032 4480
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 13636 4743 13688 4752
rect 13636 4709 13645 4743
rect 13645 4709 13679 4743
rect 13679 4709 13688 4743
rect 13636 4700 13688 4709
rect 13820 4632 13872 4684
rect 14464 4564 14516 4616
rect 14740 4564 14792 4616
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 17960 4768 18012 4820
rect 19064 4811 19116 4820
rect 19064 4777 19073 4811
rect 19073 4777 19107 4811
rect 19107 4777 19116 4811
rect 19064 4768 19116 4777
rect 19340 4768 19392 4820
rect 20904 4811 20956 4820
rect 20904 4777 20913 4811
rect 20913 4777 20947 4811
rect 20947 4777 20956 4811
rect 20904 4768 20956 4777
rect 16396 4564 16448 4616
rect 18144 4564 18196 4616
rect 18788 4564 18840 4616
rect 18880 4607 18932 4616
rect 18880 4573 18889 4607
rect 18889 4573 18923 4607
rect 18923 4573 18932 4607
rect 18880 4564 18932 4573
rect 19432 4564 19484 4616
rect 14464 4428 14516 4480
rect 17408 4496 17460 4548
rect 22008 4632 22060 4684
rect 23112 4811 23164 4820
rect 23112 4777 23121 4811
rect 23121 4777 23155 4811
rect 23155 4777 23164 4811
rect 23112 4768 23164 4777
rect 23388 4811 23440 4820
rect 23388 4777 23397 4811
rect 23397 4777 23431 4811
rect 23431 4777 23440 4811
rect 23388 4768 23440 4777
rect 24860 4811 24912 4820
rect 24860 4777 24869 4811
rect 24869 4777 24903 4811
rect 24903 4777 24912 4811
rect 24860 4768 24912 4777
rect 27528 4768 27580 4820
rect 23296 4700 23348 4752
rect 22652 4632 22704 4684
rect 25044 4675 25096 4684
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 26608 4700 26660 4752
rect 27344 4632 27396 4684
rect 29368 4811 29420 4820
rect 29368 4777 29377 4811
rect 29377 4777 29411 4811
rect 29411 4777 29420 4811
rect 29368 4768 29420 4777
rect 29920 4811 29972 4820
rect 29920 4777 29929 4811
rect 29929 4777 29963 4811
rect 29963 4777 29972 4811
rect 29920 4768 29972 4777
rect 33968 4768 34020 4820
rect 34980 4811 35032 4820
rect 34980 4777 34989 4811
rect 34989 4777 35023 4811
rect 35023 4777 35032 4811
rect 34980 4768 35032 4777
rect 35164 4768 35216 4820
rect 37096 4811 37148 4820
rect 37096 4777 37105 4811
rect 37105 4777 37139 4811
rect 37139 4777 37148 4811
rect 37096 4768 37148 4777
rect 37832 4768 37884 4820
rect 39396 4811 39448 4820
rect 39396 4777 39405 4811
rect 39405 4777 39439 4811
rect 39439 4777 39448 4811
rect 39396 4768 39448 4777
rect 31392 4700 31444 4752
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 23572 4607 23624 4616
rect 23572 4573 23581 4607
rect 23581 4573 23615 4607
rect 23615 4573 23624 4607
rect 23572 4564 23624 4573
rect 25228 4564 25280 4616
rect 26332 4564 26384 4616
rect 27528 4607 27580 4616
rect 27528 4573 27537 4607
rect 27537 4573 27571 4607
rect 27571 4573 27580 4607
rect 27528 4564 27580 4573
rect 24860 4496 24912 4548
rect 26792 4496 26844 4548
rect 27436 4496 27488 4548
rect 28448 4607 28500 4616
rect 28448 4573 28457 4607
rect 28457 4573 28491 4607
rect 28491 4573 28500 4607
rect 28448 4564 28500 4573
rect 28632 4564 28684 4616
rect 32588 4632 32640 4684
rect 30104 4607 30156 4616
rect 30104 4573 30113 4607
rect 30113 4573 30147 4607
rect 30147 4573 30156 4607
rect 30104 4564 30156 4573
rect 35992 4564 36044 4616
rect 38568 4607 38620 4616
rect 38568 4573 38577 4607
rect 38577 4573 38611 4607
rect 38611 4573 38620 4607
rect 38568 4564 38620 4573
rect 38752 4564 38804 4616
rect 36268 4496 36320 4548
rect 38476 4496 38528 4548
rect 38936 4496 38988 4548
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 21548 4428 21600 4480
rect 21732 4428 21784 4480
rect 25320 4428 25372 4480
rect 27620 4428 27672 4480
rect 28632 4428 28684 4480
rect 28724 4428 28776 4480
rect 34796 4471 34848 4480
rect 34796 4437 34805 4471
rect 34805 4437 34839 4471
rect 34839 4437 34848 4471
rect 34796 4428 34848 4437
rect 36452 4428 36504 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 5724 4224 5776 4276
rect 1216 4156 1268 4208
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 8208 4224 8260 4276
rect 8300 4224 8352 4276
rect 10876 4224 10928 4276
rect 11520 4224 11572 4276
rect 14648 4267 14700 4276
rect 14648 4233 14657 4267
rect 14657 4233 14691 4267
rect 14691 4233 14700 4267
rect 14648 4224 14700 4233
rect 17224 4224 17276 4276
rect 19432 4224 19484 4276
rect 20260 4224 20312 4276
rect 21916 4224 21968 4276
rect 24492 4224 24544 4276
rect 27436 4224 27488 4276
rect 30104 4224 30156 4276
rect 8760 4156 8812 4208
rect 10508 4156 10560 4208
rect 10232 4088 10284 4140
rect 10600 4088 10652 4140
rect 22376 4156 22428 4208
rect 25688 4156 25740 4208
rect 14372 4088 14424 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17224 4088 17276 4140
rect 17500 4088 17552 4140
rect 25228 4131 25280 4140
rect 25228 4097 25237 4131
rect 25237 4097 25271 4131
rect 25271 4097 25280 4131
rect 25228 4088 25280 4097
rect 27620 4088 27672 4140
rect 28448 4088 28500 4140
rect 29092 4088 29144 4140
rect 30288 4088 30340 4140
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 3792 3952 3844 3961
rect 7288 4020 7340 4072
rect 10048 3952 10100 4004
rect 5908 3884 5960 3936
rect 9956 3884 10008 3936
rect 14464 4063 14516 4072
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 14740 4020 14792 4072
rect 15384 3952 15436 4004
rect 16948 4020 17000 4072
rect 26884 4020 26936 4072
rect 28264 4020 28316 4072
rect 37280 4063 37332 4072
rect 37280 4029 37289 4063
rect 37289 4029 37323 4063
rect 37323 4029 37332 4063
rect 37280 4020 37332 4029
rect 21364 3952 21416 4004
rect 21548 3952 21600 4004
rect 22928 3952 22980 4004
rect 16580 3884 16632 3936
rect 17684 3927 17736 3936
rect 17684 3893 17693 3927
rect 17693 3893 17727 3927
rect 17727 3893 17736 3927
rect 17684 3884 17736 3893
rect 19156 3884 19208 3936
rect 23480 3884 23532 3936
rect 27712 3995 27764 4004
rect 27712 3961 27721 3995
rect 27721 3961 27755 3995
rect 27755 3961 27764 3995
rect 27712 3952 27764 3961
rect 38844 4131 38896 4140
rect 38844 4097 38853 4131
rect 38853 4097 38887 4131
rect 38887 4097 38896 4131
rect 38844 4088 38896 4097
rect 39488 4088 39540 4140
rect 29000 3884 29052 3936
rect 30472 3884 30524 3936
rect 39028 3995 39080 4004
rect 39028 3961 39037 3995
rect 39037 3961 39071 3995
rect 39071 3961 39080 3995
rect 39028 3952 39080 3961
rect 39396 3995 39448 4004
rect 39396 3961 39405 3995
rect 39405 3961 39439 3995
rect 39439 3961 39448 3995
rect 39396 3952 39448 3961
rect 32312 3927 32364 3936
rect 32312 3893 32321 3927
rect 32321 3893 32355 3927
rect 32355 3893 32364 3927
rect 32312 3884 32364 3893
rect 38660 3927 38712 3936
rect 38660 3893 38669 3927
rect 38669 3893 38703 3927
rect 38703 3893 38712 3927
rect 38660 3884 38712 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 16028 3680 16080 3732
rect 4436 3612 4488 3664
rect 17684 3612 17736 3664
rect 5448 3476 5500 3528
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 15476 3476 15528 3528
rect 5816 3451 5868 3460
rect 5816 3417 5825 3451
rect 5825 3417 5859 3451
rect 5859 3417 5868 3451
rect 5816 3408 5868 3417
rect 5908 3408 5960 3460
rect 6828 3408 6880 3460
rect 16672 3408 16724 3460
rect 26608 3612 26660 3664
rect 26976 3680 27028 3732
rect 32404 3680 32456 3732
rect 39580 3680 39632 3732
rect 27068 3612 27120 3664
rect 30380 3612 30432 3664
rect 38936 3612 38988 3664
rect 39948 3612 40000 3664
rect 18880 3476 18932 3528
rect 20444 3544 20496 3596
rect 21364 3544 21416 3596
rect 20352 3476 20404 3528
rect 22376 3476 22428 3528
rect 26516 3476 26568 3528
rect 30288 3544 30340 3596
rect 33876 3544 33928 3596
rect 36544 3544 36596 3596
rect 29184 3476 29236 3528
rect 36820 3476 36872 3528
rect 38752 3476 38804 3528
rect 39764 3476 39816 3528
rect 19340 3408 19392 3460
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 14280 3340 14332 3392
rect 20168 3340 20220 3392
rect 22192 3340 22244 3392
rect 23296 3340 23348 3392
rect 24676 3340 24728 3392
rect 27068 3408 27120 3460
rect 34612 3408 34664 3460
rect 26884 3340 26936 3392
rect 27344 3340 27396 3392
rect 29276 3340 29328 3392
rect 29460 3340 29512 3392
rect 33876 3340 33928 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 16948 3136 17000 3188
rect 16580 3068 16632 3120
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 20168 3136 20220 3188
rect 22008 3136 22060 3188
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 20444 3068 20496 3120
rect 5356 2932 5408 2984
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 16672 2864 16724 2916
rect 21916 3043 21968 3052
rect 21916 3009 21926 3043
rect 21926 3009 21960 3043
rect 21960 3009 21968 3043
rect 21916 3000 21968 3009
rect 22192 2932 22244 2984
rect 22928 3043 22980 3052
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 22928 3000 22980 3009
rect 23296 3043 23348 3052
rect 23296 3009 23335 3043
rect 23335 3009 23348 3043
rect 23296 3000 23348 3009
rect 23480 3043 23532 3052
rect 23480 3009 23489 3043
rect 23489 3009 23523 3043
rect 23523 3009 23532 3043
rect 23480 3000 23532 3009
rect 24032 3000 24084 3052
rect 25320 3136 25372 3188
rect 25872 3136 25924 3188
rect 26700 3136 26752 3188
rect 26516 3068 26568 3120
rect 27344 3068 27396 3120
rect 22284 2864 22336 2916
rect 22560 2932 22612 2984
rect 23572 2932 23624 2984
rect 24676 2975 24728 2984
rect 24676 2941 24685 2975
rect 24685 2941 24719 2975
rect 24719 2941 24728 2975
rect 24676 2932 24728 2941
rect 26332 3043 26384 3052
rect 26332 3009 26341 3043
rect 26341 3009 26375 3043
rect 26375 3009 26384 3043
rect 29092 3136 29144 3188
rect 29184 3179 29236 3188
rect 29184 3145 29193 3179
rect 29193 3145 29227 3179
rect 29227 3145 29236 3179
rect 29184 3136 29236 3145
rect 29460 3179 29512 3188
rect 29460 3145 29469 3179
rect 29469 3145 29503 3179
rect 29503 3145 29512 3179
rect 29460 3136 29512 3145
rect 29828 3136 29880 3188
rect 30288 3136 30340 3188
rect 32496 3136 32548 3188
rect 34612 3179 34664 3188
rect 34612 3145 34621 3179
rect 34621 3145 34655 3179
rect 34655 3145 34664 3179
rect 34612 3136 34664 3145
rect 35900 3136 35952 3188
rect 35164 3068 35216 3120
rect 35348 3068 35400 3120
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 26332 3000 26384 3009
rect 29276 3043 29328 3052
rect 29276 3009 29285 3043
rect 29285 3009 29319 3043
rect 29319 3009 29328 3043
rect 29276 3000 29328 3009
rect 27712 2932 27764 2984
rect 30564 3043 30616 3052
rect 30564 3009 30573 3043
rect 30573 3009 30607 3043
rect 30607 3009 30616 3043
rect 30564 3000 30616 3009
rect 31760 3000 31812 3052
rect 31852 2932 31904 2984
rect 34152 3000 34204 3052
rect 35256 2932 35308 2984
rect 38476 3043 38528 3052
rect 38476 3009 38485 3043
rect 38485 3009 38519 3043
rect 38519 3009 38528 3043
rect 38476 3000 38528 3009
rect 38844 3043 38896 3052
rect 38844 3009 38853 3043
rect 38853 3009 38887 3043
rect 38887 3009 38896 3043
rect 38844 3000 38896 3009
rect 38936 3000 38988 3052
rect 23480 2864 23532 2916
rect 25044 2864 25096 2916
rect 34520 2864 34572 2916
rect 22376 2796 22428 2848
rect 22560 2839 22612 2848
rect 22560 2805 22569 2839
rect 22569 2805 22603 2839
rect 22603 2805 22612 2839
rect 22560 2796 22612 2805
rect 23020 2796 23072 2848
rect 26884 2796 26936 2848
rect 40132 2864 40184 2916
rect 38660 2839 38712 2848
rect 38660 2805 38669 2839
rect 38669 2805 38703 2839
rect 38703 2805 38712 2839
rect 38660 2796 38712 2805
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 1308 2388 1360 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4528 2388 4580 2440
rect 22560 2592 22612 2644
rect 39396 2635 39448 2644
rect 39396 2601 39405 2635
rect 39405 2601 39439 2635
rect 39439 2601 39448 2635
rect 39396 2592 39448 2601
rect 7564 2524 7616 2576
rect 23480 2524 23532 2576
rect 30748 2524 30800 2576
rect 38568 2524 38620 2576
rect 6368 2456 6420 2508
rect 2780 2252 2832 2304
rect 4252 2252 4304 2304
rect 5724 2252 5776 2304
rect 9404 2388 9456 2440
rect 11612 2388 11664 2440
rect 37004 2456 37056 2508
rect 38476 2431 38528 2440
rect 38476 2397 38485 2431
rect 38485 2397 38519 2431
rect 38519 2397 38528 2431
rect 38476 2388 38528 2397
rect 39672 2456 39724 2508
rect 39212 2431 39264 2440
rect 39212 2397 39221 2431
rect 39221 2397 39255 2431
rect 39255 2397 39264 2431
rect 39212 2388 39264 2397
rect 21456 2320 21508 2372
rect 6184 2252 6236 2304
rect 7196 2252 7248 2304
rect 8668 2252 8720 2304
rect 23848 2252 23900 2304
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2252 40000 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 1032 1980 1084 2032
rect 6184 1980 6236 2032
rect 11428 2048 11480 2100
rect 32312 2048 32364 2100
rect 30656 1980 30708 2032
rect 27896 1912 27948 1964
rect 1676 1844 1728 1896
rect 14372 1844 14424 1896
rect 3792 1776 3844 1828
rect 38476 1776 38528 1828
rect 23388 824 23440 876
rect 27712 824 27764 876
rect 20444 348 20496 400
rect 35256 348 35308 400
rect 18972 280 19024 332
rect 34796 280 34848 332
rect 16028 212 16080 264
rect 33416 212 33468 264
rect 11980 144 12032 196
rect 33692 144 33744 196
rect 14648 76 14700 128
rect 37372 76 37424 128
rect 10232 8 10284 60
rect 31760 8 31812 60
<< metal2 >>
rect 1860 11212 1912 11218
rect 3238 11194 3294 11250
rect 3514 11194 3570 11250
rect 3790 11194 3846 11250
rect 4066 11194 4122 11250
rect 4342 11194 4398 11250
rect 4618 11194 4674 11250
rect 4894 11194 4950 11250
rect 5170 11194 5226 11250
rect 5446 11194 5502 11250
rect 5722 11194 5778 11250
rect 5998 11194 6054 11250
rect 6274 11194 6330 11250
rect 6550 11194 6606 11250
rect 6826 11194 6882 11250
rect 7102 11194 7158 11250
rect 7378 11194 7434 11250
rect 7654 11194 7710 11250
rect 7930 11194 7986 11250
rect 8206 11194 8262 11250
rect 8482 11194 8538 11250
rect 8758 11194 8814 11250
rect 9034 11194 9090 11250
rect 9310 11194 9366 11250
rect 9586 11194 9642 11250
rect 9862 11194 9918 11250
rect 10138 11194 10194 11250
rect 10414 11194 10470 11250
rect 10690 11194 10746 11250
rect 10966 11194 11022 11250
rect 11242 11194 11298 11250
rect 11518 11194 11574 11250
rect 11794 11194 11850 11250
rect 12070 11194 12126 11250
rect 12346 11194 12402 11250
rect 12622 11194 12678 11250
rect 12898 11194 12954 11250
rect 13174 11194 13230 11250
rect 13450 11194 13506 11250
rect 13726 11194 13782 11250
rect 14002 11194 14058 11250
rect 14278 11194 14334 11250
rect 14554 11194 14610 11250
rect 14830 11194 14886 11250
rect 15106 11194 15162 11250
rect 15382 11194 15438 11250
rect 15658 11194 15714 11250
rect 15934 11194 15990 11250
rect 16210 11194 16266 11250
rect 16486 11194 16542 11250
rect 16762 11194 16818 11250
rect 17038 11194 17094 11250
rect 17314 11194 17370 11250
rect 17590 11194 17646 11250
rect 17866 11194 17922 11250
rect 18142 11194 18198 11250
rect 18418 11194 18474 11250
rect 18694 11194 18750 11250
rect 18970 11194 19026 11250
rect 19246 11194 19302 11250
rect 19522 11194 19578 11250
rect 19798 11194 19854 11250
rect 20074 11194 20130 11250
rect 20350 11194 20406 11250
rect 20626 11194 20682 11250
rect 20902 11194 20958 11250
rect 21178 11194 21234 11250
rect 21454 11194 21510 11250
rect 21730 11194 21786 11250
rect 22006 11194 22062 11250
rect 22282 11194 22338 11250
rect 22558 11194 22614 11250
rect 22834 11194 22890 11250
rect 23110 11194 23166 11250
rect 23386 11194 23442 11250
rect 23662 11194 23718 11250
rect 23938 11194 23994 11250
rect 24214 11194 24270 11250
rect 24490 11194 24546 11250
rect 24766 11194 24822 11250
rect 25042 11194 25098 11250
rect 25318 11194 25374 11250
rect 25594 11212 25650 11250
rect 25594 11194 25596 11212
rect 1860 11154 1912 11160
rect 1030 9616 1086 9625
rect 1030 9551 1086 9560
rect 662 9344 718 9353
rect 662 9279 718 9288
rect 294 9208 350 9217
rect 294 9143 350 9152
rect 204 6316 256 6322
rect 204 6258 256 6264
rect 216 6089 244 6258
rect 202 6080 258 6089
rect 202 6015 258 6024
rect 308 3913 336 9143
rect 478 8936 534 8945
rect 478 8871 534 8880
rect 388 8424 440 8430
rect 388 8366 440 8372
rect 400 7993 428 8366
rect 386 7984 442 7993
rect 386 7919 442 7928
rect 388 4548 440 4554
rect 388 4490 440 4496
rect 294 3904 350 3913
rect 294 3839 350 3848
rect 400 2553 428 4490
rect 492 3641 520 8871
rect 572 8356 624 8362
rect 572 8298 624 8304
rect 584 4729 612 8298
rect 676 7342 704 9279
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 756 7880 808 7886
rect 756 7822 808 7828
rect 768 7721 796 7822
rect 848 7812 900 7818
rect 848 7754 900 7760
rect 754 7712 810 7721
rect 754 7647 810 7656
rect 860 7449 888 7754
rect 952 7478 980 8735
rect 1044 8022 1072 9551
rect 1490 9480 1546 9489
rect 1490 9415 1546 9424
rect 1122 9072 1178 9081
rect 1122 9007 1178 9016
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1032 8016 1084 8022
rect 1032 7958 1084 7964
rect 1136 7954 1164 9007
rect 1308 8560 1360 8566
rect 1306 8528 1308 8537
rect 1360 8528 1362 8537
rect 1216 8492 1268 8498
rect 1306 8463 1362 8472
rect 1216 8434 1268 8440
rect 1228 8265 1256 8434
rect 1412 8378 1440 9007
rect 1320 8350 1440 8378
rect 1504 8362 1532 9415
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1492 8356 1544 8362
rect 1214 8256 1270 8265
rect 1214 8191 1270 8200
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 940 7472 992 7478
rect 846 7440 902 7449
rect 756 7404 808 7410
rect 940 7414 992 7420
rect 846 7375 902 7384
rect 756 7346 808 7352
rect 664 7336 716 7342
rect 664 7278 716 7284
rect 768 7177 796 7346
rect 754 7168 810 7177
rect 754 7103 810 7112
rect 1124 6996 1176 7002
rect 1124 6938 1176 6944
rect 754 6896 810 6905
rect 754 6831 810 6840
rect 1032 6860 1084 6866
rect 768 6798 796 6831
rect 1032 6802 1084 6808
rect 756 6792 808 6798
rect 756 6734 808 6740
rect 848 6724 900 6730
rect 848 6666 900 6672
rect 860 6633 888 6666
rect 846 6624 902 6633
rect 846 6559 902 6568
rect 1044 6361 1072 6802
rect 1030 6352 1086 6361
rect 1030 6287 1086 6296
rect 848 6248 900 6254
rect 848 6190 900 6196
rect 860 5817 888 6190
rect 846 5808 902 5817
rect 846 5743 902 5752
rect 756 5704 808 5710
rect 756 5646 808 5652
rect 768 5545 796 5646
rect 848 5636 900 5642
rect 848 5578 900 5584
rect 754 5536 810 5545
rect 754 5471 810 5480
rect 860 5273 888 5578
rect 846 5264 902 5273
rect 756 5228 808 5234
rect 846 5199 902 5208
rect 756 5170 808 5176
rect 768 5001 796 5170
rect 754 4992 810 5001
rect 754 4927 810 4936
rect 570 4720 626 4729
rect 570 4655 626 4664
rect 478 3632 534 3641
rect 478 3567 534 3576
rect 1030 3360 1086 3369
rect 1030 3295 1086 3304
rect 386 2544 442 2553
rect 386 2479 442 2488
rect 1044 2038 1072 3295
rect 1032 2032 1084 2038
rect 1136 2009 1164 6938
rect 1320 4457 1348 8350
rect 1492 8298 1544 8304
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1596 7313 1624 7686
rect 1582 7304 1638 7313
rect 1582 7239 1638 7248
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5914 1624 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1688 5302 1716 8366
rect 1872 7886 1900 11154
rect 2778 9888 2834 9897
rect 2504 9852 2556 9858
rect 2778 9823 2834 9832
rect 2504 9794 2556 9800
rect 2516 8634 2544 9794
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2792 7886 2820 9823
rect 3252 9466 3280 11194
rect 3252 9438 3464 9466
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8634 2912 8774
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3330 8528 3386 8537
rect 3330 8463 3386 8472
rect 3344 8090 3372 8463
rect 3436 8090 3464 9438
rect 3528 8362 3556 11194
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3620 8498 3648 9046
rect 3804 8634 3832 11194
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 4080 8090 4108 11194
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2424 7478 2452 7686
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2700 7002 2728 7686
rect 2884 7342 2912 7754
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 6390 2636 6598
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2778 6216 2834 6225
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2516 5914 2544 6190
rect 2688 6180 2740 6186
rect 2778 6151 2780 6160
rect 2688 6122 2740 6128
rect 2832 6151 2834 6160
rect 2780 6122 2832 6128
rect 2700 6066 2728 6122
rect 2700 6038 2820 6066
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 2792 5098 2820 6038
rect 3148 5704 3200 5710
rect 3146 5672 3148 5681
rect 3200 5672 3202 5681
rect 3146 5607 3202 5616
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 3620 4593 3648 7822
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3896 6361 3924 7210
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6662 4016 7142
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3882 6352 3938 6361
rect 3882 6287 3938 6296
rect 4172 5574 4200 9318
rect 4356 8634 4384 11194
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4540 8498 4568 8910
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4632 8090 4660 11194
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4724 8498 4752 9114
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4816 8430 4844 9386
rect 4908 8634 4936 11194
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5092 8498 5120 9454
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 5184 8090 5212 11194
rect 5356 8492 5408 8498
rect 5460 8480 5488 11194
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5644 8498 5672 9590
rect 5408 8452 5488 8480
rect 5632 8492 5684 8498
rect 5356 8434 5408 8440
rect 5632 8434 5684 8440
rect 5736 8362 5764 11194
rect 5908 8628 5960 8634
rect 6012 8616 6040 11194
rect 6184 9308 6236 9314
rect 6184 9250 6236 9256
rect 6092 9240 6144 9246
rect 6092 9182 6144 9188
rect 5960 8588 6040 8616
rect 5908 8570 5960 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5828 8401 5856 8434
rect 5814 8392 5870 8401
rect 5724 8356 5776 8362
rect 5814 8327 5870 8336
rect 5724 8298 5776 8304
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 3606 4584 3662 4593
rect 3516 4548 3568 4554
rect 3606 4519 3662 4528
rect 3516 4490 3568 4496
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 1216 4208 1268 4214
rect 1216 4150 1268 4156
rect 1032 1974 1084 1980
rect 1122 2000 1178 2009
rect 1122 1935 1178 1944
rect 1228 1465 1256 4150
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3528 3097 3556 4490
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1214 1456 1270 1465
rect 1214 1391 1270 1400
rect 1320 56 1348 2382
rect 1688 1902 1716 2382
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 1676 1896 1728 1902
rect 1676 1838 1728 1844
rect 2792 56 2820 2246
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3804 1834 3832 3946
rect 4448 3670 4476 7822
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5092 5778 5120 6190
rect 5262 5808 5318 5817
rect 5080 5772 5132 5778
rect 5262 5743 5264 5752
rect 5080 5714 5132 5720
rect 5316 5743 5318 5752
rect 5264 5714 5316 5720
rect 5092 4690 5120 5714
rect 5276 4690 5304 5714
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4540 2446 4568 4422
rect 5368 2990 5396 6734
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5460 4146 5488 6394
rect 5552 6390 5580 7482
rect 5828 7342 5856 7686
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5920 6934 5948 7754
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5644 5846 5672 6394
rect 6104 6236 6132 9182
rect 6012 6208 6132 6236
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5828 5166 5856 6054
rect 6012 5710 6040 6208
rect 6196 6118 6224 9250
rect 6288 8634 6316 11194
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6564 8090 6592 11194
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6748 7857 6776 8774
rect 6840 8634 6868 11194
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 7116 8090 7144 11194
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 6920 7880 6972 7886
rect 6734 7848 6790 7857
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6460 7812 6512 7818
rect 6920 7822 6972 7828
rect 6734 7783 6790 7792
rect 6460 7754 6512 7760
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6288 5794 6316 7754
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6196 5766 6316 5794
rect 6000 5704 6052 5710
rect 5998 5672 6000 5681
rect 6092 5704 6144 5710
rect 6052 5672 6054 5681
rect 6092 5646 6144 5652
rect 5998 5607 6054 5616
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4690 5856 5102
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5736 4282 5764 4626
rect 6012 4622 6040 5607
rect 6104 5574 6132 5646
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6104 5234 6132 5510
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6104 4622 6132 5170
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3534 5488 4082
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5814 3496 5870 3505
rect 5920 3466 5948 3878
rect 5814 3431 5816 3440
rect 5868 3431 5870 3440
rect 5908 3460 5960 3466
rect 5816 3402 5868 3408
rect 5908 3402 5960 3408
rect 5356 2984 5408 2990
rect 6196 2961 6224 5766
rect 6276 5704 6328 5710
rect 6274 5672 6276 5681
rect 6328 5672 6330 5681
rect 6274 5607 6330 5616
rect 5356 2926 5408 2932
rect 6182 2952 6238 2961
rect 6182 2887 6238 2896
rect 6380 2514 6408 7686
rect 6472 2553 6500 7754
rect 6932 7274 6960 7822
rect 7300 7449 7328 8910
rect 7392 8634 7420 11194
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8634 7604 8774
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6564 5817 6592 6258
rect 6840 5914 6868 6734
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6736 5840 6788 5846
rect 6550 5808 6606 5817
rect 6736 5782 6788 5788
rect 6550 5743 6606 5752
rect 6748 5574 6776 5782
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6840 3466 6868 5850
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4826 7236 4966
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7300 4078 7328 7142
rect 7484 6905 7512 7822
rect 7470 6896 7526 6905
rect 7470 6831 7526 6840
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4690 7512 4966
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 7576 2582 7604 8434
rect 7668 8090 7696 11194
rect 7944 8362 7972 11194
rect 8022 9752 8078 9761
rect 8022 9687 8078 9696
rect 8036 8498 8064 9687
rect 8116 8628 8168 8634
rect 8220 8616 8248 11194
rect 8390 11112 8446 11121
rect 8390 11047 8446 11056
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8168 8588 8248 8616
rect 8116 8570 8168 8576
rect 8312 8566 8340 8774
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7654 7984 7710 7993
rect 7654 7919 7710 7928
rect 7668 4185 7696 7919
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8036 7750 8064 7822
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7760 6798 7788 7346
rect 7852 7313 7880 7482
rect 7838 7304 7894 7313
rect 7838 7239 7894 7248
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7852 5817 7880 7142
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8312 6118 8340 8298
rect 8404 7410 8432 11047
rect 8496 8634 8524 11194
rect 8666 9208 8722 9217
rect 8576 9172 8628 9178
rect 8666 9143 8722 9152
rect 8576 9114 8628 9120
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8496 6984 8524 7822
rect 8588 7274 8616 9114
rect 8680 7886 8708 9143
rect 8772 8294 8800 11194
rect 9048 8820 9076 11194
rect 8864 8792 9076 8820
rect 9324 8820 9352 11194
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9324 8792 9444 8820
rect 8864 8634 8892 8792
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8942 8528 8998 8537
rect 8852 8492 8904 8498
rect 8942 8463 8998 8472
rect 8852 8434 8904 8440
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8772 7732 8800 8026
rect 8680 7704 8800 7732
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8496 6956 8616 6984
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7838 5808 7894 5817
rect 7838 5743 7894 5752
rect 8404 5234 8432 6598
rect 8496 6322 8524 6802
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8312 4690 8340 4966
rect 8404 4758 8432 5170
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8496 4622 8524 5170
rect 8484 4616 8536 4622
rect 8298 4584 8354 4593
rect 8208 4548 8260 4554
rect 8484 4558 8536 4564
rect 8298 4519 8354 4528
rect 8208 4490 8260 4496
rect 8220 4282 8248 4490
rect 8312 4282 8340 4519
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 7654 4176 7710 4185
rect 7654 4111 7710 4120
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 8588 2961 8616 6956
rect 8680 3641 8708 7704
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8772 4690 8800 5170
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8772 4214 8800 4626
rect 8864 4593 8892 8434
rect 8956 7818 8984 8463
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8090 9076 8230
rect 9416 8090 9444 8792
rect 9508 8498 9536 9658
rect 9600 8634 9628 11194
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9876 8090 9904 11194
rect 10048 9784 10100 9790
rect 10048 9726 10100 9732
rect 10060 8498 10088 9726
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10152 8362 10180 11194
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8498 10272 8842
rect 10428 8634 10456 11194
rect 10508 9308 10560 9314
rect 10508 9250 10560 9256
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10520 8498 10548 9250
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10612 8537 10640 9046
rect 10704 8634 10732 11194
rect 10980 8634 11008 11194
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10598 8528 10654 8537
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10508 8492 10560 8498
rect 10598 8463 10654 8472
rect 10508 8434 10560 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9128 8016 9180 8022
rect 9126 7984 9128 7993
rect 9180 7984 9182 7993
rect 9126 7919 9182 7928
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9416 6497 9444 7822
rect 9692 7002 9720 7822
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6934 9812 7210
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9402 6488 9458 6497
rect 9402 6423 9458 6432
rect 9404 6384 9456 6390
rect 9456 6344 9536 6372
rect 9404 6326 9456 6332
rect 9220 6180 9272 6186
rect 9220 6122 9272 6128
rect 9128 6112 9180 6118
rect 9232 6089 9260 6122
rect 9128 6054 9180 6060
rect 9218 6080 9274 6089
rect 9140 5556 9168 6054
rect 9218 6015 9274 6024
rect 9140 5528 9444 5556
rect 9508 5545 9536 6344
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5710 9720 6054
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 8850 4584 8906 4593
rect 8850 4519 8906 4528
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8666 3632 8722 3641
rect 8666 3567 8722 3576
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 8574 2952 8630 2961
rect 8574 2887 8630 2896
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7564 2576 7616 2582
rect 6458 2544 6514 2553
rect 6368 2508 6420 2514
rect 7564 2518 7616 2524
rect 6458 2479 6514 2488
rect 6368 2450 6420 2456
rect 9416 2446 9444 5528
rect 9494 5536 9550 5545
rect 9494 5471 9550 5480
rect 9968 3942 9996 6870
rect 10060 4010 10088 7686
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 6322 10180 7142
rect 10244 7002 10272 7822
rect 10336 7818 10364 8434
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10784 8016 10836 8022
rect 11072 7993 11100 8366
rect 10784 7958 10836 7964
rect 11058 7984 11114 7993
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10152 5846 10180 6258
rect 10704 5846 10732 6326
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10140 5704 10192 5710
rect 10138 5672 10140 5681
rect 10192 5672 10194 5681
rect 10138 5607 10194 5616
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4146 10272 5102
rect 10336 4826 10364 5578
rect 10428 5114 10456 5578
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 5234 10640 5510
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10428 5086 10548 5114
rect 10520 5030 10548 5086
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10428 4826 10456 4966
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10612 4690 10640 5170
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4214 10548 4422
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10612 4146 10640 4490
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10796 4049 10824 7958
rect 10876 7948 10928 7954
rect 11058 7919 11114 7928
rect 10876 7890 10928 7896
rect 10888 7478 10916 7890
rect 10876 7472 10928 7478
rect 11164 7449 11192 8774
rect 11256 8090 11284 11194
rect 11532 8634 11560 11194
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11348 8294 11376 8434
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11808 8090 11836 11194
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 10876 7414 10928 7420
rect 11150 7440 11206 7449
rect 11150 7375 11206 7384
rect 10874 7304 10930 7313
rect 10874 7239 10876 7248
rect 10928 7239 10930 7248
rect 10876 7210 10928 7216
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 5778 11008 6598
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4282 10916 4558
rect 10980 4554 11008 5170
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10782 4040 10838 4049
rect 10048 4004 10100 4010
rect 10782 3975 10838 3984
rect 10048 3946 10100 3952
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 3792 1828 3844 1834
rect 3792 1770 3844 1776
rect 4264 56 4292 2246
rect 5736 56 5764 2246
rect 6196 2038 6224 2246
rect 6184 2032 6236 2038
rect 6184 1974 6236 1980
rect 7208 56 7236 2246
rect 8680 56 8708 2246
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 11440 2106 11468 6870
rect 11532 6798 11560 6870
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11716 6730 11744 6802
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11624 5710 11652 6666
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11532 5098 11560 5646
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4282 11560 5034
rect 11992 4486 12020 9454
rect 12084 8634 12112 11194
rect 12164 9308 12216 9314
rect 12164 9250 12216 9256
rect 12176 9042 12204 9250
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12360 8634 12388 11194
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12636 8090 12664 11194
rect 12912 8634 12940 11194
rect 13188 8634 13216 11194
rect 13268 9240 13320 9246
rect 13268 9182 13320 9188
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13280 8566 13308 9182
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13372 8498 13400 9114
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 12728 8362 12756 8434
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7478 12204 7822
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 12452 6866 12480 7210
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12636 6798 12664 7754
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12714 6760 12770 6769
rect 12714 6695 12770 6704
rect 12728 6662 12756 6695
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12268 4622 12296 5102
rect 12820 5098 12848 8434
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12912 7750 12940 7958
rect 13464 7818 13492 11194
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 8974 13676 9318
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13636 8628 13688 8634
rect 13740 8616 13768 11194
rect 13820 9308 13872 9314
rect 13820 9250 13872 9256
rect 13688 8588 13768 8616
rect 13636 8570 13688 8576
rect 13832 8566 13860 9250
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13924 8498 13952 8910
rect 14016 8634 14044 11194
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13464 6458 13492 7346
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13464 5846 13492 6122
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13556 5273 13584 8434
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13648 7426 13676 8298
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 8090 14320 11194
rect 14568 8634 14596 11194
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14370 8120 14426 8129
rect 14280 8084 14332 8090
rect 14370 8055 14426 8064
rect 14280 8026 14332 8032
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13740 7857 13768 7958
rect 14188 7880 14240 7886
rect 13726 7848 13782 7857
rect 14240 7840 14320 7868
rect 14188 7822 14240 7828
rect 13726 7783 13782 7792
rect 13648 7398 13860 7426
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13542 5264 13598 5273
rect 13542 5199 13598 5208
rect 13648 5137 13676 7142
rect 13740 6866 13768 7278
rect 13832 6866 13860 7398
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13740 6662 13768 6802
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 5778 13768 6598
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13832 6089 13860 6258
rect 13818 6080 13874 6089
rect 13818 6015 13874 6024
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13728 5772 13780 5778
rect 13780 5732 13860 5760
rect 13728 5714 13780 5720
rect 13726 5672 13782 5681
rect 13726 5607 13728 5616
rect 13780 5607 13782 5616
rect 13728 5578 13780 5584
rect 13634 5128 13690 5137
rect 12808 5092 12860 5098
rect 13634 5063 13690 5072
rect 12808 5034 12860 5040
rect 13636 4752 13688 4758
rect 13634 4720 13636 4729
rect 13688 4720 13690 4729
rect 13832 4690 13860 5732
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13634 4655 13690 4664
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 10152 66 10272 82
rect 10152 60 10284 66
rect 10152 56 10232 60
rect 1306 0 1362 56
rect 2778 0 2834 56
rect 4250 0 4306 56
rect 5722 0 5778 56
rect 7194 0 7250 56
rect 8666 0 8722 56
rect 10138 54 10232 56
rect 10138 0 10194 54
rect 11624 56 11652 2382
rect 11992 202 12020 3470
rect 14292 3398 14320 7840
rect 14384 7721 14412 8055
rect 14370 7712 14426 7721
rect 14370 7647 14426 7656
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14384 4146 14412 5578
rect 14476 4622 14504 8434
rect 14660 8294 14688 8842
rect 14556 8288 14608 8294
rect 14554 8256 14556 8265
rect 14648 8288 14700 8294
rect 14608 8256 14610 8265
rect 14648 8230 14700 8236
rect 14554 8191 14610 8200
rect 14844 8090 14872 11194
rect 15120 9602 15148 11194
rect 14936 9574 15148 9602
rect 14936 8634 14964 9574
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 11194
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14648 7880 14700 7886
rect 14646 7848 14648 7857
rect 14700 7848 14702 7857
rect 14646 7783 14702 7792
rect 15028 7732 15056 8570
rect 15488 8090 15516 9386
rect 15672 8634 15700 11194
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15764 8498 15792 8774
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15948 8090 15976 11194
rect 16120 8900 16172 8906
rect 16120 8842 16172 8848
rect 16132 8498 16160 8842
rect 16224 8634 16252 11194
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16408 8537 16436 9590
rect 16500 8634 16528 11194
rect 16776 8634 16804 11194
rect 17052 9314 17080 11194
rect 17040 9308 17092 9314
rect 17040 9250 17092 9256
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16210 8528 16266 8537
rect 16120 8492 16172 8498
rect 16210 8463 16266 8472
rect 16394 8528 16450 8537
rect 17328 8498 17356 11194
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 16394 8463 16450 8472
rect 17316 8492 17368 8498
rect 16120 8434 16172 8440
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 14936 7704 15056 7732
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14844 6254 14872 6598
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14568 5710 14596 5850
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14554 5536 14610 5545
rect 14554 5471 14610 5480
rect 14568 4865 14596 5471
rect 14936 5370 14964 7704
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15396 7426 15424 7822
rect 15488 7546 15516 7822
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15580 7585 15608 7686
rect 15566 7576 15622 7585
rect 15476 7540 15528 7546
rect 15566 7511 15622 7520
rect 15476 7482 15528 7488
rect 15292 7404 15344 7410
rect 15396 7398 15516 7426
rect 15292 7346 15344 7352
rect 15304 7177 15332 7346
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15290 7168 15346 7177
rect 15290 7103 15346 7112
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15016 6384 15068 6390
rect 15014 6352 15016 6361
rect 15068 6352 15070 6361
rect 15120 6338 15148 6394
rect 15198 6352 15254 6361
rect 15120 6310 15198 6338
rect 15014 6287 15070 6296
rect 15198 6287 15254 6296
rect 15396 5642 15424 7278
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14554 4856 14610 4865
rect 14554 4791 14610 4800
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 12176 2961 12204 3334
rect 12162 2952 12218 2961
rect 12162 2887 12218 2896
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13082 2000 13138 2009
rect 13082 1935 13138 1944
rect 11980 196 12032 202
rect 11980 138 12032 144
rect 13096 56 13124 1935
rect 14384 1902 14412 4082
rect 14476 4078 14504 4422
rect 14660 4282 14688 4966
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14752 4078 14780 4558
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 15396 4010 15424 4558
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15488 3534 15516 7398
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5778 15884 6054
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 16040 3738 16068 8366
rect 16224 6458 16252 8463
rect 17316 8434 17368 8440
rect 17222 8120 17278 8129
rect 17222 8055 17278 8064
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16316 7410 16344 7958
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16408 6497 16436 7822
rect 16672 7744 16724 7750
rect 17236 7721 17264 8055
rect 17512 7818 17540 9862
rect 17604 8090 17632 11194
rect 17684 9308 17736 9314
rect 17684 9250 17736 9256
rect 17696 8362 17724 9250
rect 17776 9240 17828 9246
rect 17776 9182 17828 9188
rect 17788 8566 17816 9182
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17788 8265 17816 8366
rect 17774 8256 17830 8265
rect 17774 8191 17830 8200
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17696 7750 17724 7822
rect 17684 7744 17736 7750
rect 16672 7686 16724 7692
rect 17222 7712 17278 7721
rect 16684 7342 16712 7686
rect 17684 7686 17736 7692
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17222 7647 17278 7656
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16500 7002 16528 7142
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16684 6662 16712 7278
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16394 6488 16450 6497
rect 16212 6452 16264 6458
rect 16394 6423 16450 6432
rect 16212 6394 16264 6400
rect 16396 4616 16448 4622
rect 16684 4604 16712 6598
rect 17696 6322 17724 7686
rect 17788 6662 17816 7686
rect 17880 7410 17908 11194
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 18064 8498 18092 9522
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17972 8362 18000 8434
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 18156 7410 18184 11194
rect 18432 8498 18460 11194
rect 18708 8498 18736 11194
rect 18984 8498 19012 11194
rect 19260 8498 19288 11194
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 18340 8350 18552 8378
rect 18340 7818 18368 8350
rect 18524 8294 18552 8350
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18144 7200 18196 7206
rect 18340 7177 18368 7754
rect 18432 7290 18460 8230
rect 18432 7262 18552 7290
rect 18524 7206 18552 7262
rect 18420 7200 18472 7206
rect 18144 7142 18196 7148
rect 18326 7168 18382 7177
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 16960 5914 16988 6258
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 16448 4576 16712 4604
rect 16396 4558 16448 4564
rect 16684 4146 16712 4576
rect 17420 4554 17448 5578
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17972 4826 18000 5199
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 18156 4622 18184 7142
rect 18420 7142 18472 7148
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18326 7103 18382 7112
rect 18432 5574 18460 7142
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18616 5030 18644 8230
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18878 4856 18934 4865
rect 19076 4826 19104 5034
rect 18878 4791 18934 4800
rect 19064 4820 19116 4826
rect 18892 4622 18920 4791
rect 19064 4762 19116 4768
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17236 4146 17264 4218
rect 17512 4146 17540 4422
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 16592 3126 16620 3878
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16684 3058 16712 3402
rect 16960 3194 16988 4014
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16684 2922 16712 2994
rect 17236 2990 17264 4082
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17696 3670 17724 3878
rect 17684 3664 17736 3670
rect 17684 3606 17736 3612
rect 18800 3516 18828 4558
rect 19168 3942 19196 8230
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5846 19288 6054
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19352 4826 19380 8298
rect 19444 6186 19472 8774
rect 19536 8498 19564 11194
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19536 8090 19564 8230
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19536 7274 19564 7822
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19628 5574 19656 8570
rect 19812 8498 19840 11194
rect 20088 9217 20116 11194
rect 20364 11121 20392 11194
rect 20350 11112 20406 11121
rect 20350 11047 20406 11056
rect 20640 9926 20668 11194
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20074 9208 20130 9217
rect 20074 9143 20130 9152
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 20732 8430 20760 8842
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20536 8288 20588 8294
rect 20640 8265 20668 8366
rect 20916 8294 20944 11194
rect 21192 9874 21220 11194
rect 21192 9846 21404 9874
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21192 9217 21220 9318
rect 21178 9208 21234 9217
rect 21178 9143 21234 9152
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21376 8498 21404 9846
rect 21468 8498 21496 11194
rect 21744 8566 21772 11194
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 20904 8288 20956 8294
rect 20536 8230 20588 8236
rect 20626 8256 20682 8265
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7750 19748 7822
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 6458 19748 7686
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19812 6390 19840 7958
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20350 7576 20406 7585
rect 20350 7511 20406 7520
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20364 7041 20392 7511
rect 20456 7410 20484 7822
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20350 7032 20406 7041
rect 20350 6967 20406 6976
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 20456 6322 20484 6394
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19444 4622 19472 5238
rect 20548 5166 20576 8230
rect 20904 8230 20956 8236
rect 20626 8191 20682 8200
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20640 7177 20668 8026
rect 20732 7818 20760 8026
rect 21008 7954 21036 8298
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 21100 7750 21128 7822
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20626 7168 20682 7177
rect 20626 7103 20682 7112
rect 20718 6488 20774 6497
rect 20628 6452 20680 6458
rect 20718 6423 20774 6432
rect 20628 6394 20680 6400
rect 20640 6322 20668 6394
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20640 5710 20668 6258
rect 20732 5953 20760 6423
rect 20916 6186 20944 7210
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20718 5944 20774 5953
rect 20718 5879 20774 5888
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 20810 5400 20866 5409
rect 21010 5403 21318 5412
rect 20810 5335 20866 5344
rect 20824 5166 20852 5335
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 21376 5030 21404 8298
rect 21652 7970 21680 8502
rect 22020 8430 22048 11194
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 22112 8362 22140 8774
rect 22296 8566 22324 11194
rect 22572 8634 22600 11194
rect 22652 9444 22704 9450
rect 22652 9386 22704 9392
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22284 8560 22336 8566
rect 22190 8528 22246 8537
rect 22480 8537 22508 8570
rect 22284 8502 22336 8508
rect 22466 8528 22522 8537
rect 22190 8463 22246 8472
rect 22466 8463 22522 8472
rect 22100 8356 22152 8362
rect 22100 8298 22152 8304
rect 22204 8022 22232 8463
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22192 8016 22244 8022
rect 21652 7942 21772 7970
rect 22192 7958 22244 7964
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 20812 5024 20864 5030
rect 20810 4992 20812 5001
rect 20904 5024 20956 5030
rect 20864 4992 20866 5001
rect 20904 4966 20956 4972
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 19950 4924 20258 4933
rect 20810 4927 20866 4936
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20916 4826 20944 4966
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19444 4282 19472 4558
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20272 4282 20300 4422
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 18880 3528 18932 3534
rect 18800 3488 18880 3516
rect 18880 3470 18932 3476
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19352 3194 19380 3402
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19444 2990 19472 4218
rect 20272 4026 20300 4218
rect 20272 3998 20392 4026
rect 19950 3836 20258 3845
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20364 3534 20392 3998
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 21376 3602 21404 3946
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 20180 3194 20208 3334
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20456 3126 20484 3538
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 20444 3120 20496 3126
rect 20444 3062 20496 3068
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 20456 2825 20484 3062
rect 20442 2816 20498 2825
rect 19950 2748 20258 2757
rect 20442 2751 20498 2760
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 21468 2378 21496 7686
rect 21546 7576 21602 7585
rect 21652 7546 21680 7822
rect 21546 7511 21602 7520
rect 21640 7540 21692 7546
rect 21560 6458 21588 7511
rect 21640 7482 21692 7488
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21546 5264 21602 5273
rect 21546 5199 21602 5208
rect 21560 5166 21588 5199
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21548 5024 21600 5030
rect 21546 4992 21548 5001
rect 21600 4992 21602 5001
rect 21546 4927 21602 4936
rect 21744 4486 21772 7942
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21836 7274 21864 7754
rect 22296 7750 22324 8230
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21836 6458 21864 6734
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21928 6202 21956 6598
rect 22112 6458 22140 6802
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 21928 6174 22048 6202
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 21928 5778 21956 6054
rect 22020 5778 22048 6174
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 22020 4690 22048 5102
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 21824 4616 21876 4622
rect 21876 4576 21956 4604
rect 21824 4558 21876 4564
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21732 4480 21784 4486
rect 21732 4422 21784 4428
rect 21560 4010 21588 4422
rect 21928 4282 21956 4576
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21928 3058 21956 4218
rect 22388 4214 22416 8230
rect 22480 8022 22508 8230
rect 22468 8016 22520 8022
rect 22468 7958 22520 7964
rect 22664 4690 22692 9386
rect 22848 8566 22876 11194
rect 23124 9654 23152 11194
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23018 9208 23074 9217
rect 23018 9143 23074 9152
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 22192 3392 22244 3398
rect 22192 3334 22244 3340
rect 22006 3224 22062 3233
rect 22006 3159 22008 3168
rect 22060 3159 22062 3168
rect 22008 3130 22060 3136
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 22204 2990 22232 3334
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 22296 2666 22324 2858
rect 22388 2854 22416 3470
rect 22940 3058 22968 3946
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 22560 2984 22612 2990
rect 22480 2944 22560 2972
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22480 2666 22508 2944
rect 22560 2926 22612 2932
rect 23032 2854 23060 9143
rect 23400 8566 23428 11194
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23492 8498 23520 9590
rect 23676 8634 23704 11194
rect 23952 9874 23980 11194
rect 23952 9846 24164 9874
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23202 8392 23258 8401
rect 23308 8362 23520 8378
rect 23202 8327 23258 8336
rect 23296 8356 23520 8362
rect 23216 7342 23244 8327
rect 23348 8350 23520 8356
rect 23296 8298 23348 8304
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 7886 23428 8230
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23112 7336 23164 7342
rect 23112 7278 23164 7284
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23124 4826 23152 7278
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23308 5710 23336 6598
rect 23388 6384 23440 6390
rect 23388 6326 23440 6332
rect 23400 5914 23428 6326
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23400 4826 23428 4966
rect 23112 4820 23164 4826
rect 23112 4762 23164 4768
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23308 3398 23336 4694
rect 23492 4026 23520 8350
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23584 4622 23612 8298
rect 23664 8288 23716 8294
rect 23716 8248 23796 8276
rect 23664 8230 23716 8236
rect 23768 5234 23796 8248
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7449 23888 7686
rect 23846 7440 23902 7449
rect 23846 7375 23902 7384
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 23860 5574 23888 6734
rect 23952 6322 23980 8298
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23492 3998 23612 4026
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23308 3058 23336 3334
rect 23492 3058 23520 3878
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23480 3052 23532 3058
rect 23480 2994 23532 3000
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 23020 2848 23072 2854
rect 23308 2825 23336 2994
rect 23584 2990 23612 3998
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23020 2790 23072 2796
rect 23294 2816 23350 2825
rect 22296 2638 22508 2666
rect 22572 2650 22600 2790
rect 23294 2751 23350 2760
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 23492 2582 23520 2858
rect 23952 2774 23980 5646
rect 24044 3058 24072 8774
rect 24136 8498 24164 9846
rect 24228 8566 24256 11194
rect 24504 10062 24532 11194
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24780 9874 24808 11194
rect 24584 9852 24636 9858
rect 24780 9846 24900 9874
rect 24584 9794 24636 9800
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24400 9308 24452 9314
rect 24400 9250 24452 9256
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24320 8412 24348 8774
rect 24228 8384 24348 8412
rect 24228 8294 24256 8384
rect 24216 8288 24268 8294
rect 24412 8242 24440 9250
rect 24216 8230 24268 8236
rect 24320 8214 24440 8242
rect 24320 6798 24348 8214
rect 24398 8120 24454 8129
rect 24398 8055 24400 8064
rect 24452 8055 24454 8064
rect 24400 8026 24452 8032
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24228 6118 24256 6258
rect 24216 6112 24268 6118
rect 24216 6054 24268 6060
rect 24320 5778 24348 6394
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24412 5846 24440 6054
rect 24400 5840 24452 5846
rect 24400 5782 24452 5788
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24136 5302 24164 5510
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24504 4282 24532 9522
rect 24596 6662 24624 9794
rect 24766 8936 24822 8945
rect 24766 8871 24822 8880
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24688 6730 24716 8298
rect 24780 7478 24808 8871
rect 24872 8634 24900 9846
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24964 8514 24992 8910
rect 24872 8486 24992 8514
rect 24768 7472 24820 7478
rect 24768 7414 24820 7420
rect 24766 7168 24822 7177
rect 24766 7103 24822 7112
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24596 5710 24624 6598
rect 24780 5710 24808 7103
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24872 5522 24900 8486
rect 25056 8430 25084 11194
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25148 8498 25176 9998
rect 25332 8566 25360 11194
rect 25648 11194 25650 11212
rect 25870 11194 25926 11250
rect 26146 11194 26202 11250
rect 26422 11194 26478 11250
rect 26698 11194 26754 11250
rect 26974 11194 27030 11250
rect 27250 11194 27306 11250
rect 27526 11194 27582 11250
rect 27802 11194 27858 11250
rect 28078 11194 28134 11250
rect 28354 11194 28410 11250
rect 28630 11194 28686 11250
rect 28906 11194 28962 11250
rect 29182 11194 29238 11250
rect 29458 11194 29514 11250
rect 29734 11194 29790 11250
rect 30010 11194 30066 11250
rect 30286 11194 30342 11250
rect 30562 11194 30618 11250
rect 30838 11194 30894 11250
rect 31114 11194 31170 11250
rect 31390 11194 31446 11250
rect 31666 11194 31722 11250
rect 31942 11194 31998 11250
rect 32218 11194 32274 11250
rect 32494 11194 32550 11250
rect 32770 11194 32826 11250
rect 33046 11194 33102 11250
rect 33322 11194 33378 11250
rect 33598 11194 33654 11250
rect 33874 11194 33930 11250
rect 34150 11194 34206 11250
rect 34426 11194 34482 11250
rect 34702 11194 34758 11250
rect 34978 11194 35034 11250
rect 35254 11194 35310 11250
rect 35530 11194 35586 11250
rect 35806 11194 35862 11250
rect 36082 11194 36138 11250
rect 36358 11194 36414 11250
rect 36634 11194 36690 11250
rect 36910 11194 36966 11250
rect 37186 11194 37242 11250
rect 37462 11194 37518 11250
rect 37738 11194 37794 11250
rect 25596 11154 25648 11160
rect 25686 9072 25742 9081
rect 25686 9007 25742 9016
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24952 8288 25004 8294
rect 24952 8230 25004 8236
rect 25134 8256 25190 8265
rect 24780 5494 24900 5522
rect 24780 5166 24808 5494
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 24872 4826 24900 5306
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24964 4570 24992 8230
rect 25134 8191 25190 8200
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25056 5302 25084 6598
rect 25148 5302 25176 8191
rect 25318 6896 25374 6905
rect 25318 6831 25374 6840
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25240 6662 25268 6734
rect 25332 6662 25360 6831
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25424 6254 25452 8570
rect 25502 7848 25558 7857
rect 25502 7783 25558 7792
rect 25516 7750 25544 7783
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25516 6798 25544 7346
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25608 6390 25636 8570
rect 25700 7546 25728 9007
rect 25884 8430 25912 11194
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25976 8634 26004 8910
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 26160 8276 26188 11194
rect 26436 10198 26464 11194
rect 26424 10192 26476 10198
rect 26424 10134 26476 10140
rect 26424 8560 26476 8566
rect 26424 8502 26476 8508
rect 25884 8248 26188 8276
rect 26332 8288 26384 8294
rect 25780 8016 25832 8022
rect 25780 7958 25832 7964
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25412 6248 25464 6254
rect 25412 6190 25464 6196
rect 25502 5944 25558 5953
rect 25502 5879 25558 5888
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 25136 5296 25188 5302
rect 25136 5238 25188 5244
rect 25056 4690 25084 5238
rect 25136 5160 25188 5166
rect 25136 5102 25188 5108
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24872 4554 24992 4570
rect 24860 4548 24992 4554
rect 24912 4542 24992 4548
rect 24860 4490 24912 4496
rect 24492 4276 24544 4282
rect 24492 4218 24544 4224
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24688 2990 24716 3334
rect 25042 3224 25098 3233
rect 25042 3159 25098 3168
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 25056 2922 25084 3159
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 23860 2746 23980 2774
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 23860 2310 23888 2746
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 14372 1896 14424 1902
rect 14372 1838 14424 1844
rect 23388 876 23440 882
rect 23388 818 23440 824
rect 20444 400 20496 406
rect 20444 342 20496 348
rect 18972 332 19024 338
rect 18972 274 19024 280
rect 16028 264 16080 270
rect 16028 206 16080 212
rect 14648 128 14700 134
rect 14568 76 14648 82
rect 14568 70 14700 76
rect 14568 56 14688 70
rect 16040 56 16068 206
rect 17498 96 17554 105
rect 10232 2 10284 8
rect 11610 0 11666 56
rect 13082 0 13138 56
rect 14554 54 14688 56
rect 14554 0 14610 54
rect 16026 0 16082 56
rect 18984 56 19012 274
rect 20456 56 20484 342
rect 21914 232 21970 241
rect 21914 167 21970 176
rect 21928 56 21956 167
rect 23400 56 23428 818
rect 24872 56 24992 82
rect 17498 0 17554 40
rect 18970 0 19026 56
rect 20442 0 20498 56
rect 21914 0 21970 56
rect 23386 0 23442 56
rect 24858 54 24992 56
rect 24858 0 24914 54
rect 24964 42 24992 54
rect 25148 42 25176 5102
rect 25516 5030 25544 5879
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25240 4146 25268 4558
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 25332 3194 25360 4422
rect 25700 4214 25728 7346
rect 25792 6186 25820 7958
rect 25884 7410 25912 8248
rect 26332 8230 26384 8236
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25964 6928 26016 6934
rect 25964 6870 26016 6876
rect 25976 6662 26004 6870
rect 25964 6656 26016 6662
rect 25964 6598 26016 6604
rect 25872 6384 25924 6390
rect 25872 6326 25924 6332
rect 25780 6180 25832 6186
rect 25780 6122 25832 6128
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25884 3194 25912 6326
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 25976 5234 26004 5646
rect 26160 5574 26188 5646
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 26344 4622 26372 8230
rect 26436 6322 26464 8502
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26528 8090 26556 8366
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26620 7585 26648 8230
rect 26606 7576 26662 7585
rect 26606 7511 26662 7520
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26528 5930 26556 7278
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26436 5902 26556 5930
rect 26436 5370 26464 5902
rect 26620 5710 26648 6598
rect 26712 6254 26740 11194
rect 26988 9674 27016 11194
rect 26896 9646 27016 9674
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 26620 5574 26648 5646
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 26620 4758 26648 5510
rect 26608 4752 26660 4758
rect 26608 4694 26660 4700
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26804 4554 26832 8774
rect 26896 6905 26924 9646
rect 27264 8922 27292 11194
rect 27264 8894 27384 8922
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26882 6896 26938 6905
rect 26882 6831 26938 6840
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27356 6186 27384 8894
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27448 7342 27476 8298
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27448 6866 27476 7278
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27344 6180 27396 6186
rect 27344 6122 27396 6128
rect 27448 5710 27476 6598
rect 27540 6322 27568 11194
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27528 6180 27580 6186
rect 27528 6122 27580 6128
rect 26884 5704 26936 5710
rect 27344 5704 27396 5710
rect 26936 5664 27344 5692
rect 26884 5646 26936 5652
rect 27344 5646 27396 5652
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 26792 4548 26844 4554
rect 26792 4490 26844 4496
rect 26896 4162 26924 5306
rect 27356 4690 27384 5646
rect 27434 5400 27490 5409
rect 27434 5335 27490 5344
rect 27448 5001 27476 5335
rect 27540 5302 27568 6122
rect 27528 5296 27580 5302
rect 27528 5238 27580 5244
rect 27434 4992 27490 5001
rect 27434 4927 27490 4936
rect 27528 4820 27580 4826
rect 27528 4762 27580 4768
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 27540 4622 27568 4762
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27436 4548 27488 4554
rect 27436 4490 27488 4496
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27448 4282 27476 4490
rect 27632 4486 27660 8298
rect 27724 6390 27752 8842
rect 27816 8498 27844 11194
rect 28092 9874 28120 11194
rect 28092 9846 28212 9874
rect 27894 8528 27950 8537
rect 27804 8492 27856 8498
rect 28184 8498 28212 9846
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 27894 8463 27950 8472
rect 28172 8492 28224 8498
rect 27804 8434 27856 8440
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27816 6633 27844 6734
rect 27908 6662 27936 8463
rect 28172 8434 28224 8440
rect 28276 7818 28304 9114
rect 28368 8498 28396 11194
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28460 7342 28488 7686
rect 28172 7336 28224 7342
rect 28172 7278 28224 7284
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 27988 6860 28040 6866
rect 27988 6802 28040 6808
rect 28000 6730 28028 6802
rect 28184 6798 28212 7278
rect 28356 7200 28408 7206
rect 28354 7168 28356 7177
rect 28448 7200 28500 7206
rect 28408 7168 28410 7177
rect 28448 7142 28500 7148
rect 28354 7103 28410 7112
rect 28460 6934 28488 7142
rect 28448 6928 28500 6934
rect 28262 6896 28318 6905
rect 28448 6870 28500 6876
rect 28262 6831 28318 6840
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 27988 6724 28040 6730
rect 27988 6666 28040 6672
rect 27896 6656 27948 6662
rect 27802 6624 27858 6633
rect 27896 6598 27948 6604
rect 27802 6559 27858 6568
rect 27908 6497 27936 6598
rect 27894 6488 27950 6497
rect 27894 6423 27950 6432
rect 27712 6384 27764 6390
rect 27712 6326 27764 6332
rect 27988 6384 28040 6390
rect 27988 6326 28040 6332
rect 27804 6180 27856 6186
rect 27804 6122 27856 6128
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 26804 4134 26924 4162
rect 27632 4146 27660 4422
rect 27620 4140 27672 4146
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 26608 3664 26660 3670
rect 26608 3606 26660 3612
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25872 3188 25924 3194
rect 25872 3130 25924 3136
rect 26528 3126 26556 3470
rect 26620 3210 26648 3606
rect 26620 3194 26740 3210
rect 26620 3188 26752 3194
rect 26620 3182 26700 3188
rect 26700 3130 26752 3136
rect 26516 3120 26568 3126
rect 26516 3062 26568 3068
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 26344 2009 26372 2994
rect 26804 2774 26832 4134
rect 27620 4082 27672 4088
rect 26884 4072 26936 4078
rect 26936 4020 27016 4026
rect 26884 4014 27016 4020
rect 26896 3998 27016 4014
rect 27724 4010 27752 4966
rect 27816 4185 27844 6122
rect 27896 5568 27948 5574
rect 27896 5510 27948 5516
rect 27802 4176 27858 4185
rect 27802 4111 27858 4120
rect 26988 3738 27016 3998
rect 27712 4004 27764 4010
rect 27712 3946 27764 3952
rect 26976 3732 27028 3738
rect 26976 3674 27028 3680
rect 27068 3664 27120 3670
rect 27068 3606 27120 3612
rect 27080 3466 27108 3606
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 26896 2854 26924 3334
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27356 3126 27384 3334
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27712 2984 27764 2990
rect 27712 2926 27764 2932
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 26712 2746 26832 2774
rect 26330 2000 26386 2009
rect 26330 1935 26386 1944
rect 26344 56 26464 82
rect 24964 14 25176 42
rect 26330 54 26464 56
rect 26330 0 26386 54
rect 26436 42 26464 54
rect 26712 42 26740 2746
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 27724 882 27752 2926
rect 27908 1970 27936 5510
rect 27896 1964 27948 1970
rect 27896 1906 27948 1912
rect 27712 876 27764 882
rect 27712 818 27764 824
rect 27816 56 27936 82
rect 26436 14 26740 42
rect 27802 54 27936 56
rect 27802 0 27858 54
rect 27908 42 27936 54
rect 28000 42 28028 6326
rect 28080 5840 28132 5846
rect 28080 5782 28132 5788
rect 28092 5370 28120 5782
rect 28080 5364 28132 5370
rect 28080 5306 28132 5312
rect 28276 4078 28304 6831
rect 28448 4616 28500 4622
rect 28552 4604 28580 8570
rect 28644 8412 28672 11194
rect 28722 9752 28778 9761
rect 28722 9687 28778 9696
rect 28736 8514 28764 9687
rect 28920 8634 28948 11194
rect 29196 9874 29224 11194
rect 29104 9846 29224 9874
rect 29000 9240 29052 9246
rect 29000 9182 29052 9188
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28736 8486 28856 8514
rect 28724 8424 28776 8430
rect 28644 8384 28724 8412
rect 28724 8366 28776 8372
rect 28828 7936 28856 8486
rect 28736 7908 28856 7936
rect 28736 7206 28764 7908
rect 28816 7812 28868 7818
rect 28816 7754 28868 7760
rect 28724 7200 28776 7206
rect 28724 7142 28776 7148
rect 28632 6928 28684 6934
rect 28632 6870 28684 6876
rect 28644 6633 28672 6870
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28630 6624 28686 6633
rect 28630 6559 28686 6568
rect 28736 6497 28764 6734
rect 28722 6488 28778 6497
rect 28722 6423 28778 6432
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28500 4576 28580 4604
rect 28632 4616 28684 4622
rect 28448 4558 28500 4564
rect 28632 4558 28684 4564
rect 28460 4146 28488 4558
rect 28644 4486 28672 4558
rect 28736 4486 28764 5170
rect 28632 4480 28684 4486
rect 28632 4422 28684 4428
rect 28724 4480 28776 4486
rect 28724 4422 28776 4428
rect 28448 4140 28500 4146
rect 28448 4082 28500 4088
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 28828 377 28856 7754
rect 28906 7168 28962 7177
rect 28906 7103 28962 7112
rect 28920 6866 28948 7103
rect 28908 6860 28960 6866
rect 28908 6802 28960 6808
rect 29012 3942 29040 9182
rect 29104 8498 29132 9846
rect 29184 9444 29236 9450
rect 29184 9386 29236 9392
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 29196 8294 29224 9386
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29472 7886 29500 11194
rect 29748 8566 29776 11194
rect 29828 9172 29880 9178
rect 29828 9114 29880 9120
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29104 7478 29132 7686
rect 29196 7546 29224 7754
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29092 7472 29144 7478
rect 29092 7414 29144 7420
rect 29092 4140 29144 4146
rect 29092 4082 29144 4088
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29104 3194 29132 4082
rect 29184 3528 29236 3534
rect 29184 3470 29236 3476
rect 29196 3194 29224 3470
rect 29288 3398 29316 7482
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29748 5710 29776 6054
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29380 4826 29408 5646
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29460 3392 29512 3398
rect 29460 3334 29512 3340
rect 29472 3194 29500 3334
rect 29840 3194 29868 9114
rect 29920 7472 29972 7478
rect 29918 7440 29920 7449
rect 29972 7440 29974 7449
rect 29918 7375 29974 7384
rect 29918 7032 29974 7041
rect 29918 6967 29974 6976
rect 29932 4826 29960 6967
rect 30024 5574 30052 11194
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30208 7954 30236 8230
rect 30196 7948 30248 7954
rect 30196 7890 30248 7896
rect 30012 5568 30064 5574
rect 30012 5510 30064 5516
rect 29920 4820 29972 4826
rect 29920 4762 29972 4768
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 30116 4282 30144 4558
rect 30104 4276 30156 4282
rect 30104 4218 30156 4224
rect 30300 4146 30328 11194
rect 30380 9104 30432 9110
rect 30380 9046 30432 9052
rect 30392 8634 30420 9046
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30392 3670 30420 7142
rect 30484 3942 30512 7686
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30300 3194 30328 3538
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29460 3188 29512 3194
rect 29460 3130 29512 3136
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 30288 3188 30340 3194
rect 30288 3130 30340 3136
rect 30576 3058 30604 11194
rect 30852 6798 30880 11194
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 29276 3052 29328 3058
rect 29276 2994 29328 3000
rect 30564 3052 30616 3058
rect 30564 2994 30616 3000
rect 28814 368 28870 377
rect 28814 303 28870 312
rect 29288 56 29316 2994
rect 30668 2038 30696 6258
rect 30760 5846 30788 6258
rect 30840 6112 30892 6118
rect 30840 6054 30892 6060
rect 30852 5846 30880 6054
rect 30748 5840 30800 5846
rect 30748 5782 30800 5788
rect 30840 5840 30892 5846
rect 30840 5782 30892 5788
rect 31128 5778 31156 11194
rect 31116 5772 31168 5778
rect 31116 5714 31168 5720
rect 31404 4758 31432 11194
rect 31680 9058 31708 11194
rect 31680 9030 31892 9058
rect 31392 4752 31444 4758
rect 31392 4694 31444 4700
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 30748 2576 30800 2582
rect 30748 2518 30800 2524
rect 30656 2032 30708 2038
rect 30656 1974 30708 1980
rect 30760 56 30788 2518
rect 31772 66 31800 2994
rect 31864 2990 31892 9030
rect 31956 8294 31984 11194
rect 32232 8634 32260 11194
rect 32508 8634 32536 11194
rect 32588 10192 32640 10198
rect 32588 10134 32640 10140
rect 32220 8628 32272 8634
rect 32220 8570 32272 8576
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 31956 7274 31984 7686
rect 31944 7268 31996 7274
rect 31944 7210 31996 7216
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32324 2106 32352 3878
rect 32416 3738 32444 8366
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32508 3194 32536 8434
rect 32600 7954 32628 10134
rect 32680 8900 32732 8906
rect 32680 8842 32732 8848
rect 32692 8498 32720 8842
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32784 8362 32812 11194
rect 33060 9602 33088 11194
rect 32876 9574 33088 9602
rect 33336 9602 33364 11194
rect 33336 9574 33548 9602
rect 32876 8634 32904 9574
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33520 8634 33548 9574
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33612 8362 33640 11194
rect 33888 9194 33916 11194
rect 33888 9166 34008 9194
rect 33784 8900 33836 8906
rect 33784 8842 33836 8848
rect 33692 8492 33744 8498
rect 33692 8434 33744 8440
rect 32772 8356 32824 8362
rect 32772 8298 32824 8304
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 33508 7744 33560 7750
rect 33508 7686 33560 7692
rect 32588 4684 32640 4690
rect 32588 4626 32640 4632
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32312 2100 32364 2106
rect 32312 2042 32364 2048
rect 31760 60 31812 66
rect 27908 14 28028 42
rect 29274 0 29330 56
rect 30746 0 30802 56
rect 32232 56 32352 82
rect 31760 2 31812 8
rect 32218 54 32352 56
rect 32218 0 32274 54
rect 32324 42 32352 54
rect 32600 42 32628 4626
rect 32784 1737 32812 7686
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33428 7206 33456 7686
rect 33416 7200 33468 7206
rect 33416 7142 33468 7148
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 32862 5400 32918 5409
rect 33010 5403 33318 5412
rect 32862 5335 32918 5344
rect 32876 4185 32904 5335
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 32862 4176 32918 4185
rect 32862 4111 32918 4120
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 32770 1728 32826 1737
rect 32770 1663 32826 1672
rect 33428 270 33456 5170
rect 33520 2417 33548 7686
rect 33704 5370 33732 8434
rect 33692 5364 33744 5370
rect 33692 5306 33744 5312
rect 33796 5098 33824 8842
rect 33980 8634 34008 9166
rect 34060 8832 34112 8838
rect 34060 8774 34112 8780
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34072 6186 34100 8774
rect 34164 8566 34192 11194
rect 34244 8968 34296 8974
rect 34244 8910 34296 8916
rect 34152 8560 34204 8566
rect 34152 8502 34204 8508
rect 34256 8430 34284 8910
rect 34244 8424 34296 8430
rect 34244 8366 34296 8372
rect 34440 8090 34468 11194
rect 34716 8362 34744 11194
rect 34992 8922 35020 11194
rect 34992 8894 35112 8922
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 34704 8356 34756 8362
rect 34704 8298 34756 8304
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34060 6180 34112 6186
rect 34060 6122 34112 6128
rect 34152 5568 34204 5574
rect 34152 5510 34204 5516
rect 33784 5092 33836 5098
rect 33784 5034 33836 5040
rect 33968 5024 34020 5030
rect 33968 4966 34020 4972
rect 33980 4826 34008 4966
rect 33968 4820 34020 4826
rect 33968 4762 34020 4768
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 33888 3398 33916 3538
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 34164 3058 34192 5510
rect 34992 4826 35020 8434
rect 35084 8430 35112 8894
rect 35268 8566 35296 11194
rect 35440 9104 35492 9110
rect 35440 9046 35492 9052
rect 35256 8560 35308 8566
rect 35256 8502 35308 8508
rect 35452 8498 35480 9046
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35072 8424 35124 8430
rect 35072 8366 35124 8372
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35072 7744 35124 7750
rect 35072 7686 35124 7692
rect 35084 6934 35112 7686
rect 35072 6928 35124 6934
rect 35072 6870 35124 6876
rect 35176 4826 35204 7822
rect 34980 4820 35032 4826
rect 34980 4762 35032 4768
rect 35164 4820 35216 4826
rect 35164 4762 35216 4768
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 34624 3194 34652 3402
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 34520 2916 34572 2922
rect 34520 2858 34572 2864
rect 33506 2408 33562 2417
rect 33506 2343 33562 2352
rect 33416 264 33468 270
rect 33416 206 33468 212
rect 33692 196 33744 202
rect 33692 138 33744 144
rect 33704 56 33732 138
rect 34532 105 34560 2858
rect 34808 338 34836 4422
rect 35360 3126 35388 8434
rect 35544 8090 35572 11194
rect 35624 8900 35676 8906
rect 35624 8842 35676 8848
rect 35636 8498 35664 8842
rect 35820 8634 35848 11194
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35624 8492 35676 8498
rect 35624 8434 35676 8440
rect 35900 8288 35952 8294
rect 35900 8230 35952 8236
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35912 3194 35940 8230
rect 36096 8090 36124 11194
rect 36176 8832 36228 8838
rect 36176 8774 36228 8780
rect 36188 8498 36216 8774
rect 36176 8492 36228 8498
rect 36176 8434 36228 8440
rect 36372 8430 36400 11194
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36360 8424 36412 8430
rect 36360 8366 36412 8372
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36452 7880 36504 7886
rect 36452 7822 36504 7828
rect 35992 4616 36044 4622
rect 35992 4558 36044 4564
rect 35900 3188 35952 3194
rect 35900 3130 35952 3136
rect 35164 3120 35216 3126
rect 35164 3062 35216 3068
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 34796 332 34848 338
rect 34796 274 34848 280
rect 34518 96 34574 105
rect 32324 14 32628 42
rect 33690 0 33746 56
rect 35176 56 35204 3062
rect 35256 2984 35308 2990
rect 35256 2926 35308 2932
rect 35268 406 35296 2926
rect 35256 400 35308 406
rect 35256 342 35308 348
rect 36004 241 36032 4558
rect 36268 4548 36320 4554
rect 36268 4490 36320 4496
rect 35990 232 36046 241
rect 35990 167 36046 176
rect 34518 31 34574 40
rect 35162 0 35218 56
rect 36280 42 36308 4490
rect 36464 4486 36492 7822
rect 36452 4480 36504 4486
rect 36452 4422 36504 4428
rect 36556 3602 36584 8434
rect 36648 8090 36676 11194
rect 36924 8634 36952 11194
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 36820 8560 36872 8566
rect 36820 8502 36872 8508
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 36740 2961 36768 7822
rect 36832 3534 36860 8502
rect 37096 8492 37148 8498
rect 37096 8434 37148 8440
rect 37004 8016 37056 8022
rect 37004 7958 37056 7964
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 36726 2952 36782 2961
rect 36726 2887 36782 2896
rect 37016 2514 37044 7958
rect 37108 4826 37136 8434
rect 37200 8362 37228 11194
rect 37280 9784 37332 9790
rect 37280 9726 37332 9732
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37292 8072 37320 9726
rect 37476 8566 37504 11194
rect 37648 9716 37700 9722
rect 37648 9658 37700 9664
rect 37556 9036 37608 9042
rect 37556 8978 37608 8984
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37464 8424 37516 8430
rect 37464 8366 37516 8372
rect 37200 8044 37320 8072
rect 37200 5522 37228 8044
rect 37278 7984 37334 7993
rect 37278 7919 37334 7928
rect 37292 6662 37320 7919
rect 37372 7472 37424 7478
rect 37372 7414 37424 7420
rect 37280 6656 37332 6662
rect 37280 6598 37332 6604
rect 37384 5794 37412 7414
rect 37292 5766 37412 5794
rect 37292 5710 37320 5766
rect 37280 5704 37332 5710
rect 37280 5646 37332 5652
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 37200 5494 37320 5522
rect 37096 4820 37148 4826
rect 37096 4762 37148 4768
rect 37292 4078 37320 5494
rect 37280 4072 37332 4078
rect 37280 4014 37332 4020
rect 37004 2508 37056 2514
rect 37004 2450 37056 2456
rect 37384 134 37412 5646
rect 37476 5030 37504 8366
rect 37568 6798 37596 8978
rect 37660 7970 37688 9658
rect 37752 8090 37780 11194
rect 38382 9888 38438 9897
rect 38382 9823 38438 9832
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37660 7942 37780 7970
rect 37648 7812 37700 7818
rect 37648 7754 37700 7760
rect 37556 6792 37608 6798
rect 37556 6734 37608 6740
rect 37556 6656 37608 6662
rect 37556 6598 37608 6604
rect 37568 6458 37596 6598
rect 37660 6458 37688 7754
rect 37556 6452 37608 6458
rect 37556 6394 37608 6400
rect 37648 6452 37700 6458
rect 37648 6394 37700 6400
rect 37556 6248 37608 6254
rect 37556 6190 37608 6196
rect 37464 5024 37516 5030
rect 37464 4966 37516 4972
rect 37568 3369 37596 6190
rect 37752 6118 37780 7942
rect 37740 6112 37792 6118
rect 37740 6054 37792 6060
rect 37844 5914 37872 8910
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38120 7313 38148 7346
rect 38304 7342 38332 7822
rect 38396 7546 38424 9823
rect 39670 9616 39726 9625
rect 39670 9551 39726 9560
rect 38844 9376 38896 9382
rect 38658 9344 38714 9353
rect 38844 9318 38896 9324
rect 38658 9279 38714 9288
rect 38476 8492 38528 8498
rect 38476 8434 38528 8440
rect 38384 7540 38436 7546
rect 38384 7482 38436 7488
rect 38292 7336 38344 7342
rect 38106 7304 38162 7313
rect 38292 7278 38344 7284
rect 38106 7239 38162 7248
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38198 6896 38254 6905
rect 38488 6882 38516 8434
rect 38672 7546 38700 9279
rect 38752 9172 38804 9178
rect 38752 9114 38804 9120
rect 38764 8566 38792 9114
rect 38752 8560 38804 8566
rect 38752 8502 38804 8508
rect 38856 8498 38884 9318
rect 39578 8800 39634 8809
rect 39010 8732 39318 8741
rect 39578 8735 39634 8744
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 38934 8528 38990 8537
rect 38844 8492 38896 8498
rect 38934 8463 38990 8472
rect 38844 8434 38896 8440
rect 38948 7546 38976 8463
rect 39028 8356 39080 8362
rect 39028 8298 39080 8304
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 39040 8265 39068 8298
rect 39026 8256 39082 8265
rect 39026 8191 39082 8200
rect 39408 7993 39436 8298
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 39396 7744 39448 7750
rect 39396 7686 39448 7692
rect 39486 7712 39542 7721
rect 39010 7644 39318 7653
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 38660 7540 38712 7546
rect 38660 7482 38712 7488
rect 38936 7540 38988 7546
rect 38936 7482 38988 7488
rect 39408 7449 39436 7686
rect 39486 7647 39542 7656
rect 39394 7440 39450 7449
rect 38568 7404 38620 7410
rect 38568 7346 38620 7352
rect 38844 7404 38896 7410
rect 39394 7375 39450 7384
rect 38844 7346 38896 7352
rect 38198 6831 38254 6840
rect 38304 6854 38516 6882
rect 38212 6798 38240 6831
rect 38016 6792 38068 6798
rect 38016 6734 38068 6740
rect 38200 6792 38252 6798
rect 38200 6734 38252 6740
rect 38028 6118 38056 6734
rect 38016 6112 38068 6118
rect 38016 6054 38068 6060
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 37740 5228 37792 5234
rect 37740 5170 37792 5176
rect 37554 3360 37610 3369
rect 37554 3295 37610 3304
rect 37752 2774 37780 5170
rect 37830 5128 37886 5137
rect 38304 5098 38332 6854
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38384 6656 38436 6662
rect 38384 6598 38436 6604
rect 38396 6390 38424 6598
rect 38384 6384 38436 6390
rect 38384 6326 38436 6332
rect 38488 6225 38516 6734
rect 38474 6216 38530 6225
rect 38474 6151 38530 6160
rect 38476 6112 38528 6118
rect 38476 6054 38528 6060
rect 38488 5914 38516 6054
rect 38476 5908 38528 5914
rect 38476 5850 38528 5856
rect 38580 5681 38608 7346
rect 38856 7002 38884 7346
rect 39304 7268 39356 7274
rect 39304 7210 39356 7216
rect 38844 6996 38896 7002
rect 38844 6938 38896 6944
rect 39316 6905 39344 7210
rect 39302 6896 39358 6905
rect 39302 6831 39358 6840
rect 38842 6760 38898 6769
rect 38842 6695 38898 6704
rect 38660 6656 38712 6662
rect 38660 6598 38712 6604
rect 38672 6361 38700 6598
rect 38750 6488 38806 6497
rect 38750 6423 38806 6432
rect 38658 6352 38714 6361
rect 38658 6287 38714 6296
rect 38764 6202 38792 6423
rect 38856 6322 38884 6695
rect 39500 6662 39528 7647
rect 39592 7546 39620 8735
rect 39580 7540 39632 7546
rect 39580 7482 39632 7488
rect 39578 7168 39634 7177
rect 39578 7103 39634 7112
rect 39488 6656 39540 6662
rect 39394 6624 39450 6633
rect 39488 6598 39540 6604
rect 39010 6556 39318 6565
rect 39394 6559 39450 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 38844 6316 38896 6322
rect 38844 6258 38896 6264
rect 38936 6316 38988 6322
rect 38936 6258 38988 6264
rect 38764 6174 38884 6202
rect 38660 6112 38712 6118
rect 38658 6080 38660 6089
rect 38712 6080 38714 6089
rect 38658 6015 38714 6024
rect 38660 5840 38712 5846
rect 38660 5782 38712 5788
rect 38566 5672 38622 5681
rect 38566 5607 38622 5616
rect 37830 5063 37886 5072
rect 38292 5092 38344 5098
rect 37844 4826 37872 5063
rect 38292 5034 38344 5040
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 38568 4616 38620 4622
rect 38474 4584 38530 4593
rect 38568 4558 38620 4564
rect 38474 4519 38476 4528
rect 38528 4519 38530 4528
rect 38476 4490 38528 4496
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38474 3088 38530 3097
rect 38474 3023 38476 3032
rect 38528 3023 38530 3032
rect 38476 2994 38528 3000
rect 37752 2746 37872 2774
rect 37372 128 37424 134
rect 36556 56 36676 82
rect 37372 70 37424 76
rect 36556 54 36690 56
rect 36556 42 36584 54
rect 36280 14 36584 42
rect 36634 0 36690 54
rect 37844 42 37872 2746
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38580 2582 38608 4558
rect 38672 4060 38700 5782
rect 38856 5710 38884 6174
rect 38844 5704 38896 5710
rect 38844 5646 38896 5652
rect 38948 5386 38976 6258
rect 39408 5914 39436 6559
rect 39592 6458 39620 7103
rect 39580 6452 39632 6458
rect 39580 6394 39632 6400
rect 39488 6384 39540 6390
rect 39488 6326 39540 6332
rect 39396 5908 39448 5914
rect 39396 5850 39448 5856
rect 39210 5808 39266 5817
rect 39210 5743 39266 5752
rect 39394 5808 39450 5817
rect 39394 5743 39450 5752
rect 39224 5710 39252 5743
rect 39212 5704 39264 5710
rect 39212 5646 39264 5652
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 38764 5358 38976 5386
rect 39408 5370 39436 5743
rect 39396 5364 39448 5370
rect 38764 5166 38792 5358
rect 39396 5306 39448 5312
rect 38936 5296 38988 5302
rect 38936 5238 38988 5244
rect 39210 5264 39266 5273
rect 38844 5228 38896 5234
rect 38844 5170 38896 5176
rect 38752 5160 38804 5166
rect 38752 5102 38804 5108
rect 38856 4729 38884 5170
rect 38842 4720 38898 4729
rect 38842 4655 38898 4664
rect 38752 4616 38804 4622
rect 38752 4558 38804 4564
rect 38764 4185 38792 4558
rect 38948 4554 38976 5238
rect 39210 5199 39212 5208
rect 39264 5199 39266 5208
rect 39394 5264 39450 5273
rect 39394 5199 39450 5208
rect 39212 5170 39264 5176
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39408 4826 39436 5199
rect 39396 4820 39448 4826
rect 39396 4762 39448 4768
rect 39394 4720 39450 4729
rect 39394 4655 39450 4664
rect 38936 4548 38988 4554
rect 38936 4490 38988 4496
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 38750 4176 38806 4185
rect 39026 4176 39082 4185
rect 38750 4111 38806 4120
rect 38844 4140 38896 4146
rect 39026 4111 39082 4120
rect 38844 4082 38896 4088
rect 38672 4032 38792 4060
rect 38856 4049 38884 4082
rect 38660 3936 38712 3942
rect 38660 3878 38712 3884
rect 38672 3641 38700 3878
rect 38658 3632 38714 3641
rect 38658 3567 38714 3576
rect 38764 3534 38792 4032
rect 38842 4040 38898 4049
rect 39040 4010 39068 4111
rect 39408 4010 39436 4655
rect 39500 4146 39528 6326
rect 39684 6186 39712 9551
rect 40038 9072 40094 9081
rect 40038 9007 40094 9016
rect 39764 8016 39816 8022
rect 39764 7958 39816 7964
rect 39672 6180 39724 6186
rect 39672 6122 39724 6128
rect 39578 4448 39634 4457
rect 39578 4383 39634 4392
rect 39488 4140 39540 4146
rect 39488 4082 39540 4088
rect 38842 3975 38898 3984
rect 39028 4004 39080 4010
rect 39028 3946 39080 3952
rect 39396 4004 39448 4010
rect 39396 3946 39448 3952
rect 39394 3904 39450 3913
rect 39394 3839 39450 3848
rect 38936 3664 38988 3670
rect 38936 3606 38988 3612
rect 38752 3528 38804 3534
rect 38752 3470 38804 3476
rect 38842 3496 38898 3505
rect 38842 3431 38898 3440
rect 38856 3058 38884 3431
rect 38948 3058 38976 3606
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39408 3194 39436 3839
rect 39592 3738 39620 4383
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39776 3534 39804 7958
rect 39856 7200 39908 7206
rect 39856 7142 39908 7148
rect 39764 3528 39816 3534
rect 39764 3470 39816 3476
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39394 3088 39450 3097
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 38936 3052 38988 3058
rect 39394 3023 39450 3032
rect 38936 2994 38988 3000
rect 38660 2848 38712 2854
rect 39028 2848 39080 2854
rect 38660 2790 38712 2796
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 38568 2576 38620 2582
rect 38672 2553 38700 2790
rect 39026 2751 39082 2760
rect 39408 2650 39436 3023
rect 39868 2774 39896 7142
rect 40052 6730 40080 9007
rect 40132 7812 40184 7818
rect 40132 7754 40184 7760
rect 40040 6724 40092 6730
rect 40040 6666 40092 6672
rect 39948 5840 40000 5846
rect 39948 5782 40000 5788
rect 39960 5545 39988 5782
rect 39946 5536 40002 5545
rect 39946 5471 40002 5480
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 39960 3369 39988 3606
rect 39946 3360 40002 3369
rect 39946 3295 40002 3304
rect 40144 2922 40172 7754
rect 40132 2916 40184 2922
rect 40132 2858 40184 2864
rect 39684 2746 39896 2774
rect 39396 2644 39448 2650
rect 39396 2586 39448 2592
rect 38568 2518 38620 2524
rect 38658 2544 38714 2553
rect 39684 2514 39712 2746
rect 38658 2479 38714 2488
rect 39672 2508 39724 2514
rect 39672 2450 39724 2456
rect 38476 2440 38528 2446
rect 39212 2440 39264 2446
rect 38476 2382 38528 2388
rect 39210 2408 39212 2417
rect 39264 2408 39266 2417
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 37936 2009 37964 2246
rect 37922 2000 37978 2009
rect 37922 1935 37978 1944
rect 38304 1737 38332 2246
rect 38488 1834 38516 2382
rect 39210 2343 39266 2352
rect 38660 2304 38712 2310
rect 39948 2304 40000 2310
rect 38660 2246 38712 2252
rect 39946 2272 39948 2281
rect 40000 2272 40002 2281
rect 38476 1828 38528 1834
rect 38476 1770 38528 1776
rect 38290 1728 38346 1737
rect 38290 1663 38346 1672
rect 38672 1465 38700 2246
rect 39010 2204 39318 2213
rect 39946 2207 40002 2216
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38658 1456 38714 1465
rect 38658 1391 38714 1400
rect 39578 368 39634 377
rect 39578 303 39634 312
rect 38028 56 38148 82
rect 39592 56 39620 303
rect 38028 54 38162 56
rect 38028 42 38056 54
rect 37844 14 38056 42
rect 38106 0 38162 54
rect 39578 0 39634 56
<< via2 >>
rect 1030 9560 1086 9616
rect 662 9288 718 9344
rect 294 9152 350 9208
rect 202 6024 258 6080
rect 478 8880 534 8936
rect 386 7928 442 7984
rect 294 3848 350 3904
rect 938 8744 994 8800
rect 754 7656 810 7712
rect 1490 9424 1546 9480
rect 1122 9016 1178 9072
rect 1398 9016 1454 9072
rect 1306 8508 1308 8528
rect 1308 8508 1360 8528
rect 1360 8508 1362 8528
rect 1306 8472 1362 8508
rect 1214 8200 1270 8256
rect 846 7384 902 7440
rect 754 7112 810 7168
rect 754 6840 810 6896
rect 846 6568 902 6624
rect 1030 6296 1086 6352
rect 846 5752 902 5808
rect 754 5480 810 5536
rect 846 5208 902 5264
rect 754 4936 810 4992
rect 570 4664 626 4720
rect 478 3576 534 3632
rect 1030 3304 1086 3360
rect 386 2488 442 2544
rect 1582 7248 1638 7304
rect 2778 9832 2834 9888
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3330 8472 3386 8528
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2778 6180 2834 6216
rect 2778 6160 2780 6180
rect 2780 6160 2832 6180
rect 2832 6160 2834 6180
rect 3146 5652 3148 5672
rect 3148 5652 3200 5672
rect 3200 5652 3202 5672
rect 3146 5616 3202 5652
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 3882 6296 3938 6352
rect 5814 8336 5870 8392
rect 3606 4528 3662 4584
rect 1306 4392 1362 4448
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 1122 1944 1178 2000
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3514 3032 3570 3088
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1214 1400 1270 1456
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 5262 5772 5318 5808
rect 5262 5752 5264 5772
rect 5264 5752 5316 5772
rect 5316 5752 5318 5772
rect 6734 7792 6790 7848
rect 5998 5652 6000 5672
rect 6000 5652 6052 5672
rect 6052 5652 6054 5672
rect 5998 5616 6054 5652
rect 5814 3460 5870 3496
rect 5814 3440 5816 3460
rect 5816 3440 5868 3460
rect 5868 3440 5870 3460
rect 6274 5652 6276 5672
rect 6276 5652 6328 5672
rect 6328 5652 6330 5672
rect 6274 5616 6330 5652
rect 6182 2896 6238 2952
rect 7286 7384 7342 7440
rect 6550 5752 6606 5808
rect 7470 6840 7526 6896
rect 8022 9696 8078 9752
rect 8390 11056 8446 11112
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7654 7928 7710 7984
rect 7838 7248 7894 7304
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 8666 9152 8722 9208
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 8942 8472 8998 8528
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7838 5752 7894 5808
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 8298 4528 8354 4584
rect 7654 4120 7710 4176
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 10598 8472 10654 8528
rect 9126 7964 9128 7984
rect 9128 7964 9180 7984
rect 9180 7964 9182 7984
rect 9126 7928 9182 7964
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9402 6432 9458 6488
rect 9218 6024 9274 6080
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 8850 4528 8906 4584
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 8666 3576 8722 3632
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 8574 2896 8630 2952
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 6458 2488 6514 2544
rect 9494 5480 9550 5536
rect 10138 5652 10140 5672
rect 10140 5652 10192 5672
rect 10192 5652 10194 5672
rect 10138 5616 10194 5652
rect 11058 7928 11114 7984
rect 11150 7384 11206 7440
rect 10874 7268 10930 7304
rect 10874 7248 10876 7268
rect 10876 7248 10928 7268
rect 10928 7248 10930 7268
rect 10782 3984 10838 4040
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 12714 6704 12770 6760
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14370 8064 14426 8120
rect 13726 7792 13782 7848
rect 13542 5208 13598 5264
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 13818 6024 13874 6080
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13726 5636 13782 5672
rect 13726 5616 13728 5636
rect 13728 5616 13780 5636
rect 13780 5616 13782 5636
rect 13634 5072 13690 5128
rect 13634 4700 13636 4720
rect 13636 4700 13688 4720
rect 13688 4700 13690 4720
rect 13634 4664 13690 4700
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14370 7656 14426 7712
rect 14554 8236 14556 8256
rect 14556 8236 14608 8256
rect 14608 8236 14610 8256
rect 14554 8200 14610 8236
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14646 7828 14648 7848
rect 14648 7828 14700 7848
rect 14700 7828 14702 7848
rect 14646 7792 14702 7828
rect 16210 8472 16266 8528
rect 16394 8472 16450 8528
rect 14554 5480 14610 5536
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 15566 7520 15622 7576
rect 15290 7112 15346 7168
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 15014 6332 15016 6352
rect 15016 6332 15068 6352
rect 15068 6332 15070 6352
rect 15014 6296 15070 6332
rect 15198 6296 15254 6352
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 14554 4800 14610 4856
rect 12162 2896 12218 2952
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 13082 1944 13138 2000
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 17222 8064 17278 8120
rect 17774 8200 17830 8256
rect 17222 7656 17278 7712
rect 16394 6432 16450 6488
rect 17958 5208 18014 5264
rect 18326 7112 18382 7168
rect 18878 4800 18934 4856
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 20350 11056 20406 11112
rect 20074 9152 20130 9208
rect 21178 9152 21234 9208
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 20350 7520 20406 7576
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20350 6976 20406 7032
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 20626 8200 20682 8256
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 20626 7112 20682 7168
rect 20718 6432 20774 6488
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 20718 5888 20774 5944
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 20810 5344 20866 5400
rect 22190 8472 22246 8528
rect 22466 8472 22522 8528
rect 20810 4972 20812 4992
rect 20812 4972 20864 4992
rect 20864 4972 20866 4992
rect 20810 4936 20866 4972
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20442 2760 20498 2816
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 21546 7520 21602 7576
rect 21546 5208 21602 5264
rect 21546 4972 21548 4992
rect 21548 4972 21600 4992
rect 21600 4972 21602 4992
rect 21546 4936 21602 4972
rect 23018 9152 23074 9208
rect 22006 3188 22062 3224
rect 22006 3168 22008 3188
rect 22008 3168 22060 3188
rect 22060 3168 22062 3188
rect 23202 8336 23258 8392
rect 23846 7384 23902 7440
rect 23294 2760 23350 2816
rect 24398 8084 24454 8120
rect 24398 8064 24400 8084
rect 24400 8064 24452 8084
rect 24452 8064 24454 8084
rect 24766 8880 24822 8936
rect 24766 7112 24822 7168
rect 25686 9016 25742 9072
rect 25134 8200 25190 8256
rect 25318 6840 25374 6896
rect 25502 7792 25558 7848
rect 25502 5888 25558 5944
rect 25042 3168 25098 3224
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 17498 40 17554 96
rect 21914 176 21970 232
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 26606 7520 26662 7576
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 26882 6840 26938 6896
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27434 5344 27490 5400
rect 27434 4936 27490 4992
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27894 8472 27950 8528
rect 28354 7148 28356 7168
rect 28356 7148 28408 7168
rect 28408 7148 28410 7168
rect 28354 7112 28410 7148
rect 28262 6840 28318 6896
rect 27802 6568 27858 6624
rect 27894 6432 27950 6488
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 27802 4120 27858 4176
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 26330 1944 26386 2000
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 28722 9696 28778 9752
rect 28630 6568 28686 6624
rect 28722 6432 28778 6488
rect 28906 7112 28962 7168
rect 29918 7420 29920 7440
rect 29920 7420 29972 7440
rect 29972 7420 29974 7440
rect 29918 7384 29974 7420
rect 29918 6976 29974 7032
rect 28814 312 28870 368
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 32862 5344 32918 5400
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 32862 4120 32918 4176
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 32770 1672 32826 1728
rect 33506 2352 33562 2408
rect 34518 40 34574 96
rect 35990 176 36046 232
rect 36726 2896 36782 2952
rect 37278 7928 37334 7984
rect 38382 9832 38438 9888
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 39670 9560 39726 9616
rect 38658 9288 38714 9344
rect 38106 7248 38162 7304
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 38198 6840 38254 6896
rect 39578 8744 39634 8800
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 38934 8472 38990 8528
rect 39026 8200 39082 8256
rect 39394 7928 39450 7984
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 39486 7656 39542 7712
rect 39394 7384 39450 7440
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37554 3304 37610 3360
rect 37830 5072 37886 5128
rect 38474 6160 38530 6216
rect 39302 6840 39358 6896
rect 38842 6704 38898 6760
rect 38750 6432 38806 6488
rect 38658 6296 38714 6352
rect 39578 7112 39634 7168
rect 39394 6568 39450 6624
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 38658 6060 38660 6080
rect 38660 6060 38712 6080
rect 38712 6060 38714 6080
rect 38658 6024 38714 6060
rect 38566 5616 38622 5672
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 38474 4548 38530 4584
rect 38474 4528 38476 4548
rect 38476 4528 38528 4548
rect 38528 4528 38530 4548
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 38474 3052 38530 3088
rect 38474 3032 38476 3052
rect 38476 3032 38528 3052
rect 38528 3032 38530 3052
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 39210 5752 39266 5808
rect 39394 5752 39450 5808
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 38842 4664 38898 4720
rect 39210 5228 39266 5264
rect 39210 5208 39212 5228
rect 39212 5208 39264 5228
rect 39264 5208 39266 5228
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 39394 4664 39450 4720
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 38750 4120 38806 4176
rect 39026 4120 39082 4176
rect 38658 3576 38714 3632
rect 38842 3984 38898 4040
rect 40038 9016 40094 9072
rect 39578 4392 39634 4448
rect 39394 3848 39450 3904
rect 38842 3440 38898 3496
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39394 3032 39450 3088
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 39946 5480 40002 5536
rect 39946 3304 40002 3360
rect 38658 2488 38714 2544
rect 39210 2388 39212 2408
rect 39212 2388 39264 2408
rect 39264 2388 39266 2408
rect 37922 1944 37978 2000
rect 39210 2352 39266 2388
rect 39946 2252 39948 2272
rect 39948 2252 40000 2272
rect 40000 2252 40002 2272
rect 38290 1672 38346 1728
rect 39946 2216 40002 2252
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38658 1400 38714 1456
rect 39578 312 39634 368
<< metal3 >>
rect 8385 11114 8451 11117
rect 20345 11114 20411 11117
rect 8385 11112 20411 11114
rect 8385 11056 8390 11112
rect 8446 11056 20350 11112
rect 20406 11056 20411 11112
rect 8385 11054 20411 11056
rect 8385 11051 8451 11054
rect 20345 11051 20411 11054
rect 0 9890 120 9920
rect 2773 9890 2839 9893
rect 0 9888 2839 9890
rect 0 9832 2778 9888
rect 2834 9832 2839 9888
rect 0 9830 2839 9832
rect 0 9800 120 9830
rect 2773 9827 2839 9830
rect 38377 9890 38443 9893
rect 40880 9890 41000 9920
rect 38377 9888 41000 9890
rect 38377 9832 38382 9888
rect 38438 9832 41000 9888
rect 38377 9830 41000 9832
rect 38377 9827 38443 9830
rect 40880 9800 41000 9830
rect 8017 9754 8083 9757
rect 28717 9754 28783 9757
rect 8017 9752 28783 9754
rect 8017 9696 8022 9752
rect 8078 9696 28722 9752
rect 28778 9696 28783 9752
rect 8017 9694 28783 9696
rect 8017 9691 8083 9694
rect 28717 9691 28783 9694
rect 0 9618 120 9648
rect 1025 9618 1091 9621
rect 0 9616 1091 9618
rect 0 9560 1030 9616
rect 1086 9560 1091 9616
rect 0 9558 1091 9560
rect 0 9528 120 9558
rect 1025 9555 1091 9558
rect 39665 9618 39731 9621
rect 40880 9618 41000 9648
rect 39665 9616 41000 9618
rect 39665 9560 39670 9616
rect 39726 9560 41000 9616
rect 39665 9558 41000 9560
rect 39665 9555 39731 9558
rect 40880 9528 41000 9558
rect 1485 9482 1551 9485
rect 37222 9482 37228 9484
rect 1485 9480 37228 9482
rect 1485 9424 1490 9480
rect 1546 9424 37228 9480
rect 1485 9422 37228 9424
rect 1485 9419 1551 9422
rect 37222 9420 37228 9422
rect 37292 9420 37298 9484
rect 0 9346 120 9376
rect 657 9346 723 9349
rect 24710 9346 24716 9348
rect 0 9344 723 9346
rect 0 9288 662 9344
rect 718 9288 723 9344
rect 0 9286 723 9288
rect 0 9256 120 9286
rect 657 9283 723 9286
rect 2730 9286 24716 9346
rect 289 9210 355 9213
rect 2730 9210 2790 9286
rect 24710 9284 24716 9286
rect 24780 9284 24786 9348
rect 38653 9346 38719 9349
rect 40880 9346 41000 9376
rect 38653 9344 41000 9346
rect 38653 9288 38658 9344
rect 38714 9288 41000 9344
rect 38653 9286 41000 9288
rect 38653 9283 38719 9286
rect 40880 9256 41000 9286
rect 289 9208 2790 9210
rect 289 9152 294 9208
rect 350 9152 2790 9208
rect 289 9150 2790 9152
rect 8661 9210 8727 9213
rect 20069 9210 20135 9213
rect 8661 9208 20135 9210
rect 8661 9152 8666 9208
rect 8722 9152 20074 9208
rect 20130 9152 20135 9208
rect 8661 9150 20135 9152
rect 289 9147 355 9150
rect 8661 9147 8727 9150
rect 20069 9147 20135 9150
rect 21173 9210 21239 9213
rect 23013 9210 23079 9213
rect 21173 9208 23079 9210
rect 21173 9152 21178 9208
rect 21234 9152 23018 9208
rect 23074 9152 23079 9208
rect 21173 9150 23079 9152
rect 21173 9147 21239 9150
rect 23013 9147 23079 9150
rect 0 9074 120 9104
rect 1117 9074 1183 9077
rect 0 9072 1183 9074
rect 0 9016 1122 9072
rect 1178 9016 1183 9072
rect 0 9014 1183 9016
rect 0 8984 120 9014
rect 1117 9011 1183 9014
rect 1393 9074 1459 9077
rect 25681 9074 25747 9077
rect 1393 9072 25747 9074
rect 1393 9016 1398 9072
rect 1454 9016 25686 9072
rect 25742 9016 25747 9072
rect 1393 9014 25747 9016
rect 1393 9011 1459 9014
rect 25681 9011 25747 9014
rect 40033 9074 40099 9077
rect 40880 9074 41000 9104
rect 40033 9072 41000 9074
rect 40033 9016 40038 9072
rect 40094 9016 41000 9072
rect 40033 9014 41000 9016
rect 40033 9011 40099 9014
rect 40880 8984 41000 9014
rect 473 8938 539 8941
rect 24761 8938 24827 8941
rect 473 8936 24827 8938
rect 473 8880 478 8936
rect 534 8880 24766 8936
rect 24822 8880 24827 8936
rect 473 8878 24827 8880
rect 473 8875 539 8878
rect 24761 8875 24827 8878
rect 0 8802 120 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 120 8742
rect 933 8739 999 8742
rect 39573 8802 39639 8805
rect 40880 8802 41000 8832
rect 39573 8800 41000 8802
rect 39573 8744 39578 8800
rect 39634 8744 41000 8800
rect 39573 8742 41000 8744
rect 39573 8739 39639 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 0 8530 120 8560
rect 1301 8530 1367 8533
rect 0 8528 1367 8530
rect 0 8472 1306 8528
rect 1362 8472 1367 8528
rect 0 8470 1367 8472
rect 0 8440 120 8470
rect 1301 8467 1367 8470
rect 3325 8530 3391 8533
rect 8937 8530 9003 8533
rect 3325 8528 9003 8530
rect 3325 8472 3330 8528
rect 3386 8472 8942 8528
rect 8998 8472 9003 8528
rect 3325 8470 9003 8472
rect 3325 8467 3391 8470
rect 8937 8467 9003 8470
rect 10593 8530 10659 8533
rect 16205 8530 16271 8533
rect 10593 8528 16271 8530
rect 10593 8472 10598 8528
rect 10654 8472 16210 8528
rect 16266 8472 16271 8528
rect 10593 8470 16271 8472
rect 10593 8467 10659 8470
rect 16205 8467 16271 8470
rect 16389 8530 16455 8533
rect 22185 8530 22251 8533
rect 16389 8528 22251 8530
rect 16389 8472 16394 8528
rect 16450 8472 22190 8528
rect 22246 8472 22251 8528
rect 16389 8470 22251 8472
rect 16389 8467 16455 8470
rect 22185 8467 22251 8470
rect 22461 8530 22527 8533
rect 27889 8530 27955 8533
rect 22461 8528 27955 8530
rect 22461 8472 22466 8528
rect 22522 8472 27894 8528
rect 27950 8472 27955 8528
rect 22461 8470 27955 8472
rect 22461 8467 22527 8470
rect 27889 8467 27955 8470
rect 38929 8530 38995 8533
rect 40880 8530 41000 8560
rect 38929 8528 41000 8530
rect 38929 8472 38934 8528
rect 38990 8472 41000 8528
rect 38929 8470 41000 8472
rect 38929 8467 38995 8470
rect 40880 8440 41000 8470
rect 5809 8394 5875 8397
rect 23197 8394 23263 8397
rect 5809 8392 23263 8394
rect 5809 8336 5814 8392
rect 5870 8336 23202 8392
rect 23258 8336 23263 8392
rect 5809 8334 23263 8336
rect 5809 8331 5875 8334
rect 23197 8331 23263 8334
rect 0 8258 120 8288
rect 1209 8258 1275 8261
rect 0 8256 1275 8258
rect 0 8200 1214 8256
rect 1270 8200 1275 8256
rect 0 8198 1275 8200
rect 0 8168 120 8198
rect 1209 8195 1275 8198
rect 14549 8258 14615 8261
rect 17769 8258 17835 8261
rect 14549 8256 17835 8258
rect 14549 8200 14554 8256
rect 14610 8200 17774 8256
rect 17830 8200 17835 8256
rect 14549 8198 17835 8200
rect 14549 8195 14615 8198
rect 17769 8195 17835 8198
rect 20621 8258 20687 8261
rect 25129 8258 25195 8261
rect 20621 8256 25195 8258
rect 20621 8200 20626 8256
rect 20682 8200 25134 8256
rect 25190 8200 25195 8256
rect 20621 8198 25195 8200
rect 20621 8195 20687 8198
rect 25129 8195 25195 8198
rect 39021 8258 39087 8261
rect 40880 8258 41000 8288
rect 39021 8256 41000 8258
rect 39021 8200 39026 8256
rect 39082 8200 41000 8256
rect 39021 8198 41000 8200
rect 39021 8195 39087 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 14365 8122 14431 8125
rect 17217 8122 17283 8125
rect 24393 8122 24459 8125
rect 14365 8120 17283 8122
rect 14365 8064 14370 8120
rect 14426 8064 17222 8120
rect 17278 8064 17283 8120
rect 14365 8062 17283 8064
rect 14365 8059 14431 8062
rect 17217 8059 17283 8062
rect 20486 8120 24459 8122
rect 20486 8064 24398 8120
rect 24454 8064 24459 8120
rect 20486 8062 24459 8064
rect 0 7986 120 8016
rect 381 7986 447 7989
rect 0 7984 447 7986
rect 0 7928 386 7984
rect 442 7928 447 7984
rect 0 7926 447 7928
rect 0 7896 120 7926
rect 381 7923 447 7926
rect 7649 7986 7715 7989
rect 9121 7986 9187 7989
rect 7649 7984 9187 7986
rect 7649 7928 7654 7984
rect 7710 7928 9126 7984
rect 9182 7928 9187 7984
rect 7649 7926 9187 7928
rect 7649 7923 7715 7926
rect 9121 7923 9187 7926
rect 11053 7986 11119 7989
rect 20486 7986 20546 8062
rect 24393 8059 24459 8062
rect 37273 7986 37339 7989
rect 11053 7984 20546 7986
rect 11053 7928 11058 7984
rect 11114 7928 20546 7984
rect 11053 7926 20546 7928
rect 20670 7984 37339 7986
rect 20670 7928 37278 7984
rect 37334 7928 37339 7984
rect 20670 7926 37339 7928
rect 11053 7923 11119 7926
rect 6729 7850 6795 7853
rect 13721 7850 13787 7853
rect 6729 7848 13787 7850
rect 6729 7792 6734 7848
rect 6790 7792 13726 7848
rect 13782 7792 13787 7848
rect 6729 7790 13787 7792
rect 6729 7787 6795 7790
rect 13721 7787 13787 7790
rect 14641 7850 14707 7853
rect 20670 7850 20730 7926
rect 37273 7923 37339 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 25497 7850 25563 7853
rect 14641 7848 20730 7850
rect 14641 7792 14646 7848
rect 14702 7792 20730 7848
rect 14641 7790 20730 7792
rect 20854 7848 25563 7850
rect 20854 7792 25502 7848
rect 25558 7792 25563 7848
rect 20854 7790 25563 7792
rect 14641 7787 14707 7790
rect 0 7714 120 7744
rect 749 7714 815 7717
rect 14365 7714 14431 7717
rect 0 7712 815 7714
rect 0 7656 754 7712
rect 810 7656 815 7712
rect 0 7654 815 7656
rect 0 7624 120 7654
rect 749 7651 815 7654
rect 9446 7712 14431 7714
rect 9446 7656 14370 7712
rect 14426 7656 14431 7712
rect 9446 7654 14431 7656
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 0 7442 120 7472
rect 841 7442 907 7445
rect 0 7440 907 7442
rect 0 7384 846 7440
rect 902 7384 907 7440
rect 0 7382 907 7384
rect 0 7352 120 7382
rect 841 7379 907 7382
rect 7281 7442 7347 7445
rect 9446 7442 9506 7654
rect 14365 7651 14431 7654
rect 17217 7714 17283 7717
rect 20854 7714 20914 7790
rect 25497 7787 25563 7790
rect 17217 7712 20914 7714
rect 17217 7656 17222 7712
rect 17278 7656 20914 7712
rect 17217 7654 20914 7656
rect 39481 7714 39547 7717
rect 40880 7714 41000 7744
rect 39481 7712 41000 7714
rect 39481 7656 39486 7712
rect 39542 7656 41000 7712
rect 39481 7654 41000 7656
rect 17217 7651 17283 7654
rect 39481 7651 39547 7654
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 15561 7578 15627 7581
rect 20345 7578 20411 7581
rect 15561 7576 20411 7578
rect 15561 7520 15566 7576
rect 15622 7520 20350 7576
rect 20406 7520 20411 7576
rect 15561 7518 20411 7520
rect 15561 7515 15627 7518
rect 20345 7515 20411 7518
rect 21541 7578 21607 7581
rect 26601 7578 26667 7581
rect 21541 7576 26667 7578
rect 21541 7520 21546 7576
rect 21602 7520 26606 7576
rect 26662 7520 26667 7576
rect 21541 7518 26667 7520
rect 21541 7515 21607 7518
rect 26601 7515 26667 7518
rect 7281 7440 9506 7442
rect 7281 7384 7286 7440
rect 7342 7384 9506 7440
rect 7281 7382 9506 7384
rect 11145 7442 11211 7445
rect 23841 7442 23907 7445
rect 11145 7440 23907 7442
rect 11145 7384 11150 7440
rect 11206 7384 23846 7440
rect 23902 7384 23907 7440
rect 11145 7382 23907 7384
rect 7281 7379 7347 7382
rect 11145 7379 11211 7382
rect 23841 7379 23907 7382
rect 24710 7380 24716 7444
rect 24780 7442 24786 7444
rect 29913 7442 29979 7445
rect 24780 7440 29979 7442
rect 24780 7384 29918 7440
rect 29974 7384 29979 7440
rect 24780 7382 29979 7384
rect 24780 7380 24786 7382
rect 29913 7379 29979 7382
rect 39389 7442 39455 7445
rect 40880 7442 41000 7472
rect 39389 7440 41000 7442
rect 39389 7384 39394 7440
rect 39450 7384 41000 7440
rect 39389 7382 41000 7384
rect 39389 7379 39455 7382
rect 40880 7352 41000 7382
rect 1577 7306 1643 7309
rect 7833 7306 7899 7309
rect 1577 7304 7899 7306
rect 1577 7248 1582 7304
rect 1638 7248 7838 7304
rect 7894 7248 7899 7304
rect 1577 7246 7899 7248
rect 1577 7243 1643 7246
rect 7833 7243 7899 7246
rect 10869 7306 10935 7309
rect 38101 7306 38167 7309
rect 10869 7304 38167 7306
rect 10869 7248 10874 7304
rect 10930 7248 38106 7304
rect 38162 7248 38167 7304
rect 10869 7246 38167 7248
rect 10869 7243 10935 7246
rect 38101 7243 38167 7246
rect 0 7170 120 7200
rect 749 7170 815 7173
rect 0 7168 815 7170
rect 0 7112 754 7168
rect 810 7112 815 7168
rect 0 7110 815 7112
rect 0 7080 120 7110
rect 749 7107 815 7110
rect 15285 7170 15351 7173
rect 18321 7170 18387 7173
rect 15285 7168 18387 7170
rect 15285 7112 15290 7168
rect 15346 7112 18326 7168
rect 18382 7112 18387 7168
rect 15285 7110 18387 7112
rect 15285 7107 15351 7110
rect 18321 7107 18387 7110
rect 20621 7170 20687 7173
rect 24761 7170 24827 7173
rect 20621 7168 24827 7170
rect 20621 7112 20626 7168
rect 20682 7112 24766 7168
rect 24822 7112 24827 7168
rect 20621 7110 24827 7112
rect 20621 7107 20687 7110
rect 24761 7107 24827 7110
rect 28349 7170 28415 7173
rect 28901 7170 28967 7173
rect 28349 7168 28967 7170
rect 28349 7112 28354 7168
rect 28410 7112 28906 7168
rect 28962 7112 28967 7168
rect 28349 7110 28967 7112
rect 28349 7107 28415 7110
rect 28901 7107 28967 7110
rect 39573 7170 39639 7173
rect 40880 7170 41000 7200
rect 39573 7168 41000 7170
rect 39573 7112 39578 7168
rect 39634 7112 41000 7168
rect 39573 7110 41000 7112
rect 39573 7107 39639 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 20345 7034 20411 7037
rect 29913 7034 29979 7037
rect 20345 7032 25882 7034
rect 20345 6976 20350 7032
rect 20406 6976 25882 7032
rect 20345 6974 25882 6976
rect 20345 6971 20411 6974
rect 0 6898 120 6928
rect 749 6898 815 6901
rect 0 6896 815 6898
rect 0 6840 754 6896
rect 810 6840 815 6896
rect 0 6838 815 6840
rect 0 6808 120 6838
rect 749 6835 815 6838
rect 7465 6898 7531 6901
rect 25313 6898 25379 6901
rect 7465 6896 25379 6898
rect 7465 6840 7470 6896
rect 7526 6840 25318 6896
rect 25374 6840 25379 6896
rect 7465 6838 25379 6840
rect 25822 6898 25882 6974
rect 26374 7032 29979 7034
rect 26374 6976 29918 7032
rect 29974 6976 29979 7032
rect 26374 6974 29979 6976
rect 26374 6898 26434 6974
rect 29913 6971 29979 6974
rect 25822 6838 26434 6898
rect 26877 6898 26943 6901
rect 28257 6898 28323 6901
rect 26877 6896 28323 6898
rect 26877 6840 26882 6896
rect 26938 6840 28262 6896
rect 28318 6840 28323 6896
rect 26877 6838 28323 6840
rect 7465 6835 7531 6838
rect 25313 6835 25379 6838
rect 26877 6835 26943 6838
rect 28257 6835 28323 6838
rect 37222 6836 37228 6900
rect 37292 6898 37298 6900
rect 38193 6898 38259 6901
rect 37292 6896 38259 6898
rect 37292 6840 38198 6896
rect 38254 6840 38259 6896
rect 37292 6838 38259 6840
rect 37292 6836 37298 6838
rect 38193 6835 38259 6838
rect 39297 6898 39363 6901
rect 40880 6898 41000 6928
rect 39297 6896 41000 6898
rect 39297 6840 39302 6896
rect 39358 6840 41000 6896
rect 39297 6838 41000 6840
rect 39297 6835 39363 6838
rect 40880 6808 41000 6838
rect 12709 6762 12775 6765
rect 38837 6762 38903 6765
rect 12709 6760 38903 6762
rect 12709 6704 12714 6760
rect 12770 6704 38842 6760
rect 38898 6704 38903 6760
rect 12709 6702 38903 6704
rect 12709 6699 12775 6702
rect 38837 6699 38903 6702
rect 0 6626 120 6656
rect 841 6626 907 6629
rect 0 6624 907 6626
rect 0 6568 846 6624
rect 902 6568 907 6624
rect 0 6566 907 6568
rect 0 6536 120 6566
rect 841 6563 907 6566
rect 27797 6626 27863 6629
rect 28625 6626 28691 6629
rect 27797 6624 28691 6626
rect 27797 6568 27802 6624
rect 27858 6568 28630 6624
rect 28686 6568 28691 6624
rect 27797 6566 28691 6568
rect 27797 6563 27863 6566
rect 28625 6563 28691 6566
rect 39389 6626 39455 6629
rect 40880 6626 41000 6656
rect 39389 6624 41000 6626
rect 39389 6568 39394 6624
rect 39450 6568 41000 6624
rect 39389 6566 41000 6568
rect 39389 6563 39455 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 9397 6492 9463 6493
rect 9397 6488 9444 6492
rect 9508 6490 9514 6492
rect 16389 6490 16455 6493
rect 20713 6490 20779 6493
rect 9397 6432 9402 6488
rect 9397 6428 9444 6432
rect 9508 6430 9554 6490
rect 16389 6488 20779 6490
rect 16389 6432 16394 6488
rect 16450 6432 20718 6488
rect 20774 6432 20779 6488
rect 16389 6430 20779 6432
rect 9508 6428 9514 6430
rect 9397 6427 9463 6428
rect 16389 6427 16455 6430
rect 20713 6427 20779 6430
rect 27889 6490 27955 6493
rect 28717 6490 28783 6493
rect 38745 6490 38811 6493
rect 27889 6488 28783 6490
rect 27889 6432 27894 6488
rect 27950 6432 28722 6488
rect 28778 6432 28783 6488
rect 27889 6430 28783 6432
rect 27889 6427 27955 6430
rect 28717 6427 28783 6430
rect 35206 6488 38811 6490
rect 35206 6432 38750 6488
rect 38806 6432 38811 6488
rect 35206 6430 38811 6432
rect 0 6354 120 6384
rect 1025 6354 1091 6357
rect 0 6352 1091 6354
rect 0 6296 1030 6352
rect 1086 6296 1091 6352
rect 0 6294 1091 6296
rect 0 6264 120 6294
rect 1025 6291 1091 6294
rect 3877 6354 3943 6357
rect 15009 6354 15075 6357
rect 3877 6352 15075 6354
rect 3877 6296 3882 6352
rect 3938 6296 15014 6352
rect 15070 6296 15075 6352
rect 3877 6294 15075 6296
rect 3877 6291 3943 6294
rect 15009 6291 15075 6294
rect 15193 6354 15259 6357
rect 35206 6354 35266 6430
rect 38745 6427 38811 6430
rect 15193 6352 35266 6354
rect 15193 6296 15198 6352
rect 15254 6296 35266 6352
rect 15193 6294 35266 6296
rect 38653 6354 38719 6357
rect 40880 6354 41000 6384
rect 38653 6352 41000 6354
rect 38653 6296 38658 6352
rect 38714 6296 41000 6352
rect 38653 6294 41000 6296
rect 15193 6291 15259 6294
rect 38653 6291 38719 6294
rect 40880 6264 41000 6294
rect 2773 6218 2839 6221
rect 38469 6218 38535 6221
rect 2773 6216 38535 6218
rect 2773 6160 2778 6216
rect 2834 6160 38474 6216
rect 38530 6160 38535 6216
rect 2773 6158 38535 6160
rect 2773 6155 2839 6158
rect 38469 6155 38535 6158
rect 0 6082 120 6112
rect 197 6082 263 6085
rect 0 6080 263 6082
rect 0 6024 202 6080
rect 258 6024 263 6080
rect 0 6022 263 6024
rect 0 5992 120 6022
rect 197 6019 263 6022
rect 9213 6082 9279 6085
rect 13813 6082 13879 6085
rect 9213 6080 13879 6082
rect 9213 6024 9218 6080
rect 9274 6024 13818 6080
rect 13874 6024 13879 6080
rect 9213 6022 13879 6024
rect 9213 6019 9279 6022
rect 13813 6019 13879 6022
rect 38653 6082 38719 6085
rect 40880 6082 41000 6112
rect 38653 6080 41000 6082
rect 38653 6024 38658 6080
rect 38714 6024 41000 6080
rect 38653 6022 41000 6024
rect 38653 6019 38719 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 20713 5946 20779 5949
rect 25497 5946 25563 5949
rect 20713 5944 25563 5946
rect 20713 5888 20718 5944
rect 20774 5888 25502 5944
rect 25558 5888 25563 5944
rect 20713 5886 25563 5888
rect 20713 5883 20779 5886
rect 25497 5883 25563 5886
rect 0 5810 120 5840
rect 841 5810 907 5813
rect 0 5808 907 5810
rect 0 5752 846 5808
rect 902 5752 907 5808
rect 0 5750 907 5752
rect 0 5720 120 5750
rect 841 5747 907 5750
rect 5257 5810 5323 5813
rect 6545 5810 6611 5813
rect 5257 5808 6611 5810
rect 5257 5752 5262 5808
rect 5318 5752 6550 5808
rect 6606 5752 6611 5808
rect 5257 5750 6611 5752
rect 5257 5747 5323 5750
rect 6545 5747 6611 5750
rect 7833 5810 7899 5813
rect 39205 5810 39271 5813
rect 7833 5808 39271 5810
rect 7833 5752 7838 5808
rect 7894 5752 39210 5808
rect 39266 5752 39271 5808
rect 7833 5750 39271 5752
rect 7833 5747 7899 5750
rect 39205 5747 39271 5750
rect 39389 5810 39455 5813
rect 40880 5810 41000 5840
rect 39389 5808 41000 5810
rect 39389 5752 39394 5808
rect 39450 5752 41000 5808
rect 39389 5750 41000 5752
rect 39389 5747 39455 5750
rect 40880 5720 41000 5750
rect 3141 5674 3207 5677
rect 5993 5674 6059 5677
rect 3141 5672 6059 5674
rect 3141 5616 3146 5672
rect 3202 5616 5998 5672
rect 6054 5616 6059 5672
rect 3141 5614 6059 5616
rect 3141 5611 3207 5614
rect 5993 5611 6059 5614
rect 6269 5674 6335 5677
rect 10133 5674 10199 5677
rect 6269 5672 10199 5674
rect 6269 5616 6274 5672
rect 6330 5616 10138 5672
rect 10194 5616 10199 5672
rect 6269 5614 10199 5616
rect 6269 5611 6335 5614
rect 10133 5611 10199 5614
rect 13721 5674 13787 5677
rect 38561 5674 38627 5677
rect 13721 5672 38627 5674
rect 13721 5616 13726 5672
rect 13782 5616 38566 5672
rect 38622 5616 38627 5672
rect 13721 5614 38627 5616
rect 13721 5611 13787 5614
rect 38561 5611 38627 5614
rect 0 5538 120 5568
rect 749 5538 815 5541
rect 0 5536 815 5538
rect 0 5480 754 5536
rect 810 5480 815 5536
rect 0 5478 815 5480
rect 0 5448 120 5478
rect 749 5475 815 5478
rect 9489 5538 9555 5541
rect 14549 5538 14615 5541
rect 9489 5536 14615 5538
rect 9489 5480 9494 5536
rect 9550 5480 14554 5536
rect 14610 5480 14615 5536
rect 9489 5478 14615 5480
rect 9489 5475 9555 5478
rect 14549 5475 14615 5478
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 39941 5475 40007 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 20805 5402 20871 5405
rect 27429 5402 27495 5405
rect 32857 5402 32923 5405
rect 17726 5400 20871 5402
rect 17726 5344 20810 5400
rect 20866 5344 20871 5400
rect 17726 5342 20871 5344
rect 0 5266 120 5296
rect 841 5266 907 5269
rect 0 5264 907 5266
rect 0 5208 846 5264
rect 902 5208 907 5264
rect 0 5206 907 5208
rect 0 5176 120 5206
rect 841 5203 907 5206
rect 13537 5266 13603 5269
rect 17726 5266 17786 5342
rect 20805 5339 20871 5342
rect 21406 5342 26802 5402
rect 13537 5264 17786 5266
rect 13537 5208 13542 5264
rect 13598 5208 17786 5264
rect 13537 5206 17786 5208
rect 17953 5266 18019 5269
rect 21406 5266 21466 5342
rect 17953 5264 21466 5266
rect 17953 5208 17958 5264
rect 18014 5208 21466 5264
rect 17953 5206 21466 5208
rect 21541 5266 21607 5269
rect 26742 5266 26802 5342
rect 27429 5400 32923 5402
rect 27429 5344 27434 5400
rect 27490 5344 32862 5400
rect 32918 5344 32923 5400
rect 27429 5342 32923 5344
rect 27429 5339 27495 5342
rect 32857 5339 32923 5342
rect 39205 5266 39271 5269
rect 21541 5264 26618 5266
rect 21541 5208 21546 5264
rect 21602 5208 26618 5264
rect 21541 5206 26618 5208
rect 26742 5264 39271 5266
rect 26742 5208 39210 5264
rect 39266 5208 39271 5264
rect 26742 5206 39271 5208
rect 13537 5203 13603 5206
rect 17953 5203 18019 5206
rect 21541 5203 21607 5206
rect 13629 5130 13695 5133
rect 26558 5130 26618 5206
rect 39205 5203 39271 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 37825 5130 37891 5133
rect 13629 5128 26434 5130
rect 13629 5072 13634 5128
rect 13690 5072 26434 5128
rect 13629 5070 26434 5072
rect 26558 5128 37891 5130
rect 26558 5072 37830 5128
rect 37886 5072 37891 5128
rect 26558 5070 37891 5072
rect 13629 5067 13695 5070
rect 0 4994 120 5024
rect 749 4994 815 4997
rect 0 4992 815 4994
rect 0 4936 754 4992
rect 810 4936 815 4992
rect 0 4934 815 4936
rect 0 4904 120 4934
rect 749 4931 815 4934
rect 20805 4994 20871 4997
rect 21541 4994 21607 4997
rect 20805 4992 21607 4994
rect 20805 4936 20810 4992
rect 20866 4936 21546 4992
rect 21602 4936 21607 4992
rect 20805 4934 21607 4936
rect 26374 4994 26434 5070
rect 37825 5067 37891 5070
rect 27429 4994 27495 4997
rect 26374 4992 27495 4994
rect 26374 4936 27434 4992
rect 27490 4936 27495 4992
rect 26374 4934 27495 4936
rect 20805 4931 20871 4934
rect 21541 4931 21607 4934
rect 27429 4931 27495 4934
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 14549 4858 14615 4861
rect 18873 4858 18939 4861
rect 14549 4856 18939 4858
rect 14549 4800 14554 4856
rect 14610 4800 18878 4856
rect 18934 4800 18939 4856
rect 14549 4798 18939 4800
rect 14549 4795 14615 4798
rect 18873 4795 18939 4798
rect 0 4722 120 4752
rect 565 4722 631 4725
rect 0 4720 631 4722
rect 0 4664 570 4720
rect 626 4664 631 4720
rect 0 4662 631 4664
rect 0 4632 120 4662
rect 565 4659 631 4662
rect 13629 4722 13695 4725
rect 38837 4722 38903 4725
rect 13629 4720 38903 4722
rect 13629 4664 13634 4720
rect 13690 4664 38842 4720
rect 38898 4664 38903 4720
rect 13629 4662 38903 4664
rect 13629 4659 13695 4662
rect 38837 4659 38903 4662
rect 39389 4722 39455 4725
rect 40880 4722 41000 4752
rect 39389 4720 41000 4722
rect 39389 4664 39394 4720
rect 39450 4664 41000 4720
rect 39389 4662 41000 4664
rect 39389 4659 39455 4662
rect 40880 4632 41000 4662
rect 3601 4586 3667 4589
rect 8293 4586 8359 4589
rect 3601 4584 8359 4586
rect 3601 4528 3606 4584
rect 3662 4528 8298 4584
rect 8354 4528 8359 4584
rect 3601 4526 8359 4528
rect 3601 4523 3667 4526
rect 8293 4523 8359 4526
rect 8845 4586 8911 4589
rect 38469 4586 38535 4589
rect 8845 4584 38535 4586
rect 8845 4528 8850 4584
rect 8906 4528 38474 4584
rect 38530 4528 38535 4584
rect 8845 4526 38535 4528
rect 8845 4523 8911 4526
rect 38469 4523 38535 4526
rect 0 4450 120 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 120 4390
rect 1301 4387 1367 4390
rect 39573 4450 39639 4453
rect 40880 4450 41000 4480
rect 39573 4448 41000 4450
rect 39573 4392 39578 4448
rect 39634 4392 41000 4448
rect 39573 4390 41000 4392
rect 39573 4387 39639 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 0 4178 120 4208
rect 7649 4178 7715 4181
rect 0 4176 7715 4178
rect 0 4120 7654 4176
rect 7710 4120 7715 4176
rect 0 4118 7715 4120
rect 0 4088 120 4118
rect 7649 4115 7715 4118
rect 9438 4116 9444 4180
rect 9508 4178 9514 4180
rect 27797 4178 27863 4181
rect 9508 4176 27863 4178
rect 9508 4120 27802 4176
rect 27858 4120 27863 4176
rect 9508 4118 27863 4120
rect 9508 4116 9514 4118
rect 27797 4115 27863 4118
rect 32857 4178 32923 4181
rect 38745 4178 38811 4181
rect 32857 4176 38811 4178
rect 32857 4120 32862 4176
rect 32918 4120 38750 4176
rect 38806 4120 38811 4176
rect 32857 4118 38811 4120
rect 32857 4115 32923 4118
rect 38745 4115 38811 4118
rect 39021 4178 39087 4181
rect 40880 4178 41000 4208
rect 39021 4176 41000 4178
rect 39021 4120 39026 4176
rect 39082 4120 41000 4176
rect 39021 4118 41000 4120
rect 39021 4115 39087 4118
rect 40880 4088 41000 4118
rect 10777 4042 10843 4045
rect 38837 4042 38903 4045
rect 10777 4040 38903 4042
rect 10777 3984 10782 4040
rect 10838 3984 38842 4040
rect 38898 3984 38903 4040
rect 10777 3982 38903 3984
rect 10777 3979 10843 3982
rect 38837 3979 38903 3982
rect 0 3906 120 3936
rect 289 3906 355 3909
rect 0 3904 355 3906
rect 0 3848 294 3904
rect 350 3848 355 3904
rect 0 3846 355 3848
rect 0 3816 120 3846
rect 289 3843 355 3846
rect 39389 3906 39455 3909
rect 40880 3906 41000 3936
rect 39389 3904 41000 3906
rect 39389 3848 39394 3904
rect 39450 3848 41000 3904
rect 39389 3846 41000 3848
rect 39389 3843 39455 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 0 3634 120 3664
rect 473 3634 539 3637
rect 0 3632 539 3634
rect 0 3576 478 3632
rect 534 3576 539 3632
rect 0 3574 539 3576
rect 0 3544 120 3574
rect 473 3571 539 3574
rect 8661 3634 8727 3637
rect 38653 3634 38719 3637
rect 40880 3634 41000 3664
rect 8661 3632 35266 3634
rect 8661 3576 8666 3632
rect 8722 3576 35266 3632
rect 8661 3574 35266 3576
rect 8661 3571 8727 3574
rect 5809 3498 5875 3501
rect 35206 3498 35266 3574
rect 38653 3632 41000 3634
rect 38653 3576 38658 3632
rect 38714 3576 41000 3632
rect 38653 3574 41000 3576
rect 38653 3571 38719 3574
rect 40880 3544 41000 3574
rect 38837 3498 38903 3501
rect 5809 3496 35082 3498
rect 5809 3440 5814 3496
rect 5870 3440 35082 3496
rect 5809 3438 35082 3440
rect 35206 3496 38903 3498
rect 35206 3440 38842 3496
rect 38898 3440 38903 3496
rect 35206 3438 38903 3440
rect 5809 3435 5875 3438
rect 0 3362 120 3392
rect 1025 3362 1091 3365
rect 0 3360 1091 3362
rect 0 3304 1030 3360
rect 1086 3304 1091 3360
rect 0 3302 1091 3304
rect 35022 3362 35082 3438
rect 38837 3435 38903 3438
rect 37549 3362 37615 3365
rect 35022 3360 37615 3362
rect 35022 3304 37554 3360
rect 37610 3304 37615 3360
rect 35022 3302 37615 3304
rect 0 3272 120 3302
rect 1025 3299 1091 3302
rect 37549 3299 37615 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 22001 3226 22067 3229
rect 25037 3226 25103 3229
rect 22001 3224 25103 3226
rect 22001 3168 22006 3224
rect 22062 3168 25042 3224
rect 25098 3168 25103 3224
rect 22001 3166 25103 3168
rect 22001 3163 22067 3166
rect 25037 3163 25103 3166
rect 0 3090 120 3120
rect 3509 3090 3575 3093
rect 38469 3090 38535 3093
rect 0 3030 3434 3090
rect 0 3000 120 3030
rect 3374 2954 3434 3030
rect 3509 3088 38535 3090
rect 3509 3032 3514 3088
rect 3570 3032 38474 3088
rect 38530 3032 38535 3088
rect 3509 3030 38535 3032
rect 3509 3027 3575 3030
rect 38469 3027 38535 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 6177 2954 6243 2957
rect 8569 2954 8635 2957
rect 1350 2894 2790 2954
rect 3374 2952 6243 2954
rect 3374 2896 6182 2952
rect 6238 2896 6243 2952
rect 3374 2894 6243 2896
rect 0 2818 120 2848
rect 1350 2818 1410 2894
rect 0 2758 1410 2818
rect 2730 2818 2790 2894
rect 6177 2891 6243 2894
rect 6318 2952 8635 2954
rect 6318 2896 8574 2952
rect 8630 2896 8635 2952
rect 6318 2894 8635 2896
rect 6318 2818 6378 2894
rect 8569 2891 8635 2894
rect 12157 2954 12223 2957
rect 36721 2954 36787 2957
rect 12157 2952 36787 2954
rect 12157 2896 12162 2952
rect 12218 2896 36726 2952
rect 36782 2896 36787 2952
rect 12157 2894 36787 2896
rect 12157 2891 12223 2894
rect 36721 2891 36787 2894
rect 2730 2758 6378 2818
rect 20437 2818 20503 2821
rect 23289 2818 23355 2821
rect 20437 2816 23355 2818
rect 20437 2760 20442 2816
rect 20498 2760 23294 2816
rect 23350 2760 23355 2816
rect 20437 2758 23355 2760
rect 0 2728 120 2758
rect 20437 2755 20503 2758
rect 23289 2755 23355 2758
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 39021 2755 39087 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 0 2546 120 2576
rect 381 2546 447 2549
rect 0 2544 447 2546
rect 0 2488 386 2544
rect 442 2488 447 2544
rect 0 2486 447 2488
rect 0 2456 120 2486
rect 381 2483 447 2486
rect 6453 2546 6519 2549
rect 38653 2546 38719 2549
rect 40880 2546 41000 2576
rect 6453 2544 35450 2546
rect 6453 2488 6458 2544
rect 6514 2488 35450 2544
rect 6453 2486 35450 2488
rect 6453 2483 6519 2486
rect 33501 2410 33567 2413
rect 2730 2408 33567 2410
rect 2730 2352 33506 2408
rect 33562 2352 33567 2408
rect 2730 2350 33567 2352
rect 35390 2410 35450 2486
rect 38653 2544 41000 2546
rect 38653 2488 38658 2544
rect 38714 2488 41000 2544
rect 38653 2486 41000 2488
rect 38653 2483 38719 2486
rect 40880 2456 41000 2486
rect 39205 2410 39271 2413
rect 35390 2408 39271 2410
rect 35390 2352 39210 2408
rect 39266 2352 39271 2408
rect 35390 2350 39271 2352
rect 0 2274 120 2304
rect 2730 2274 2790 2350
rect 33501 2347 33567 2350
rect 39205 2347 39271 2350
rect 0 2214 2790 2274
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 0 2184 120 2214
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 1117 2002 1183 2005
rect 0 2000 1183 2002
rect 0 1944 1122 2000
rect 1178 1944 1183 2000
rect 0 1942 1183 1944
rect 0 1912 120 1942
rect 1117 1939 1183 1942
rect 13077 2002 13143 2005
rect 26325 2002 26391 2005
rect 13077 2000 26391 2002
rect 13077 1944 13082 2000
rect 13138 1944 26330 2000
rect 26386 1944 26391 2000
rect 13077 1942 26391 1944
rect 13077 1939 13143 1942
rect 26325 1939 26391 1942
rect 37917 2002 37983 2005
rect 40880 2002 41000 2032
rect 37917 2000 41000 2002
rect 37917 1944 37922 2000
rect 37978 1944 41000 2000
rect 37917 1942 41000 1944
rect 37917 1939 37983 1942
rect 40880 1912 41000 1942
rect 0 1730 120 1760
rect 32765 1730 32831 1733
rect 0 1728 32831 1730
rect 0 1672 32770 1728
rect 32826 1672 32831 1728
rect 0 1670 32831 1672
rect 0 1640 120 1670
rect 32765 1667 32831 1670
rect 38285 1730 38351 1733
rect 40880 1730 41000 1760
rect 38285 1728 41000 1730
rect 38285 1672 38290 1728
rect 38346 1672 41000 1728
rect 38285 1670 41000 1672
rect 38285 1667 38351 1670
rect 40880 1640 41000 1670
rect 0 1458 120 1488
rect 1209 1458 1275 1461
rect 0 1456 1275 1458
rect 0 1400 1214 1456
rect 1270 1400 1275 1456
rect 0 1398 1275 1400
rect 0 1368 120 1398
rect 1209 1395 1275 1398
rect 38653 1458 38719 1461
rect 40880 1458 41000 1488
rect 38653 1456 41000 1458
rect 38653 1400 38658 1456
rect 38714 1400 41000 1456
rect 38653 1398 41000 1400
rect 38653 1395 38719 1398
rect 40880 1368 41000 1398
rect 28809 370 28875 373
rect 39573 370 39639 373
rect 28809 368 39639 370
rect 28809 312 28814 368
rect 28870 312 39578 368
rect 39634 312 39639 368
rect 28809 310 39639 312
rect 28809 307 28875 310
rect 39573 307 39639 310
rect 21909 234 21975 237
rect 35985 234 36051 237
rect 21909 232 36051 234
rect 21909 176 21914 232
rect 21970 176 35990 232
rect 36046 176 36051 232
rect 21909 174 36051 176
rect 21909 171 21975 174
rect 35985 171 36051 174
rect 17493 98 17559 101
rect 34513 98 34579 101
rect 17493 96 34579 98
rect 17493 40 17498 96
rect 17554 40 34518 96
rect 34574 40 34579 96
rect 17493 38 34579 40
rect 17493 35 17559 38
rect 34513 35 34579 38
<< via3 >>
rect 37228 9420 37292 9484
rect 24716 9284 24780 9348
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 24716 7380 24780 7444
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 37228 6836 37292 6900
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 9444 6488 9508 6492
rect 9444 6432 9458 6488
rect 9458 6432 9508 6488
rect 9444 6428 9508 6432
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 9444 4116 9508 4180
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9446 4181 9506 6427
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 9443 4180 9509 4181
rect 9443 4116 9444 4180
rect 9508 4116 9509 4180
rect 9443 4115 9509 4116
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19944 0 20264 2688
rect 21004 8736 21324 11250
rect 24715 9348 24781 9349
rect 24715 9284 24716 9348
rect 24780 9284 24781 9348
rect 24715 9283 24781 9284
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 21004 6560 21324 7584
rect 24718 7445 24778 9283
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 24715 7444 24781 7445
rect 24715 7380 24716 7444
rect 24780 7380 24781 7444
rect 24715 7379 24781 7380
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 37227 9484 37293 9485
rect 37227 9420 37228 9484
rect 37292 9420 37293 9484
rect 37227 9419 37293 9420
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 37230 6901 37290 9419
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37227 6900 37293 6901
rect 37227 6836 37228 6900
rect 37292 6836 37293 6900
rect 37227 6835 37293 6836
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__inv_1  _030_
timestamp -3599
transform -1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _031_
timestamp -3599
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _032_
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp -3599
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _034_
timestamp -3599
transform -1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _035_
timestamp -3599
transform 1 0 5060 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _036_
timestamp -3599
transform -1 0 10856 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _037_
timestamp -3599
transform 1 0 10856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _038_
timestamp -3599
transform 1 0 10120 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _039_
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _040_
timestamp -3599
transform 1 0 9292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _041_
timestamp -3599
transform -1 0 21712 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _042_
timestamp -3599
transform -1 0 22172 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _043_
timestamp -3599
transform -1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _044_
timestamp -3599
transform 1 0 23000 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _045_
timestamp -3599
transform 1 0 20424 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _046_
timestamp -3599
transform 1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _047_
timestamp -3599
transform 1 0 27508 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _048_
timestamp -3599
transform 1 0 25944 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _049_
timestamp -3599
transform -1 0 27140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _050_
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _051_
timestamp -3599
transform 1 0 27140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _052_
timestamp -3599
transform 1 0 28704 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _053_
timestamp -3599
transform -1 0 23092 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _054_
timestamp -3599
transform -1 0 23552 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _055_
timestamp -3599
transform -1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _056_
timestamp -3599
transform 1 0 24104 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _057_
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _058_
timestamp -3599
transform 1 0 22540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _059_
timestamp -3599
transform 1 0 5060 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2b_1  _060_
timestamp -3599
transform -1 0 8556 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _061_
timestamp -3599
transform 1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _062_
timestamp -3599
transform 1 0 9200 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _063_
timestamp -3599
transform -1 0 8648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _064_
timestamp -3599
transform 1 0 6992 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _065_
timestamp -3599
transform 1 0 17480 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _066_
timestamp -3599
transform 1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp -3599
transform 1 0 14904 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp -3599
transform -1 0 15088 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dlxtp_1  _069_
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _070_
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _071_
timestamp -3599
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _072_
timestamp -3599
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _073_
timestamp -3599
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _074_
timestamp -3599
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _075_
timestamp -3599
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _076_
timestamp -3599
transform 1 0 17204 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _077_
timestamp -3599
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _078_
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _079_
timestamp -3599
transform 1 0 25208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _080_
timestamp -3599
transform 1 0 25024 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _081_
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _082_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _083_
timestamp -3599
transform 1 0 17940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _084_
timestamp -3599
transform 1 0 17848 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _085_
timestamp -3599
transform -1 0 13432 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _086_
timestamp -3599
transform -1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _087_
timestamp -3599
transform -1 0 10580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp -3599
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp -3599
transform -1 0 33120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp -3599
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp -3599
transform -1 0 33396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _093_
timestamp -3599
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _094_
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _095_
timestamp -3599
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp -3599
transform -1 0 30912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp -3599
transform 1 0 29072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp -3599
transform 1 0 30176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp -3599
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp -3599
transform -1 0 38456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp -3599
transform -1 0 38456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform 1 0 13432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_
timestamp -3599
transform 1 0 13432 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp -3599
transform 1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp -3599
transform -1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp -3599
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp -3599
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp -3599
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _110_
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp -3599
transform -1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp -3599
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _113_
timestamp -3599
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp -3599
transform 1 0 23552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _115_
timestamp -3599
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _116_
timestamp -3599
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _117_
timestamp -3599
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp -3599
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp -3599
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp -3599
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _121_
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp -3599
transform -1 0 26680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp -3599
transform 1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp -3599
transform -1 0 33488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp -3599
transform 1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp -3599
transform 1 0 34960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp -3599
transform 1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp -3599
transform 1 0 35696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp -3599
transform -1 0 29808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp -3599
transform -1 0 32752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp -3599
transform -1 0 34132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp -3599
transform 1 0 37628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp -3599
transform -1 0 29532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp -3599
transform 1 0 38364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp -3599
transform -1 0 37168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp -3599
transform 1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _137_
timestamp -3599
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp -3599
transform -1 0 33856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp -3599
transform -1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp -3599
transform -1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp -3599
transform -1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _142_
timestamp -3599
transform -1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp -3599
transform -1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp -3599
transform -1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp -3599
transform -1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp -3599
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp -3599
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp -3599
transform 1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp -3599
transform -1 0 22448 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp -3599
transform -1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp -3599
transform -1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp -3599
transform 1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _154_
timestamp -3599
transform -1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp -3599
transform -1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp -3599
transform -1 0 25208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp -3599
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp -3599
transform -1 0 24104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp -3599
transform -1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _160_
timestamp -3599
transform -1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp -3599
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp -3599
transform -1 0 39008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp -3599
transform -1 0 32568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp -3599
transform -1 0 37628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _165_
timestamp -3599
transform -1 0 35328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp -3599
transform -1 0 37628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp -3599
transform -1 0 32200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp -3599
transform -1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp -3599
transform -1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _170_
timestamp -3599
transform -1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp -3599
transform -1 0 29808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _172_
timestamp -3599
transform -1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp -3599
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp -3599
transform -1 0 22356 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _175_
timestamp -3599
transform -1 0 30176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp -3599
transform -1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _177_
timestamp -3599
transform -1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _178_
timestamp -3599
transform -1 0 34132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp -3599
transform -1 0 38364 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _180_
timestamp -3599
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp -3599
transform -1 0 37536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _182_
timestamp -3599
transform -1 0 30636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _183_
timestamp -3599
transform -1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _184_
timestamp -3599
transform -1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _185_
timestamp -3599
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp -3599
transform 1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _187_
timestamp -3599
transform -1 0 27968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp -3599
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _189_
timestamp -3599
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _191_
timestamp -3599
transform -1 0 27416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp -3599
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _193_
timestamp -3599
transform 1 0 32200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 38180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 32844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 33580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 29072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 29992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform 1 0 37996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 26220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 36156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 34960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 24840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout7
timestamp -3599
transform -1 0 17020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout8
timestamp -3599
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13
timestamp -3599
transform 1 0 2300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39
timestamp 1636964856
transform 1 0 4692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp -3599
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65
timestamp -3599
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71
timestamp 1636964856
transform 1 0 7636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp -3599
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89
timestamp 1636964856
transform 1 0 9292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101
timestamp -3599
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118
timestamp 1636964856
transform 1 0 11960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp -3599
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp -3599
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636964856
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636964856
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp -3599
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636964856
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp -3599
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636964856
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636964856
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636964856
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636964856
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_187
timestamp -3599
transform 1 0 18308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_195
timestamp -3599
transform 1 0 19044 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_211
timestamp -3599
transform 1 0 20516 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_219
timestamp -3599
transform 1 0 21252 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_247
timestamp -3599
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_265
timestamp -3599
transform 1 0 25484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp -3599
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_289
timestamp -3599
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_294
timestamp -3599
transform 1 0 28152 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_302
timestamp -3599
transform 1 0 28888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_312
timestamp -3599
transform 1 0 29808 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1636964856
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp -3599
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_342
timestamp 1636964856
transform 1 0 32568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_354
timestamp -3599
transform 1 0 33672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp -3599
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_363
timestamp -3599
transform 1 0 34500 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_367
timestamp 1636964856
transform 1 0 34868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_379
timestamp -3599
transform 1 0 35972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp -3599
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_401
timestamp -3599
transform 1 0 37996 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_41
timestamp -3599
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp -3599
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_52
timestamp 1636964856
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_64
timestamp 1636964856
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_76
timestamp -3599
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp -3599
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp -3599
transform 1 0 11868 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636964856
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636964856
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636964856
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636964856
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636964856
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636964856
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp -3599
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636964856
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636964856
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636964856
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636964856
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp -3599
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -3599
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636964856
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636964856
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636964856
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636964856
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp -3599
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636964856
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_401
timestamp -3599
transform 1 0 37996 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_409
timestamp -3599
transform 1 0 38732 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_23
timestamp -3599
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_30
timestamp 1636964856
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp -3599
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp -3599
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_93
timestamp -3599
transform 1 0 9660 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_137
timestamp -3599
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_152
timestamp 1636964856
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp -3599
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_173
timestamp -3599
transform 1 0 17020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_179
timestamp -3599
transform 1 0 17572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_183
timestamp 1636964856
transform 1 0 17940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_195
timestamp 1636964856
transform 1 0 19044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1636964856
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp -3599
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636964856
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636964856
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_261
timestamp -3599
transform 1 0 25116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_265
timestamp 1636964856
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp -3599
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_286
timestamp -3599
transform 1 0 27416 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_292
timestamp 1636964856
transform 1 0 27968 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1636964856
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1636964856
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp -3599
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_342
timestamp 1636964856
transform 1 0 32568 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_354
timestamp 1636964856
transform 1 0 33672 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_366
timestamp 1636964856
transform 1 0 34776 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_378
timestamp 1636964856
transform 1 0 35880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp -3599
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_397
timestamp -3599
transform 1 0 37628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_15
timestamp -3599
transform 1 0 2484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp -3599
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp -3599
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_107
timestamp 1636964856
transform 1 0 10948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_122
timestamp 1636964856
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp -3599
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_156
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_160
timestamp -3599
transform 1 0 15824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp -3599
transform 1 0 17296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_187
timestamp -3599
transform 1 0 18308 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp -3599
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_257
timestamp -3599
transform 1 0 24748 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_272
timestamp 1636964856
transform 1 0 26128 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_284
timestamp -3599
transform 1 0 27232 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_312
timestamp -3599
transform 1 0 29808 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_316
timestamp 1636964856
transform 1 0 30176 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_328
timestamp 1636964856
transform 1 0 31280 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_340
timestamp 1636964856
transform 1 0 32384 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_352
timestamp -3599
transform 1 0 33488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp -3599
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_371
timestamp -3599
transform 1 0 35236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_375
timestamp -3599
transform 1 0 35604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_379
timestamp -3599
transform 1 0 35972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_387
timestamp -3599
transform 1 0 36708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_392
timestamp -3599
transform 1 0 37168 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_400
timestamp -3599
transform 1 0 37904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_412
timestamp -3599
transform 1 0 39008 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_6
timestamp 1636964856
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_18
timestamp 1636964856
transform 1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_37
timestamp 1636964856
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp -3599
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_75
timestamp -3599
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_86
timestamp 1636964856
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_98
timestamp -3599
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp -3599
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636964856
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636964856
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636964856
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp -3599
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp -3599
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636964856
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636964856
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636964856
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp -3599
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636964856
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636964856
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636964856
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp -3599
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_344
timestamp -3599
transform 1 0 32752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_348
timestamp -3599
transform 1 0 33120 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_355
timestamp 1636964856
transform 1 0 33764 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_367
timestamp 1636964856
transform 1 0 34868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_379
timestamp 1636964856
transform 1 0 35972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp -3599
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_9
timestamp 1636964856
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_21
timestamp -3599
transform 1 0 3036 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp -3599
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_64
timestamp 1636964856
transform 1 0 6992 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp -3599
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636964856
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_105
timestamp -3599
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_114
timestamp -3599
transform 1 0 11592 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp -3599
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636964856
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636964856
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_165
timestamp -3599
transform 1 0 16284 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_171
timestamp -3599
transform 1 0 16836 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_181
timestamp 1636964856
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp -3599
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_205
timestamp -3599
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636964856
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636964856
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_233
timestamp -3599
transform 1 0 22540 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_241
timestamp -3599
transform 1 0 23276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp -3599
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_269
timestamp -3599
transform 1 0 25852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_291
timestamp -3599
transform 1 0 27876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_299
timestamp -3599
transform 1 0 28612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp -3599
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_312
timestamp 1636964856
transform 1 0 29808 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_324
timestamp 1636964856
transform 1 0 30912 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_336
timestamp 1636964856
transform 1 0 32016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_348
timestamp 1636964856
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp -3599
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636964856
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636964856
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_401
timestamp -3599
transform 1 0 37996 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_9
timestamp -3599
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1636964856
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_43
timestamp -3599
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp -3599
transform 1 0 5796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_62
timestamp 1636964856
transform 1 0 6808 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_74
timestamp 1636964856
transform 1 0 7912 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_86
timestamp -3599
transform 1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp -3599
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1636964856
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636964856
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636964856
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_137
timestamp -3599
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp -3599
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_175
timestamp -3599
transform 1 0 17204 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp -3599
transform 1 0 19320 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_231
timestamp 1636964856
transform 1 0 22356 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_243
timestamp 1636964856
transform 1 0 23460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_255
timestamp 1636964856
transform 1 0 24564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1636964856
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp -3599
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636964856
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_320
timestamp -3599
transform 1 0 30544 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_324
timestamp 1636964856
transform 1 0 30912 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_349
timestamp -3599
transform 1 0 33212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_355
timestamp -3599
transform 1 0 33764 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_359
timestamp 1636964856
transform 1 0 34132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_371
timestamp 1636964856
transform 1 0 35236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_383
timestamp -3599
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_400
timestamp -3599
transform 1 0 37904 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_12
timestamp 1636964856
transform 1 0 2208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp -3599
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636964856
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636964856
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_127
timestamp 1636964856
transform 1 0 12788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636964856
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636964856
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636964856
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp -3599
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636964856
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636964856
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636964856
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636964856
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp -3599
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_261
timestamp -3599
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_274
timestamp 1636964856
transform 1 0 26312 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636964856
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636964856
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636964856
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636964856
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_389
timestamp -3599
transform 1 0 36892 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_396
timestamp -3599
transform 1 0 37536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_400
timestamp -3599
transform 1 0 37904 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_12
timestamp 1636964856
transform 1 0 2208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1636964856
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1636964856
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_84
timestamp -3599
transform 1 0 8832 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_90
timestamp -3599
transform 1 0 9384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp -3599
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -3599
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_125
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp -3599
transform 1 0 13340 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_149
timestamp -3599
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_159
timestamp -3599
transform 1 0 15732 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_189
timestamp 1636964856
transform 1 0 18492 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_201
timestamp 1636964856
transform 1 0 19596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_213
timestamp -3599
transform 1 0 20700 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp -3599
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636964856
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636964856
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636964856
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp -3599
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_268
timestamp 1636964856
transform 1 0 25760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_305
timestamp -3599
transform 1 0 29164 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_313
timestamp -3599
transform 1 0 29900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_319
timestamp 1636964856
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp -3599
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp -3599
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636964856
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636964856
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1636964856
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636964856
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp -3599
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp -3599
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_397
timestamp -3599
transform 1 0 37628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp -3599
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp -3599
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp -3599
transform 1 0 8096 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp -3599
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_94
timestamp -3599
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp -3599
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp -3599
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_134
timestamp -3599
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_148
timestamp -3599
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp -3599
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_166
timestamp -3599
transform 1 0 16376 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_174
timestamp -3599
transform 1 0 17112 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp -3599
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_205
timestamp -3599
transform 1 0 19964 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_209
timestamp -3599
transform 1 0 20332 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_232
timestamp -3599
transform 1 0 22448 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp -3599
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_256
timestamp -3599
transform 1 0 24656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_264
timestamp -3599
transform 1 0 25392 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_268
timestamp 1636964856
transform 1 0 25760 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_280
timestamp -3599
transform 1 0 26864 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_285
timestamp 1636964856
transform 1 0 27324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_297
timestamp -3599
transform 1 0 28428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_301
timestamp -3599
transform 1 0 28796 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_312
timestamp 1636964856
transform 1 0 29808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_332
timestamp -3599
transform 1 0 31648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_338
timestamp -3599
transform 1 0 32200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_342
timestamp -3599
transform 1 0 32568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp -3599
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp -3599
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_372
timestamp -3599
transform 1 0 35328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_379
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_399
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_410
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp -3599
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp -3599
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_207
timestamp 1636964856
transform 1 0 20148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_271
timestamp -3599
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -3599
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp -3599
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_306
timestamp -3599
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_323
timestamp 1636964856
transform 1 0 30820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp -3599
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp -3599
transform 1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -3599
transform -1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -3599
transform 1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input13
timestamp -3599
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -3599
transform 1 0 2576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -3599
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp -3599
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp -3599
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -3599
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input22
timestamp -3599
transform 1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp -3599
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp -3599
transform -1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp -3599
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp -3599
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp -3599
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp -3599
transform -1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -3599
transform -1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -3599
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp -3599
transform -1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp -3599
transform -1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -3599
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp -3599
transform 1 0 19320 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp -3599
transform -1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp -3599
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp -3599
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp -3599
transform -1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp -3599
transform 1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp -3599
transform 1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp -3599
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp -3599
transform -1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp -3599
transform -1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp -3599
transform -1 0 28428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp -3599
transform -1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input50
timestamp -3599
transform -1 0 29256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp -3599
transform 1 0 28704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp -3599
transform -1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp -3599
transform -1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp -3599
transform -1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp -3599
transform 1 0 38456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp -3599
transform 1 0 38456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp -3599
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 38456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 38456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 35972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 36524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform -1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform -1 0 34408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform -1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform -1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform -1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform -1 0 3680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform -1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform -1 0 5060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform -1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform -1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform -1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform -1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform -1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform -1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform -1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform 1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform -1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform -1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform -1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform -1 0 13892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform -1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform -1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform -1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform -1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform -1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform -1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output163
timestamp -3599
transform -1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_WARMBOOT_164
timestamp -3599
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 2778 0 2834 56 0 FreeSans 224 0 0 0 BOOT_top
port 0 nsew signal output
flabel metal2 s 17590 11194 17646 11250 0 FreeSans 224 0 0 0 Co
port 1 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 2 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 3 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 4 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 5 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 6 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 7 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 8 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 9 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 10 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 11 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 12 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 13 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 14 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 15 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 16 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 17 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 18 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 19 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 20 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 21 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 22 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 23 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 24 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 25 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 26 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 27 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 28 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 29 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 30 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 31 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 32 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 33 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 34 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 35 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 36 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 37 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 38 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 39 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 40 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 41 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 42 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 43 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 44 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 45 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 46 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 47 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 48 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 49 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 50 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 51 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 52 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 53 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 54 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 55 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 56 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 57 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 58 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 59 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 60 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 61 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 62 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 63 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 64 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 65 nsew signal output
flabel metal2 s 11610 0 11666 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 66 nsew signal input
flabel metal2 s 26330 0 26386 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 67 nsew signal input
flabel metal2 s 27802 0 27858 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 68 nsew signal input
flabel metal2 s 29274 0 29330 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 69 nsew signal input
flabel metal2 s 30746 0 30802 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 70 nsew signal input
flabel metal2 s 32218 0 32274 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 71 nsew signal input
flabel metal2 s 33690 0 33746 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 72 nsew signal input
flabel metal2 s 35162 0 35218 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 73 nsew signal input
flabel metal2 s 36634 0 36690 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 74 nsew signal input
flabel metal2 s 38106 0 38162 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 75 nsew signal input
flabel metal2 s 39578 0 39634 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 76 nsew signal input
flabel metal2 s 13082 0 13138 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 77 nsew signal input
flabel metal2 s 14554 0 14610 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 78 nsew signal input
flabel metal2 s 16026 0 16082 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 79 nsew signal input
flabel metal2 s 17498 0 17554 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 80 nsew signal input
flabel metal2 s 18970 0 19026 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 81 nsew signal input
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 82 nsew signal input
flabel metal2 s 21914 0 21970 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 83 nsew signal input
flabel metal2 s 23386 0 23442 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 84 nsew signal input
flabel metal2 s 24858 0 24914 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 85 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 86 nsew signal output
flabel metal2 s 35254 11194 35310 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 87 nsew signal output
flabel metal2 s 35530 11194 35586 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 88 nsew signal output
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 89 nsew signal output
flabel metal2 s 36082 11194 36138 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 90 nsew signal output
flabel metal2 s 36358 11194 36414 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 91 nsew signal output
flabel metal2 s 36634 11194 36690 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 92 nsew signal output
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 93 nsew signal output
flabel metal2 s 37186 11194 37242 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 94 nsew signal output
flabel metal2 s 37462 11194 37518 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 95 nsew signal output
flabel metal2 s 37738 11194 37794 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 96 nsew signal output
flabel metal2 s 32770 11194 32826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 97 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 98 nsew signal output
flabel metal2 s 33322 11194 33378 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 99 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 100 nsew signal output
flabel metal2 s 33874 11194 33930 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 101 nsew signal output
flabel metal2 s 34150 11194 34206 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 102 nsew signal output
flabel metal2 s 34426 11194 34482 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 103 nsew signal output
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 104 nsew signal output
flabel metal2 s 34978 11194 35034 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 105 nsew signal output
flabel metal2 s 3238 11194 3294 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 106 nsew signal output
flabel metal2 s 3514 11194 3570 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 107 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 108 nsew signal output
flabel metal2 s 4066 11194 4122 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 109 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 110 nsew signal output
flabel metal2 s 4618 11194 4674 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 111 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 112 nsew signal output
flabel metal2 s 5170 11194 5226 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 113 nsew signal output
flabel metal2 s 5446 11194 5502 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 114 nsew signal output
flabel metal2 s 5722 11194 5778 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 115 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 116 nsew signal output
flabel metal2 s 6274 11194 6330 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 117 nsew signal output
flabel metal2 s 6550 11194 6606 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 118 nsew signal output
flabel metal2 s 6826 11194 6882 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 119 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 120 nsew signal output
flabel metal2 s 7378 11194 7434 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 121 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 122 nsew signal output
flabel metal2 s 7930 11194 7986 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 123 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 124 nsew signal output
flabel metal2 s 8482 11194 8538 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 125 nsew signal output
flabel metal2 s 8758 11194 8814 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 126 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 127 nsew signal output
flabel metal2 s 11794 11194 11850 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 128 nsew signal output
flabel metal2 s 12070 11194 12126 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 129 nsew signal output
flabel metal2 s 12346 11194 12402 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 130 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 131 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 132 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 133 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 134 nsew signal output
flabel metal2 s 9586 11194 9642 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 135 nsew signal output
flabel metal2 s 9862 11194 9918 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 136 nsew signal output
flabel metal2 s 10138 11194 10194 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 137 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 138 nsew signal output
flabel metal2 s 10690 11194 10746 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 139 nsew signal output
flabel metal2 s 10966 11194 11022 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 140 nsew signal output
flabel metal2 s 11242 11194 11298 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 141 nsew signal output
flabel metal2 s 13174 11194 13230 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 142 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 143 nsew signal output
flabel metal2 s 16210 11194 16266 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 144 nsew signal output
flabel metal2 s 16486 11194 16542 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 145 nsew signal output
flabel metal2 s 16762 11194 16818 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 146 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 147 nsew signal output
flabel metal2 s 17314 11194 17370 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 148 nsew signal output
flabel metal2 s 13450 11194 13506 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 149 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 150 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 151 nsew signal output
flabel metal2 s 14278 11194 14334 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 152 nsew signal output
flabel metal2 s 14554 11194 14610 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 153 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 154 nsew signal output
flabel metal2 s 15106 11194 15162 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 155 nsew signal output
flabel metal2 s 15382 11194 15438 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 156 nsew signal output
flabel metal2 s 15658 11194 15714 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 157 nsew signal output
flabel metal2 s 1306 0 1362 56 0 FreeSans 224 0 0 0 RESET_top
port 158 nsew signal input
flabel metal2 s 17866 11194 17922 11250 0 FreeSans 224 0 0 0 S1END[0]
port 159 nsew signal input
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 S1END[1]
port 160 nsew signal input
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 S1END[2]
port 161 nsew signal input
flabel metal2 s 18694 11194 18750 11250 0 FreeSans 224 0 0 0 S1END[3]
port 162 nsew signal input
flabel metal2 s 21178 11194 21234 11250 0 FreeSans 224 0 0 0 S2END[0]
port 163 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S2END[1]
port 164 nsew signal input
flabel metal2 s 21730 11194 21786 11250 0 FreeSans 224 0 0 0 S2END[2]
port 165 nsew signal input
flabel metal2 s 22006 11194 22062 11250 0 FreeSans 224 0 0 0 S2END[3]
port 166 nsew signal input
flabel metal2 s 22282 11194 22338 11250 0 FreeSans 224 0 0 0 S2END[4]
port 167 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2END[5]
port 168 nsew signal input
flabel metal2 s 22834 11194 22890 11250 0 FreeSans 224 0 0 0 S2END[6]
port 169 nsew signal input
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 S2END[7]
port 170 nsew signal input
flabel metal2 s 18970 11194 19026 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 171 nsew signal input
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 172 nsew signal input
flabel metal2 s 19522 11194 19578 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 173 nsew signal input
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 174 nsew signal input
flabel metal2 s 20074 11194 20130 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 175 nsew signal input
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 176 nsew signal input
flabel metal2 s 20626 11194 20682 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 177 nsew signal input
flabel metal2 s 20902 11194 20958 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 178 nsew signal input
flabel metal2 s 23386 11194 23442 11250 0 FreeSans 224 0 0 0 S4END[0]
port 179 nsew signal input
flabel metal2 s 26146 11194 26202 11250 0 FreeSans 224 0 0 0 S4END[10]
port 180 nsew signal input
flabel metal2 s 26422 11194 26478 11250 0 FreeSans 224 0 0 0 S4END[11]
port 181 nsew signal input
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 S4END[12]
port 182 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S4END[13]
port 183 nsew signal input
flabel metal2 s 27250 11194 27306 11250 0 FreeSans 224 0 0 0 S4END[14]
port 184 nsew signal input
flabel metal2 s 27526 11194 27582 11250 0 FreeSans 224 0 0 0 S4END[15]
port 185 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S4END[1]
port 186 nsew signal input
flabel metal2 s 23938 11194 23994 11250 0 FreeSans 224 0 0 0 S4END[2]
port 187 nsew signal input
flabel metal2 s 24214 11194 24270 11250 0 FreeSans 224 0 0 0 S4END[3]
port 188 nsew signal input
flabel metal2 s 24490 11194 24546 11250 0 FreeSans 224 0 0 0 S4END[4]
port 189 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S4END[5]
port 190 nsew signal input
flabel metal2 s 25042 11194 25098 11250 0 FreeSans 224 0 0 0 S4END[6]
port 191 nsew signal input
flabel metal2 s 25318 11194 25374 11250 0 FreeSans 224 0 0 0 S4END[7]
port 192 nsew signal input
flabel metal2 s 25594 11194 25650 11250 0 FreeSans 224 0 0 0 S4END[8]
port 193 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S4END[9]
port 194 nsew signal input
flabel metal2 s 4250 0 4306 56 0 FreeSans 224 0 0 0 SLOT_top0
port 195 nsew signal output
flabel metal2 s 5722 0 5778 56 0 FreeSans 224 0 0 0 SLOT_top1
port 196 nsew signal output
flabel metal2 s 7194 0 7250 56 0 FreeSans 224 0 0 0 SLOT_top2
port 197 nsew signal output
flabel metal2 s 8666 0 8722 56 0 FreeSans 224 0 0 0 SLOT_top3
port 198 nsew signal output
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 199 nsew signal input
flabel metal2 s 30562 11194 30618 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 200 nsew signal input
flabel metal2 s 30838 11194 30894 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 201 nsew signal input
flabel metal2 s 31114 11194 31170 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 202 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 203 nsew signal input
flabel metal2 s 31666 11194 31722 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 204 nsew signal input
flabel metal2 s 31942 11194 31998 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 205 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 206 nsew signal input
flabel metal2 s 28354 11194 28410 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 207 nsew signal input
flabel metal2 s 28630 11194 28686 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 208 nsew signal input
flabel metal2 s 28906 11194 28962 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 209 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 210 nsew signal input
flabel metal2 s 29458 11194 29514 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 211 nsew signal input
flabel metal2 s 29734 11194 29790 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 212 nsew signal input
flabel metal2 s 30010 11194 30066 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 213 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 214 nsew signal input
flabel metal2 s 10138 0 10194 56 0 FreeSans 224 0 0 0 UserCLK
port 215 nsew signal input
flabel metal2 s 32218 11194 32274 11250 0 FreeSans 224 0 0 0 UserCLKo
port 216 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 217 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 218 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal2 2806 1160 2806 1160 0 BOOT_top
rlabel metal3 666 1428 666 1428 0 FrameData[0]
rlabel metal1 9752 7990 9752 7990 0 FrameData[10]
rlabel metal3 712 4420 712 4420 0 FrameData[11]
rlabel metal3 344 4692 344 4692 0 FrameData[12]
rlabel metal3 436 4964 436 4964 0 FrameData[13]
rlabel metal3 482 5236 482 5236 0 FrameData[14]
rlabel metal3 436 5508 436 5508 0 FrameData[15]
rlabel metal3 482 5780 482 5780 0 FrameData[16]
rlabel metal3 160 6052 160 6052 0 FrameData[17]
rlabel metal3 574 6324 574 6324 0 FrameData[18]
rlabel metal3 482 6596 482 6596 0 FrameData[19]
rlabel metal1 32844 7854 32844 7854 0 FrameData[1]
rlabel metal3 436 6868 436 6868 0 FrameData[20]
rlabel metal3 436 7140 436 7140 0 FrameData[21]
rlabel metal3 482 7412 482 7412 0 FrameData[22]
rlabel metal3 436 7684 436 7684 0 FrameData[23]
rlabel metal3 252 7956 252 7956 0 FrameData[24]
rlabel metal3 666 8228 666 8228 0 FrameData[25]
rlabel metal3 712 8500 712 8500 0 FrameData[26]
rlabel metal3 528 8772 528 8772 0 FrameData[27]
rlabel metal3 620 9044 620 9044 0 FrameData[28]
rlabel metal3 390 9316 390 9316 0 FrameData[29]
rlabel metal3 620 1972 620 1972 0 FrameData[2]
rlabel metal3 574 9588 574 9588 0 FrameData[30]
rlabel metal2 2806 8857 2806 8857 0 FrameData[31]
rlabel metal1 33304 7854 33304 7854 0 FrameData[3]
rlabel metal3 252 2516 252 2516 0 FrameData[4]
rlabel metal3 735 2788 735 2788 0 FrameData[5]
rlabel metal3 3404 2992 3404 2992 0 FrameData[6]
rlabel metal3 574 3332 574 3332 0 FrameData[7]
rlabel metal3 298 3604 298 3604 0 FrameData[8]
rlabel metal3 206 3876 206 3876 0 FrameData[9]
rlabel metal3 39798 1428 39798 1428 0 FrameData_O[0]
rlabel metal3 39982 4148 39982 4148 0 FrameData_O[10]
rlabel metal1 39514 3706 39514 3706 0 FrameData_O[11]
rlabel metal2 39422 4335 39422 4335 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal2 39422 5015 39422 5015 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal2 39422 5559 39422 5559 0 FrameData_O[16]
rlabel metal3 39798 6052 39798 6052 0 FrameData_O[17]
rlabel metal3 39798 6324 39798 6324 0 FrameData_O[18]
rlabel metal2 39422 6239 39422 6239 0 FrameData_O[19]
rlabel metal3 39614 1700 39614 1700 0 FrameData_O[1]
rlabel metal3 40120 6868 40120 6868 0 FrameData_O[20]
rlabel metal1 39514 6426 39514 6426 0 FrameData_O[21]
rlabel metal3 40166 7412 40166 7412 0 FrameData_O[22]
rlabel metal1 39468 6630 39468 6630 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal3 39982 8228 39982 8228 0 FrameData_O[25]
rlabel metal1 39008 7514 39008 7514 0 FrameData_O[26]
rlabel metal1 39514 7514 39514 7514 0 FrameData_O[27]
rlabel metal1 39054 6664 39054 6664 0 FrameData_O[28]
rlabel metal2 38686 8415 38686 8415 0 FrameData_O[29]
rlabel metal3 39430 1972 39430 1972 0 FrameData_O[2]
rlabel metal1 39376 6154 39376 6154 0 FrameData_O[30]
rlabel metal1 38364 7514 38364 7514 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 39798 2516 39798 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal3 39798 3604 39798 3604 0 FrameData_O[8]
rlabel metal2 39422 3519 39422 3519 0 FrameData_O[9]
rlabel metal2 11638 1228 11638 1228 0 FrameStrobe[0]
rlabel metal2 26358 55 26358 55 0 FrameStrobe[10]
rlabel metal1 37858 6324 37858 6324 0 FrameStrobe[11]
rlabel metal2 29302 1534 29302 1534 0 FrameStrobe[12]
rlabel metal2 38594 3570 38594 3570 0 FrameStrobe[13]
rlabel metal2 32246 55 32246 55 0 FrameStrobe[14]
rlabel metal2 33718 106 33718 106 0 FrameStrobe[15]
rlabel metal2 35190 1568 35190 1568 0 FrameStrobe[16]
rlabel metal2 36662 55 36662 55 0 FrameStrobe[17]
rlabel metal2 38134 55 38134 55 0 FrameStrobe[18]
rlabel metal2 39606 191 39606 191 0 FrameStrobe[19]
rlabel metal2 13110 1007 13110 1007 0 FrameStrobe[1]
rlabel metal2 14582 55 14582 55 0 FrameStrobe[2]
rlabel metal2 16054 140 16054 140 0 FrameStrobe[3]
rlabel via2 17526 55 17526 55 0 FrameStrobe[4]
rlabel metal2 18998 174 18998 174 0 FrameStrobe[5]
rlabel metal2 20470 208 20470 208 0 FrameStrobe[6]
rlabel metal2 21942 123 21942 123 0 FrameStrobe[7]
rlabel metal2 23414 446 23414 446 0 FrameStrobe[8]
rlabel metal2 24886 55 24886 55 0 FrameStrobe[9]
rlabel metal1 32660 8602 32660 8602 0 FrameStrobe_O[0]
rlabel metal1 36386 8296 36386 8296 0 FrameStrobe_O[10]
rlabel metal1 35650 8058 35650 8058 0 FrameStrobe_O[11]
rlabel metal1 36294 8602 36294 8602 0 FrameStrobe_O[12]
rlabel metal1 36202 8058 36202 8058 0 FrameStrobe_O[13]
rlabel metal1 37306 8262 37306 8262 0 FrameStrobe_O[14]
rlabel metal1 36800 8058 36800 8058 0 FrameStrobe_O[15]
rlabel metal1 37398 8602 37398 8602 0 FrameStrobe_O[16]
rlabel metal1 37720 8330 37720 8330 0 FrameStrobe_O[17]
rlabel metal1 38594 8568 38594 8568 0 FrameStrobe_O[18]
rlabel metal1 38226 8058 38226 8058 0 FrameStrobe_O[19]
rlabel metal1 32982 8330 32982 8330 0 FrameStrobe_O[1]
rlabel metal1 33166 8602 33166 8602 0 FrameStrobe_O[2]
rlabel metal1 33718 8602 33718 8602 0 FrameStrobe_O[3]
rlabel metal1 33902 8330 33902 8330 0 FrameStrobe_O[4]
rlabel metal1 34408 8602 34408 8602 0 FrameStrobe_O[5]
rlabel metal1 35190 8568 35190 8568 0 FrameStrobe_O[6]
rlabel metal1 34638 8058 34638 8058 0 FrameStrobe_O[7]
rlabel metal1 35190 8330 35190 8330 0 FrameStrobe_O[8]
rlabel metal1 36018 8364 36018 8364 0 FrameStrobe_O[9]
rlabel metal2 14490 4250 14490 4250 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q
rlabel metal1 15502 7276 15502 7276 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 16698 5746 16698 5746 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q
rlabel metal1 17664 4658 17664 4658 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q
rlabel metal1 5980 4250 5980 4250 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q
rlabel metal1 6072 4658 6072 4658 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
rlabel metal1 8170 5202 8170 5202 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q
rlabel metal1 19826 3536 19826 3536 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 21896 4590 21896 4590 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 20976 3026 20976 3026 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 26634 5202 26634 5202 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q
rlabel via1 27352 5678 27352 5678 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
rlabel metal1 29578 5644 29578 5644 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q
rlabel viali 22017 7854 22017 7854 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 20470 6358 20470 6358 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
rlabel metal1 18906 7752 18906 7752 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q
rlabel metal1 11362 5712 11362 5712 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q
rlabel via1 10166 5678 10166 5678 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
rlabel via1 10148 6289 10148 6289 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
rlabel metal1 15226 3978 15226 3978 0 Inst_S_WARMBOOT_switch_matrix.N1BEG0
rlabel metal1 15226 7514 15226 7514 0 Inst_S_WARMBOOT_switch_matrix.N1BEG1
rlabel metal2 16974 6086 16974 6086 0 Inst_S_WARMBOOT_switch_matrix.N1BEG2
rlabel metal1 17710 4114 17710 4114 0 Inst_S_WARMBOOT_switch_matrix.N1BEG3
rlabel metal2 3450 8755 3450 8755 0 N1BEG[0]
rlabel metal1 3312 8330 3312 8330 0 N1BEG[1]
rlabel metal1 3634 8602 3634 8602 0 N1BEG[2]
rlabel metal1 4186 8058 4186 8058 0 N1BEG[3]
rlabel metal1 4278 8602 4278 8602 0 N2BEG[0]
rlabel metal1 4738 8058 4738 8058 0 N2BEG[1]
rlabel metal1 4738 8602 4738 8602 0 N2BEG[2]
rlabel metal1 5290 8058 5290 8058 0 N2BEG[3]
rlabel metal1 4922 8364 4922 8364 0 N2BEG[4]
rlabel metal1 5520 8330 5520 8330 0 N2BEG[5]
rlabel metal1 5796 8602 5796 8602 0 N2BEG[6]
rlabel metal1 6164 8602 6164 8602 0 N2BEG[7]
rlabel metal1 6670 8058 6670 8058 0 N2BEGb[0]
rlabel metal1 6808 8602 6808 8602 0 N2BEGb[1]
rlabel metal1 7222 8058 7222 8058 0 N2BEGb[2]
rlabel metal1 7268 8602 7268 8602 0 N2BEGb[3]
rlabel metal1 7774 8058 7774 8058 0 N2BEGb[4]
rlabel metal1 7728 8330 7728 8330 0 N2BEGb[5]
rlabel metal1 8004 8602 8004 8602 0 N2BEGb[6]
rlabel metal1 8372 8602 8372 8602 0 N2BEGb[7]
rlabel metal2 9062 8160 9062 8160 0 N4BEG[0]
rlabel metal1 11362 8602 11362 8602 0 N4BEG[10]
rlabel metal1 11914 8058 11914 8058 0 N4BEG[11]
rlabel metal1 12052 8602 12052 8602 0 N4BEG[12]
rlabel metal1 12328 8602 12328 8602 0 N4BEG[13]
rlabel metal1 12742 8058 12742 8058 0 N4BEG[14]
rlabel metal1 12788 8602 12788 8602 0 N4BEG[15]
rlabel metal1 8740 8602 8740 8602 0 N4BEG[1]
rlabel metal1 9476 8058 9476 8058 0 N4BEG[2]
rlabel metal1 9476 8602 9476 8602 0 N4BEG[3]
rlabel metal1 9982 8058 9982 8058 0 N4BEG[4]
rlabel metal1 9936 8330 9936 8330 0 N4BEG[5]
rlabel metal1 10258 8602 10258 8602 0 N4BEG[6]
rlabel metal1 10626 8602 10626 8602 0 N4BEG[7]
rlabel metal1 10948 8602 10948 8602 0 N4BEG[8]
rlabel metal1 11362 8058 11362 8058 0 N4BEG[9]
rlabel metal1 13110 8602 13110 8602 0 NN4BEG[0]
rlabel metal1 16054 8058 16054 8058 0 NN4BEG[10]
rlabel metal1 16100 8602 16100 8602 0 NN4BEG[11]
rlabel metal1 16468 8602 16468 8602 0 NN4BEG[12]
rlabel metal1 16882 8602 16882 8602 0 NN4BEG[13]
rlabel metal1 17802 8330 17802 8330 0 NN4BEG[14]
rlabel metal1 17526 8398 17526 8398 0 NN4BEG[15]
rlabel metal1 13662 7752 13662 7752 0 NN4BEG[1]
rlabel metal1 13524 8602 13524 8602 0 NN4BEG[2]
rlabel metal1 13892 8602 13892 8602 0 NN4BEG[3]
rlabel metal1 14398 8058 14398 8058 0 NN4BEG[4]
rlabel metal1 14536 8602 14536 8602 0 NN4BEG[5]
rlabel metal1 14950 8058 14950 8058 0 NN4BEG[6]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[7]
rlabel metal1 15364 8602 15364 8602 0 NN4BEG[8]
rlabel metal1 15640 8602 15640 8602 0 NN4BEG[9]
rlabel metal2 1334 1228 1334 1228 0 RESET_top
rlabel metal2 17894 9292 17894 9292 0 S1END[0]
rlabel metal2 18170 9292 18170 9292 0 S1END[1]
rlabel metal2 18446 9836 18446 9836 0 S1END[2]
rlabel metal2 18722 9836 18722 9836 0 S1END[3]
rlabel metal2 21206 10533 21206 10533 0 S2END[0]
rlabel metal2 21482 9836 21482 9836 0 S2END[1]
rlabel metal2 21758 9870 21758 9870 0 S2END[2]
rlabel metal2 22034 9802 22034 9802 0 S2END[3]
rlabel metal2 22310 9870 22310 9870 0 S2END[4]
rlabel metal2 22586 9904 22586 9904 0 S2END[5]
rlabel metal2 22862 9870 22862 9870 0 S2END[6]
rlabel metal2 23138 10414 23138 10414 0 S2END[7]
rlabel metal2 18998 9836 18998 9836 0 S2MID[0]
rlabel metal2 19274 9836 19274 9836 0 S2MID[1]
rlabel metal2 19550 9836 19550 9836 0 S2MID[2]
rlabel metal2 19826 9836 19826 9836 0 S2MID[3]
rlabel metal2 20102 10193 20102 10193 0 S2MID[4]
rlabel metal2 20378 11145 20378 11145 0 S2MID[5]
rlabel metal2 20654 10550 20654 10550 0 S2MID[6]
rlabel metal2 20930 9734 20930 9734 0 S2MID[7]
rlabel metal2 23414 9870 23414 9870 0 S4END[0]
rlabel metal2 26174 9734 26174 9734 0 S4END[10]
rlabel metal2 32614 9044 32614 9044 0 S4END[11]
rlabel metal1 37490 6256 37490 6256 0 S4END[12]
rlabel metal1 32118 4114 32118 4114 0 S4END[13]
rlabel metal2 38962 4896 38962 4896 0 S4END[14]
rlabel metal2 27554 8748 27554 8748 0 S4END[15]
rlabel metal2 23690 9904 23690 9904 0 S4END[1]
rlabel metal2 23966 10533 23966 10533 0 S4END[2]
rlabel metal2 24242 9870 24242 9870 0 S4END[3]
rlabel metal2 24518 10618 24518 10618 0 S4END[4]
rlabel metal2 24794 10533 24794 10533 0 S4END[5]
rlabel metal2 25070 9802 25070 9802 0 S4END[6]
rlabel metal2 25346 9870 25346 9870 0 S4END[7]
rlabel metal2 1886 9520 1886 9520 0 S4END[8]
rlabel metal1 31947 7854 31947 7854 0 S4END[9]
rlabel metal2 4278 1160 4278 1160 0 SLOT_top0
rlabel metal2 5750 1160 5750 1160 0 SLOT_top1
rlabel metal2 7222 1160 7222 1160 0 SLOT_top2
rlabel metal2 8694 1160 8694 1160 0 SLOT_top3
rlabel metal2 27830 9836 27830 9836 0 SS4END[0]
rlabel metal2 30590 7116 30590 7116 0 SS4END[10]
rlabel metal2 30866 8986 30866 8986 0 SS4END[11]
rlabel metal1 38778 5712 38778 5712 0 SS4END[12]
rlabel metal1 38318 4658 38318 4658 0 SS4END[13]
rlabel metal2 31878 6001 31878 6001 0 SS4END[14]
rlabel metal2 31970 9734 31970 9734 0 SS4END[15]
rlabel metal2 28106 10533 28106 10533 0 SS4END[1]
rlabel metal2 28382 9836 28382 9836 0 SS4END[2]
rlabel metal2 28658 9802 28658 9802 0 SS4END[3]
rlabel metal2 28934 9904 28934 9904 0 SS4END[4]
rlabel metal2 29210 10533 29210 10533 0 SS4END[5]
rlabel metal2 29486 9530 29486 9530 0 SS4END[6]
rlabel metal2 29762 9870 29762 9870 0 SS4END[7]
rlabel metal2 34178 4284 34178 4284 0 SS4END[8]
rlabel metal2 30314 7660 30314 7660 0 SS4END[9]
rlabel metal1 32016 3026 32016 3026 0 UserCLK
rlabel metal1 32292 8602 32292 8602 0 UserCLKo
rlabel metal1 9913 6222 9913 6222 0 _000_
rlabel metal1 21298 7514 21298 7514 0 _001_
rlabel metal1 29440 5746 29440 5746 0 _002_
rlabel metal1 22816 2958 22816 2958 0 _003_
rlabel metal2 7498 4828 7498 4828 0 _004_
rlabel metal2 9706 5882 9706 5882 0 _005_
rlabel metal1 10580 4998 10580 4998 0 _006_
rlabel metal1 10741 5678 10741 5678 0 _007_
rlabel metal1 10258 4794 10258 4794 0 _008_
rlabel metal2 10718 6086 10718 6086 0 _009_
rlabel metal2 19826 7174 19826 7174 0 _010_
rlabel metal1 21298 7786 21298 7786 0 _011_
rlabel metal1 20840 7854 20840 7854 0 _012_
rlabel metal2 20746 7922 20746 7922 0 _013_
rlabel metal1 21252 7854 21252 7854 0 _014_
rlabel metal2 29394 5236 29394 5236 0 _015_
rlabel metal1 27186 5610 27186 5610 0 _016_
rlabel metal1 27602 5678 27602 5678 0 _017_
rlabel metal2 27462 6154 27462 6154 0 _018_
rlabel metal1 28382 5678 28382 5678 0 _019_
rlabel metal2 21574 4216 21574 4216 0 _020_
rlabel metal1 22688 3094 22688 3094 0 _021_
rlabel metal1 22315 2992 22315 2992 0 _022_
rlabel metal1 22126 3128 22126 3128 0 _023_
rlabel metal1 22632 3026 22632 3026 0 _024_
rlabel metal1 7176 4658 7176 4658 0 _025_
rlabel metal1 8188 4250 8188 4250 0 _026_
rlabel metal1 8231 4590 8231 4590 0 _027_
rlabel metal1 8326 4488 8326 4488 0 _028_
rlabel metal1 7222 4522 7222 4522 0 _029_
rlabel metal2 7222 4896 7222 4896 0 net1
rlabel metal1 2070 6698 2070 6698 0 net10
rlabel metal2 32706 8670 32706 8670 0 net100
rlabel metal1 38088 5882 38088 5882 0 net101
rlabel metal1 33580 5338 33580 5338 0 net102
rlabel metal1 36156 3162 36156 3162 0 net103
rlabel metal2 35006 6630 35006 6630 0 net104
rlabel metal1 38226 3128 38226 3128 0 net105
rlabel metal1 35466 4794 35466 4794 0 net106
rlabel metal2 35466 8772 35466 8772 0 net107
rlabel metal1 33258 5066 33258 5066 0 net108
rlabel metal1 13570 4488 13570 4488 0 net109
rlabel metal1 19550 4556 19550 4556 0 net11
rlabel metal1 15410 8058 15410 8058 0 net110
rlabel metal2 3634 8772 3634 8772 0 net111
rlabel metal2 17710 3774 17710 3774 0 net112
rlabel metal2 14398 7888 14398 7888 0 net113
rlabel metal2 12926 7854 12926 7854 0 net114
rlabel metal2 8602 8194 8602 8194 0 net115
rlabel metal1 5566 7888 5566 7888 0 net116
rlabel metal1 12052 4454 12052 4454 0 net117
rlabel metal2 16422 9061 16422 9061 0 net118
rlabel metal2 5842 8415 5842 8415 0 net119
rlabel metal1 1886 7752 1886 7752 0 net12
rlabel metal1 7590 8874 7590 8874 0 net120
rlabel metal1 10120 3910 10120 3910 0 net121
rlabel metal3 20516 8024 20516 8024 0 net122
rlabel metal2 7498 7361 7498 7361 0 net123
rlabel metal1 15548 2550 15548 2550 0 net124
rlabel metal1 10304 3978 10304 3978 0 net125
rlabel metal2 11178 8109 11178 8109 0 net126
rlabel metal2 8050 9095 8050 9095 0 net127
rlabel metal1 8418 8500 8418 8500 0 net128
rlabel metal2 27830 5151 27830 5151 0 net129
rlabel metal1 23805 7378 23805 7378 0 net13
rlabel metal2 20654 8313 20654 8313 0 net130
rlabel metal1 14674 7310 14674 7310 0 net131
rlabel metal1 7544 6086 7544 6086 0 net132
rlabel metal2 13846 7123 13846 7123 0 net133
rlabel metal2 20378 7276 20378 7276 0 net134
rlabel via2 21574 4981 21574 4981 0 net135
rlabel via2 38502 4539 38502 4539 0 net136
rlabel metal2 32338 2992 32338 2992 0 net137
rlabel metal1 37582 6086 37582 6086 0 net138
rlabel metal2 35098 7310 35098 7310 0 net139
rlabel metal2 1702 6834 1702 6834 0 net14
rlabel metal2 37306 4777 37306 4777 0 net140
rlabel metal2 14674 8568 14674 8568 0 net141
rlabel metal2 10350 8126 10350 8126 0 net142
rlabel metal2 6210 7684 6210 7684 0 net143
rlabel metal2 21850 6596 21850 6596 0 net144
rlabel metal2 13386 8806 13386 8806 0 net145
rlabel metal2 16422 7157 16422 7157 0 net146
rlabel metal2 20930 4896 20930 4896 0 net147
rlabel metal2 14950 6528 14950 6528 0 net148
rlabel metal1 19872 5542 19872 5542 0 net149
rlabel metal2 2530 9214 2530 9214 0 net15
rlabel metal2 18078 9010 18078 9010 0 net150
rlabel metal1 20010 4794 20010 4794 0 net151
rlabel metal2 14306 5610 14306 5610 0 net152
rlabel metal2 21574 5185 21574 5185 0 net153
rlabel metal2 13938 8704 13938 8704 0 net154
rlabel metal3 20700 7888 20700 7888 0 net155
rlabel metal1 16882 4012 16882 4012 0 net156
rlabel metal1 18814 3536 18814 3536 0 net157
rlabel metal1 26726 3672 26726 3672 0 net158
rlabel metal2 13846 8908 13846 8908 0 net159
rlabel metal2 16330 7684 16330 7684 0 net16
rlabel metal1 19504 6154 19504 6154 0 net160
rlabel metal1 4646 2516 4646 2516 0 net161
rlabel metal1 6210 1972 6210 1972 0 net162
rlabel metal1 21344 7718 21344 7718 0 net163
rlabel metal1 9338 2414 9338 2414 0 net164
rlabel metal1 32476 3162 32476 3162 0 net165
rlabel metal1 17572 8058 17572 8058 0 net166
rlabel metal1 18262 6324 18262 6324 0 net17
rlabel metal1 17618 7888 17618 7888 0 net18
rlabel metal1 13340 5610 13340 5610 0 net19
rlabel metal2 5658 6120 5658 6120 0 net2
rlabel metal2 2714 7344 2714 7344 0 net20
rlabel metal1 9568 7378 9568 7378 0 net21
rlabel metal1 17894 2278 17894 2278 0 net22
rlabel metal2 1702 2142 1702 2142 0 net23
rlabel metal1 18032 4590 18032 4590 0 net24
rlabel metal1 18308 5542 18308 5542 0 net25
rlabel metal2 18538 8313 18538 8313 0 net26
rlabel metal2 14674 4624 14674 4624 0 net27
rlabel metal1 24288 3026 24288 3026 0 net28
rlabel metal1 27876 6630 27876 6630 0 net29
rlabel metal2 1610 5984 1610 5984 0 net3
rlabel metal1 22862 7718 22862 7718 0 net30
rlabel metal1 10718 4148 10718 4148 0 net31
rlabel metal1 24104 2958 24104 2958 0 net32
rlabel metal1 27692 6834 27692 6834 0 net33
rlabel metal1 23460 7854 23460 7854 0 net34
rlabel metal2 23782 6732 23782 6732 0 net35
rlabel metal2 19182 6086 19182 6086 0 net36
rlabel metal1 25392 5678 25392 5678 0 net37
rlabel metal2 21022 8126 21022 8126 0 net38
rlabel metal2 20562 6698 20562 6698 0 net39
rlabel metal2 2714 6103 2714 6103 0 net4
rlabel metal2 23598 6460 23598 6460 0 net40
rlabel metal1 27738 4556 27738 4556 0 net41
rlabel metal1 21482 6324 21482 6324 0 net42
rlabel metal2 24702 7514 24702 7514 0 net43
rlabel metal1 23322 4556 23322 4556 0 net44
rlabel metal1 26956 4590 26956 4590 0 net45
rlabel metal1 22034 6256 22034 6256 0 net46
rlabel metal2 23414 6120 23414 6120 0 net47
rlabel metal1 21643 4658 21643 4658 0 net48
rlabel metal1 27508 4114 27508 4114 0 net49
rlabel metal2 5474 5270 5474 5270 0 net5
rlabel via1 20641 6290 20641 6290 0 net50
rlabel metal2 21942 5916 21942 5916 0 net51
rlabel metal1 21114 4692 21114 4692 0 net52
rlabel metal2 28520 4590 28520 4590 0 net53
rlabel metal1 20930 6222 20930 6222 0 net54
rlabel metal1 17066 9044 17066 9044 0 net55
rlabel metal1 3864 2414 3864 2414 0 net56
rlabel metal2 3818 2890 3818 2890 0 net57
rlabel metal2 38870 4063 38870 4063 0 net58
rlabel metal1 39514 3502 39514 3502 0 net59
rlabel metal2 2622 6494 2622 6494 0 net6
rlabel metal1 39376 4114 39376 4114 0 net60
rlabel via2 13662 4709 13662 4709 0 net61
rlabel metal2 13662 6137 13662 6137 0 net62
rlabel metal2 15180 6324 15180 6324 0 net63
rlabel metal1 17066 4794 17066 4794 0 net64
rlabel metal3 35052 3400 35052 3400 0 net65
rlabel metal2 38502 6477 38502 6477 0 net66
rlabel metal2 39238 5729 39238 5729 0 net67
rlabel metal1 37582 2482 37582 2482 0 net68
rlabel metal1 19550 2856 19550 2856 0 net69
rlabel metal1 17848 6290 17848 6290 0 net7
rlabel metal2 19090 4930 19090 4930 0 net70
rlabel metal2 19366 3298 19366 3298 0 net71
rlabel metal1 39238 6800 39238 6800 0 net72
rlabel metal2 38778 8840 38778 8840 0 net73
rlabel metal2 38870 8908 38870 8908 0 net74
rlabel metal2 16514 7072 16514 7072 0 net75
rlabel metal2 19274 5950 19274 5950 0 net76
rlabel metal2 22034 5967 22034 5967 0 net77
rlabel via2 13754 5627 13754 5627 0 net78
rlabel metal1 14237 2482 14237 2482 0 net79
rlabel metal2 2530 6052 2530 6052 0 net8
rlabel metal2 12742 6681 12742 6681 0 net80
rlabel metal2 38134 7327 38134 7327 0 net81
rlabel metal1 39284 2482 39284 2482 0 net82
rlabel via2 38502 3043 38502 3043 0 net83
rlabel metal3 35236 3536 35236 3536 0 net84
rlabel metal3 35420 2448 35420 2448 0 net85
rlabel metal2 38686 4930 38686 4930 0 net86
rlabel metal1 31878 3944 31878 3944 0 net87
rlabel metal2 38962 3332 38962 3332 0 net88
rlabel metal1 16928 3162 16928 3162 0 net89
rlabel metal1 1886 6868 1886 6868 0 net9
rlabel metal2 34086 7480 34086 7480 0 net90
rlabel metal2 37674 7106 37674 7106 0 net91
rlabel metal2 33902 3468 33902 3468 0 net92
rlabel metal1 37444 4454 37444 4454 0 net93
rlabel metal2 37122 6630 37122 6630 0 net94
rlabel metal2 36754 5389 36754 5389 0 net95
rlabel metal2 36846 6018 36846 6018 0 net96
rlabel metal1 33902 4794 33902 4794 0 net97
rlabel metal1 33810 4998 33810 4998 0 net98
rlabel metal2 38318 7582 38318 7582 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
