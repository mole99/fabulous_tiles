module S_term_IHP_SRAM (UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    S1END,
    S2END,
    S2MID,
    S4END);
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;

 sg13g2_buf_1 _00_ (.A(FrameData[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _01_ (.A(FrameData[1]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _02_ (.A(FrameData[2]),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _03_ (.A(FrameData[3]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _04_ (.A(FrameData[4]),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _05_ (.A(FrameData[5]),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _06_ (.A(FrameData[6]),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _07_ (.A(FrameData[7]),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _08_ (.A(FrameData[8]),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _09_ (.A(FrameData[9]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10_ (.A(FrameData[10]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _11_ (.A(FrameData[11]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _12_ (.A(FrameData[12]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _13_ (.A(FrameData[13]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _14_ (.A(FrameData[14]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _15_ (.A(FrameData[15]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _16_ (.A(FrameData[16]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _17_ (.A(FrameData[17]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _18_ (.A(FrameData[18]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _19_ (.A(FrameData[19]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _20_ (.A(FrameData[20]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _21_ (.A(FrameData[21]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _22_ (.A(FrameData[22]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _23_ (.A(FrameData[23]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _24_ (.A(FrameData[24]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _25_ (.A(FrameData[25]),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _26_ (.A(FrameData[26]),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _27_ (.A(FrameData[27]),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _28_ (.A(FrameData[28]),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _29_ (.A(FrameData[29]),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _30_ (.A(FrameData[30]),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _31_ (.A(FrameData[31]),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _32_ (.A(FrameStrobe[0]),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _33_ (.A(FrameStrobe[1]),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _34_ (.A(FrameStrobe[2]),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _35_ (.A(FrameStrobe[3]),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _36_ (.A(FrameStrobe[4]),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _37_ (.A(FrameStrobe[5]),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _38_ (.A(FrameStrobe[6]),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _39_ (.A(FrameStrobe[7]),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _40_ (.A(FrameStrobe[8]),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _41_ (.A(FrameStrobe[9]),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _42_ (.A(FrameStrobe[10]),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _43_ (.A(FrameStrobe[11]),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _44_ (.A(FrameStrobe[12]),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _45_ (.A(FrameStrobe[13]),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _46_ (.A(FrameStrobe[14]),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _47_ (.A(FrameStrobe[15]),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _48_ (.A(FrameStrobe[16]),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _49_ (.A(FrameStrobe[17]),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _50_ (.A(FrameStrobe[18]),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _51_ (.A(FrameStrobe[19]),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _52_ (.A(S1END[3]),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _53_ (.A(S1END[2]),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _54_ (.A(S1END[1]),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _55_ (.A(S1END[0]),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _56_ (.A(S2MID[7]),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _57_ (.A(S2MID[6]),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _58_ (.A(S2MID[5]),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _59_ (.A(S2MID[4]),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _60_ (.A(S2MID[3]),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _61_ (.A(S2MID[2]),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _62_ (.A(S2MID[1]),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _63_ (.A(S2MID[0]),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _64_ (.A(S2END[7]),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _65_ (.A(S2END[6]),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _66_ (.A(S2END[5]),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _67_ (.A(S2END[4]),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _68_ (.A(S2END[3]),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _69_ (.A(S2END[2]),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _70_ (.A(S2END[1]),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _71_ (.A(S2END[0]),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _72_ (.A(S4END[15]),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _73_ (.A(S4END[14]),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _74_ (.A(S4END[13]),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _75_ (.A(S4END[12]),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _76_ (.A(S4END[11]),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _77_ (.A(S4END[10]),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _78_ (.A(S4END[9]),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _79_ (.A(S4END[8]),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _80_ (.A(S4END[7]),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _81_ (.A(S4END[6]),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _82_ (.A(S4END[5]),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _83_ (.A(S4END[4]),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _84_ (.A(S4END[3]),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _85_ (.A(S4END[2]),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _86_ (.A(S4END[1]),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _87_ (.A(S4END[0]),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _88_ (.A(UserCLK),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output53 (.A(net53),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output54 (.A(net54),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output55 (.A(net55),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output56 (.A(net56),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output57 (.A(net57),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output58 (.A(net58),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output59 (.A(net59),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output60 (.A(net60),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output61 (.A(net61),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output62 (.A(net62),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output63 (.A(net63),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output64 (.A(net64),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output65 (.A(net65),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output66 (.A(net66),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output67 (.A(net67),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output68 (.A(net68),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output69 (.A(net69),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output70 (.A(net70),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output71 (.A(net71),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output72 (.A(net72),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output73 (.A(net73),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output74 (.A(net74),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output75 (.A(net75),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output76 (.A(net76),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output77 (.A(net77),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output78 (.A(net78),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output79 (.A(net79),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output80 (.A(net80),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output81 (.A(net81),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output82 (.A(net82),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output83 (.A(net83),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output84 (.A(net84),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output85 (.A(net85),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output86 (.A(net86),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output87 (.A(net87),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output88 (.A(net88),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output89 (.A(net89),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_200 (.VDD(VPWR),
    .VSS(VGND));
endmodule
