VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_term_single2
  CLASS BLOCK ;
  FOREIGN S_term_single2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 266.400 BY 59.220 ;
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2.740 0.450 3.140 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 19.540 0.450 19.940 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 21.220 0.450 21.620 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.900 0.450 23.300 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 24.580 0.450 24.980 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 26.260 0.450 26.660 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.940 0.450 28.340 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 29.620 0.450 30.020 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 31.300 0.450 31.700 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.980 0.450 33.380 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 34.660 0.450 35.060 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 4.420 0.450 4.820 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 36.340 0.450 36.740 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.020 0.450 38.420 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 39.700 0.450 40.100 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 41.380 0.450 41.780 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 43.060 0.450 43.460 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 44.740 0.450 45.140 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 46.420 0.450 46.820 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.100 0.450 48.500 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 49.780 0.450 50.180 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 51.460 0.450 51.860 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 6.100 0.450 6.500 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 53.140 0.450 53.540 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 54.820 0.450 55.220 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 7.780 0.450 8.180 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 9.460 0.450 9.860 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 11.140 0.450 11.540 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 12.820 0.450 13.220 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 14.500 0.450 14.900 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 16.180 0.450 16.580 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 17.860 0.450 18.260 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 2.740 266.400 3.140 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 19.540 266.400 19.940 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 21.220 266.400 21.620 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 22.900 266.400 23.300 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 24.580 266.400 24.980 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 26.260 266.400 26.660 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 27.940 266.400 28.340 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 29.620 266.400 30.020 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 31.300 266.400 31.700 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 32.980 266.400 33.380 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 34.660 266.400 35.060 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 4.420 266.400 4.820 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 36.340 266.400 36.740 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 38.020 266.400 38.420 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 39.700 266.400 40.100 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 41.380 266.400 41.780 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 43.060 266.400 43.460 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 44.740 266.400 45.140 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 46.420 266.400 46.820 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 48.100 266.400 48.500 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 49.780 266.400 50.180 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 51.460 266.400 51.860 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 6.100 266.400 6.500 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 53.140 266.400 53.540 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 54.820 266.400 55.220 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 7.780 266.400 8.180 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 9.460 266.400 9.860 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 11.140 266.400 11.540 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 12.820 266.400 13.220 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 14.500 266.400 14.900 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 16.180 266.400 16.580 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.950 17.860 266.400 18.260 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 20.440 0.000 20.840 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 145.240 0.000 145.640 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 157.720 0.000 158.120 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 170.200 0.000 170.600 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 182.680 0.000 183.080 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 195.160 0.000 195.560 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 207.640 0.000 208.040 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 220.120 0.000 220.520 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 232.600 0.000 233.000 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 245.080 0.000 245.480 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 257.560 0.000 257.960 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 0.000 108.200 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 120.280 0.000 120.680 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 0.000 133.160 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 215.320 58.820 215.720 59.220 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 234.520 58.820 234.920 59.220 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 236.440 58.820 236.840 59.220 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 238.360 58.820 238.760 59.220 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 240.280 58.820 240.680 59.220 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 242.200 58.820 242.600 59.220 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 244.120 58.820 244.520 59.220 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.040 58.820 246.440 59.220 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 247.960 58.820 248.360 59.220 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 249.880 58.820 250.280 59.220 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 251.800 58.820 252.200 59.220 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 217.240 58.820 217.640 59.220 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 219.160 58.820 219.560 59.220 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 221.080 58.820 221.480 59.220 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 223.000 58.820 223.400 59.220 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 224.920 58.820 225.320 59.220 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 226.840 58.820 227.240 59.220 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 228.760 58.820 229.160 59.220 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 230.680 58.820 231.080 59.220 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 232.600 58.820 233.000 59.220 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 13.720 58.820 14.120 59.220 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 15.640 58.820 16.040 59.220 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 17.560 58.820 17.960 59.220 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 19.480 58.820 19.880 59.220 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 21.400 58.820 21.800 59.220 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 23.320 58.820 23.720 59.220 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 25.240 58.820 25.640 59.220 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 27.160 58.820 27.560 59.220 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 29.080 58.820 29.480 59.220 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 31.000 58.820 31.400 59.220 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 32.920 58.820 33.320 59.220 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 34.840 58.820 35.240 59.220 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 36.760 58.820 37.160 59.220 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 38.680 58.820 39.080 59.220 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 40.600 58.820 41.000 59.220 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 42.520 58.820 42.920 59.220 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 44.440 58.820 44.840 59.220 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 46.360 58.820 46.760 59.220 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 48.280 58.820 48.680 59.220 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 50.200 58.820 50.600 59.220 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 52.120 58.820 52.520 59.220 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 71.320 58.820 71.720 59.220 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 73.240 58.820 73.640 59.220 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 75.160 58.820 75.560 59.220 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 77.080 58.820 77.480 59.220 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 79.000 58.820 79.400 59.220 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 80.920 58.820 81.320 59.220 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 54.040 58.820 54.440 59.220 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 55.960 58.820 56.360 59.220 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 57.880 58.820 58.280 59.220 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 59.800 58.820 60.200 59.220 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 61.720 58.820 62.120 59.220 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 63.640 58.820 64.040 59.220 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 65.560 58.820 65.960 59.220 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 67.480 58.820 67.880 59.220 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 69.400 58.820 69.800 59.220 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 82.840 58.820 83.240 59.220 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 102.040 58.820 102.440 59.220 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 103.960 58.820 104.360 59.220 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 105.880 58.820 106.280 59.220 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.800 58.820 108.200 59.220 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 109.720 58.820 110.120 59.220 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 111.640 58.820 112.040 59.220 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 84.760 58.820 85.160 59.220 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 86.680 58.820 87.080 59.220 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 88.600 58.820 89.000 59.220 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 90.520 58.820 90.920 59.220 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 92.440 58.820 92.840 59.220 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 94.360 58.820 94.760 59.220 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 96.280 58.820 96.680 59.220 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 98.200 58.820 98.600 59.220 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 100.120 58.820 100.520 59.220 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 113.560 58.820 113.960 59.220 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 115.480 58.820 115.880 59.220 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 117.400 58.820 117.800 59.220 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 119.320 58.820 119.720 59.220 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 136.600 58.820 137.000 59.220 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 138.520 58.820 138.920 59.220 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 140.440 58.820 140.840 59.220 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 142.360 58.820 142.760 59.220 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 144.280 58.820 144.680 59.220 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 146.200 58.820 146.600 59.220 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 148.120 58.820 148.520 59.220 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 150.040 58.820 150.440 59.220 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 121.240 58.820 121.640 59.220 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 123.160 58.820 123.560 59.220 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 125.080 58.820 125.480 59.220 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 127.000 58.820 127.400 59.220 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 128.920 58.820 129.320 59.220 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 130.840 58.820 131.240 59.220 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 132.760 58.820 133.160 59.220 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 134.680 58.820 135.080 59.220 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 151.960 58.820 152.360 59.220 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 171.160 58.820 171.560 59.220 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 173.080 58.820 173.480 59.220 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 175.000 58.820 175.400 59.220 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 176.920 58.820 177.320 59.220 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 178.840 58.820 179.240 59.220 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 180.760 58.820 181.160 59.220 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 153.880 58.820 154.280 59.220 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 155.800 58.820 156.200 59.220 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 157.720 58.820 158.120 59.220 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 159.640 58.820 160.040 59.220 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 161.560 58.820 161.960 59.220 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 163.480 58.820 163.880 59.220 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 165.400 58.820 165.800 59.220 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 167.320 58.820 167.720 59.220 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 169.240 58.820 169.640 59.220 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 182.680 58.820 183.080 59.220 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 201.880 58.820 202.280 59.220 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 203.800 58.820 204.200 59.220 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 205.720 58.820 206.120 59.220 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 207.640 58.820 208.040 59.220 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 209.560 58.820 209.960 59.220 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 211.480 58.820 211.880 59.220 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 184.600 58.820 185.000 59.220 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 186.520 58.820 186.920 59.220 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 188.440 58.820 188.840 59.220 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 190.360 58.820 190.760 59.220 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 192.280 58.820 192.680 59.220 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 194.200 58.820 194.600 59.220 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 196.120 58.820 196.520 59.220 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 198.040 58.820 198.440 59.220 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 199.960 58.820 200.360 59.220 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 7.960 0.000 8.360 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.654800 ;
    PORT
      LAYER Metal3 ;
        RECT 213.400 58.820 213.800 59.220 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 24.460 0.000 26.660 59.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 100.060 0.000 102.260 59.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 175.660 0.000 177.860 59.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 251.260 0.000 253.460 59.220 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 18.260 0.000 20.460 59.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 93.860 0.000 96.060 59.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 169.460 0.000 171.660 59.220 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 245.060 0.000 247.260 59.220 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 5.760 7.410 260.640 49.290 ;
      LAYER Metal1 ;
        RECT 5.760 7.340 260.640 49.360 ;
      LAYER Metal2 ;
        RECT 0.380 55.430 266.065 58.900 ;
        RECT 0.660 54.610 265.740 55.430 ;
        RECT 0.380 53.750 266.065 54.610 ;
        RECT 0.660 52.930 265.740 53.750 ;
        RECT 0.380 52.070 266.065 52.930 ;
        RECT 0.660 51.250 265.740 52.070 ;
        RECT 0.380 50.390 266.065 51.250 ;
        RECT 0.660 49.570 265.740 50.390 ;
        RECT 0.380 48.710 266.065 49.570 ;
        RECT 0.660 47.890 265.740 48.710 ;
        RECT 0.380 47.030 266.065 47.890 ;
        RECT 0.660 46.210 265.740 47.030 ;
        RECT 0.380 45.350 266.065 46.210 ;
        RECT 0.660 44.530 265.740 45.350 ;
        RECT 0.380 43.670 266.065 44.530 ;
        RECT 0.660 42.850 265.740 43.670 ;
        RECT 0.380 41.990 266.065 42.850 ;
        RECT 0.660 41.170 265.740 41.990 ;
        RECT 0.380 40.310 266.065 41.170 ;
        RECT 0.660 39.490 265.740 40.310 ;
        RECT 0.380 38.630 266.065 39.490 ;
        RECT 0.660 37.810 265.740 38.630 ;
        RECT 0.380 36.950 266.065 37.810 ;
        RECT 0.660 36.130 265.740 36.950 ;
        RECT 0.380 35.270 266.065 36.130 ;
        RECT 0.660 34.450 265.740 35.270 ;
        RECT 0.380 33.590 266.065 34.450 ;
        RECT 0.660 32.770 265.740 33.590 ;
        RECT 0.380 31.910 266.065 32.770 ;
        RECT 0.660 31.090 265.740 31.910 ;
        RECT 0.380 30.230 266.065 31.090 ;
        RECT 0.660 29.410 265.740 30.230 ;
        RECT 0.380 28.550 266.065 29.410 ;
        RECT 0.660 27.730 265.740 28.550 ;
        RECT 0.380 26.870 266.065 27.730 ;
        RECT 0.660 26.050 265.740 26.870 ;
        RECT 0.380 25.190 266.065 26.050 ;
        RECT 0.660 24.370 265.740 25.190 ;
        RECT 0.380 23.510 266.065 24.370 ;
        RECT 0.660 22.690 265.740 23.510 ;
        RECT 0.380 21.830 266.065 22.690 ;
        RECT 0.660 21.010 265.740 21.830 ;
        RECT 0.380 20.150 266.065 21.010 ;
        RECT 0.660 19.330 265.740 20.150 ;
        RECT 0.380 18.470 266.065 19.330 ;
        RECT 0.660 17.650 265.740 18.470 ;
        RECT 0.380 16.790 266.065 17.650 ;
        RECT 0.660 15.970 265.740 16.790 ;
        RECT 0.380 15.110 266.065 15.970 ;
        RECT 0.660 14.290 265.740 15.110 ;
        RECT 0.380 13.430 266.065 14.290 ;
        RECT 0.660 12.610 265.740 13.430 ;
        RECT 0.380 11.750 266.065 12.610 ;
        RECT 0.660 10.930 265.740 11.750 ;
        RECT 0.380 10.070 266.065 10.930 ;
        RECT 0.660 9.250 265.740 10.070 ;
        RECT 0.380 8.390 266.065 9.250 ;
        RECT 0.660 7.570 265.740 8.390 ;
        RECT 0.380 6.710 266.065 7.570 ;
        RECT 0.660 5.890 265.740 6.710 ;
        RECT 0.380 5.030 266.065 5.890 ;
        RECT 0.660 4.210 265.740 5.030 ;
        RECT 0.380 3.350 266.065 4.210 ;
        RECT 0.660 2.840 265.740 3.350 ;
      LAYER Metal3 ;
        RECT 1.340 58.610 13.510 58.945 ;
        RECT 14.330 58.610 15.430 58.945 ;
        RECT 16.250 58.610 17.350 58.945 ;
        RECT 18.170 58.610 19.270 58.945 ;
        RECT 20.090 58.610 21.190 58.945 ;
        RECT 22.010 58.610 23.110 58.945 ;
        RECT 23.930 58.610 25.030 58.945 ;
        RECT 25.850 58.610 26.950 58.945 ;
        RECT 27.770 58.610 28.870 58.945 ;
        RECT 29.690 58.610 30.790 58.945 ;
        RECT 31.610 58.610 32.710 58.945 ;
        RECT 33.530 58.610 34.630 58.945 ;
        RECT 35.450 58.610 36.550 58.945 ;
        RECT 37.370 58.610 38.470 58.945 ;
        RECT 39.290 58.610 40.390 58.945 ;
        RECT 41.210 58.610 42.310 58.945 ;
        RECT 43.130 58.610 44.230 58.945 ;
        RECT 45.050 58.610 46.150 58.945 ;
        RECT 46.970 58.610 48.070 58.945 ;
        RECT 48.890 58.610 49.990 58.945 ;
        RECT 50.810 58.610 51.910 58.945 ;
        RECT 52.730 58.610 53.830 58.945 ;
        RECT 54.650 58.610 55.750 58.945 ;
        RECT 56.570 58.610 57.670 58.945 ;
        RECT 58.490 58.610 59.590 58.945 ;
        RECT 60.410 58.610 61.510 58.945 ;
        RECT 62.330 58.610 63.430 58.945 ;
        RECT 64.250 58.610 65.350 58.945 ;
        RECT 66.170 58.610 67.270 58.945 ;
        RECT 68.090 58.610 69.190 58.945 ;
        RECT 70.010 58.610 71.110 58.945 ;
        RECT 71.930 58.610 73.030 58.945 ;
        RECT 73.850 58.610 74.950 58.945 ;
        RECT 75.770 58.610 76.870 58.945 ;
        RECT 77.690 58.610 78.790 58.945 ;
        RECT 79.610 58.610 80.710 58.945 ;
        RECT 81.530 58.610 82.630 58.945 ;
        RECT 83.450 58.610 84.550 58.945 ;
        RECT 85.370 58.610 86.470 58.945 ;
        RECT 87.290 58.610 88.390 58.945 ;
        RECT 89.210 58.610 90.310 58.945 ;
        RECT 91.130 58.610 92.230 58.945 ;
        RECT 93.050 58.610 94.150 58.945 ;
        RECT 94.970 58.610 96.070 58.945 ;
        RECT 96.890 58.610 97.990 58.945 ;
        RECT 98.810 58.610 99.910 58.945 ;
        RECT 100.730 58.610 101.830 58.945 ;
        RECT 102.650 58.610 103.750 58.945 ;
        RECT 104.570 58.610 105.670 58.945 ;
        RECT 106.490 58.610 107.590 58.945 ;
        RECT 108.410 58.610 109.510 58.945 ;
        RECT 110.330 58.610 111.430 58.945 ;
        RECT 112.250 58.610 113.350 58.945 ;
        RECT 114.170 58.610 115.270 58.945 ;
        RECT 116.090 58.610 117.190 58.945 ;
        RECT 118.010 58.610 119.110 58.945 ;
        RECT 119.930 58.610 121.030 58.945 ;
        RECT 121.850 58.610 122.950 58.945 ;
        RECT 123.770 58.610 124.870 58.945 ;
        RECT 125.690 58.610 126.790 58.945 ;
        RECT 127.610 58.610 128.710 58.945 ;
        RECT 129.530 58.610 130.630 58.945 ;
        RECT 131.450 58.610 132.550 58.945 ;
        RECT 133.370 58.610 134.470 58.945 ;
        RECT 135.290 58.610 136.390 58.945 ;
        RECT 137.210 58.610 138.310 58.945 ;
        RECT 139.130 58.610 140.230 58.945 ;
        RECT 141.050 58.610 142.150 58.945 ;
        RECT 142.970 58.610 144.070 58.945 ;
        RECT 144.890 58.610 145.990 58.945 ;
        RECT 146.810 58.610 147.910 58.945 ;
        RECT 148.730 58.610 149.830 58.945 ;
        RECT 150.650 58.610 151.750 58.945 ;
        RECT 152.570 58.610 153.670 58.945 ;
        RECT 154.490 58.610 155.590 58.945 ;
        RECT 156.410 58.610 157.510 58.945 ;
        RECT 158.330 58.610 159.430 58.945 ;
        RECT 160.250 58.610 161.350 58.945 ;
        RECT 162.170 58.610 163.270 58.945 ;
        RECT 164.090 58.610 165.190 58.945 ;
        RECT 166.010 58.610 167.110 58.945 ;
        RECT 167.930 58.610 169.030 58.945 ;
        RECT 169.850 58.610 170.950 58.945 ;
        RECT 171.770 58.610 172.870 58.945 ;
        RECT 173.690 58.610 174.790 58.945 ;
        RECT 175.610 58.610 176.710 58.945 ;
        RECT 177.530 58.610 178.630 58.945 ;
        RECT 179.450 58.610 180.550 58.945 ;
        RECT 181.370 58.610 182.470 58.945 ;
        RECT 183.290 58.610 184.390 58.945 ;
        RECT 185.210 58.610 186.310 58.945 ;
        RECT 187.130 58.610 188.230 58.945 ;
        RECT 189.050 58.610 190.150 58.945 ;
        RECT 190.970 58.610 192.070 58.945 ;
        RECT 192.890 58.610 193.990 58.945 ;
        RECT 194.810 58.610 195.910 58.945 ;
        RECT 196.730 58.610 197.830 58.945 ;
        RECT 198.650 58.610 199.750 58.945 ;
        RECT 200.570 58.610 201.670 58.945 ;
        RECT 202.490 58.610 203.590 58.945 ;
        RECT 204.410 58.610 205.510 58.945 ;
        RECT 206.330 58.610 207.430 58.945 ;
        RECT 208.250 58.610 209.350 58.945 ;
        RECT 210.170 58.610 211.270 58.945 ;
        RECT 212.090 58.610 213.190 58.945 ;
        RECT 214.010 58.610 215.110 58.945 ;
        RECT 215.930 58.610 217.030 58.945 ;
        RECT 217.850 58.610 218.950 58.945 ;
        RECT 219.770 58.610 220.870 58.945 ;
        RECT 221.690 58.610 222.790 58.945 ;
        RECT 223.610 58.610 224.710 58.945 ;
        RECT 225.530 58.610 226.630 58.945 ;
        RECT 227.450 58.610 228.550 58.945 ;
        RECT 229.370 58.610 230.470 58.945 ;
        RECT 231.290 58.610 232.390 58.945 ;
        RECT 233.210 58.610 234.310 58.945 ;
        RECT 235.130 58.610 236.230 58.945 ;
        RECT 237.050 58.610 238.150 58.945 ;
        RECT 238.970 58.610 240.070 58.945 ;
        RECT 240.890 58.610 241.990 58.945 ;
        RECT 242.810 58.610 243.910 58.945 ;
        RECT 244.730 58.610 245.830 58.945 ;
        RECT 246.650 58.610 247.750 58.945 ;
        RECT 248.570 58.610 249.670 58.945 ;
        RECT 250.490 58.610 251.590 58.945 ;
        RECT 252.410 58.610 266.020 58.945 ;
        RECT 1.340 0.610 266.020 58.610 ;
        RECT 1.340 0.100 7.750 0.610 ;
        RECT 8.570 0.100 20.230 0.610 ;
        RECT 21.050 0.100 32.710 0.610 ;
        RECT 33.530 0.100 45.190 0.610 ;
        RECT 46.010 0.100 57.670 0.610 ;
        RECT 58.490 0.100 70.150 0.610 ;
        RECT 70.970 0.100 82.630 0.610 ;
        RECT 83.450 0.100 95.110 0.610 ;
        RECT 95.930 0.100 107.590 0.610 ;
        RECT 108.410 0.100 120.070 0.610 ;
        RECT 120.890 0.100 132.550 0.610 ;
        RECT 133.370 0.100 145.030 0.610 ;
        RECT 145.850 0.100 157.510 0.610 ;
        RECT 158.330 0.100 169.990 0.610 ;
        RECT 170.810 0.100 182.470 0.610 ;
        RECT 183.290 0.100 194.950 0.610 ;
        RECT 195.770 0.100 207.430 0.610 ;
        RECT 208.250 0.100 219.910 0.610 ;
        RECT 220.730 0.100 232.390 0.610 ;
        RECT 233.210 0.100 244.870 0.610 ;
        RECT 245.690 0.100 257.350 0.610 ;
        RECT 258.170 0.100 266.020 0.610 ;
      LAYER Metal4 ;
        RECT 1.295 0.320 257.425 58.900 ;
  END
END S_term_single2
END LIBRARY

