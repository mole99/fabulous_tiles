module S_term_IHP_SRAM (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    S1END,
    S2END,
    S2MID,
    S4END);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;

 sg13g2_buf_1 _00_ (.A(FrameData[0]),
    .X(net1));
 sg13g2_buf_1 _01_ (.A(FrameData[1]),
    .X(net12));
 sg13g2_buf_1 _02_ (.A(FrameData[2]),
    .X(net23));
 sg13g2_buf_1 _03_ (.A(FrameData[3]),
    .X(net26));
 sg13g2_buf_1 _04_ (.A(FrameData[4]),
    .X(net27));
 sg13g2_buf_1 _05_ (.A(FrameData[5]),
    .X(net28));
 sg13g2_buf_1 _06_ (.A(FrameData[6]),
    .X(net29));
 sg13g2_buf_1 _07_ (.A(FrameData[7]),
    .X(net30));
 sg13g2_buf_1 _08_ (.A(FrameData[8]),
    .X(net31));
 sg13g2_buf_1 _09_ (.A(FrameData[9]),
    .X(net32));
 sg13g2_buf_1 _10_ (.A(FrameData[10]),
    .X(net2));
 sg13g2_buf_1 _11_ (.A(FrameData[11]),
    .X(net3));
 sg13g2_buf_1 _12_ (.A(FrameData[12]),
    .X(net4));
 sg13g2_buf_1 _13_ (.A(FrameData[13]),
    .X(net5));
 sg13g2_buf_1 _14_ (.A(FrameData[14]),
    .X(net6));
 sg13g2_buf_1 _15_ (.A(FrameData[15]),
    .X(net7));
 sg13g2_buf_1 _16_ (.A(FrameData[16]),
    .X(net8));
 sg13g2_buf_1 _17_ (.A(FrameData[17]),
    .X(net9));
 sg13g2_buf_1 _18_ (.A(FrameData[18]),
    .X(net10));
 sg13g2_buf_1 _19_ (.A(FrameData[19]),
    .X(net11));
 sg13g2_buf_1 _20_ (.A(FrameData[20]),
    .X(net13));
 sg13g2_buf_1 _21_ (.A(FrameData[21]),
    .X(net14));
 sg13g2_buf_1 _22_ (.A(FrameData[22]),
    .X(net15));
 sg13g2_buf_1 _23_ (.A(FrameData[23]),
    .X(net16));
 sg13g2_buf_1 _24_ (.A(FrameData[24]),
    .X(net17));
 sg13g2_buf_1 _25_ (.A(FrameData[25]),
    .X(net18));
 sg13g2_buf_1 _26_ (.A(FrameData[26]),
    .X(net19));
 sg13g2_buf_1 _27_ (.A(FrameData[27]),
    .X(net20));
 sg13g2_buf_1 _28_ (.A(FrameData[28]),
    .X(net21));
 sg13g2_buf_1 _29_ (.A(FrameData[29]),
    .X(net22));
 sg13g2_buf_1 _30_ (.A(FrameData[30]),
    .X(net24));
 sg13g2_buf_1 _31_ (.A(FrameData[31]),
    .X(net25));
 sg13g2_buf_1 _32_ (.A(FrameStrobe[0]),
    .X(net33));
 sg13g2_buf_1 _33_ (.A(FrameStrobe[1]),
    .X(net44));
 sg13g2_buf_1 _34_ (.A(FrameStrobe[2]),
    .X(net45));
 sg13g2_buf_1 _35_ (.A(FrameStrobe[3]),
    .X(net46));
 sg13g2_buf_1 _36_ (.A(FrameStrobe[4]),
    .X(net47));
 sg13g2_buf_1 _37_ (.A(FrameStrobe[5]),
    .X(net48));
 sg13g2_buf_1 _38_ (.A(FrameStrobe[6]),
    .X(net49));
 sg13g2_buf_1 _39_ (.A(FrameStrobe[7]),
    .X(net50));
 sg13g2_buf_1 _40_ (.A(FrameStrobe[8]),
    .X(net51));
 sg13g2_buf_1 _41_ (.A(FrameStrobe[9]),
    .X(net52));
 sg13g2_buf_1 _42_ (.A(FrameStrobe[10]),
    .X(net34));
 sg13g2_buf_1 _43_ (.A(FrameStrobe[11]),
    .X(net35));
 sg13g2_buf_1 _44_ (.A(FrameStrobe[12]),
    .X(net36));
 sg13g2_buf_1 _45_ (.A(FrameStrobe[13]),
    .X(net37));
 sg13g2_buf_1 _46_ (.A(FrameStrobe[14]),
    .X(net38));
 sg13g2_buf_1 _47_ (.A(FrameStrobe[15]),
    .X(net39));
 sg13g2_buf_1 _48_ (.A(FrameStrobe[16]),
    .X(net40));
 sg13g2_buf_1 _49_ (.A(FrameStrobe[17]),
    .X(net41));
 sg13g2_buf_1 _50_ (.A(FrameStrobe[18]),
    .X(net42));
 sg13g2_buf_1 _51_ (.A(FrameStrobe[19]),
    .X(net43));
 sg13g2_buf_1 _52_ (.A(S1END[3]),
    .X(net53));
 sg13g2_buf_1 _53_ (.A(S1END[2]),
    .X(net54));
 sg13g2_buf_1 _54_ (.A(S1END[1]),
    .X(net55));
 sg13g2_buf_1 _55_ (.A(S1END[0]),
    .X(net56));
 sg13g2_buf_1 _56_ (.A(S2MID[7]),
    .X(net57));
 sg13g2_buf_1 _57_ (.A(S2MID[6]),
    .X(net58));
 sg13g2_buf_1 _58_ (.A(S2MID[5]),
    .X(net59));
 sg13g2_buf_1 _59_ (.A(S2MID[4]),
    .X(net60));
 sg13g2_buf_1 _60_ (.A(S2MID[3]),
    .X(net61));
 sg13g2_buf_1 _61_ (.A(S2MID[2]),
    .X(net62));
 sg13g2_buf_1 _62_ (.A(S2MID[1]),
    .X(net63));
 sg13g2_buf_1 _63_ (.A(S2MID[0]),
    .X(net64));
 sg13g2_buf_1 _64_ (.A(S2END[7]),
    .X(net65));
 sg13g2_buf_1 _65_ (.A(S2END[6]),
    .X(net66));
 sg13g2_buf_1 _66_ (.A(S2END[5]),
    .X(net67));
 sg13g2_buf_1 _67_ (.A(S2END[4]),
    .X(net68));
 sg13g2_buf_1 _68_ (.A(S2END[3]),
    .X(net69));
 sg13g2_buf_1 _69_ (.A(S2END[2]),
    .X(net70));
 sg13g2_buf_1 _70_ (.A(S2END[1]),
    .X(net71));
 sg13g2_buf_1 _71_ (.A(S2END[0]),
    .X(net72));
 sg13g2_buf_1 _72_ (.A(S4END[15]),
    .X(net73));
 sg13g2_buf_1 _73_ (.A(S4END[14]),
    .X(net80));
 sg13g2_buf_1 _74_ (.A(S4END[13]),
    .X(net81));
 sg13g2_buf_1 _75_ (.A(S4END[12]),
    .X(net82));
 sg13g2_buf_1 _76_ (.A(S4END[11]),
    .X(net83));
 sg13g2_buf_1 _77_ (.A(S4END[10]),
    .X(net84));
 sg13g2_buf_1 _78_ (.A(S4END[9]),
    .X(net85));
 sg13g2_buf_1 _79_ (.A(S4END[8]),
    .X(net86));
 sg13g2_buf_1 _80_ (.A(S4END[7]),
    .X(net87));
 sg13g2_buf_1 _81_ (.A(S4END[6]),
    .X(net88));
 sg13g2_buf_1 _82_ (.A(S4END[5]),
    .X(net74));
 sg13g2_buf_1 _83_ (.A(S4END[4]),
    .X(net75));
 sg13g2_buf_1 _84_ (.A(S4END[3]),
    .X(net76));
 sg13g2_buf_1 _85_ (.A(S4END[2]),
    .X(net77));
 sg13g2_buf_1 _86_ (.A(S4END[1]),
    .X(net78));
 sg13g2_buf_1 _87_ (.A(S4END[0]),
    .X(net79));
 sg13g2_buf_1 _88_ (.A(UserCLK),
    .X(net89));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output53 (.A(net53),
    .X(N1BEG[0]));
 sg13g2_buf_1 output54 (.A(net54),
    .X(N1BEG[1]));
 sg13g2_buf_1 output55 (.A(net55),
    .X(N1BEG[2]));
 sg13g2_buf_1 output56 (.A(net56),
    .X(N1BEG[3]));
 sg13g2_buf_1 output57 (.A(net57),
    .X(N2BEG[0]));
 sg13g2_buf_1 output58 (.A(net58),
    .X(N2BEG[1]));
 sg13g2_buf_1 output59 (.A(net59),
    .X(N2BEG[2]));
 sg13g2_buf_1 output60 (.A(net60),
    .X(N2BEG[3]));
 sg13g2_buf_1 output61 (.A(net61),
    .X(N2BEG[4]));
 sg13g2_buf_1 output62 (.A(net62),
    .X(N2BEG[5]));
 sg13g2_buf_1 output63 (.A(net63),
    .X(N2BEG[6]));
 sg13g2_buf_1 output64 (.A(net64),
    .X(N2BEG[7]));
 sg13g2_buf_1 output65 (.A(net65),
    .X(N2BEGb[0]));
 sg13g2_buf_1 output66 (.A(net66),
    .X(N2BEGb[1]));
 sg13g2_buf_1 output67 (.A(net67),
    .X(N2BEGb[2]));
 sg13g2_buf_1 output68 (.A(net68),
    .X(N2BEGb[3]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(N2BEGb[4]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(N2BEGb[5]));
 sg13g2_buf_1 output71 (.A(net71),
    .X(N2BEGb[6]));
 sg13g2_buf_1 output72 (.A(net72),
    .X(N2BEGb[7]));
 sg13g2_buf_1 output73 (.A(net73),
    .X(N4BEG[0]));
 sg13g2_buf_1 output74 (.A(net74),
    .X(N4BEG[10]));
 sg13g2_buf_1 output75 (.A(net75),
    .X(N4BEG[11]));
 sg13g2_buf_1 output76 (.A(net76),
    .X(N4BEG[12]));
 sg13g2_buf_1 output77 (.A(net77),
    .X(N4BEG[13]));
 sg13g2_buf_1 output78 (.A(net78),
    .X(N4BEG[14]));
 sg13g2_buf_1 output79 (.A(net79),
    .X(N4BEG[15]));
 sg13g2_buf_1 output80 (.A(net80),
    .X(N4BEG[1]));
 sg13g2_buf_1 output81 (.A(net81),
    .X(N4BEG[2]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(N4BEG[3]));
 sg13g2_buf_1 output83 (.A(net83),
    .X(N4BEG[4]));
 sg13g2_buf_1 output84 (.A(net84),
    .X(N4BEG[5]));
 sg13g2_buf_1 output85 (.A(net85),
    .X(N4BEG[6]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(N4BEG[7]));
 sg13g2_buf_1 output87 (.A(net87),
    .X(N4BEG[8]));
 sg13g2_buf_1 output88 (.A(net88),
    .X(N4BEG[9]));
 sg13g2_buf_1 output89 (.A(net89),
    .X(UserCLKo));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_fill_1 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_fill_2 FILLER_0_172 ();
 sg13g2_fill_2 FILLER_0_182 ();
 sg13g2_fill_1 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_60 ();
 sg13g2_decap_8 FILLER_1_67 ();
 sg13g2_decap_8 FILLER_1_74 ();
 sg13g2_decap_8 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_88 ();
 sg13g2_decap_8 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_102 ();
 sg13g2_decap_8 FILLER_1_109 ();
 sg13g2_decap_8 FILLER_1_116 ();
 sg13g2_decap_8 FILLER_1_123 ();
 sg13g2_decap_8 FILLER_1_130 ();
 sg13g2_decap_8 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_144 ();
 sg13g2_decap_8 FILLER_1_151 ();
 sg13g2_decap_8 FILLER_1_158 ();
 sg13g2_fill_1 FILLER_1_165 ();
 sg13g2_decap_4 FILLER_1_170 ();
 sg13g2_fill_2 FILLER_1_174 ();
 sg13g2_fill_1 FILLER_1_180 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_57 ();
 sg13g2_decap_8 FILLER_2_64 ();
 sg13g2_decap_4 FILLER_2_71 ();
 sg13g2_fill_1 FILLER_2_75 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_4 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_103 ();
 sg13g2_fill_2 FILLER_2_110 ();
 sg13g2_fill_1 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_117 ();
 sg13g2_fill_2 FILLER_2_124 ();
 sg13g2_fill_1 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_fill_1 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_4 FILLER_2_154 ();
 sg13g2_fill_2 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_fill_2 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_115 ();
 sg13g2_decap_8 FILLER_3_122 ();
 sg13g2_decap_8 FILLER_3_129 ();
 sg13g2_decap_8 FILLER_3_136 ();
 sg13g2_fill_2 FILLER_3_143 ();
 sg13g2_decap_8 FILLER_3_149 ();
 sg13g2_decap_8 FILLER_3_156 ();
 sg13g2_decap_8 FILLER_3_163 ();
 sg13g2_decap_8 FILLER_3_170 ();
 sg13g2_decap_4 FILLER_3_177 ();
 sg13g2_fill_2 FILLER_3_181 ();
 sg13g2_fill_2 FILLER_3_195 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_4 FILLER_4_21 ();
 sg13g2_fill_1 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_30 ();
 sg13g2_decap_4 FILLER_4_37 ();
 sg13g2_decap_8 FILLER_4_45 ();
 sg13g2_decap_4 FILLER_4_52 ();
 sg13g2_fill_1 FILLER_4_56 ();
 sg13g2_fill_2 FILLER_4_65 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_decap_8 FILLER_4_76 ();
 sg13g2_decap_8 FILLER_4_83 ();
 sg13g2_decap_8 FILLER_4_90 ();
 sg13g2_decap_8 FILLER_4_97 ();
 sg13g2_decap_8 FILLER_4_104 ();
 sg13g2_decap_8 FILLER_4_111 ();
 sg13g2_decap_8 FILLER_4_118 ();
 sg13g2_decap_4 FILLER_4_125 ();
 sg13g2_fill_2 FILLER_4_129 ();
 sg13g2_decap_8 FILLER_4_135 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_4 FILLER_4_149 ();
 sg13g2_fill_1 FILLER_4_153 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_fill_2 FILLER_4_179 ();
 sg13g2_fill_1 FILLER_4_181 ();
 sg13g2_fill_2 FILLER_4_190 ();
 sg13g2_fill_1 FILLER_4_192 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_fill_2 FILLER_5_32 ();
 sg13g2_fill_1 FILLER_5_34 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_50 ();
 sg13g2_decap_8 FILLER_5_57 ();
 sg13g2_decap_8 FILLER_5_64 ();
 sg13g2_fill_2 FILLER_5_71 ();
 sg13g2_fill_1 FILLER_5_73 ();
 sg13g2_decap_4 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_82 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_fill_2 FILLER_5_95 ();
 sg13g2_fill_1 FILLER_5_97 ();
 sg13g2_decap_8 FILLER_5_106 ();
 sg13g2_decap_8 FILLER_5_117 ();
 sg13g2_decap_8 FILLER_5_124 ();
 sg13g2_decap_8 FILLER_5_131 ();
 sg13g2_decap_4 FILLER_5_138 ();
 sg13g2_fill_1 FILLER_5_142 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_179 ();
 sg13g2_fill_2 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_26 ();
 sg13g2_decap_8 FILLER_6_37 ();
 sg13g2_decap_8 FILLER_6_44 ();
 sg13g2_decap_8 FILLER_6_51 ();
 sg13g2_decap_8 FILLER_6_58 ();
 sg13g2_decap_8 FILLER_6_65 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_4 FILLER_6_79 ();
 sg13g2_decap_8 FILLER_6_87 ();
 sg13g2_decap_8 FILLER_6_94 ();
 sg13g2_decap_8 FILLER_6_101 ();
 sg13g2_decap_8 FILLER_6_108 ();
 sg13g2_decap_4 FILLER_6_115 ();
 sg13g2_fill_1 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_128 ();
 sg13g2_decap_4 FILLER_6_135 ();
 sg13g2_fill_1 FILLER_6_139 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_fill_2 FILLER_6_195 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_12 ();
 sg13g2_decap_8 FILLER_7_19 ();
 sg13g2_decap_8 FILLER_7_26 ();
 sg13g2_decap_4 FILLER_7_37 ();
 sg13g2_fill_1 FILLER_7_41 ();
 sg13g2_decap_8 FILLER_7_50 ();
 sg13g2_decap_8 FILLER_7_57 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_decap_8 FILLER_7_71 ();
 sg13g2_decap_8 FILLER_7_78 ();
 sg13g2_decap_4 FILLER_7_85 ();
 sg13g2_fill_2 FILLER_7_89 ();
 sg13g2_decap_8 FILLER_7_99 ();
 sg13g2_decap_4 FILLER_7_106 ();
 sg13g2_fill_1 FILLER_7_110 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_decap_8 FILLER_7_137 ();
 sg13g2_decap_4 FILLER_7_144 ();
 sg13g2_fill_2 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_154 ();
 sg13g2_fill_2 FILLER_7_159 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_fill_2 FILLER_7_194 ();
 sg13g2_fill_1 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_13 ();
 sg13g2_decap_8 FILLER_8_20 ();
 sg13g2_decap_8 FILLER_8_27 ();
 sg13g2_decap_8 FILLER_8_34 ();
 sg13g2_decap_8 FILLER_8_41 ();
 sg13g2_decap_8 FILLER_8_48 ();
 sg13g2_decap_8 FILLER_8_55 ();
 sg13g2_decap_8 FILLER_8_62 ();
 sg13g2_decap_8 FILLER_8_69 ();
 sg13g2_decap_8 FILLER_8_76 ();
 sg13g2_decap_8 FILLER_8_83 ();
 sg13g2_fill_1 FILLER_8_90 ();
 sg13g2_decap_8 FILLER_8_99 ();
 sg13g2_decap_8 FILLER_8_106 ();
 sg13g2_decap_8 FILLER_8_113 ();
 sg13g2_decap_8 FILLER_8_120 ();
 sg13g2_decap_8 FILLER_8_127 ();
 sg13g2_decap_8 FILLER_8_134 ();
 sg13g2_decap_8 FILLER_8_141 ();
 sg13g2_decap_8 FILLER_8_148 ();
 sg13g2_fill_2 FILLER_8_155 ();
 sg13g2_fill_1 FILLER_9_20 ();
 sg13g2_decap_8 FILLER_9_69 ();
 sg13g2_decap_8 FILLER_9_76 ();
 sg13g2_decap_8 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_decap_8 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_104 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_200 ();
 sg13g2_fill_1 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_8 FILLER_10_92 ();
 sg13g2_decap_8 FILLER_10_99 ();
 sg13g2_decap_4 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_decap_4 FILLER_10_115 ();
 sg13g2_fill_2 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_8 FILLER_10_132 ();
 sg13g2_fill_1 FILLER_10_143 ();
 sg13g2_fill_1 FILLER_10_200 ();
endmodule
