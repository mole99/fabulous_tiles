module S_term_single2 (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;

 sg13g2_buf_1 _000_ (.A(FrameData[0]),
    .X(net1));
 sg13g2_buf_1 _001_ (.A(FrameData[1]),
    .X(net12));
 sg13g2_buf_1 _002_ (.A(FrameData[2]),
    .X(net23));
 sg13g2_buf_1 _003_ (.A(FrameData[3]),
    .X(net26));
 sg13g2_buf_1 _004_ (.A(FrameData[4]),
    .X(net27));
 sg13g2_buf_1 _005_ (.A(FrameData[5]),
    .X(net28));
 sg13g2_buf_1 _006_ (.A(FrameData[6]),
    .X(net29));
 sg13g2_buf_1 _007_ (.A(FrameData[7]),
    .X(net30));
 sg13g2_buf_1 _008_ (.A(FrameData[8]),
    .X(net31));
 sg13g2_buf_1 _009_ (.A(FrameData[9]),
    .X(net32));
 sg13g2_buf_1 _010_ (.A(FrameData[10]),
    .X(net2));
 sg13g2_buf_1 _011_ (.A(FrameData[11]),
    .X(net3));
 sg13g2_buf_1 _012_ (.A(FrameData[12]),
    .X(net4));
 sg13g2_buf_1 _013_ (.A(FrameData[13]),
    .X(net5));
 sg13g2_buf_1 _014_ (.A(FrameData[14]),
    .X(net6));
 sg13g2_buf_1 _015_ (.A(FrameData[15]),
    .X(net7));
 sg13g2_buf_1 _016_ (.A(FrameData[16]),
    .X(net8));
 sg13g2_buf_1 _017_ (.A(FrameData[17]),
    .X(net9));
 sg13g2_buf_1 _018_ (.A(FrameData[18]),
    .X(net10));
 sg13g2_buf_1 _019_ (.A(FrameData[19]),
    .X(net11));
 sg13g2_buf_1 _020_ (.A(FrameData[20]),
    .X(net13));
 sg13g2_buf_1 _021_ (.A(FrameData[21]),
    .X(net14));
 sg13g2_buf_1 _022_ (.A(FrameData[22]),
    .X(net15));
 sg13g2_buf_1 _023_ (.A(FrameData[23]),
    .X(net16));
 sg13g2_buf_1 _024_ (.A(FrameData[24]),
    .X(net17));
 sg13g2_buf_1 _025_ (.A(FrameData[25]),
    .X(net18));
 sg13g2_buf_1 _026_ (.A(FrameData[26]),
    .X(net19));
 sg13g2_buf_1 _027_ (.A(FrameData[27]),
    .X(net20));
 sg13g2_buf_1 _028_ (.A(FrameData[28]),
    .X(net21));
 sg13g2_buf_1 _029_ (.A(FrameData[29]),
    .X(net22));
 sg13g2_buf_1 _030_ (.A(FrameData[30]),
    .X(net24));
 sg13g2_buf_1 _031_ (.A(FrameData[31]),
    .X(net25));
 sg13g2_buf_1 _032_ (.A(FrameStrobe[0]),
    .X(net33));
 sg13g2_buf_1 _033_ (.A(FrameStrobe[1]),
    .X(net44));
 sg13g2_buf_1 _034_ (.A(FrameStrobe[2]),
    .X(net45));
 sg13g2_buf_1 _035_ (.A(FrameStrobe[3]),
    .X(net46));
 sg13g2_buf_1 _036_ (.A(FrameStrobe[4]),
    .X(net47));
 sg13g2_buf_1 _037_ (.A(FrameStrobe[5]),
    .X(net48));
 sg13g2_buf_1 _038_ (.A(FrameStrobe[6]),
    .X(net49));
 sg13g2_buf_1 _039_ (.A(FrameStrobe[7]),
    .X(net50));
 sg13g2_buf_1 _040_ (.A(FrameStrobe[8]),
    .X(net51));
 sg13g2_buf_1 _041_ (.A(FrameStrobe[9]),
    .X(net52));
 sg13g2_buf_1 _042_ (.A(FrameStrobe[10]),
    .X(net34));
 sg13g2_buf_1 _043_ (.A(FrameStrobe[11]),
    .X(net35));
 sg13g2_buf_1 _044_ (.A(FrameStrobe[12]),
    .X(net36));
 sg13g2_buf_1 _045_ (.A(FrameStrobe[13]),
    .X(net37));
 sg13g2_buf_1 _046_ (.A(FrameStrobe[14]),
    .X(net38));
 sg13g2_buf_1 _047_ (.A(FrameStrobe[15]),
    .X(net39));
 sg13g2_buf_1 _048_ (.A(FrameStrobe[16]),
    .X(net40));
 sg13g2_buf_1 _049_ (.A(FrameStrobe[17]),
    .X(net41));
 sg13g2_buf_1 _050_ (.A(FrameStrobe[18]),
    .X(net42));
 sg13g2_buf_1 _051_ (.A(FrameStrobe[19]),
    .X(net43));
 sg13g2_buf_1 _052_ (.A(S1END[3]),
    .X(net53));
 sg13g2_buf_1 _053_ (.A(S1END[2]),
    .X(net54));
 sg13g2_buf_1 _054_ (.A(S1END[1]),
    .X(net55));
 sg13g2_buf_1 _055_ (.A(S1END[0]),
    .X(net56));
 sg13g2_buf_1 _056_ (.A(S2MID[7]),
    .X(net57));
 sg13g2_buf_1 _057_ (.A(S2MID[6]),
    .X(net58));
 sg13g2_buf_1 _058_ (.A(S2MID[5]),
    .X(net59));
 sg13g2_buf_1 _059_ (.A(S2MID[4]),
    .X(net60));
 sg13g2_buf_1 _060_ (.A(S2MID[3]),
    .X(net61));
 sg13g2_buf_1 _061_ (.A(S2MID[2]),
    .X(net62));
 sg13g2_buf_1 _062_ (.A(S2MID[1]),
    .X(net63));
 sg13g2_buf_1 _063_ (.A(S2MID[0]),
    .X(net64));
 sg13g2_buf_1 _064_ (.A(S2END[7]),
    .X(net65));
 sg13g2_buf_1 _065_ (.A(S2END[6]),
    .X(net66));
 sg13g2_buf_1 _066_ (.A(S2END[5]),
    .X(net67));
 sg13g2_buf_1 _067_ (.A(S2END[4]),
    .X(net68));
 sg13g2_buf_1 _068_ (.A(S2END[3]),
    .X(net69));
 sg13g2_buf_1 _069_ (.A(S2END[2]),
    .X(net70));
 sg13g2_buf_1 _070_ (.A(S2END[1]),
    .X(net71));
 sg13g2_buf_1 _071_ (.A(S2END[0]),
    .X(net72));
 sg13g2_buf_1 _072_ (.A(S4END[15]),
    .X(net73));
 sg13g2_buf_1 _073_ (.A(S4END[14]),
    .X(net80));
 sg13g2_buf_1 _074_ (.A(S4END[13]),
    .X(net81));
 sg13g2_buf_1 _075_ (.A(S4END[12]),
    .X(net82));
 sg13g2_buf_1 _076_ (.A(S4END[11]),
    .X(net83));
 sg13g2_buf_1 _077_ (.A(S4END[10]),
    .X(net84));
 sg13g2_buf_1 _078_ (.A(S4END[9]),
    .X(net85));
 sg13g2_buf_1 _079_ (.A(S4END[8]),
    .X(net86));
 sg13g2_buf_1 _080_ (.A(S4END[7]),
    .X(net87));
 sg13g2_buf_1 _081_ (.A(S4END[6]),
    .X(net88));
 sg13g2_buf_1 _082_ (.A(S4END[5]),
    .X(net74));
 sg13g2_buf_1 _083_ (.A(S4END[4]),
    .X(net75));
 sg13g2_buf_1 _084_ (.A(S4END[3]),
    .X(net76));
 sg13g2_buf_1 _085_ (.A(S4END[2]),
    .X(net77));
 sg13g2_buf_1 _086_ (.A(S4END[1]),
    .X(net78));
 sg13g2_buf_1 _087_ (.A(S4END[0]),
    .X(net79));
 sg13g2_buf_1 _088_ (.A(SS4END[15]),
    .X(net89));
 sg13g2_buf_1 _089_ (.A(SS4END[14]),
    .X(net96));
 sg13g2_buf_1 _090_ (.A(SS4END[13]),
    .X(net97));
 sg13g2_buf_1 _091_ (.A(SS4END[12]),
    .X(net98));
 sg13g2_buf_1 _092_ (.A(SS4END[11]),
    .X(net99));
 sg13g2_buf_1 _093_ (.A(SS4END[10]),
    .X(net100));
 sg13g2_buf_1 _094_ (.A(SS4END[9]),
    .X(net101));
 sg13g2_buf_1 _095_ (.A(SS4END[8]),
    .X(net102));
 sg13g2_buf_1 _096_ (.A(SS4END[7]),
    .X(net103));
 sg13g2_buf_1 _097_ (.A(SS4END[6]),
    .X(net104));
 sg13g2_buf_1 _098_ (.A(SS4END[5]),
    .X(net90));
 sg13g2_buf_1 _099_ (.A(SS4END[4]),
    .X(net91));
 sg13g2_buf_1 _100_ (.A(SS4END[3]),
    .X(net92));
 sg13g2_buf_1 _101_ (.A(SS4END[2]),
    .X(net93));
 sg13g2_buf_1 _102_ (.A(SS4END[1]),
    .X(net94));
 sg13g2_buf_1 _103_ (.A(SS4END[0]),
    .X(net95));
 sg13g2_buf_1 _104_ (.A(UserCLK),
    .X(net105));
 sg13g2_buf_1 output1 (.A(net1),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output27 (.A(net27),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output28 (.A(net28),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output29 (.A(net29),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output30 (.A(net30),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output31 (.A(net31),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output32 (.A(net32),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output53 (.A(net53),
    .X(N1BEG[0]));
 sg13g2_buf_1 output54 (.A(net54),
    .X(N1BEG[1]));
 sg13g2_buf_1 output55 (.A(net55),
    .X(N1BEG[2]));
 sg13g2_buf_1 output56 (.A(net56),
    .X(N1BEG[3]));
 sg13g2_buf_1 output57 (.A(net57),
    .X(N2BEG[0]));
 sg13g2_buf_1 output58 (.A(net58),
    .X(N2BEG[1]));
 sg13g2_buf_1 output59 (.A(net59),
    .X(N2BEG[2]));
 sg13g2_buf_1 output60 (.A(net60),
    .X(N2BEG[3]));
 sg13g2_buf_1 output61 (.A(net61),
    .X(N2BEG[4]));
 sg13g2_buf_1 output62 (.A(net62),
    .X(N2BEG[5]));
 sg13g2_buf_1 output63 (.A(net63),
    .X(N2BEG[6]));
 sg13g2_buf_1 output64 (.A(net64),
    .X(N2BEG[7]));
 sg13g2_buf_1 output65 (.A(net65),
    .X(N2BEGb[0]));
 sg13g2_buf_1 output66 (.A(net66),
    .X(N2BEGb[1]));
 sg13g2_buf_1 output67 (.A(net67),
    .X(N2BEGb[2]));
 sg13g2_buf_1 output68 (.A(net68),
    .X(N2BEGb[3]));
 sg13g2_buf_1 output69 (.A(net69),
    .X(N2BEGb[4]));
 sg13g2_buf_1 output70 (.A(net70),
    .X(N2BEGb[5]));
 sg13g2_buf_1 output71 (.A(net71),
    .X(N2BEGb[6]));
 sg13g2_buf_1 output72 (.A(net72),
    .X(N2BEGb[7]));
 sg13g2_buf_1 output73 (.A(net73),
    .X(N4BEG[0]));
 sg13g2_buf_1 output74 (.A(net74),
    .X(N4BEG[10]));
 sg13g2_buf_1 output75 (.A(net75),
    .X(N4BEG[11]));
 sg13g2_buf_1 output76 (.A(net76),
    .X(N4BEG[12]));
 sg13g2_buf_1 output77 (.A(net77),
    .X(N4BEG[13]));
 sg13g2_buf_1 output78 (.A(net78),
    .X(N4BEG[14]));
 sg13g2_buf_1 output79 (.A(net79),
    .X(N4BEG[15]));
 sg13g2_buf_1 output80 (.A(net80),
    .X(N4BEG[1]));
 sg13g2_buf_1 output81 (.A(net81),
    .X(N4BEG[2]));
 sg13g2_buf_1 output82 (.A(net82),
    .X(N4BEG[3]));
 sg13g2_buf_1 output83 (.A(net83),
    .X(N4BEG[4]));
 sg13g2_buf_1 output84 (.A(net84),
    .X(N4BEG[5]));
 sg13g2_buf_1 output85 (.A(net85),
    .X(N4BEG[6]));
 sg13g2_buf_1 output86 (.A(net86),
    .X(N4BEG[7]));
 sg13g2_buf_1 output87 (.A(net87),
    .X(N4BEG[8]));
 sg13g2_buf_1 output88 (.A(net88),
    .X(N4BEG[9]));
 sg13g2_buf_1 output89 (.A(net89),
    .X(NN4BEG[0]));
 sg13g2_buf_1 output90 (.A(net90),
    .X(NN4BEG[10]));
 sg13g2_buf_1 output91 (.A(net91),
    .X(NN4BEG[11]));
 sg13g2_buf_1 output92 (.A(net92),
    .X(NN4BEG[12]));
 sg13g2_buf_1 output93 (.A(net93),
    .X(NN4BEG[13]));
 sg13g2_buf_1 output94 (.A(net94),
    .X(NN4BEG[14]));
 sg13g2_buf_1 output95 (.A(net95),
    .X(NN4BEG[15]));
 sg13g2_buf_1 output96 (.A(net96),
    .X(NN4BEG[1]));
 sg13g2_buf_1 output97 (.A(net97),
    .X(NN4BEG[2]));
 sg13g2_buf_1 output98 (.A(net98),
    .X(NN4BEG[3]));
 sg13g2_buf_1 output99 (.A(net99),
    .X(NN4BEG[4]));
 sg13g2_buf_1 output100 (.A(net100),
    .X(NN4BEG[5]));
 sg13g2_buf_1 output101 (.A(net101),
    .X(NN4BEG[6]));
 sg13g2_buf_1 output102 (.A(net102),
    .X(NN4BEG[7]));
 sg13g2_buf_1 output103 (.A(net103),
    .X(NN4BEG[8]));
 sg13g2_buf_1 output104 (.A(net104),
    .X(NN4BEG[9]));
 sg13g2_buf_1 output105 (.A(net105),
    .X(UserCLKo));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_4 FILLER_1_245 ();
 sg13g2_fill_1 FILLER_1_249 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_decap_8 FILLER_1_261 ();
 sg13g2_decap_8 FILLER_1_268 ();
 sg13g2_decap_8 FILLER_1_275 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_decap_8 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_decap_8 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_1_436 ();
 sg13g2_decap_8 FILLER_1_443 ();
 sg13g2_decap_8 FILLER_1_450 ();
 sg13g2_decap_8 FILLER_1_457 ();
 sg13g2_decap_8 FILLER_1_464 ();
 sg13g2_decap_8 FILLER_1_471 ();
 sg13g2_decap_8 FILLER_1_478 ();
 sg13g2_decap_8 FILLER_1_485 ();
 sg13g2_decap_8 FILLER_1_492 ();
 sg13g2_decap_8 FILLER_1_499 ();
 sg13g2_decap_8 FILLER_1_506 ();
 sg13g2_decap_4 FILLER_1_513 ();
 sg13g2_fill_2 FILLER_1_517 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_4 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_218 ();
 sg13g2_fill_2 FILLER_2_225 ();
 sg13g2_fill_1 FILLER_2_227 ();
 sg13g2_decap_8 FILLER_2_232 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_fill_2 FILLER_2_244 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_286 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_300 ();
 sg13g2_decap_8 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_2_412 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_8 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_2_433 ();
 sg13g2_decap_8 FILLER_2_440 ();
 sg13g2_decap_8 FILLER_2_447 ();
 sg13g2_decap_8 FILLER_2_454 ();
 sg13g2_decap_8 FILLER_2_461 ();
 sg13g2_decap_8 FILLER_2_468 ();
 sg13g2_decap_8 FILLER_2_475 ();
 sg13g2_decap_8 FILLER_2_482 ();
 sg13g2_decap_8 FILLER_2_489 ();
 sg13g2_decap_8 FILLER_2_496 ();
 sg13g2_decap_8 FILLER_2_503 ();
 sg13g2_decap_8 FILLER_2_510 ();
 sg13g2_decap_4 FILLER_2_517 ();
 sg13g2_fill_2 FILLER_2_521 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_4 FILLER_3_196 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_fill_1 FILLER_3_221 ();
 sg13g2_decap_4 FILLER_3_234 ();
 sg13g2_decap_8 FILLER_3_262 ();
 sg13g2_decap_8 FILLER_3_269 ();
 sg13g2_decap_8 FILLER_3_276 ();
 sg13g2_decap_8 FILLER_3_283 ();
 sg13g2_decap_8 FILLER_3_290 ();
 sg13g2_decap_8 FILLER_3_297 ();
 sg13g2_decap_8 FILLER_3_304 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_332 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_3_409 ();
 sg13g2_decap_8 FILLER_3_416 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_3_430 ();
 sg13g2_decap_8 FILLER_3_437 ();
 sg13g2_decap_8 FILLER_3_444 ();
 sg13g2_decap_8 FILLER_3_451 ();
 sg13g2_decap_8 FILLER_3_458 ();
 sg13g2_decap_8 FILLER_3_465 ();
 sg13g2_decap_8 FILLER_3_472 ();
 sg13g2_decap_8 FILLER_3_479 ();
 sg13g2_decap_8 FILLER_3_486 ();
 sg13g2_decap_8 FILLER_3_493 ();
 sg13g2_decap_8 FILLER_3_500 ();
 sg13g2_decap_8 FILLER_3_507 ();
 sg13g2_decap_8 FILLER_3_514 ();
 sg13g2_fill_2 FILLER_3_521 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_fill_2 FILLER_4_315 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_fill_2 FILLER_4_322 ();
 sg13g2_fill_1 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_4 FILLER_4_518 ();
 sg13g2_fill_1 FILLER_4_522 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_4 FILLER_5_270 ();
 sg13g2_fill_1 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_279 ();
 sg13g2_decap_8 FILLER_5_286 ();
 sg13g2_decap_4 FILLER_5_293 ();
 sg13g2_fill_1 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_fill_1 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_321 ();
 sg13g2_decap_4 FILLER_5_328 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_fill_2 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_475 ();
 sg13g2_decap_8 FILLER_5_482 ();
 sg13g2_decap_8 FILLER_5_489 ();
 sg13g2_decap_4 FILLER_5_496 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_4 FILLER_5_518 ();
 sg13g2_fill_1 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_4 FILLER_6_224 ();
 sg13g2_fill_1 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_237 ();
 sg13g2_decap_4 FILLER_6_244 ();
 sg13g2_fill_2 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_258 ();
 sg13g2_decap_8 FILLER_6_265 ();
 sg13g2_decap_8 FILLER_6_272 ();
 sg13g2_decap_8 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_293 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_8 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_335 ();
 sg13g2_decap_8 FILLER_6_342 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_4 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_404 ();
 sg13g2_decap_8 FILLER_6_411 ();
 sg13g2_decap_8 FILLER_6_418 ();
 sg13g2_fill_2 FILLER_6_425 ();
 sg13g2_fill_1 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_432 ();
 sg13g2_decap_8 FILLER_6_439 ();
 sg13g2_decap_8 FILLER_6_446 ();
 sg13g2_decap_8 FILLER_6_453 ();
 sg13g2_decap_8 FILLER_6_460 ();
 sg13g2_decap_8 FILLER_6_467 ();
 sg13g2_decap_8 FILLER_6_474 ();
 sg13g2_decap_8 FILLER_6_481 ();
 sg13g2_decap_8 FILLER_6_488 ();
 sg13g2_decap_4 FILLER_6_495 ();
 sg13g2_fill_2 FILLER_6_499 ();
 sg13g2_decap_8 FILLER_6_505 ();
 sg13g2_decap_8 FILLER_6_512 ();
 sg13g2_decap_4 FILLER_6_519 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_fill_2 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_100 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_fill_2 FILLER_7_114 ();
 sg13g2_fill_1 FILLER_7_116 ();
 sg13g2_decap_4 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_125 ();
 sg13g2_decap_4 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_139 ();
 sg13g2_decap_8 FILLER_7_148 ();
 sg13g2_decap_8 FILLER_7_155 ();
 sg13g2_fill_2 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_277 ();
 sg13g2_fill_2 FILLER_7_284 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_fill_2 FILLER_7_375 ();
 sg13g2_fill_2 FILLER_7_381 ();
 sg13g2_fill_1 FILLER_7_383 ();
 sg13g2_decap_4 FILLER_7_388 ();
 sg13g2_fill_1 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_8 FILLER_7_404 ();
 sg13g2_decap_8 FILLER_7_411 ();
 sg13g2_decap_8 FILLER_7_418 ();
 sg13g2_decap_8 FILLER_7_425 ();
 sg13g2_decap_8 FILLER_7_432 ();
 sg13g2_decap_8 FILLER_7_439 ();
 sg13g2_decap_8 FILLER_7_446 ();
 sg13g2_decap_8 FILLER_7_453 ();
 sg13g2_decap_8 FILLER_7_460 ();
 sg13g2_decap_8 FILLER_7_467 ();
 sg13g2_decap_8 FILLER_7_474 ();
 sg13g2_decap_8 FILLER_7_481 ();
 sg13g2_decap_8 FILLER_7_488 ();
 sg13g2_decap_8 FILLER_7_495 ();
 sg13g2_decap_8 FILLER_7_502 ();
 sg13g2_decap_8 FILLER_7_509 ();
 sg13g2_decap_8 FILLER_7_516 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_fill_1 FILLER_8_32 ();
 sg13g2_decap_4 FILLER_8_37 ();
 sg13g2_fill_1 FILLER_8_41 ();
 sg13g2_decap_4 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_50 ();
 sg13g2_decap_8 FILLER_8_55 ();
 sg13g2_decap_8 FILLER_8_62 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_fill_2 FILLER_8_109 ();
 sg13g2_fill_1 FILLER_8_111 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_fill_2 FILLER_8_144 ();
 sg13g2_fill_1 FILLER_8_146 ();
 sg13g2_fill_2 FILLER_8_183 ();
 sg13g2_fill_1 FILLER_8_185 ();
 sg13g2_decap_4 FILLER_8_194 ();
 sg13g2_fill_1 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_208 ();
 sg13g2_decap_8 FILLER_8_215 ();
 sg13g2_decap_8 FILLER_8_222 ();
 sg13g2_decap_8 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_236 ();
 sg13g2_decap_8 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_250 ();
 sg13g2_decap_8 FILLER_8_257 ();
 sg13g2_decap_8 FILLER_8_264 ();
 sg13g2_decap_8 FILLER_8_271 ();
 sg13g2_decap_4 FILLER_8_278 ();
 sg13g2_fill_1 FILLER_8_282 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_fill_1 FILLER_8_348 ();
 sg13g2_fill_1 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_fill_1 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_fill_2 FILLER_9_210 ();
 sg13g2_fill_1 FILLER_9_212 ();
 sg13g2_fill_1 FILLER_9_217 ();
 sg13g2_fill_2 FILLER_9_226 ();
 sg13g2_fill_2 FILLER_9_232 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_fill_1 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_324 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_decap_8 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_422 ();
 sg13g2_decap_8 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_9_436 ();
 sg13g2_decap_8 FILLER_9_443 ();
 sg13g2_decap_8 FILLER_9_450 ();
 sg13g2_decap_8 FILLER_9_457 ();
 sg13g2_decap_8 FILLER_9_464 ();
 sg13g2_decap_8 FILLER_9_471 ();
 sg13g2_decap_8 FILLER_9_478 ();
 sg13g2_decap_8 FILLER_9_485 ();
 sg13g2_decap_8 FILLER_9_492 ();
 sg13g2_decap_8 FILLER_9_499 ();
 sg13g2_fill_1 FILLER_9_506 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_16 ();
 sg13g2_decap_8 FILLER_10_225 ();
 sg13g2_decap_8 FILLER_10_232 ();
 sg13g2_decap_8 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_246 ();
 sg13g2_decap_8 FILLER_10_253 ();
 sg13g2_decap_8 FILLER_10_260 ();
 sg13g2_decap_8 FILLER_10_267 ();
 sg13g2_decap_8 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_281 ();
 sg13g2_decap_8 FILLER_10_288 ();
 sg13g2_decap_8 FILLER_10_295 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_decap_8 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_10_414 ();
 sg13g2_decap_8 FILLER_10_421 ();
 sg13g2_decap_4 FILLER_10_428 ();
 sg13g2_fill_1 FILLER_10_432 ();
 sg13g2_fill_2 FILLER_10_517 ();
endmodule
