magic
tech sky130A
magscale 1 2
timestamp 1740331796
<< viali >>
rect 1593 42313 1627 42347
rect 2145 42313 2179 42347
rect 2605 42313 2639 42347
rect 2973 42313 3007 42347
rect 3433 42313 3467 42347
rect 3893 42313 3927 42347
rect 4353 42313 4387 42347
rect 4813 42313 4847 42347
rect 5273 42313 5307 42347
rect 5641 42313 5675 42347
rect 6009 42313 6043 42347
rect 6745 42313 6779 42347
rect 7297 42313 7331 42347
rect 7665 42313 7699 42347
rect 8401 42313 8435 42347
rect 9505 42313 9539 42347
rect 1777 42177 1811 42211
rect 1961 42177 1995 42211
rect 2421 42177 2455 42211
rect 3157 42177 3191 42211
rect 3617 42177 3651 42211
rect 4077 42177 4111 42211
rect 4537 42177 4571 42211
rect 4997 42177 5031 42211
rect 5457 42177 5491 42211
rect 5825 42177 5859 42211
rect 6193 42177 6227 42211
rect 6561 42177 6595 42211
rect 7481 42177 7515 42211
rect 7849 42177 7883 42211
rect 8585 42177 8619 42211
rect 9229 42177 9263 42211
rect 9321 42177 9355 42211
rect 9045 42041 9079 42075
rect 7021 41973 7055 42007
rect 8125 41973 8159 42007
rect 1409 41769 1443 41803
rect 6561 41769 6595 41803
rect 6745 41769 6779 41803
rect 7481 41769 7515 41803
rect 8585 41769 8619 41803
rect 9321 41769 9355 41803
rect 8125 41701 8159 41735
rect 1593 41565 1627 41599
rect 6285 41565 6319 41599
rect 6377 41565 6411 41599
rect 6929 41565 6963 41599
rect 7205 41565 7239 41599
rect 7297 41565 7331 41599
rect 7573 41565 7607 41599
rect 8033 41565 8067 41599
rect 8309 41565 8343 41599
rect 8769 41565 8803 41599
rect 9137 41565 9171 41599
rect 9505 41565 9539 41599
rect 6193 41429 6227 41463
rect 7021 41429 7055 41463
rect 7849 41429 7883 41463
rect 9689 41429 9723 41463
rect 6745 41225 6779 41259
rect 7389 41225 7423 41259
rect 7941 41225 7975 41259
rect 8217 41225 8251 41259
rect 8677 41225 8711 41259
rect 9229 41225 9263 41259
rect 9505 41225 9539 41259
rect 1501 41089 1535 41123
rect 6929 41089 6963 41123
rect 7021 41089 7055 41123
rect 7573 41089 7607 41123
rect 7665 41089 7699 41123
rect 8125 41089 8159 41123
rect 8401 41089 8435 41123
rect 8861 41089 8895 41123
rect 9413 41089 9447 41123
rect 9689 41089 9723 41123
rect 1685 40953 1719 40987
rect 7849 40953 7883 40987
rect 8585 40885 8619 40919
rect 9045 40885 9079 40919
rect 7389 40681 7423 40715
rect 8585 40681 8619 40715
rect 8953 40681 8987 40715
rect 7573 40477 7607 40511
rect 8769 40477 8803 40511
rect 9137 40477 9171 40511
rect 1501 40409 1535 40443
rect 1685 40409 1719 40443
rect 7941 40409 7975 40443
rect 6837 40341 6871 40375
rect 7757 40341 7791 40375
rect 8309 40341 8343 40375
rect 9321 40341 9355 40375
rect 9597 40341 9631 40375
rect 8953 40001 8987 40035
rect 9137 40001 9171 40035
rect 9505 40001 9539 40035
rect 8769 39865 8803 39899
rect 9321 39865 9355 39899
rect 7389 39797 7423 39831
rect 8677 39797 8711 39831
rect 9689 39797 9723 39831
rect 9321 39525 9355 39559
rect 5181 39389 5215 39423
rect 5457 39389 5491 39423
rect 9137 39389 9171 39423
rect 9505 39389 9539 39423
rect 1501 39321 1535 39355
rect 1685 39321 1719 39355
rect 4445 39253 4479 39287
rect 9689 39253 9723 39287
rect 9321 39049 9355 39083
rect 1501 38913 1535 38947
rect 3893 38913 3927 38947
rect 4445 38913 4479 38947
rect 4721 38913 4755 38947
rect 5733 38913 5767 38947
rect 6377 38913 6411 38947
rect 8769 38913 8803 38947
rect 9137 38913 9171 38947
rect 9505 38913 9539 38947
rect 1685 38777 1719 38811
rect 8953 38777 8987 38811
rect 4077 38709 4111 38743
rect 5457 38709 5491 38743
rect 5917 38709 5951 38743
rect 6561 38709 6595 38743
rect 9689 38709 9723 38743
rect 6009 38505 6043 38539
rect 4813 38437 4847 38471
rect 9321 38437 9355 38471
rect 4353 38369 4387 38403
rect 5206 38369 5240 38403
rect 5365 38369 5399 38403
rect 6469 38369 6503 38403
rect 1961 38301 1995 38335
rect 2237 38301 2271 38335
rect 4169 38301 4203 38335
rect 5089 38301 5123 38335
rect 6193 38301 6227 38335
rect 6745 38301 6779 38335
rect 8493 38301 8527 38335
rect 9137 38301 9171 38335
rect 9505 38301 9539 38335
rect 1501 38233 1535 38267
rect 1593 38165 1627 38199
rect 2973 38165 3007 38199
rect 6377 38165 6411 38199
rect 7481 38165 7515 38199
rect 8677 38165 8711 38199
rect 9689 38165 9723 38199
rect 4353 37961 4387 37995
rect 9321 37961 9355 37995
rect 1409 37825 1443 37859
rect 1685 37825 1719 37859
rect 4721 37825 4755 37859
rect 5641 37825 5675 37859
rect 6377 37825 6411 37859
rect 8677 37825 8711 37859
rect 8769 37825 8803 37859
rect 9137 37825 9171 37859
rect 9505 37825 9539 37859
rect 2513 37757 2547 37791
rect 2697 37757 2731 37791
rect 3157 37757 3191 37791
rect 3433 37757 3467 37791
rect 3550 37757 3584 37791
rect 3709 37757 3743 37791
rect 4445 37757 4479 37791
rect 5825 37689 5859 37723
rect 8953 37689 8987 37723
rect 2421 37621 2455 37655
rect 5457 37621 5491 37655
rect 7665 37621 7699 37655
rect 8493 37621 8527 37655
rect 9689 37621 9723 37655
rect 5549 37417 5583 37451
rect 7021 37417 7055 37451
rect 7573 37281 7607 37315
rect 1685 37213 1719 37247
rect 1777 37213 1811 37247
rect 2145 37213 2179 37247
rect 2421 37213 2455 37247
rect 4261 37213 4295 37247
rect 4537 37213 4571 37247
rect 7849 37213 7883 37247
rect 9137 37213 9171 37247
rect 9505 37213 9539 37247
rect 1501 37145 1535 37179
rect 5733 37145 5767 37179
rect 1961 37077 1995 37111
rect 2329 37077 2363 37111
rect 2605 37077 2639 37111
rect 5273 37077 5307 37111
rect 8585 37077 8619 37111
rect 9321 37077 9355 37111
rect 9689 37077 9723 37111
rect 5825 36873 5859 36907
rect 7205 36873 7239 36907
rect 2053 36737 2087 36771
rect 3985 36737 4019 36771
rect 4528 36737 4562 36771
rect 6009 36737 6043 36771
rect 7849 36737 7883 36771
rect 8861 36737 8895 36771
rect 9137 36737 9171 36771
rect 9505 36737 9539 36771
rect 1777 36669 1811 36703
rect 4261 36669 4295 36703
rect 7987 36669 8021 36703
rect 8125 36669 8159 36703
rect 8401 36669 8435 36703
rect 9045 36669 9079 36703
rect 9321 36601 9355 36635
rect 2789 36533 2823 36567
rect 4169 36533 4203 36567
rect 5641 36533 5675 36567
rect 9689 36533 9723 36567
rect 4261 36329 4295 36363
rect 2053 36125 2087 36159
rect 2329 36125 2363 36159
rect 7573 36125 7607 36159
rect 7849 36125 7883 36159
rect 9137 36125 9171 36159
rect 9505 36125 9539 36159
rect 1501 36057 1535 36091
rect 1685 36057 1719 36091
rect 5549 36057 5583 36091
rect 5733 36057 5767 36091
rect 7481 36057 7515 36091
rect 3065 35989 3099 36023
rect 7021 35989 7055 36023
rect 8585 35989 8619 36023
rect 9321 35989 9355 36023
rect 9689 35989 9723 36023
rect 1961 35785 1995 35819
rect 4353 35785 4387 35819
rect 6561 35785 6595 35819
rect 7665 35785 7699 35819
rect 1501 35649 1535 35683
rect 1777 35649 1811 35683
rect 2237 35649 2271 35683
rect 2513 35649 2547 35683
rect 3709 35649 3743 35683
rect 6377 35649 6411 35683
rect 8309 35649 8343 35683
rect 8585 35649 8619 35683
rect 2697 35581 2731 35615
rect 3157 35581 3191 35615
rect 3433 35581 3467 35615
rect 3571 35581 3605 35615
rect 8468 35581 8502 35615
rect 8861 35581 8895 35615
rect 9321 35581 9355 35615
rect 9505 35581 9539 35615
rect 1685 35513 1719 35547
rect 2421 35445 2455 35479
rect 1961 35241 1995 35275
rect 8217 35241 8251 35275
rect 8677 35173 8711 35207
rect 1777 35037 1811 35071
rect 5365 35037 5399 35071
rect 5641 35037 5675 35071
rect 5733 35037 5767 35071
rect 7205 35037 7239 35071
rect 7481 35037 7515 35071
rect 8493 35037 8527 35071
rect 8953 35037 8987 35071
rect 9321 35037 9355 35071
rect 6000 34969 6034 35003
rect 4629 34901 4663 34935
rect 7113 34901 7147 34935
rect 9137 34901 9171 34935
rect 9505 34901 9539 34935
rect 1593 34697 1627 34731
rect 5181 34697 5215 34731
rect 6561 34697 6595 34731
rect 1869 34629 1903 34663
rect 8033 34629 8067 34663
rect 1501 34561 1535 34595
rect 3249 34561 3283 34595
rect 4813 34561 4847 34595
rect 5917 34561 5951 34595
rect 6377 34561 6411 34595
rect 7205 34561 7239 34595
rect 2053 34493 2087 34527
rect 2973 34493 3007 34527
rect 5089 34493 5123 34527
rect 6193 34493 6227 34527
rect 6929 34493 6963 34527
rect 9321 34425 9355 34459
rect 3985 34357 4019 34391
rect 4077 34357 4111 34391
rect 7941 34357 7975 34391
rect 1593 34085 1627 34119
rect 4445 34085 4479 34119
rect 8677 34085 8711 34119
rect 1685 34017 1719 34051
rect 4997 34017 5031 34051
rect 7113 34017 7147 34051
rect 1409 33949 1443 33983
rect 1961 33949 1995 33983
rect 3433 33949 3467 33983
rect 3801 33949 3835 33983
rect 3985 33949 4019 33983
rect 4721 33949 4755 33983
rect 4838 33949 4872 33983
rect 5641 33949 5675 33983
rect 5733 33949 5767 33983
rect 7389 33949 7423 33983
rect 8217 33949 8251 33983
rect 8493 33949 8527 33983
rect 9137 33949 9171 33983
rect 9505 33949 9539 33983
rect 2697 33813 2731 33847
rect 3617 33813 3651 33847
rect 5917 33813 5951 33847
rect 8125 33813 8159 33847
rect 8401 33813 8435 33847
rect 9321 33813 9355 33847
rect 9689 33813 9723 33847
rect 1593 33609 1627 33643
rect 9413 33609 9447 33643
rect 2421 33541 2455 33575
rect 1501 33473 1535 33507
rect 1869 33473 1903 33507
rect 8769 33473 8803 33507
rect 3065 33405 3099 33439
rect 3224 33405 3258 33439
rect 3341 33405 3375 33439
rect 3617 33405 3651 33439
rect 4077 33405 4111 33439
rect 4261 33405 4295 33439
rect 7573 33405 7607 33439
rect 7757 33405 7791 33439
rect 8217 33405 8251 33439
rect 8493 33405 8527 33439
rect 8631 33405 8665 33439
rect 2053 33337 2087 33371
rect 9505 33337 9539 33371
rect 1593 33065 1627 33099
rect 2697 33065 2731 33099
rect 6837 32997 6871 33031
rect 7573 32997 7607 33031
rect 9321 32997 9355 33031
rect 5825 32929 5859 32963
rect 7849 32929 7883 32963
rect 7987 32929 8021 32963
rect 1409 32861 1443 32895
rect 1685 32861 1719 32895
rect 1961 32861 1995 32895
rect 6101 32861 6135 32895
rect 6929 32861 6963 32895
rect 7113 32861 7147 32895
rect 8125 32861 8159 32895
rect 9045 32861 9079 32895
rect 9137 32861 9171 32895
rect 9505 32861 9539 32895
rect 8769 32725 8803 32759
rect 8953 32725 8987 32759
rect 9689 32725 9723 32759
rect 6193 32521 6227 32555
rect 8677 32521 8711 32555
rect 1501 32385 1535 32419
rect 3433 32385 3467 32419
rect 4905 32385 4939 32419
rect 5457 32385 5491 32419
rect 6561 32385 6595 32419
rect 7113 32385 7147 32419
rect 8217 32385 8251 32419
rect 8493 32385 8527 32419
rect 8769 32385 8803 32419
rect 9137 32385 9171 32419
rect 9505 32385 9539 32419
rect 5181 32317 5215 32351
rect 6837 32317 6871 32351
rect 7849 32249 7883 32283
rect 8953 32249 8987 32283
rect 1593 32181 1627 32215
rect 3617 32181 3651 32215
rect 5089 32181 5123 32215
rect 6745 32181 6779 32215
rect 8401 32181 8435 32215
rect 9321 32181 9355 32215
rect 9689 32181 9723 32215
rect 1777 31977 1811 32011
rect 4353 31977 4387 32011
rect 5549 31909 5583 31943
rect 9321 31909 9355 31943
rect 9689 31909 9723 31943
rect 1685 31841 1719 31875
rect 2559 31841 2593 31875
rect 2697 31841 2731 31875
rect 2973 31841 3007 31875
rect 4997 31841 5031 31875
rect 7297 31841 7331 31875
rect 1501 31773 1535 31807
rect 2421 31773 2455 31807
rect 3433 31773 3467 31807
rect 3617 31773 3651 31807
rect 5135 31773 5169 31807
rect 5273 31773 5307 31807
rect 6009 31773 6043 31807
rect 6193 31773 6227 31807
rect 7573 31773 7607 31807
rect 8585 31773 8619 31807
rect 9137 31773 9171 31807
rect 9505 31773 9539 31807
rect 8309 31637 8343 31671
rect 8769 31637 8803 31671
rect 2513 31433 2547 31467
rect 3525 31433 3559 31467
rect 3709 31433 3743 31467
rect 9505 31433 9539 31467
rect 1501 31297 1535 31331
rect 1777 31297 1811 31331
rect 3341 31297 3375 31331
rect 4512 31297 4546 31331
rect 5641 31297 5675 31331
rect 7849 31297 7883 31331
rect 8585 31297 8619 31331
rect 8861 31297 8895 31331
rect 9781 31297 9815 31331
rect 4353 31229 4387 31263
rect 4629 31229 4663 31263
rect 5365 31229 5399 31263
rect 5549 31229 5583 31263
rect 7665 31229 7699 31263
rect 8309 31229 8343 31263
rect 8702 31229 8736 31263
rect 4905 31161 4939 31195
rect 5825 31093 5859 31127
rect 9597 31093 9631 31127
rect 2513 30889 2547 30923
rect 3617 30889 3651 30923
rect 3985 30889 4019 30923
rect 7665 30889 7699 30923
rect 9321 30889 9355 30923
rect 8217 30821 8251 30855
rect 6285 30753 6319 30787
rect 1501 30685 1535 30719
rect 1777 30685 1811 30719
rect 2605 30685 2639 30719
rect 2881 30685 2915 30719
rect 3801 30685 3835 30719
rect 6561 30685 6595 30719
rect 7481 30685 7515 30719
rect 8401 30685 8435 30719
rect 8493 30685 8527 30719
rect 9137 30685 9171 30719
rect 9505 30685 9539 30719
rect 7297 30549 7331 30583
rect 8677 30549 8711 30583
rect 9689 30549 9723 30583
rect 1685 30277 1719 30311
rect 9045 30277 9079 30311
rect 1501 30209 1535 30243
rect 3157 30209 3191 30243
rect 6377 30209 6411 30243
rect 7389 30209 7423 30243
rect 8125 30209 8159 30243
rect 8401 30209 8435 30243
rect 9137 30209 9171 30243
rect 9505 30209 9539 30243
rect 2881 30141 2915 30175
rect 7205 30141 7239 30175
rect 8263 30141 8297 30175
rect 3893 30073 3927 30107
rect 7849 30073 7883 30107
rect 9321 30073 9355 30107
rect 1593 30005 1627 30039
rect 6561 30005 6595 30039
rect 9689 30005 9723 30039
rect 1593 29801 1627 29835
rect 6469 29801 6503 29835
rect 7573 29801 7607 29835
rect 8953 29801 8987 29835
rect 1777 29733 1811 29767
rect 8033 29733 8067 29767
rect 8309 29733 8343 29767
rect 5273 29665 5307 29699
rect 5825 29665 5859 29699
rect 6561 29665 6595 29699
rect 9413 29665 9447 29699
rect 9505 29665 9539 29699
rect 1409 29597 1443 29631
rect 1961 29597 1995 29631
rect 4629 29597 4663 29631
rect 4813 29597 4847 29631
rect 5549 29597 5583 29631
rect 5666 29597 5700 29631
rect 6837 29597 6871 29631
rect 7849 29597 7883 29631
rect 8125 29597 8159 29631
rect 8493 29597 8527 29631
rect 8677 29461 8711 29495
rect 9321 29461 9355 29495
rect 1593 29257 1627 29291
rect 5181 29257 5215 29291
rect 1409 29121 1443 29155
rect 2053 29121 2087 29155
rect 4445 29121 4479 29155
rect 7389 29121 7423 29155
rect 8125 29121 8159 29155
rect 9137 29121 9171 29155
rect 9505 29121 9539 29155
rect 1777 29053 1811 29087
rect 4169 29053 4203 29087
rect 7205 29053 7239 29087
rect 8242 29053 8276 29087
rect 8401 29053 8435 29087
rect 7849 28985 7883 29019
rect 9321 28985 9355 29019
rect 9689 28985 9723 29019
rect 2789 28917 2823 28951
rect 9045 28917 9079 28951
rect 1593 28713 1627 28747
rect 3617 28713 3651 28747
rect 4997 28713 5031 28747
rect 7481 28713 7515 28747
rect 9321 28645 9355 28679
rect 6469 28577 6503 28611
rect 1501 28509 1535 28543
rect 1777 28509 1811 28543
rect 2053 28509 2087 28543
rect 3433 28509 3467 28543
rect 3985 28509 4019 28543
rect 4261 28509 4295 28543
rect 5549 28509 5583 28543
rect 6745 28509 6779 28543
rect 8585 28509 8619 28543
rect 9137 28509 9171 28543
rect 9505 28509 9539 28543
rect 5733 28441 5767 28475
rect 2789 28373 2823 28407
rect 5365 28373 5399 28407
rect 5825 28373 5859 28407
rect 8769 28373 8803 28407
rect 9689 28373 9723 28407
rect 2421 28169 2455 28203
rect 7481 28169 7515 28203
rect 8125 28169 8159 28203
rect 9413 28169 9447 28203
rect 1409 28033 1443 28067
rect 5733 28033 5767 28067
rect 6009 28033 6043 28067
rect 6469 28033 6503 28067
rect 6745 28033 6779 28067
rect 8309 28033 8343 28067
rect 8401 28033 8435 28067
rect 8677 28033 8711 28067
rect 9505 28033 9539 28067
rect 3065 27965 3099 27999
rect 3224 27965 3258 27999
rect 3341 27965 3375 27999
rect 4077 27965 4111 27999
rect 4261 27965 4295 27999
rect 3617 27897 3651 27931
rect 1593 27829 1627 27863
rect 4997 27829 5031 27863
rect 9689 27829 9723 27863
rect 4445 27625 4479 27659
rect 8769 27557 8803 27591
rect 9321 27557 9355 27591
rect 2329 27421 2363 27455
rect 2605 27421 2639 27455
rect 4261 27421 4295 27455
rect 4537 27421 4571 27455
rect 4813 27421 4847 27455
rect 8309 27421 8343 27455
rect 8585 27421 8619 27455
rect 9137 27421 9171 27455
rect 9505 27421 9539 27455
rect 8125 27353 8159 27387
rect 1593 27285 1627 27319
rect 5549 27285 5583 27319
rect 9689 27285 9723 27319
rect 2973 27081 3007 27115
rect 9321 27081 9355 27115
rect 1409 26945 1443 26979
rect 2145 26945 2179 26979
rect 4813 26945 4847 26979
rect 5181 26945 5215 26979
rect 6745 26945 6779 26979
rect 8493 26945 8527 26979
rect 8769 26945 8803 26979
rect 9137 26945 9171 26979
rect 9505 26945 9539 26979
rect 1869 26877 1903 26911
rect 3617 26877 3651 26911
rect 3776 26877 3810 26911
rect 3893 26877 3927 26911
rect 4629 26877 4663 26911
rect 4905 26877 4939 26911
rect 2881 26809 2915 26843
rect 4169 26809 4203 26843
rect 8677 26809 8711 26843
rect 8953 26809 8987 26843
rect 1593 26741 1627 26775
rect 5917 26741 5951 26775
rect 6929 26741 6963 26775
rect 9689 26741 9723 26775
rect 1593 26537 1627 26571
rect 3249 26537 3283 26571
rect 4629 26537 4663 26571
rect 6929 26537 6963 26571
rect 9689 26537 9723 26571
rect 5733 26469 5767 26503
rect 8217 26469 8251 26503
rect 9321 26469 9355 26503
rect 5089 26401 5123 26435
rect 6285 26401 6319 26435
rect 1409 26333 1443 26367
rect 1777 26333 1811 26367
rect 2237 26333 2271 26367
rect 2513 26333 2547 26367
rect 4997 26333 5031 26367
rect 5273 26333 5307 26367
rect 6009 26333 6043 26367
rect 6147 26333 6181 26367
rect 7205 26333 7239 26367
rect 7481 26333 7515 26367
rect 9137 26333 9171 26367
rect 9505 26333 9539 26367
rect 4537 26265 4571 26299
rect 1961 26197 1995 26231
rect 4813 26197 4847 26231
rect 2329 25857 2363 25891
rect 2605 25857 2639 25891
rect 3249 25857 3283 25891
rect 6561 25857 6595 25891
rect 6837 25857 6871 25891
rect 7849 25857 7883 25891
rect 3525 25789 3559 25823
rect 8033 25789 8067 25823
rect 8493 25789 8527 25823
rect 8769 25789 8803 25823
rect 8907 25789 8941 25823
rect 9045 25789 9079 25823
rect 1593 25653 1627 25687
rect 7573 25653 7607 25687
rect 9689 25653 9723 25687
rect 1961 25449 1995 25483
rect 8493 25449 8527 25483
rect 9321 25381 9355 25415
rect 6377 25313 6411 25347
rect 7481 25313 7515 25347
rect 1409 25245 1443 25279
rect 1777 25245 1811 25279
rect 4813 25245 4847 25279
rect 5089 25245 5123 25279
rect 6653 25245 6687 25279
rect 7757 25245 7791 25279
rect 8585 25245 8619 25279
rect 9137 25245 9171 25279
rect 9505 25245 9539 25279
rect 1593 25109 1627 25143
rect 5825 25109 5859 25143
rect 7389 25109 7423 25143
rect 8769 25109 8803 25143
rect 9689 25109 9723 25143
rect 5641 24905 5675 24939
rect 9229 24837 9263 24871
rect 1409 24769 1443 24803
rect 2697 24769 2731 24803
rect 5457 24769 5491 24803
rect 7389 24769 7423 24803
rect 8125 24769 8159 24803
rect 8242 24769 8276 24803
rect 9505 24769 9539 24803
rect 2421 24701 2455 24735
rect 3525 24701 3559 24735
rect 3709 24701 3743 24735
rect 4445 24701 4479 24735
rect 4583 24701 4617 24735
rect 4721 24701 4755 24735
rect 7205 24701 7239 24735
rect 8401 24701 8435 24735
rect 1593 24633 1627 24667
rect 4169 24633 4203 24667
rect 7849 24633 7883 24667
rect 3433 24565 3467 24599
rect 5365 24565 5399 24599
rect 9045 24565 9079 24599
rect 9689 24565 9723 24599
rect 1593 24361 1627 24395
rect 5181 24361 5215 24395
rect 8125 24361 8159 24395
rect 9689 24361 9723 24395
rect 6377 24293 6411 24327
rect 9321 24293 9355 24327
rect 2421 24225 2455 24259
rect 5963 24225 5997 24259
rect 1409 24157 1443 24191
rect 2697 24157 2731 24191
rect 5825 24157 5859 24191
rect 6101 24157 6135 24191
rect 6837 24157 6871 24191
rect 7021 24157 7055 24191
rect 7113 24157 7147 24191
rect 7389 24157 7423 24191
rect 8585 24157 8619 24191
rect 9137 24157 9171 24191
rect 9505 24157 9539 24191
rect 3433 24021 3467 24055
rect 8769 24021 8803 24055
rect 3065 23817 3099 23851
rect 5089 23817 5123 23851
rect 8309 23817 8343 23851
rect 9689 23817 9723 23851
rect 2329 23681 2363 23715
rect 3433 23681 3467 23715
rect 4169 23681 4203 23715
rect 4445 23681 4479 23715
rect 5181 23681 5215 23715
rect 7573 23681 7607 23715
rect 8401 23681 8435 23715
rect 9137 23681 9171 23715
rect 9505 23681 9539 23715
rect 2053 23613 2087 23647
rect 3249 23613 3283 23647
rect 3893 23613 3927 23647
rect 4307 23613 4341 23647
rect 7297 23613 7331 23647
rect 8585 23545 8619 23579
rect 5365 23477 5399 23511
rect 9321 23477 9355 23511
rect 1593 23273 1627 23307
rect 2973 23273 3007 23307
rect 1869 23205 1903 23239
rect 9689 23205 9723 23239
rect 6745 23137 6779 23171
rect 7757 23137 7791 23171
rect 1409 23069 1443 23103
rect 1685 23069 1719 23103
rect 1961 23069 1995 23103
rect 2237 23069 2271 23103
rect 8033 23069 8067 23103
rect 9137 23069 9171 23103
rect 9505 23069 9539 23103
rect 6561 23001 6595 23035
rect 6193 22933 6227 22967
rect 6653 22933 6687 22967
rect 8769 22933 8803 22967
rect 9321 22933 9355 22967
rect 1593 22729 1627 22763
rect 6377 22729 6411 22763
rect 9045 22729 9079 22763
rect 9505 22729 9539 22763
rect 9137 22661 9171 22695
rect 1409 22593 1443 22627
rect 1685 22593 1719 22627
rect 1961 22593 1995 22627
rect 4261 22593 4295 22627
rect 4537 22593 4571 22627
rect 6009 22593 6043 22627
rect 7113 22593 7147 22627
rect 8401 22593 8435 22627
rect 9781 22593 9815 22627
rect 7389 22525 7423 22559
rect 8861 22525 8895 22559
rect 8585 22457 8619 22491
rect 2697 22389 2731 22423
rect 5273 22389 5307 22423
rect 6193 22389 6227 22423
rect 9597 22389 9631 22423
rect 8401 22185 8435 22219
rect 5273 22117 5307 22151
rect 1777 22049 1811 22083
rect 5549 22049 5583 22083
rect 5666 22049 5700 22083
rect 2053 21981 2087 22015
rect 4629 21981 4663 22015
rect 4813 21981 4847 22015
rect 5825 21981 5859 22015
rect 6469 21981 6503 22015
rect 6561 21981 6595 22015
rect 8217 21981 8251 22015
rect 8493 21981 8527 22015
rect 9137 21981 9171 22015
rect 9505 21981 9539 22015
rect 2789 21845 2823 21879
rect 6745 21845 6779 21879
rect 8677 21845 8711 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 2421 21641 2455 21675
rect 5457 21641 5491 21675
rect 9321 21641 9355 21675
rect 9689 21641 9723 21675
rect 1409 21505 1443 21539
rect 1685 21505 1719 21539
rect 4353 21505 4387 21539
rect 4445 21505 4479 21539
rect 4721 21505 4755 21539
rect 9505 21505 9539 21539
rect 3157 21437 3191 21471
rect 3316 21437 3350 21471
rect 3433 21437 3467 21471
rect 3709 21437 3743 21471
rect 4169 21437 4203 21471
rect 7481 21437 7515 21471
rect 7665 21437 7699 21471
rect 8401 21437 8435 21471
rect 8518 21437 8552 21471
rect 8677 21437 8711 21471
rect 8125 21369 8159 21403
rect 2513 21301 2547 21335
rect 3249 21097 3283 21131
rect 4261 21097 4295 21131
rect 5089 21097 5123 21131
rect 9689 21097 9723 21131
rect 9321 21029 9355 21063
rect 2237 20961 2271 20995
rect 7573 20961 7607 20995
rect 7966 20961 8000 20995
rect 1409 20893 1443 20927
rect 1685 20893 1719 20927
rect 2513 20893 2547 20927
rect 4077 20893 4111 20927
rect 4905 20893 4939 20927
rect 6929 20893 6963 20927
rect 7113 20893 7147 20927
rect 7849 20893 7883 20927
rect 8125 20893 8159 20927
rect 9137 20893 9171 20927
rect 9505 20893 9539 20927
rect 1593 20757 1627 20791
rect 1869 20757 1903 20791
rect 8769 20757 8803 20791
rect 7665 20553 7699 20587
rect 8677 20553 8711 20587
rect 9689 20553 9723 20587
rect 2145 20417 2179 20451
rect 6929 20417 6963 20451
rect 8493 20417 8527 20451
rect 8769 20417 8803 20451
rect 9137 20417 9171 20451
rect 9505 20417 9539 20451
rect 6653 20349 6687 20383
rect 9321 20281 9355 20315
rect 1961 20213 1995 20247
rect 8953 20213 8987 20247
rect 4537 20009 4571 20043
rect 7389 20009 7423 20043
rect 8769 20009 8803 20043
rect 9689 20009 9723 20043
rect 9321 19941 9355 19975
rect 1777 19873 1811 19907
rect 6377 19873 6411 19907
rect 1409 19805 1443 19839
rect 2053 19805 2087 19839
rect 4353 19805 4387 19839
rect 6653 19805 6687 19839
rect 7481 19805 7515 19839
rect 7757 19805 7791 19839
rect 8585 19805 8619 19839
rect 9137 19805 9171 19839
rect 9505 19805 9539 19839
rect 1593 19669 1627 19703
rect 2789 19669 2823 19703
rect 8493 19669 8527 19703
rect 2881 19465 2915 19499
rect 4997 19465 5031 19499
rect 9413 19465 9447 19499
rect 9689 19465 9723 19499
rect 1409 19329 1443 19363
rect 2053 19329 2087 19363
rect 3663 19329 3697 19363
rect 4813 19329 4847 19363
rect 6377 19329 6411 19363
rect 6653 19329 6687 19363
rect 7573 19329 7607 19363
rect 8493 19329 8527 19363
rect 9505 19329 9539 19363
rect 1777 19261 1811 19295
rect 3525 19261 3559 19295
rect 3801 19261 3835 19295
rect 4077 19261 4111 19295
rect 4537 19261 4571 19295
rect 4721 19261 4755 19295
rect 7757 19261 7791 19295
rect 8610 19261 8644 19295
rect 8769 19261 8803 19295
rect 2789 19193 2823 19227
rect 7389 19193 7423 19227
rect 8217 19193 8251 19227
rect 1593 19125 1627 19159
rect 3801 18921 3835 18955
rect 5917 18921 5951 18955
rect 8217 18921 8251 18955
rect 9689 18921 9723 18955
rect 2973 18853 3007 18887
rect 9229 18853 9263 18887
rect 1961 18785 1995 18819
rect 4583 18785 4617 18819
rect 4721 18785 4755 18819
rect 4997 18785 5031 18819
rect 5641 18785 5675 18819
rect 2237 18717 2271 18751
rect 4445 18717 4479 18751
rect 5457 18717 5491 18751
rect 5733 18717 5767 18751
rect 6929 18717 6963 18751
rect 7205 18717 7239 18751
rect 8401 18717 8435 18751
rect 8499 18717 8533 18751
rect 9413 18717 9447 18751
rect 9505 18717 9539 18751
rect 7941 18581 7975 18615
rect 8677 18581 8711 18615
rect 4721 18377 4755 18411
rect 9689 18377 9723 18411
rect 3433 18309 3467 18343
rect 1409 18241 1443 18275
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 2329 18241 2363 18275
rect 5365 18241 5399 18275
rect 6377 18241 6411 18275
rect 6653 18241 6687 18275
rect 8769 18241 8803 18275
rect 9505 18241 9539 18275
rect 7573 18173 7607 18207
rect 7757 18173 7791 18207
rect 8217 18173 8251 18207
rect 8493 18173 8527 18207
rect 8610 18173 8644 18207
rect 1869 18105 1903 18139
rect 3065 18105 3099 18139
rect 5549 18105 5583 18139
rect 1593 18037 1627 18071
rect 7389 18037 7423 18071
rect 9413 18037 9447 18071
rect 2513 17833 2547 17867
rect 6285 17833 6319 17867
rect 6745 17833 6779 17867
rect 7021 17833 7055 17867
rect 8493 17833 8527 17867
rect 8125 17765 8159 17799
rect 1685 17697 1719 17731
rect 7113 17697 7147 17731
rect 9505 17697 9539 17731
rect 9781 17697 9815 17731
rect 1409 17629 1443 17663
rect 2329 17629 2363 17663
rect 6101 17629 6135 17663
rect 6561 17629 6595 17663
rect 6837 17629 6871 17663
rect 7389 17629 7423 17663
rect 8309 17629 8343 17663
rect 8585 17629 8619 17663
rect 2513 17493 2547 17527
rect 8769 17493 8803 17527
rect 9413 17289 9447 17323
rect 9505 17221 9539 17255
rect 1409 17153 1443 17187
rect 1685 17153 1719 17187
rect 2697 17153 2731 17187
rect 3433 17153 3467 17187
rect 4353 17153 4387 17187
rect 4445 17153 4479 17187
rect 7757 17153 7791 17187
rect 8769 17153 8803 17187
rect 9689 17153 9723 17187
rect 2513 17085 2547 17119
rect 3571 17085 3605 17119
rect 3709 17085 3743 17119
rect 7573 17085 7607 17119
rect 8217 17085 8251 17119
rect 8493 17085 8527 17119
rect 8610 17085 8644 17119
rect 3157 17017 3191 17051
rect 4629 17017 4663 17051
rect 2421 16949 2455 16983
rect 2789 16745 2823 16779
rect 8217 16745 8251 16779
rect 9551 16745 9585 16779
rect 8493 16677 8527 16711
rect 1777 16609 1811 16643
rect 5549 16609 5583 16643
rect 9781 16609 9815 16643
rect 2053 16541 2087 16575
rect 5273 16541 5307 16575
rect 6745 16541 6779 16575
rect 7021 16541 7055 16575
rect 8309 16541 8343 16575
rect 8677 16473 8711 16507
rect 4537 16405 4571 16439
rect 7757 16405 7791 16439
rect 9597 16201 9631 16235
rect 9689 16133 9723 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 2421 16065 2455 16099
rect 3617 16065 3651 16099
rect 5273 16065 5307 16099
rect 5549 16065 5583 16099
rect 6653 16065 6687 16099
rect 7573 16065 7607 16099
rect 8631 16065 8665 16099
rect 2605 15997 2639 16031
rect 3341 15997 3375 16031
rect 3479 15997 3513 16031
rect 4353 15997 4387 16031
rect 4537 15997 4571 16031
rect 4997 15997 5031 16031
rect 5411 15997 5445 16031
rect 6377 15997 6411 16031
rect 7757 15997 7791 16031
rect 8217 15997 8251 16031
rect 8493 15997 8527 16031
rect 8769 15997 8803 16031
rect 3065 15929 3099 15963
rect 4261 15861 4295 15895
rect 6193 15861 6227 15895
rect 7389 15861 7423 15895
rect 9413 15861 9447 15895
rect 3065 15657 3099 15691
rect 4537 15657 4571 15691
rect 6009 15657 6043 15691
rect 7389 15657 7423 15691
rect 7849 15657 7883 15691
rect 5641 15589 5675 15623
rect 2053 15521 2087 15555
rect 4629 15521 4663 15555
rect 8493 15521 8527 15555
rect 9781 15521 9815 15555
rect 2329 15453 2363 15487
rect 4353 15453 4387 15487
rect 4905 15453 4939 15487
rect 5825 15453 5859 15487
rect 7573 15453 7607 15487
rect 7665 15453 7699 15487
rect 8769 15453 8803 15487
rect 9505 15453 9539 15487
rect 2973 15113 3007 15147
rect 7573 15113 7607 15147
rect 9689 15045 9723 15079
rect 1685 14977 1719 15011
rect 1961 14977 1995 15011
rect 2237 14977 2271 15011
rect 6745 14977 6779 15011
rect 8376 14977 8410 15011
rect 9413 14977 9447 15011
rect 6469 14909 6503 14943
rect 8217 14909 8251 14943
rect 8493 14909 8527 14943
rect 9229 14909 9263 14943
rect 8769 14841 8803 14875
rect 9505 14841 9539 14875
rect 1501 14773 1535 14807
rect 7481 14773 7515 14807
rect 4445 14569 4479 14603
rect 9321 14569 9355 14603
rect 9597 14569 9631 14603
rect 7553 14501 7587 14535
rect 1869 14433 1903 14467
rect 7113 14433 7147 14467
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 4261 14365 4295 14399
rect 4629 14365 4663 14399
rect 4905 14365 4939 14399
rect 6469 14365 6503 14399
rect 6745 14365 6779 14399
rect 6929 14365 6963 14399
rect 7849 14365 7883 14399
rect 7987 14365 8021 14399
rect 8125 14365 8159 14399
rect 9137 14365 9171 14399
rect 9689 14365 9723 14399
rect 1501 14229 1535 14263
rect 2881 14229 2915 14263
rect 5641 14229 5675 14263
rect 5733 14229 5767 14263
rect 8769 14229 8803 14263
rect 2789 14025 2823 14059
rect 4721 14025 4755 14059
rect 9597 14025 9631 14059
rect 1777 13889 1811 13923
rect 2053 13889 2087 13923
rect 3801 13889 3835 13923
rect 4077 13889 4111 13923
rect 5089 13889 5123 13923
rect 5365 13889 5399 13923
rect 7665 13889 7699 13923
rect 8401 13889 8435 13923
rect 9781 13889 9815 13923
rect 2881 13821 2915 13855
rect 3065 13821 3099 13855
rect 3525 13821 3559 13855
rect 3939 13821 3973 13855
rect 7481 13821 7515 13855
rect 8518 13821 8552 13855
rect 8677 13821 8711 13855
rect 8125 13753 8159 13787
rect 6101 13685 6135 13719
rect 9321 13685 9355 13719
rect 7757 13481 7791 13515
rect 1961 13413 1995 13447
rect 6791 13413 6825 13447
rect 8033 13413 8067 13447
rect 8309 13413 8343 13447
rect 9505 13345 9539 13379
rect 1685 13277 1719 13311
rect 1777 13277 1811 13311
rect 6720 13277 6754 13311
rect 7941 13277 7975 13311
rect 8217 13277 8251 13311
rect 8493 13277 8527 13311
rect 8769 13277 8803 13311
rect 9321 13277 9355 13311
rect 1501 13141 1535 13175
rect 8585 13141 8619 13175
rect 8953 13141 8987 13175
rect 9413 13141 9447 13175
rect 4905 12937 4939 12971
rect 9229 12937 9263 12971
rect 6929 12869 6963 12903
rect 7113 12869 7147 12903
rect 1961 12801 1995 12835
rect 2789 12801 2823 12835
rect 3709 12801 3743 12835
rect 4629 12801 4663 12835
rect 4721 12801 4755 12835
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 8309 12801 8343 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 1685 12733 1719 12767
rect 2973 12733 3007 12767
rect 3847 12733 3881 12767
rect 3985 12733 4019 12767
rect 7573 12733 7607 12767
rect 8426 12733 8460 12767
rect 8585 12733 8619 12767
rect 2697 12665 2731 12699
rect 3433 12665 3467 12699
rect 6377 12665 6411 12699
rect 8033 12665 8067 12699
rect 9321 12665 9355 12699
rect 6745 12597 6779 12631
rect 9597 12597 9631 12631
rect 1409 12393 1443 12427
rect 2697 12393 2731 12427
rect 6837 12393 6871 12427
rect 8033 12393 8067 12427
rect 2789 12325 2823 12359
rect 8309 12325 8343 12359
rect 8585 12325 8619 12359
rect 1685 12257 1719 12291
rect 4997 12257 5031 12291
rect 5641 12257 5675 12291
rect 5917 12257 5951 12291
rect 6193 12257 6227 12291
rect 1961 12189 1995 12223
rect 3893 12189 3927 12223
rect 4169 12189 4203 12223
rect 5181 12189 5215 12223
rect 6034 12189 6068 12223
rect 7113 12189 7147 12223
rect 7481 12189 7515 12223
rect 8217 12189 8251 12223
rect 8493 12189 8527 12223
rect 8769 12189 8803 12223
rect 9505 12189 9539 12223
rect 9781 12189 9815 12223
rect 2973 12121 3007 12155
rect 7205 12121 7239 12155
rect 7297 12121 7331 12155
rect 4905 12053 4939 12087
rect 6929 12053 6963 12087
rect 5181 11849 5215 11883
rect 6561 11849 6595 11883
rect 1685 11713 1719 11747
rect 2237 11713 2271 11747
rect 3985 11713 4019 11747
rect 4102 11713 4136 11747
rect 4905 11713 4939 11747
rect 4997 11713 5031 11747
rect 6469 11713 6503 11747
rect 7757 11713 7791 11747
rect 9689 11713 9723 11747
rect 1961 11645 1995 11679
rect 3065 11645 3099 11679
rect 3249 11645 3283 11679
rect 4261 11645 4295 11679
rect 7573 11645 7607 11679
rect 8493 11645 8527 11679
rect 8610 11645 8644 11679
rect 8769 11645 8803 11679
rect 9505 11645 9539 11679
rect 3709 11577 3743 11611
rect 8217 11577 8251 11611
rect 1501 11509 1535 11543
rect 2973 11509 3007 11543
rect 9413 11509 9447 11543
rect 2881 11305 2915 11339
rect 7297 11305 7331 11339
rect 8033 11305 8067 11339
rect 8493 11305 8527 11339
rect 8585 11305 8619 11339
rect 1501 11237 1535 11271
rect 6101 11237 6135 11271
rect 7757 11237 7791 11271
rect 9689 11237 9723 11271
rect 1869 11169 1903 11203
rect 6377 11169 6411 11203
rect 6653 11169 6687 11203
rect 9137 11169 9171 11203
rect 9229 11169 9263 11203
rect 1685 11101 1719 11135
rect 2145 11101 2179 11135
rect 5457 11101 5491 11135
rect 5641 11101 5675 11135
rect 6494 11101 6528 11135
rect 7941 11101 7975 11135
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 8769 11101 8803 11135
rect 9321 10965 9355 10999
rect 1501 10761 1535 10795
rect 3065 10761 3099 10795
rect 7573 10761 7607 10795
rect 9505 10761 9539 10795
rect 3801 10693 3835 10727
rect 1777 10625 1811 10659
rect 2329 10625 2363 10659
rect 3617 10625 3651 10659
rect 5365 10625 5399 10659
rect 6837 10625 6871 10659
rect 7665 10625 7699 10659
rect 8702 10625 8736 10659
rect 9781 10625 9815 10659
rect 2053 10557 2087 10591
rect 5089 10557 5123 10591
rect 6561 10557 6595 10591
rect 7849 10557 7883 10591
rect 8585 10557 8619 10591
rect 8861 10557 8895 10591
rect 1961 10489 1995 10523
rect 5181 10489 5215 10523
rect 8309 10489 8343 10523
rect 9597 10489 9631 10523
rect 3709 10421 3743 10455
rect 5273 10421 5307 10455
rect 1961 10217 1995 10251
rect 7849 10217 7883 10251
rect 4813 10149 4847 10183
rect 8493 10149 8527 10183
rect 2605 10081 2639 10115
rect 5181 10081 5215 10115
rect 6469 10081 6503 10115
rect 6837 10081 6871 10115
rect 9781 10081 9815 10115
rect 1685 10013 1719 10047
rect 1869 10013 1903 10047
rect 2881 10013 2915 10047
rect 3801 10013 3835 10047
rect 4077 10013 4111 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 7113 10013 7147 10047
rect 8401 10013 8435 10047
rect 9505 10013 9539 10047
rect 5089 9945 5123 9979
rect 5549 9945 5583 9979
rect 6285 9945 6319 9979
rect 8677 9945 8711 9979
rect 1501 9877 1535 9911
rect 3617 9877 3651 9911
rect 5917 9877 5951 9911
rect 6377 9877 6411 9911
rect 8217 9877 8251 9911
rect 8585 9877 8619 9911
rect 4721 9673 4755 9707
rect 5365 9673 5399 9707
rect 8309 9673 8343 9707
rect 4537 9605 4571 9639
rect 5871 9605 5905 9639
rect 1685 9537 1719 9571
rect 2697 9537 2731 9571
rect 2973 9537 3007 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5227 9537 5261 9571
rect 5457 9537 5491 9571
rect 5549 9537 5583 9571
rect 5733 9537 5767 9571
rect 5974 9536 6008 9570
rect 6561 9537 6595 9571
rect 6929 9537 6963 9571
rect 7573 9537 7607 9571
rect 8585 9537 8619 9571
rect 7297 9469 7331 9503
rect 9505 9469 9539 9503
rect 9781 9469 9815 9503
rect 3709 9401 3743 9435
rect 4169 9401 4203 9435
rect 5641 9401 5675 9435
rect 1501 9333 1535 9367
rect 4537 9333 4571 9367
rect 4813 9333 4847 9367
rect 6377 9333 6411 9367
rect 6561 9333 6595 9367
rect 8677 9333 8711 9367
rect 8309 9061 8343 9095
rect 9505 9061 9539 9095
rect 1685 8925 1719 8959
rect 7849 8925 7883 8959
rect 7976 8925 8010 8959
rect 8079 8925 8113 8959
rect 8217 8925 8251 8959
rect 8493 8925 8527 8959
rect 9137 8925 9171 8959
rect 8953 8857 8987 8891
rect 9689 8857 9723 8891
rect 1501 8789 1535 8823
rect 7665 8789 7699 8823
rect 8677 8789 8711 8823
rect 9321 8789 9355 8823
rect 1961 8585 1995 8619
rect 8953 8585 8987 8619
rect 1501 8517 1535 8551
rect 1869 8517 1903 8551
rect 9505 8517 9539 8551
rect 2605 8449 2639 8483
rect 7297 8449 7331 8483
rect 9413 8449 9447 8483
rect 1685 8381 1719 8415
rect 2329 8381 2363 8415
rect 7113 8381 7147 8415
rect 8033 8381 8067 8415
rect 8171 8381 8205 8415
rect 8309 8381 8343 8415
rect 9597 8381 9631 8415
rect 3341 8313 3375 8347
rect 7757 8313 7791 8347
rect 9045 8245 9079 8279
rect 2513 8041 2547 8075
rect 6929 8041 6963 8075
rect 8585 8041 8619 8075
rect 8953 8041 8987 8075
rect 5733 7973 5767 8007
rect 7757 7973 7791 8007
rect 2605 7905 2639 7939
rect 5089 7905 5123 7939
rect 6009 7905 6043 7939
rect 6126 7905 6160 7939
rect 1501 7837 1535 7871
rect 1777 7837 1811 7871
rect 2881 7837 2915 7871
rect 5273 7837 5307 7871
rect 6285 7837 6319 7871
rect 7941 7837 7975 7871
rect 8309 7837 8343 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9505 7837 9539 7871
rect 9781 7837 9815 7871
rect 8125 7769 8159 7803
rect 8677 7769 8711 7803
rect 3617 7701 3651 7735
rect 9597 7701 9631 7735
rect 1501 7497 1535 7531
rect 2053 7497 2087 7531
rect 2421 7497 2455 7531
rect 3709 7497 3743 7531
rect 6929 7497 6963 7531
rect 7113 7497 7147 7531
rect 7757 7497 7791 7531
rect 2329 7429 2363 7463
rect 7481 7429 7515 7463
rect 8493 7429 8527 7463
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 2973 7361 3007 7395
rect 4169 7361 4203 7395
rect 6469 7361 6503 7395
rect 6745 7361 6779 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 7941 7361 7975 7395
rect 8125 7361 8159 7395
rect 8401 7361 8435 7395
rect 8861 7361 8895 7395
rect 9137 7361 9171 7395
rect 9505 7361 9539 7395
rect 9781 7361 9815 7395
rect 2697 7293 2731 7327
rect 4353 7293 4387 7327
rect 4813 7293 4847 7327
rect 5089 7293 5123 7327
rect 5227 7293 5261 7327
rect 5365 7293 5399 7327
rect 6009 7293 6043 7327
rect 9225 7293 9259 7327
rect 6653 7225 6687 7259
rect 8217 7225 8251 7259
rect 9413 7225 9447 7259
rect 9597 7225 9631 7259
rect 8033 7157 8067 7191
rect 8585 7157 8619 7191
rect 9045 7157 9079 7191
rect 9321 7157 9355 7191
rect 6837 6953 6871 6987
rect 7849 6953 7883 6987
rect 7481 6885 7515 6919
rect 8033 6885 8067 6919
rect 4997 6817 5031 6851
rect 5181 6817 5215 6851
rect 5641 6817 5675 6851
rect 5917 6817 5951 6851
rect 6034 6817 6068 6851
rect 6193 6817 6227 6851
rect 8309 6817 8343 6851
rect 8677 6817 8711 6851
rect 9505 6817 9539 6851
rect 2145 6749 2179 6783
rect 2421 6749 2455 6783
rect 7389 6749 7423 6783
rect 8125 6749 8159 6783
rect 8401 6749 8435 6783
rect 8769 6749 8803 6783
rect 9781 6749 9815 6783
rect 1409 6613 1443 6647
rect 7205 6613 7239 6647
rect 7849 6613 7883 6647
rect 8585 6613 8619 6647
rect 1593 6409 1627 6443
rect 2145 6409 2179 6443
rect 7389 6409 7423 6443
rect 8585 6409 8619 6443
rect 1409 6273 1443 6307
rect 2053 6273 2087 6307
rect 2881 6273 2915 6307
rect 4353 6273 4387 6307
rect 6377 6273 6411 6307
rect 6653 6273 6687 6307
rect 7849 6273 7883 6307
rect 8826 6273 8860 6307
rect 3157 6205 3191 6239
rect 4077 6205 4111 6239
rect 7573 6205 7607 6239
rect 9505 6205 9539 6239
rect 9781 6205 9815 6239
rect 8723 6137 8757 6171
rect 1869 6069 1903 6103
rect 5089 6069 5123 6103
rect 7573 5865 7607 5899
rect 8677 5865 8711 5899
rect 3617 5797 3651 5831
rect 5733 5797 5767 5831
rect 6469 5797 6503 5831
rect 2605 5729 2639 5763
rect 4353 5729 4387 5763
rect 6561 5729 6595 5763
rect 7665 5729 7699 5763
rect 9505 5729 9539 5763
rect 2881 5661 2915 5695
rect 4169 5661 4203 5695
rect 4261 5661 4295 5695
rect 5549 5661 5583 5695
rect 6837 5661 6871 5695
rect 7941 5661 7975 5695
rect 9781 5661 9815 5695
rect 6285 5593 6319 5627
rect 3801 5525 3835 5559
rect 3709 5321 3743 5355
rect 4537 5321 4571 5355
rect 8493 5321 8527 5355
rect 9321 5321 9355 5355
rect 4445 5253 4479 5287
rect 1685 5185 1719 5219
rect 3525 5185 3559 5219
rect 5825 5185 5859 5219
rect 6101 5185 6135 5219
rect 7481 5185 7515 5219
rect 7757 5185 7791 5219
rect 9505 5185 9539 5219
rect 9781 5185 9815 5219
rect 5089 5049 5123 5083
rect 1501 4981 1535 5015
rect 9597 4981 9631 5015
rect 1685 4709 1719 4743
rect 5733 4641 5767 4675
rect 5549 4573 5583 4607
rect 1501 4505 1535 4539
rect 2605 2601 2639 2635
rect 2421 2397 2455 2431
<< metal1 >>
rect 7834 43460 7840 43512
rect 7892 43500 7898 43512
rect 8386 43500 8392 43512
rect 7892 43472 8392 43500
rect 7892 43460 7898 43472
rect 8386 43460 8392 43472
rect 8444 43460 8450 43512
rect 934 43256 940 43308
rect 992 43296 998 43308
rect 1394 43296 1400 43308
rect 992 43268 1400 43296
rect 992 43256 998 43268
rect 1394 43256 1400 43268
rect 1452 43256 1458 43308
rect 6730 42508 6736 42560
rect 6788 42548 6794 42560
rect 9214 42548 9220 42560
rect 6788 42520 9220 42548
rect 6788 42508 6794 42520
rect 9214 42508 9220 42520
rect 9272 42508 9278 42560
rect 1104 42458 10120 42480
rect 1104 42406 3010 42458
rect 3062 42406 3074 42458
rect 3126 42406 3138 42458
rect 3190 42406 3202 42458
rect 3254 42406 3266 42458
rect 3318 42406 9010 42458
rect 9062 42406 9074 42458
rect 9126 42406 9138 42458
rect 9190 42406 9202 42458
rect 9254 42406 9266 42458
rect 9318 42406 10120 42458
rect 1104 42384 10120 42406
rect 1486 42304 1492 42356
rect 1544 42344 1550 42356
rect 1581 42347 1639 42353
rect 1581 42344 1593 42347
rect 1544 42316 1593 42344
rect 1544 42304 1550 42316
rect 1581 42313 1593 42316
rect 1627 42313 1639 42347
rect 1581 42307 1639 42313
rect 1854 42304 1860 42356
rect 1912 42344 1918 42356
rect 2133 42347 2191 42353
rect 2133 42344 2145 42347
rect 1912 42316 2145 42344
rect 1912 42304 1918 42316
rect 2133 42313 2145 42316
rect 2179 42313 2191 42347
rect 2133 42307 2191 42313
rect 2314 42304 2320 42356
rect 2372 42344 2378 42356
rect 2593 42347 2651 42353
rect 2593 42344 2605 42347
rect 2372 42316 2605 42344
rect 2372 42304 2378 42316
rect 2593 42313 2605 42316
rect 2639 42313 2651 42347
rect 2593 42307 2651 42313
rect 2774 42304 2780 42356
rect 2832 42344 2838 42356
rect 2961 42347 3019 42353
rect 2961 42344 2973 42347
rect 2832 42316 2973 42344
rect 2832 42304 2838 42316
rect 2961 42313 2973 42316
rect 3007 42313 3019 42347
rect 2961 42307 3019 42313
rect 3418 42304 3424 42356
rect 3476 42304 3482 42356
rect 3694 42304 3700 42356
rect 3752 42344 3758 42356
rect 3881 42347 3939 42353
rect 3881 42344 3893 42347
rect 3752 42316 3893 42344
rect 3752 42304 3758 42316
rect 3881 42313 3893 42316
rect 3927 42313 3939 42347
rect 3881 42307 3939 42313
rect 4154 42304 4160 42356
rect 4212 42344 4218 42356
rect 4341 42347 4399 42353
rect 4341 42344 4353 42347
rect 4212 42316 4353 42344
rect 4212 42304 4218 42316
rect 4341 42313 4353 42316
rect 4387 42313 4399 42347
rect 4341 42307 4399 42313
rect 4614 42304 4620 42356
rect 4672 42344 4678 42356
rect 4801 42347 4859 42353
rect 4801 42344 4813 42347
rect 4672 42316 4813 42344
rect 4672 42304 4678 42316
rect 4801 42313 4813 42316
rect 4847 42313 4859 42347
rect 4801 42307 4859 42313
rect 5074 42304 5080 42356
rect 5132 42344 5138 42356
rect 5261 42347 5319 42353
rect 5261 42344 5273 42347
rect 5132 42316 5273 42344
rect 5132 42304 5138 42316
rect 5261 42313 5273 42316
rect 5307 42313 5319 42347
rect 5261 42307 5319 42313
rect 5534 42304 5540 42356
rect 5592 42344 5598 42356
rect 5629 42347 5687 42353
rect 5629 42344 5641 42347
rect 5592 42316 5641 42344
rect 5592 42304 5598 42316
rect 5629 42313 5641 42316
rect 5675 42313 5687 42347
rect 5629 42307 5687 42313
rect 5994 42304 6000 42356
rect 6052 42304 6058 42356
rect 6454 42304 6460 42356
rect 6512 42344 6518 42356
rect 6733 42347 6791 42353
rect 6733 42344 6745 42347
rect 6512 42316 6745 42344
rect 6512 42304 6518 42316
rect 6733 42313 6745 42316
rect 6779 42313 6791 42347
rect 6733 42307 6791 42313
rect 6914 42304 6920 42356
rect 6972 42344 6978 42356
rect 7285 42347 7343 42353
rect 7285 42344 7297 42347
rect 6972 42316 7297 42344
rect 6972 42304 6978 42316
rect 7285 42313 7297 42316
rect 7331 42313 7343 42347
rect 7285 42307 7343 42313
rect 7374 42304 7380 42356
rect 7432 42344 7438 42356
rect 7653 42347 7711 42353
rect 7653 42344 7665 42347
rect 7432 42316 7665 42344
rect 7432 42304 7438 42316
rect 7653 42313 7665 42316
rect 7699 42313 7711 42347
rect 7653 42307 7711 42313
rect 8386 42304 8392 42356
rect 8444 42304 8450 42356
rect 8754 42304 8760 42356
rect 8812 42344 8818 42356
rect 9493 42347 9551 42353
rect 9493 42344 9505 42347
rect 8812 42316 9505 42344
rect 8812 42304 8818 42316
rect 9493 42313 9505 42316
rect 9539 42313 9551 42347
rect 9493 42307 9551 42313
rect 3970 42276 3976 42288
rect 3160 42248 3976 42276
rect 1118 42168 1124 42220
rect 1176 42208 1182 42220
rect 1765 42211 1823 42217
rect 1765 42208 1777 42211
rect 1176 42180 1777 42208
rect 1176 42168 1182 42180
rect 1765 42177 1777 42180
rect 1811 42177 1823 42211
rect 1765 42171 1823 42177
rect 1949 42211 2007 42217
rect 1949 42177 1961 42211
rect 1995 42177 2007 42211
rect 1949 42171 2007 42177
rect 1964 42072 1992 42171
rect 2314 42168 2320 42220
rect 2372 42208 2378 42220
rect 3160 42217 3188 42248
rect 3970 42236 3976 42248
rect 4028 42236 4034 42288
rect 7190 42276 7196 42288
rect 4080 42248 7196 42276
rect 4080 42217 4108 42248
rect 7190 42236 7196 42248
rect 7248 42236 7254 42288
rect 8478 42236 8484 42288
rect 8536 42276 8542 42288
rect 8536 42248 9352 42276
rect 8536 42236 8542 42248
rect 2409 42211 2467 42217
rect 2409 42208 2421 42211
rect 2372 42180 2421 42208
rect 2372 42168 2378 42180
rect 2409 42177 2421 42180
rect 2455 42177 2467 42211
rect 2409 42171 2467 42177
rect 3145 42211 3203 42217
rect 3145 42177 3157 42211
rect 3191 42177 3203 42211
rect 3145 42171 3203 42177
rect 3605 42211 3663 42217
rect 3605 42177 3617 42211
rect 3651 42177 3663 42211
rect 3605 42171 3663 42177
rect 4065 42211 4123 42217
rect 4065 42177 4077 42211
rect 4111 42177 4123 42211
rect 4065 42171 4123 42177
rect 4525 42211 4583 42217
rect 4525 42177 4537 42211
rect 4571 42177 4583 42211
rect 4525 42171 4583 42177
rect 2406 42072 2412 42084
rect 1964 42044 2412 42072
rect 2406 42032 2412 42044
rect 2464 42032 2470 42084
rect 3620 42004 3648 42171
rect 4540 42072 4568 42171
rect 4982 42168 4988 42220
rect 5040 42168 5046 42220
rect 5442 42168 5448 42220
rect 5500 42168 5506 42220
rect 5813 42211 5871 42217
rect 5813 42177 5825 42211
rect 5859 42177 5871 42211
rect 5813 42171 5871 42177
rect 5828 42140 5856 42171
rect 6178 42168 6184 42220
rect 6236 42168 6242 42220
rect 6546 42168 6552 42220
rect 6604 42168 6610 42220
rect 7466 42168 7472 42220
rect 7524 42168 7530 42220
rect 7834 42168 7840 42220
rect 7892 42168 7898 42220
rect 8570 42168 8576 42220
rect 8628 42168 8634 42220
rect 9324 42217 9352 42248
rect 9217 42211 9275 42217
rect 9217 42177 9229 42211
rect 9263 42177 9275 42211
rect 9217 42171 9275 42177
rect 9309 42211 9367 42217
rect 9309 42177 9321 42211
rect 9355 42177 9367 42211
rect 9309 42171 9367 42177
rect 8754 42140 8760 42152
rect 5828 42112 8760 42140
rect 8754 42100 8760 42112
rect 8812 42100 8818 42152
rect 9232 42140 9260 42171
rect 9490 42140 9496 42152
rect 9232 42112 9496 42140
rect 9490 42100 9496 42112
rect 9548 42100 9554 42152
rect 7374 42072 7380 42084
rect 4540 42044 7380 42072
rect 7374 42032 7380 42044
rect 7432 42032 7438 42084
rect 8294 42032 8300 42084
rect 8352 42072 8358 42084
rect 9033 42075 9091 42081
rect 9033 42072 9045 42075
rect 8352 42044 9045 42072
rect 8352 42032 8358 42044
rect 9033 42041 9045 42044
rect 9079 42041 9091 42075
rect 9033 42035 9091 42041
rect 6914 42004 6920 42016
rect 3620 41976 6920 42004
rect 6914 41964 6920 41976
rect 6972 41964 6978 42016
rect 7006 41964 7012 42016
rect 7064 41964 7070 42016
rect 7282 41964 7288 42016
rect 7340 42004 7346 42016
rect 7742 42004 7748 42016
rect 7340 41976 7748 42004
rect 7340 41964 7346 41976
rect 7742 41964 7748 41976
rect 7800 42004 7806 42016
rect 8113 42007 8171 42013
rect 8113 42004 8125 42007
rect 7800 41976 8125 42004
rect 7800 41964 7806 41976
rect 8113 41973 8125 41976
rect 8159 41973 8171 42007
rect 8113 41967 8171 41973
rect 1104 41914 10120 41936
rect 1104 41862 1950 41914
rect 2002 41862 2014 41914
rect 2066 41862 2078 41914
rect 2130 41862 2142 41914
rect 2194 41862 2206 41914
rect 2258 41862 7950 41914
rect 8002 41862 8014 41914
rect 8066 41862 8078 41914
rect 8130 41862 8142 41914
rect 8194 41862 8206 41914
rect 8258 41862 10120 41914
rect 1104 41840 10120 41862
rect 1394 41760 1400 41812
rect 1452 41760 1458 41812
rect 6546 41760 6552 41812
rect 6604 41760 6610 41812
rect 6730 41760 6736 41812
rect 6788 41760 6794 41812
rect 7466 41760 7472 41812
rect 7524 41760 7530 41812
rect 7834 41760 7840 41812
rect 7892 41800 7898 41812
rect 8573 41803 8631 41809
rect 8573 41800 8585 41803
rect 7892 41772 8585 41800
rect 7892 41760 7898 41772
rect 8573 41769 8585 41772
rect 8619 41769 8631 41803
rect 8573 41763 8631 41769
rect 9309 41803 9367 41809
rect 9309 41769 9321 41803
rect 9355 41800 9367 41803
rect 10134 41800 10140 41812
rect 9355 41772 10140 41800
rect 9355 41769 9367 41772
rect 9309 41763 9367 41769
rect 10134 41760 10140 41772
rect 10192 41760 10198 41812
rect 5442 41692 5448 41744
rect 5500 41732 5506 41744
rect 8113 41735 8171 41741
rect 8113 41732 8125 41735
rect 5500 41704 8125 41732
rect 5500 41692 5506 41704
rect 8113 41701 8125 41704
rect 8159 41701 8171 41735
rect 8113 41695 8171 41701
rect 5994 41624 6000 41676
rect 6052 41664 6058 41676
rect 8386 41664 8392 41676
rect 6052 41636 6500 41664
rect 6052 41624 6058 41636
rect 1581 41599 1639 41605
rect 1581 41565 1593 41599
rect 1627 41596 1639 41599
rect 5442 41596 5448 41608
rect 1627 41568 5448 41596
rect 1627 41565 1639 41568
rect 1581 41559 1639 41565
rect 5442 41556 5448 41568
rect 5500 41556 5506 41608
rect 6273 41599 6331 41605
rect 6273 41565 6285 41599
rect 6319 41596 6331 41599
rect 6365 41599 6423 41605
rect 6365 41596 6377 41599
rect 6319 41568 6377 41596
rect 6319 41565 6331 41568
rect 6273 41559 6331 41565
rect 6365 41565 6377 41568
rect 6411 41565 6423 41599
rect 6365 41559 6423 41565
rect 4982 41488 4988 41540
rect 5040 41528 5046 41540
rect 6472 41528 6500 41636
rect 6932 41636 8392 41664
rect 6932 41605 6960 41636
rect 8386 41624 8392 41636
rect 8444 41624 8450 41676
rect 6917 41599 6975 41605
rect 6917 41565 6929 41599
rect 6963 41565 6975 41599
rect 6917 41559 6975 41565
rect 7006 41556 7012 41608
rect 7064 41596 7070 41608
rect 7193 41599 7251 41605
rect 7193 41596 7205 41599
rect 7064 41568 7205 41596
rect 7064 41556 7070 41568
rect 7193 41565 7205 41568
rect 7239 41565 7251 41599
rect 7193 41559 7251 41565
rect 7285 41599 7343 41605
rect 7285 41565 7297 41599
rect 7331 41596 7343 41599
rect 7561 41599 7619 41605
rect 7561 41596 7573 41599
rect 7331 41568 7573 41596
rect 7331 41565 7343 41568
rect 7285 41559 7343 41565
rect 7561 41565 7573 41568
rect 7607 41565 7619 41599
rect 7561 41559 7619 41565
rect 7300 41528 7328 41559
rect 8018 41556 8024 41608
rect 8076 41556 8082 41608
rect 8110 41556 8116 41608
rect 8168 41596 8174 41608
rect 8297 41599 8355 41605
rect 8297 41596 8309 41599
rect 8168 41568 8309 41596
rect 8168 41556 8174 41568
rect 8297 41565 8309 41568
rect 8343 41565 8355 41599
rect 8297 41559 8355 41565
rect 8757 41599 8815 41605
rect 8757 41565 8769 41599
rect 8803 41596 8815 41599
rect 8846 41596 8852 41608
rect 8803 41568 8852 41596
rect 8803 41565 8815 41568
rect 8757 41559 8815 41565
rect 8846 41556 8852 41568
rect 8904 41556 8910 41608
rect 9125 41599 9183 41605
rect 9125 41565 9137 41599
rect 9171 41596 9183 41599
rect 9398 41596 9404 41608
rect 9171 41568 9404 41596
rect 9171 41565 9183 41568
rect 9125 41559 9183 41565
rect 9398 41556 9404 41568
rect 9456 41556 9462 41608
rect 9493 41599 9551 41605
rect 9493 41565 9505 41599
rect 9539 41596 9551 41599
rect 9582 41596 9588 41608
rect 9539 41568 9588 41596
rect 9539 41565 9551 41568
rect 9493 41559 9551 41565
rect 9582 41556 9588 41568
rect 9640 41556 9646 41608
rect 9674 41556 9680 41608
rect 9732 41556 9738 41608
rect 9692 41528 9720 41556
rect 5040 41500 6316 41528
rect 6472 41500 7328 41528
rect 7852 41500 9720 41528
rect 5040 41488 5046 41500
rect 3786 41420 3792 41472
rect 3844 41460 3850 41472
rect 6181 41463 6239 41469
rect 6181 41460 6193 41463
rect 3844 41432 6193 41460
rect 3844 41420 3850 41432
rect 6181 41429 6193 41432
rect 6227 41429 6239 41463
rect 6288 41460 6316 41500
rect 7852 41469 7880 41500
rect 7009 41463 7067 41469
rect 7009 41460 7021 41463
rect 6288 41432 7021 41460
rect 6181 41423 6239 41429
rect 7009 41429 7021 41432
rect 7055 41429 7067 41463
rect 7009 41423 7067 41429
rect 7837 41463 7895 41469
rect 7837 41429 7849 41463
rect 7883 41429 7895 41463
rect 7837 41423 7895 41429
rect 9674 41420 9680 41472
rect 9732 41420 9738 41472
rect 1104 41370 10120 41392
rect 1104 41318 3010 41370
rect 3062 41318 3074 41370
rect 3126 41318 3138 41370
rect 3190 41318 3202 41370
rect 3254 41318 3266 41370
rect 3318 41318 9010 41370
rect 9062 41318 9074 41370
rect 9126 41318 9138 41370
rect 9190 41318 9202 41370
rect 9254 41318 9266 41370
rect 9318 41318 10120 41370
rect 1104 41296 10120 41318
rect 6178 41216 6184 41268
rect 6236 41256 6242 41268
rect 6733 41259 6791 41265
rect 6733 41256 6745 41259
rect 6236 41228 6745 41256
rect 6236 41216 6242 41228
rect 6733 41225 6745 41228
rect 6779 41225 6791 41259
rect 6733 41219 6791 41225
rect 6914 41216 6920 41268
rect 6972 41216 6978 41268
rect 7374 41216 7380 41268
rect 7432 41216 7438 41268
rect 7929 41259 7987 41265
rect 7929 41225 7941 41259
rect 7975 41225 7987 41259
rect 7929 41219 7987 41225
rect 6932 41188 6960 41216
rect 7944 41188 7972 41219
rect 8018 41216 8024 41268
rect 8076 41256 8082 41268
rect 8205 41259 8263 41265
rect 8205 41256 8217 41259
rect 8076 41228 8217 41256
rect 8076 41216 8082 41228
rect 8205 41225 8217 41228
rect 8251 41225 8263 41259
rect 8205 41219 8263 41225
rect 8665 41259 8723 41265
rect 8665 41225 8677 41259
rect 8711 41256 8723 41259
rect 8846 41256 8852 41268
rect 8711 41228 8852 41256
rect 8711 41225 8723 41228
rect 8665 41219 8723 41225
rect 8846 41216 8852 41228
rect 8904 41216 8910 41268
rect 9217 41259 9275 41265
rect 9217 41225 9229 41259
rect 9263 41256 9275 41259
rect 9398 41256 9404 41268
rect 9263 41228 9404 41256
rect 9263 41225 9275 41228
rect 9217 41219 9275 41225
rect 9398 41216 9404 41228
rect 9456 41216 9462 41268
rect 9490 41216 9496 41268
rect 9548 41216 9554 41268
rect 6932 41160 7972 41188
rect 1486 41080 1492 41132
rect 1544 41080 1550 41132
rect 6822 41080 6828 41132
rect 6880 41120 6886 41132
rect 6917 41123 6975 41129
rect 6917 41120 6929 41123
rect 6880 41092 6929 41120
rect 6880 41080 6886 41092
rect 6917 41089 6929 41092
rect 6963 41089 6975 41123
rect 6917 41083 6975 41089
rect 7006 41080 7012 41132
rect 7064 41080 7070 41132
rect 7561 41123 7619 41129
rect 7561 41089 7573 41123
rect 7607 41089 7619 41123
rect 7561 41083 7619 41089
rect 7653 41123 7711 41129
rect 7653 41089 7665 41123
rect 7699 41120 7711 41123
rect 7742 41120 7748 41132
rect 7699 41092 7748 41120
rect 7699 41089 7711 41092
rect 7653 41083 7711 41089
rect 842 41012 848 41064
rect 900 41052 906 41064
rect 7576 41052 7604 41083
rect 7742 41080 7748 41092
rect 7800 41080 7806 41132
rect 7834 41080 7840 41132
rect 7892 41120 7898 41132
rect 8113 41123 8171 41129
rect 8113 41120 8125 41123
rect 7892 41092 8125 41120
rect 7892 41080 7898 41092
rect 8113 41089 8125 41092
rect 8159 41089 8171 41123
rect 8113 41083 8171 41089
rect 8294 41080 8300 41132
rect 8352 41120 8358 41132
rect 8389 41123 8447 41129
rect 8389 41120 8401 41123
rect 8352 41092 8401 41120
rect 8352 41080 8358 41092
rect 8389 41089 8401 41092
rect 8435 41089 8447 41123
rect 8389 41083 8447 41089
rect 8849 41123 8907 41129
rect 8849 41089 8861 41123
rect 8895 41089 8907 41123
rect 8849 41083 8907 41089
rect 8864 41052 8892 41083
rect 9398 41080 9404 41132
rect 9456 41080 9462 41132
rect 9677 41123 9735 41129
rect 9677 41089 9689 41123
rect 9723 41120 9735 41123
rect 9766 41120 9772 41132
rect 9723 41092 9772 41120
rect 9723 41089 9735 41092
rect 9677 41083 9735 41089
rect 9766 41080 9772 41092
rect 9824 41080 9830 41132
rect 900 41024 7604 41052
rect 7668 41024 8892 41052
rect 900 41012 906 41024
rect 1673 40987 1731 40993
rect 1673 40953 1685 40987
rect 1719 40984 1731 40987
rect 1854 40984 1860 40996
rect 1719 40956 1860 40984
rect 1719 40953 1731 40956
rect 1673 40947 1731 40953
rect 1854 40944 1860 40956
rect 1912 40944 1918 40996
rect 3878 40944 3884 40996
rect 3936 40984 3942 40996
rect 7668 40984 7696 41024
rect 3936 40956 7696 40984
rect 7837 40987 7895 40993
rect 3936 40944 3942 40956
rect 7837 40953 7849 40987
rect 7883 40984 7895 40987
rect 8478 40984 8484 40996
rect 7883 40956 8484 40984
rect 7883 40953 7895 40956
rect 7837 40947 7895 40953
rect 8478 40944 8484 40956
rect 8536 40944 8542 40996
rect 8570 40876 8576 40928
rect 8628 40876 8634 40928
rect 9033 40919 9091 40925
rect 9033 40885 9045 40919
rect 9079 40916 9091 40919
rect 10410 40916 10416 40928
rect 9079 40888 10416 40916
rect 9079 40885 9091 40888
rect 9033 40879 9091 40885
rect 10410 40876 10416 40888
rect 10468 40876 10474 40928
rect 1104 40826 10120 40848
rect 1104 40774 1950 40826
rect 2002 40774 2014 40826
rect 2066 40774 2078 40826
rect 2130 40774 2142 40826
rect 2194 40774 2206 40826
rect 2258 40774 7950 40826
rect 8002 40774 8014 40826
rect 8066 40774 8078 40826
rect 8130 40774 8142 40826
rect 8194 40774 8206 40826
rect 8258 40774 10120 40826
rect 1104 40752 10120 40774
rect 7190 40672 7196 40724
rect 7248 40712 7254 40724
rect 7377 40715 7435 40721
rect 7377 40712 7389 40715
rect 7248 40684 7389 40712
rect 7248 40672 7254 40684
rect 7377 40681 7389 40684
rect 7423 40681 7435 40715
rect 7377 40675 7435 40681
rect 8386 40672 8392 40724
rect 8444 40712 8450 40724
rect 8573 40715 8631 40721
rect 8573 40712 8585 40715
rect 8444 40684 8585 40712
rect 8444 40672 8450 40684
rect 8573 40681 8585 40684
rect 8619 40681 8631 40715
rect 8573 40675 8631 40681
rect 8662 40672 8668 40724
rect 8720 40712 8726 40724
rect 8941 40715 8999 40721
rect 8941 40712 8953 40715
rect 8720 40684 8953 40712
rect 8720 40672 8726 40684
rect 8941 40681 8953 40684
rect 8987 40681 8999 40715
rect 8941 40675 8999 40681
rect 7374 40468 7380 40520
rect 7432 40508 7438 40520
rect 7561 40511 7619 40517
rect 7561 40508 7573 40511
rect 7432 40480 7573 40508
rect 7432 40468 7438 40480
rect 7561 40477 7573 40480
rect 7607 40477 7619 40511
rect 7561 40471 7619 40477
rect 8662 40468 8668 40520
rect 8720 40508 8726 40520
rect 8757 40511 8815 40517
rect 8757 40508 8769 40511
rect 8720 40480 8769 40508
rect 8720 40468 8726 40480
rect 8757 40477 8769 40480
rect 8803 40477 8815 40511
rect 8757 40471 8815 40477
rect 9125 40511 9183 40517
rect 9125 40477 9137 40511
rect 9171 40508 9183 40511
rect 9582 40508 9588 40520
rect 9171 40480 9588 40508
rect 9171 40477 9183 40480
rect 9125 40471 9183 40477
rect 9582 40468 9588 40480
rect 9640 40468 9646 40520
rect 1486 40400 1492 40452
rect 1544 40400 1550 40452
rect 1673 40443 1731 40449
rect 1673 40409 1685 40443
rect 1719 40440 1731 40443
rect 1762 40440 1768 40452
rect 1719 40412 1768 40440
rect 1719 40409 1731 40412
rect 1673 40403 1731 40409
rect 1762 40400 1768 40412
rect 1820 40400 1826 40452
rect 7466 40400 7472 40452
rect 7524 40440 7530 40452
rect 7834 40440 7840 40452
rect 7524 40412 7840 40440
rect 7524 40400 7530 40412
rect 7834 40400 7840 40412
rect 7892 40440 7898 40452
rect 7929 40443 7987 40449
rect 7929 40440 7941 40443
rect 7892 40412 7941 40440
rect 7892 40400 7898 40412
rect 7929 40409 7941 40412
rect 7975 40409 7987 40443
rect 7929 40403 7987 40409
rect 6822 40332 6828 40384
rect 6880 40332 6886 40384
rect 7742 40332 7748 40384
rect 7800 40332 7806 40384
rect 8294 40332 8300 40384
rect 8352 40332 8358 40384
rect 9309 40375 9367 40381
rect 9309 40341 9321 40375
rect 9355 40372 9367 40375
rect 9398 40372 9404 40384
rect 9355 40344 9404 40372
rect 9355 40341 9367 40344
rect 9309 40335 9367 40341
rect 9398 40332 9404 40344
rect 9456 40332 9462 40384
rect 9585 40375 9643 40381
rect 9585 40341 9597 40375
rect 9631 40372 9643 40375
rect 9766 40372 9772 40384
rect 9631 40344 9772 40372
rect 9631 40341 9643 40344
rect 9585 40335 9643 40341
rect 9766 40332 9772 40344
rect 9824 40332 9830 40384
rect 1104 40282 10120 40304
rect 1104 40230 3010 40282
rect 3062 40230 3074 40282
rect 3126 40230 3138 40282
rect 3190 40230 3202 40282
rect 3254 40230 3266 40282
rect 3318 40230 9010 40282
rect 9062 40230 9074 40282
rect 9126 40230 9138 40282
rect 9190 40230 9202 40282
rect 9254 40230 9266 40282
rect 9318 40230 10120 40282
rect 1104 40208 10120 40230
rect 4062 40128 4068 40180
rect 4120 40168 4126 40180
rect 4120 40140 9168 40168
rect 4120 40128 4126 40140
rect 566 40060 572 40112
rect 624 40100 630 40112
rect 624 40072 8984 40100
rect 624 40060 630 40072
rect 8956 40041 8984 40072
rect 9140 40041 9168 40140
rect 9214 40060 9220 40112
rect 9272 40100 9278 40112
rect 9272 40072 9536 40100
rect 9272 40060 9278 40072
rect 9508 40041 9536 40072
rect 8941 40035 8999 40041
rect 8941 40001 8953 40035
rect 8987 40001 8999 40035
rect 8941 39995 8999 40001
rect 9125 40035 9183 40041
rect 9125 40001 9137 40035
rect 9171 40001 9183 40035
rect 9125 39995 9183 40001
rect 9493 40035 9551 40041
rect 9493 40001 9505 40035
rect 9539 40001 9551 40035
rect 9493 39995 9551 40001
rect 8754 39856 8760 39908
rect 8812 39856 8818 39908
rect 9309 39899 9367 39905
rect 9309 39865 9321 39899
rect 9355 39896 9367 39899
rect 10594 39896 10600 39908
rect 9355 39868 10600 39896
rect 9355 39865 9367 39868
rect 9309 39859 9367 39865
rect 10594 39856 10600 39868
rect 10652 39856 10658 39908
rect 7374 39788 7380 39840
rect 7432 39788 7438 39840
rect 8662 39788 8668 39840
rect 8720 39788 8726 39840
rect 9677 39831 9735 39837
rect 9677 39797 9689 39831
rect 9723 39828 9735 39831
rect 10778 39828 10784 39840
rect 9723 39800 10784 39828
rect 9723 39797 9735 39800
rect 9677 39791 9735 39797
rect 10778 39788 10784 39800
rect 10836 39788 10842 39840
rect 1104 39738 10120 39760
rect 1104 39686 1950 39738
rect 2002 39686 2014 39738
rect 2066 39686 2078 39738
rect 2130 39686 2142 39738
rect 2194 39686 2206 39738
rect 2258 39686 7950 39738
rect 8002 39686 8014 39738
rect 8066 39686 8078 39738
rect 8130 39686 8142 39738
rect 8194 39686 8206 39738
rect 8258 39686 10120 39738
rect 1104 39664 10120 39686
rect 9309 39559 9367 39565
rect 9309 39525 9321 39559
rect 9355 39556 9367 39559
rect 10226 39556 10232 39568
rect 9355 39528 10232 39556
rect 9355 39525 9367 39528
rect 9309 39519 9367 39525
rect 10226 39516 10232 39528
rect 10284 39516 10290 39568
rect 3694 39448 3700 39500
rect 3752 39488 3758 39500
rect 3970 39488 3976 39500
rect 3752 39460 3976 39488
rect 3752 39448 3758 39460
rect 3970 39448 3976 39460
rect 4028 39448 4034 39500
rect 5166 39380 5172 39432
rect 5224 39380 5230 39432
rect 5445 39423 5503 39429
rect 5445 39389 5457 39423
rect 5491 39420 5503 39423
rect 5810 39420 5816 39432
rect 5491 39392 5816 39420
rect 5491 39389 5503 39392
rect 5445 39383 5503 39389
rect 5810 39380 5816 39392
rect 5868 39380 5874 39432
rect 9125 39423 9183 39429
rect 9125 39389 9137 39423
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 1486 39312 1492 39364
rect 1544 39312 1550 39364
rect 1673 39355 1731 39361
rect 1673 39321 1685 39355
rect 1719 39352 1731 39355
rect 2774 39352 2780 39364
rect 1719 39324 2780 39352
rect 1719 39321 1731 39324
rect 1673 39315 1731 39321
rect 2774 39312 2780 39324
rect 2832 39312 2838 39364
rect 3970 39312 3976 39364
rect 4028 39352 4034 39364
rect 9140 39352 9168 39383
rect 9490 39380 9496 39432
rect 9548 39380 9554 39432
rect 4028 39324 9168 39352
rect 4028 39312 4034 39324
rect 4430 39244 4436 39296
rect 4488 39244 4494 39296
rect 9677 39287 9735 39293
rect 9677 39253 9689 39287
rect 9723 39284 9735 39287
rect 10410 39284 10416 39296
rect 9723 39256 10416 39284
rect 9723 39253 9735 39256
rect 9677 39247 9735 39253
rect 10410 39244 10416 39256
rect 10468 39244 10474 39296
rect 1104 39194 10120 39216
rect 1104 39142 3010 39194
rect 3062 39142 3074 39194
rect 3126 39142 3138 39194
rect 3190 39142 3202 39194
rect 3254 39142 3266 39194
rect 3318 39142 9010 39194
rect 9062 39142 9074 39194
rect 9126 39142 9138 39194
rect 9190 39142 9202 39194
rect 9254 39142 9266 39194
rect 9318 39142 10120 39194
rect 1104 39120 10120 39142
rect 9309 39083 9367 39089
rect 9309 39049 9321 39083
rect 9355 39080 9367 39083
rect 10318 39080 10324 39092
rect 9355 39052 10324 39080
rect 9355 39049 9367 39052
rect 9309 39043 9367 39049
rect 10318 39040 10324 39052
rect 10376 39040 10382 39092
rect 5810 39012 5816 39024
rect 4448 38984 5816 39012
rect 750 38904 756 38956
rect 808 38944 814 38956
rect 1489 38947 1547 38953
rect 1489 38944 1501 38947
rect 808 38916 1501 38944
rect 808 38904 814 38916
rect 1489 38913 1501 38916
rect 1535 38913 1547 38947
rect 1489 38907 1547 38913
rect 3881 38947 3939 38953
rect 3881 38913 3893 38947
rect 3927 38944 3939 38947
rect 4338 38944 4344 38956
rect 3927 38916 4344 38944
rect 3927 38913 3939 38916
rect 3881 38907 3939 38913
rect 4338 38904 4344 38916
rect 4396 38904 4402 38956
rect 4448 38953 4476 38984
rect 5810 38972 5816 38984
rect 5868 38972 5874 39024
rect 4433 38947 4491 38953
rect 4433 38913 4445 38947
rect 4479 38913 4491 38947
rect 4433 38907 4491 38913
rect 4709 38947 4767 38953
rect 4709 38913 4721 38947
rect 4755 38944 4767 38947
rect 4982 38944 4988 38956
rect 4755 38916 4988 38944
rect 4755 38913 4767 38916
rect 4709 38907 4767 38913
rect 4982 38904 4988 38916
rect 5040 38904 5046 38956
rect 5718 38904 5724 38956
rect 5776 38904 5782 38956
rect 6365 38947 6423 38953
rect 6365 38913 6377 38947
rect 6411 38913 6423 38947
rect 6365 38907 6423 38913
rect 5000 38876 5028 38904
rect 6380 38876 6408 38907
rect 8754 38904 8760 38956
rect 8812 38904 8818 38956
rect 9122 38904 9128 38956
rect 9180 38904 9186 38956
rect 9490 38904 9496 38956
rect 9548 38904 9554 38956
rect 5000 38848 6408 38876
rect 1673 38811 1731 38817
rect 1673 38777 1685 38811
rect 1719 38808 1731 38811
rect 2590 38808 2596 38820
rect 1719 38780 2596 38808
rect 1719 38777 1731 38780
rect 1673 38771 1731 38777
rect 2590 38768 2596 38780
rect 2648 38768 2654 38820
rect 8941 38811 8999 38817
rect 8941 38777 8953 38811
rect 8987 38808 8999 38811
rect 10134 38808 10140 38820
rect 8987 38780 10140 38808
rect 8987 38777 8999 38780
rect 8941 38771 8999 38777
rect 10134 38768 10140 38780
rect 10192 38768 10198 38820
rect 4065 38743 4123 38749
rect 4065 38709 4077 38743
rect 4111 38740 4123 38743
rect 5258 38740 5264 38752
rect 4111 38712 5264 38740
rect 4111 38709 4123 38712
rect 4065 38703 4123 38709
rect 5258 38700 5264 38712
rect 5316 38700 5322 38752
rect 5350 38700 5356 38752
rect 5408 38740 5414 38752
rect 5445 38743 5503 38749
rect 5445 38740 5457 38743
rect 5408 38712 5457 38740
rect 5408 38700 5414 38712
rect 5445 38709 5457 38712
rect 5491 38709 5503 38743
rect 5445 38703 5503 38709
rect 5905 38743 5963 38749
rect 5905 38709 5917 38743
rect 5951 38740 5963 38743
rect 6270 38740 6276 38752
rect 5951 38712 6276 38740
rect 5951 38709 5963 38712
rect 5905 38703 5963 38709
rect 6270 38700 6276 38712
rect 6328 38700 6334 38752
rect 6549 38743 6607 38749
rect 6549 38709 6561 38743
rect 6595 38740 6607 38743
rect 8846 38740 8852 38752
rect 6595 38712 8852 38740
rect 6595 38709 6607 38712
rect 6549 38703 6607 38709
rect 8846 38700 8852 38712
rect 8904 38700 8910 38752
rect 9677 38743 9735 38749
rect 9677 38709 9689 38743
rect 9723 38740 9735 38743
rect 10502 38740 10508 38752
rect 9723 38712 10508 38740
rect 9723 38709 9735 38712
rect 9677 38703 9735 38709
rect 10502 38700 10508 38712
rect 10560 38700 10566 38752
rect 1104 38650 10120 38672
rect 1104 38598 1950 38650
rect 2002 38598 2014 38650
rect 2066 38598 2078 38650
rect 2130 38598 2142 38650
rect 2194 38598 2206 38650
rect 2258 38598 7950 38650
rect 8002 38598 8014 38650
rect 8066 38598 8078 38650
rect 8130 38598 8142 38650
rect 8194 38598 8206 38650
rect 8258 38598 10120 38650
rect 1104 38576 10120 38598
rect 3418 38496 3424 38548
rect 3476 38536 3482 38548
rect 4706 38536 4712 38548
rect 3476 38508 4712 38536
rect 3476 38496 3482 38508
rect 4706 38496 4712 38508
rect 4764 38496 4770 38548
rect 5718 38496 5724 38548
rect 5776 38536 5782 38548
rect 5997 38539 6055 38545
rect 5997 38536 6009 38539
rect 5776 38508 6009 38536
rect 5776 38496 5782 38508
rect 5997 38505 6009 38508
rect 6043 38505 6055 38539
rect 5997 38499 6055 38505
rect 4430 38428 4436 38480
rect 4488 38468 4494 38480
rect 4801 38471 4859 38477
rect 4801 38468 4813 38471
rect 4488 38440 4813 38468
rect 4488 38428 4494 38440
rect 4801 38437 4813 38440
rect 4847 38437 4859 38471
rect 4801 38431 4859 38437
rect 9309 38471 9367 38477
rect 9309 38437 9321 38471
rect 9355 38468 9367 38471
rect 10042 38468 10048 38480
rect 9355 38440 10048 38468
rect 9355 38437 9367 38440
rect 9309 38431 9367 38437
rect 10042 38428 10048 38440
rect 10100 38428 10106 38480
rect 2682 38360 2688 38412
rect 2740 38400 2746 38412
rect 4341 38403 4399 38409
rect 4341 38400 4353 38403
rect 2740 38372 4353 38400
rect 2740 38360 2746 38372
rect 4341 38369 4353 38372
rect 4387 38369 4399 38403
rect 5194 38403 5252 38409
rect 5194 38400 5206 38403
rect 4341 38363 4399 38369
rect 4448 38372 5206 38400
rect 1578 38292 1584 38344
rect 1636 38332 1642 38344
rect 1949 38335 2007 38341
rect 1949 38332 1961 38335
rect 1636 38304 1961 38332
rect 1636 38292 1642 38304
rect 1949 38301 1961 38304
rect 1995 38301 2007 38335
rect 1949 38295 2007 38301
rect 2225 38335 2283 38341
rect 2225 38301 2237 38335
rect 2271 38301 2283 38335
rect 2225 38295 2283 38301
rect 1486 38224 1492 38276
rect 1544 38224 1550 38276
rect 1854 38224 1860 38276
rect 1912 38264 1918 38276
rect 2240 38264 2268 38295
rect 2498 38292 2504 38344
rect 2556 38332 2562 38344
rect 4157 38335 4215 38341
rect 4157 38332 4169 38335
rect 2556 38304 4169 38332
rect 2556 38292 2562 38304
rect 4157 38301 4169 38304
rect 4203 38301 4215 38335
rect 4448 38332 4476 38372
rect 5194 38369 5206 38372
rect 5240 38369 5252 38403
rect 5194 38363 5252 38369
rect 5350 38360 5356 38412
rect 5408 38360 5414 38412
rect 6454 38360 6460 38412
rect 6512 38360 6518 38412
rect 7024 38372 9536 38400
rect 4157 38295 4215 38301
rect 4264 38304 4476 38332
rect 3418 38264 3424 38276
rect 1912 38236 2268 38264
rect 2746 38236 3424 38264
rect 1912 38224 1918 38236
rect 1581 38199 1639 38205
rect 1581 38165 1593 38199
rect 1627 38196 1639 38199
rect 2746 38196 2774 38236
rect 3418 38224 3424 38236
rect 3476 38224 3482 38276
rect 3510 38224 3516 38276
rect 3568 38264 3574 38276
rect 4264 38264 4292 38304
rect 5074 38292 5080 38344
rect 5132 38292 5138 38344
rect 6178 38292 6184 38344
rect 6236 38332 6242 38344
rect 6733 38335 6791 38341
rect 6733 38332 6745 38335
rect 6236 38304 6745 38332
rect 6236 38292 6242 38304
rect 6733 38301 6745 38304
rect 6779 38301 6791 38335
rect 6733 38295 6791 38301
rect 7024 38264 7052 38372
rect 8478 38292 8484 38344
rect 8536 38292 8542 38344
rect 9122 38292 9128 38344
rect 9180 38292 9186 38344
rect 9508 38341 9536 38372
rect 9493 38335 9551 38341
rect 9493 38301 9505 38335
rect 9539 38301 9551 38335
rect 9493 38295 9551 38301
rect 9950 38264 9956 38276
rect 3568 38236 4292 38264
rect 5828 38236 7052 38264
rect 8680 38236 9956 38264
rect 3568 38224 3574 38236
rect 1627 38168 2774 38196
rect 1627 38165 1639 38168
rect 1581 38159 1639 38165
rect 2866 38156 2872 38208
rect 2924 38196 2930 38208
rect 2961 38199 3019 38205
rect 2961 38196 2973 38199
rect 2924 38168 2973 38196
rect 2924 38156 2930 38168
rect 2961 38165 2973 38168
rect 3007 38165 3019 38199
rect 2961 38159 3019 38165
rect 4154 38156 4160 38208
rect 4212 38196 4218 38208
rect 5828 38196 5856 38236
rect 4212 38168 5856 38196
rect 6365 38199 6423 38205
rect 4212 38156 4218 38168
rect 6365 38165 6377 38199
rect 6411 38196 6423 38199
rect 6638 38196 6644 38208
rect 6411 38168 6644 38196
rect 6411 38165 6423 38168
rect 6365 38159 6423 38165
rect 6638 38156 6644 38168
rect 6696 38156 6702 38208
rect 7469 38199 7527 38205
rect 7469 38165 7481 38199
rect 7515 38196 7527 38199
rect 7834 38196 7840 38208
rect 7515 38168 7840 38196
rect 7515 38165 7527 38168
rect 7469 38159 7527 38165
rect 7834 38156 7840 38168
rect 7892 38156 7898 38208
rect 8680 38205 8708 38236
rect 9950 38224 9956 38236
rect 10008 38224 10014 38276
rect 8665 38199 8723 38205
rect 8665 38165 8677 38199
rect 8711 38165 8723 38199
rect 8665 38159 8723 38165
rect 9677 38199 9735 38205
rect 9677 38165 9689 38199
rect 9723 38196 9735 38199
rect 10962 38196 10968 38208
rect 9723 38168 10968 38196
rect 9723 38165 9735 38168
rect 9677 38159 9735 38165
rect 10962 38156 10968 38168
rect 11020 38156 11026 38208
rect 1104 38106 10120 38128
rect 1104 38054 3010 38106
rect 3062 38054 3074 38106
rect 3126 38054 3138 38106
rect 3190 38054 3202 38106
rect 3254 38054 3266 38106
rect 3318 38054 9010 38106
rect 9062 38054 9074 38106
rect 9126 38054 9138 38106
rect 9190 38054 9202 38106
rect 9254 38054 9266 38106
rect 9318 38054 10120 38106
rect 1104 38032 10120 38054
rect 474 37952 480 38004
rect 532 37992 538 38004
rect 3970 37992 3976 38004
rect 532 37964 3976 37992
rect 532 37952 538 37964
rect 3970 37952 3976 37964
rect 4028 37952 4034 38004
rect 4338 37952 4344 38004
rect 4396 37952 4402 38004
rect 5166 37992 5172 38004
rect 4724 37964 5172 37992
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37856 1455 37859
rect 1578 37856 1584 37868
rect 1443 37828 1584 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 1578 37816 1584 37828
rect 1636 37816 1642 37868
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37856 1731 37859
rect 1762 37856 1768 37868
rect 1719 37828 1768 37856
rect 1719 37825 1731 37828
rect 1673 37819 1731 37825
rect 1762 37816 1768 37828
rect 1820 37816 1826 37868
rect 4614 37816 4620 37868
rect 4672 37856 4678 37868
rect 4724 37865 4752 37964
rect 5166 37952 5172 37964
rect 5224 37992 5230 38004
rect 6178 37992 6184 38004
rect 5224 37964 6184 37992
rect 5224 37952 5230 37964
rect 6178 37952 6184 37964
rect 6236 37952 6242 38004
rect 9309 37995 9367 38001
rect 9309 37961 9321 37995
rect 9355 37992 9367 37995
rect 10134 37992 10140 38004
rect 9355 37964 10140 37992
rect 9355 37961 9367 37964
rect 9309 37955 9367 37961
rect 10134 37952 10140 37964
rect 10192 37952 10198 38004
rect 5902 37884 5908 37936
rect 5960 37924 5966 37936
rect 5960 37896 9168 37924
rect 5960 37884 5966 37896
rect 4709 37859 4767 37865
rect 4709 37856 4721 37859
rect 4672 37828 4721 37856
rect 4672 37816 4678 37828
rect 4709 37825 4721 37828
rect 4755 37825 4767 37859
rect 4709 37819 4767 37825
rect 5626 37816 5632 37868
rect 5684 37816 5690 37868
rect 6362 37816 6368 37868
rect 6420 37816 6426 37868
rect 8662 37816 8668 37868
rect 8720 37816 8726 37868
rect 8754 37816 8760 37868
rect 8812 37816 8818 37868
rect 9140 37865 9168 37896
rect 9125 37859 9183 37865
rect 9125 37825 9137 37859
rect 9171 37825 9183 37859
rect 9125 37819 9183 37825
rect 9493 37859 9551 37865
rect 9493 37825 9505 37859
rect 9539 37825 9551 37859
rect 9493 37819 9551 37825
rect 2498 37748 2504 37800
rect 2556 37748 2562 37800
rect 2682 37748 2688 37800
rect 2740 37748 2746 37800
rect 2866 37748 2872 37800
rect 2924 37788 2930 37800
rect 3145 37791 3203 37797
rect 3145 37788 3157 37791
rect 2924 37760 3157 37788
rect 2924 37748 2930 37760
rect 3145 37757 3157 37760
rect 3191 37757 3203 37791
rect 3145 37751 3203 37757
rect 3418 37748 3424 37800
rect 3476 37748 3482 37800
rect 3510 37748 3516 37800
rect 3568 37797 3574 37800
rect 3568 37791 3596 37797
rect 3584 37757 3596 37791
rect 3568 37751 3596 37757
rect 3697 37791 3755 37797
rect 3697 37757 3709 37791
rect 3743 37788 3755 37791
rect 3743 37760 4108 37788
rect 3743 37757 3755 37760
rect 3697 37751 3755 37757
rect 3568 37748 3574 37751
rect 2409 37655 2467 37661
rect 2409 37621 2421 37655
rect 2455 37652 2467 37655
rect 4080 37652 4108 37760
rect 4246 37748 4252 37800
rect 4304 37788 4310 37800
rect 4433 37791 4491 37797
rect 4433 37788 4445 37791
rect 4304 37760 4445 37788
rect 4304 37748 4310 37760
rect 4433 37757 4445 37760
rect 4479 37757 4491 37791
rect 4433 37751 4491 37757
rect 7006 37748 7012 37800
rect 7064 37788 7070 37800
rect 9508 37788 9536 37819
rect 7064 37760 9536 37788
rect 7064 37748 7070 37760
rect 5810 37680 5816 37732
rect 5868 37680 5874 37732
rect 8941 37723 8999 37729
rect 8941 37689 8953 37723
rect 8987 37720 8999 37723
rect 10226 37720 10232 37732
rect 8987 37692 10232 37720
rect 8987 37689 8999 37692
rect 8941 37683 8999 37689
rect 10226 37680 10232 37692
rect 10284 37680 10290 37732
rect 2455 37624 4108 37652
rect 2455 37621 2467 37624
rect 2409 37615 2467 37621
rect 4890 37612 4896 37664
rect 4948 37652 4954 37664
rect 5445 37655 5503 37661
rect 5445 37652 5457 37655
rect 4948 37624 5457 37652
rect 4948 37612 4954 37624
rect 5445 37621 5457 37624
rect 5491 37621 5503 37655
rect 5445 37615 5503 37621
rect 6914 37612 6920 37664
rect 6972 37652 6978 37664
rect 7653 37655 7711 37661
rect 7653 37652 7665 37655
rect 6972 37624 7665 37652
rect 6972 37612 6978 37624
rect 7653 37621 7665 37624
rect 7699 37621 7711 37655
rect 7653 37615 7711 37621
rect 8478 37612 8484 37664
rect 8536 37612 8542 37664
rect 9677 37655 9735 37661
rect 9677 37621 9689 37655
rect 9723 37652 9735 37655
rect 10594 37652 10600 37664
rect 9723 37624 10600 37652
rect 9723 37621 9735 37624
rect 9677 37615 9735 37621
rect 10594 37612 10600 37624
rect 10652 37612 10658 37664
rect 1104 37562 10120 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 7950 37562
rect 8002 37510 8014 37562
rect 8066 37510 8078 37562
rect 8130 37510 8142 37562
rect 8194 37510 8206 37562
rect 8258 37510 10120 37562
rect 1104 37488 10120 37510
rect 198 37408 204 37460
rect 256 37448 262 37460
rect 5537 37451 5595 37457
rect 5537 37448 5549 37451
rect 256 37420 5549 37448
rect 256 37408 262 37420
rect 5537 37417 5549 37420
rect 5583 37448 5595 37451
rect 5626 37448 5632 37460
rect 5583 37420 5632 37448
rect 5583 37417 5595 37420
rect 5537 37411 5595 37417
rect 5626 37408 5632 37420
rect 5684 37408 5690 37460
rect 6362 37408 6368 37460
rect 6420 37448 6426 37460
rect 7009 37451 7067 37457
rect 7009 37448 7021 37451
rect 6420 37420 7021 37448
rect 6420 37408 6426 37420
rect 7009 37417 7021 37420
rect 7055 37417 7067 37451
rect 7009 37411 7067 37417
rect 6086 37340 6092 37392
rect 6144 37380 6150 37392
rect 7466 37380 7472 37392
rect 6144 37352 7472 37380
rect 6144 37340 6150 37352
rect 7466 37340 7472 37352
rect 7524 37340 7530 37392
rect 5258 37272 5264 37324
rect 5316 37312 5322 37324
rect 7374 37312 7380 37324
rect 5316 37284 7380 37312
rect 5316 37272 5322 37284
rect 7374 37272 7380 37284
rect 7432 37272 7438 37324
rect 7558 37272 7564 37324
rect 7616 37272 7622 37324
rect 1670 37204 1676 37256
rect 1728 37204 1734 37256
rect 1765 37247 1823 37253
rect 1765 37213 1777 37247
rect 1811 37213 1823 37247
rect 1765 37207 1823 37213
rect 1486 37136 1492 37188
rect 1544 37136 1550 37188
rect 1578 37136 1584 37188
rect 1636 37176 1642 37188
rect 1780 37176 1808 37207
rect 1854 37204 1860 37256
rect 1912 37244 1918 37256
rect 2133 37247 2191 37253
rect 2133 37244 2145 37247
rect 1912 37216 2145 37244
rect 1912 37204 1918 37216
rect 2133 37213 2145 37216
rect 2179 37213 2191 37247
rect 2409 37247 2467 37253
rect 2409 37244 2421 37247
rect 2133 37207 2191 37213
rect 2240 37216 2421 37244
rect 1636 37148 1808 37176
rect 1636 37136 1642 37148
rect 2038 37136 2044 37188
rect 2096 37176 2102 37188
rect 2240 37176 2268 37216
rect 2409 37213 2421 37216
rect 2455 37213 2467 37247
rect 2409 37207 2467 37213
rect 4246 37204 4252 37256
rect 4304 37204 4310 37256
rect 4522 37204 4528 37256
rect 4580 37204 4586 37256
rect 4982 37204 4988 37256
rect 5040 37244 5046 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 5040 37216 7849 37244
rect 5040 37204 5046 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 7837 37207 7895 37213
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 4062 37176 4068 37188
rect 2096 37148 2268 37176
rect 2332 37148 4068 37176
rect 2096 37136 2102 37148
rect 1949 37111 2007 37117
rect 1949 37077 1961 37111
rect 1995 37108 2007 37111
rect 2222 37108 2228 37120
rect 1995 37080 2228 37108
rect 1995 37077 2007 37080
rect 1949 37071 2007 37077
rect 2222 37068 2228 37080
rect 2280 37068 2286 37120
rect 2332 37117 2360 37148
rect 4062 37136 4068 37148
rect 4120 37136 4126 37188
rect 5626 37176 5632 37188
rect 5276 37148 5632 37176
rect 2317 37111 2375 37117
rect 2317 37077 2329 37111
rect 2363 37077 2375 37111
rect 2317 37071 2375 37077
rect 2593 37111 2651 37117
rect 2593 37077 2605 37111
rect 2639 37108 2651 37111
rect 3878 37108 3884 37120
rect 2639 37080 3884 37108
rect 2639 37077 2651 37080
rect 2593 37071 2651 37077
rect 3878 37068 3884 37080
rect 3936 37068 3942 37120
rect 5276 37117 5304 37148
rect 5626 37136 5632 37148
rect 5684 37136 5690 37188
rect 5718 37136 5724 37188
rect 5776 37136 5782 37188
rect 6546 37136 6552 37188
rect 6604 37176 6610 37188
rect 9140 37176 9168 37207
rect 9398 37204 9404 37256
rect 9456 37244 9462 37256
rect 9493 37247 9551 37253
rect 9493 37244 9505 37247
rect 9456 37216 9505 37244
rect 9456 37204 9462 37216
rect 9493 37213 9505 37216
rect 9539 37213 9551 37247
rect 9493 37207 9551 37213
rect 10318 37176 10324 37188
rect 6604 37148 9168 37176
rect 9324 37148 10324 37176
rect 6604 37136 6610 37148
rect 5261 37111 5319 37117
rect 5261 37077 5273 37111
rect 5307 37077 5319 37111
rect 5261 37071 5319 37077
rect 8386 37068 8392 37120
rect 8444 37108 8450 37120
rect 9324 37117 9352 37148
rect 10318 37136 10324 37148
rect 10376 37136 10382 37188
rect 8573 37111 8631 37117
rect 8573 37108 8585 37111
rect 8444 37080 8585 37108
rect 8444 37068 8450 37080
rect 8573 37077 8585 37080
rect 8619 37077 8631 37111
rect 8573 37071 8631 37077
rect 9309 37111 9367 37117
rect 9309 37077 9321 37111
rect 9355 37077 9367 37111
rect 9309 37071 9367 37077
rect 9674 37068 9680 37120
rect 9732 37068 9738 37120
rect 1104 37018 10120 37040
rect 1104 36966 3010 37018
rect 3062 36966 3074 37018
rect 3126 36966 3138 37018
rect 3190 36966 3202 37018
rect 3254 36966 3266 37018
rect 3318 36966 9010 37018
rect 9062 36966 9074 37018
rect 9126 36966 9138 37018
rect 9190 36966 9202 37018
rect 9254 36966 9266 37018
rect 9318 36966 10120 37018
rect 1104 36944 10120 36966
rect 1578 36864 1584 36916
rect 1636 36904 1642 36916
rect 4246 36904 4252 36916
rect 1636 36876 4252 36904
rect 1636 36864 1642 36876
rect 4246 36864 4252 36876
rect 4304 36864 4310 36916
rect 5534 36864 5540 36916
rect 5592 36904 5598 36916
rect 5813 36907 5871 36913
rect 5813 36904 5825 36907
rect 5592 36876 5825 36904
rect 5592 36864 5598 36876
rect 5813 36873 5825 36876
rect 5859 36873 5871 36907
rect 5813 36867 5871 36873
rect 7193 36907 7251 36913
rect 7193 36873 7205 36907
rect 7239 36904 7251 36907
rect 8662 36904 8668 36916
rect 7239 36876 8668 36904
rect 7239 36873 7251 36876
rect 7193 36867 7251 36873
rect 8662 36864 8668 36876
rect 8720 36864 8726 36916
rect 1762 36796 1768 36848
rect 1820 36796 1826 36848
rect 3602 36796 3608 36848
rect 3660 36836 3666 36848
rect 9306 36836 9312 36848
rect 3660 36808 5764 36836
rect 3660 36796 3666 36808
rect 1780 36768 1808 36796
rect 2041 36771 2099 36777
rect 2041 36768 2053 36771
rect 1780 36740 2053 36768
rect 2041 36737 2053 36740
rect 2087 36737 2099 36771
rect 2041 36731 2099 36737
rect 3973 36771 4031 36777
rect 3973 36737 3985 36771
rect 4019 36768 4031 36771
rect 4338 36768 4344 36780
rect 4019 36740 4344 36768
rect 4019 36737 4031 36740
rect 3973 36731 4031 36737
rect 4338 36728 4344 36740
rect 4396 36728 4402 36780
rect 4522 36777 4528 36780
rect 4516 36731 4528 36777
rect 4522 36728 4528 36731
rect 4580 36728 4586 36780
rect 1670 36660 1676 36712
rect 1728 36700 1734 36712
rect 1765 36703 1823 36709
rect 1765 36700 1777 36703
rect 1728 36672 1777 36700
rect 1728 36660 1734 36672
rect 1765 36669 1777 36672
rect 1811 36669 1823 36703
rect 1765 36663 1823 36669
rect 3694 36660 3700 36712
rect 3752 36700 3758 36712
rect 3878 36700 3884 36712
rect 3752 36672 3884 36700
rect 3752 36660 3758 36672
rect 3878 36660 3884 36672
rect 3936 36660 3942 36712
rect 4246 36660 4252 36712
rect 4304 36660 4310 36712
rect 3418 36592 3424 36644
rect 3476 36632 3482 36644
rect 3476 36604 4292 36632
rect 3476 36592 3482 36604
rect 1578 36524 1584 36576
rect 1636 36564 1642 36576
rect 2038 36564 2044 36576
rect 1636 36536 2044 36564
rect 1636 36524 1642 36536
rect 2038 36524 2044 36536
rect 2096 36524 2102 36576
rect 2777 36567 2835 36573
rect 2777 36533 2789 36567
rect 2823 36564 2835 36567
rect 3694 36564 3700 36576
rect 2823 36536 3700 36564
rect 2823 36533 2835 36536
rect 2777 36527 2835 36533
rect 3694 36524 3700 36536
rect 3752 36524 3758 36576
rect 4062 36524 4068 36576
rect 4120 36564 4126 36576
rect 4157 36567 4215 36573
rect 4157 36564 4169 36567
rect 4120 36536 4169 36564
rect 4120 36524 4126 36536
rect 4157 36533 4169 36536
rect 4203 36533 4215 36567
rect 4264 36564 4292 36604
rect 5629 36567 5687 36573
rect 5629 36564 5641 36567
rect 4264 36536 5641 36564
rect 4157 36527 4215 36533
rect 5629 36533 5641 36536
rect 5675 36533 5687 36567
rect 5736 36564 5764 36808
rect 8864 36808 9312 36836
rect 5997 36771 6055 36777
rect 5997 36737 6009 36771
rect 6043 36768 6055 36771
rect 6914 36768 6920 36780
rect 6043 36740 6920 36768
rect 6043 36737 6055 36740
rect 5997 36731 6055 36737
rect 6914 36728 6920 36740
rect 6972 36728 6978 36780
rect 7834 36728 7840 36780
rect 7892 36728 7898 36780
rect 8864 36777 8892 36808
rect 9306 36796 9312 36808
rect 9364 36796 9370 36848
rect 8849 36771 8907 36777
rect 8849 36737 8861 36771
rect 8895 36737 8907 36771
rect 8849 36731 8907 36737
rect 9122 36728 9128 36780
rect 9180 36728 9186 36780
rect 9493 36771 9551 36777
rect 9493 36737 9505 36771
rect 9539 36737 9551 36771
rect 9493 36731 9551 36737
rect 7650 36660 7656 36712
rect 7708 36700 7714 36712
rect 7975 36703 8033 36709
rect 7975 36700 7987 36703
rect 7708 36672 7987 36700
rect 7708 36660 7714 36672
rect 7975 36669 7987 36672
rect 8021 36669 8033 36703
rect 7975 36663 8033 36669
rect 8110 36660 8116 36712
rect 8168 36660 8174 36712
rect 8386 36660 8392 36712
rect 8444 36660 8450 36712
rect 8754 36660 8760 36712
rect 8812 36700 8818 36712
rect 9033 36703 9091 36709
rect 9033 36700 9045 36703
rect 8812 36672 9045 36700
rect 8812 36660 8818 36672
rect 9033 36669 9045 36672
rect 9079 36669 9091 36703
rect 9508 36700 9536 36731
rect 9033 36663 9091 36669
rect 9140 36672 9536 36700
rect 9140 36564 9168 36672
rect 9309 36635 9367 36641
rect 9309 36601 9321 36635
rect 9355 36632 9367 36635
rect 10502 36632 10508 36644
rect 9355 36604 10508 36632
rect 9355 36601 9367 36604
rect 9309 36595 9367 36601
rect 10502 36592 10508 36604
rect 10560 36592 10566 36644
rect 5736 36536 9168 36564
rect 9677 36567 9735 36573
rect 5629 36527 5687 36533
rect 9677 36533 9689 36567
rect 9723 36564 9735 36567
rect 10410 36564 10416 36576
rect 9723 36536 10416 36564
rect 9723 36533 9735 36536
rect 9677 36527 9735 36533
rect 10410 36524 10416 36536
rect 10468 36524 10474 36576
rect 1104 36474 10120 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 7950 36474
rect 8002 36422 8014 36474
rect 8066 36422 8078 36474
rect 8130 36422 8142 36474
rect 8194 36422 8206 36474
rect 8258 36422 10120 36474
rect 1104 36400 10120 36422
rect 4246 36320 4252 36372
rect 4304 36320 4310 36372
rect 9398 36360 9404 36372
rect 6840 36332 9404 36360
rect 4062 36252 4068 36304
rect 4120 36292 4126 36304
rect 6730 36292 6736 36304
rect 4120 36264 6736 36292
rect 4120 36252 4126 36264
rect 6730 36252 6736 36264
rect 6788 36252 6794 36304
rect 1210 36184 1216 36236
rect 1268 36224 1274 36236
rect 1486 36224 1492 36236
rect 1268 36196 1492 36224
rect 1268 36184 1274 36196
rect 1486 36184 1492 36196
rect 1544 36184 1550 36236
rect 1670 36184 1676 36236
rect 1728 36184 1734 36236
rect 4430 36184 4436 36236
rect 4488 36224 4494 36236
rect 5994 36224 6000 36236
rect 4488 36196 6000 36224
rect 4488 36184 4494 36196
rect 5994 36184 6000 36196
rect 6052 36184 6058 36236
rect 1118 36116 1124 36168
rect 1176 36156 1182 36168
rect 1688 36156 1716 36184
rect 2041 36159 2099 36165
rect 2041 36156 2053 36159
rect 1176 36128 2053 36156
rect 1176 36116 1182 36128
rect 2041 36125 2053 36128
rect 2087 36125 2099 36159
rect 2041 36119 2099 36125
rect 2314 36116 2320 36168
rect 2372 36116 2378 36168
rect 6840 36156 6868 36332
rect 9398 36320 9404 36332
rect 9456 36320 9462 36372
rect 9490 36252 9496 36304
rect 9548 36292 9554 36304
rect 10226 36292 10232 36304
rect 9548 36264 10232 36292
rect 9548 36252 9554 36264
rect 10226 36252 10232 36264
rect 10284 36252 10290 36304
rect 8294 36184 8300 36236
rect 8352 36224 8358 36236
rect 10870 36224 10876 36236
rect 8352 36196 10876 36224
rect 8352 36184 8358 36196
rect 10870 36184 10876 36196
rect 10928 36184 10934 36236
rect 2746 36128 6868 36156
rect 1486 36048 1492 36100
rect 1544 36048 1550 36100
rect 1670 36048 1676 36100
rect 1728 36048 1734 36100
rect 290 35980 296 36032
rect 348 36020 354 36032
rect 2746 36020 2774 36128
rect 7098 36116 7104 36168
rect 7156 36156 7162 36168
rect 7561 36159 7619 36165
rect 7561 36156 7573 36159
rect 7156 36128 7573 36156
rect 7156 36116 7162 36128
rect 7561 36125 7573 36128
rect 7607 36125 7619 36159
rect 7561 36119 7619 36125
rect 7742 36116 7748 36168
rect 7800 36156 7806 36168
rect 7837 36159 7895 36165
rect 7837 36156 7849 36159
rect 7800 36128 7849 36156
rect 7800 36116 7806 36128
rect 7837 36125 7849 36128
rect 7883 36125 7895 36159
rect 7837 36119 7895 36125
rect 8846 36116 8852 36168
rect 8904 36156 8910 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 8904 36128 9137 36156
rect 8904 36116 8910 36128
rect 9125 36125 9137 36128
rect 9171 36125 9183 36159
rect 9125 36119 9183 36125
rect 9493 36159 9551 36165
rect 9493 36125 9505 36159
rect 9539 36125 9551 36159
rect 9493 36119 9551 36125
rect 5537 36091 5595 36097
rect 5537 36057 5549 36091
rect 5583 36057 5595 36091
rect 5537 36051 5595 36057
rect 348 35992 2774 36020
rect 348 35980 354 35992
rect 2866 35980 2872 36032
rect 2924 36020 2930 36032
rect 3053 36023 3111 36029
rect 3053 36020 3065 36023
rect 2924 35992 3065 36020
rect 2924 35980 2930 35992
rect 3053 35989 3065 35992
rect 3099 35989 3111 36023
rect 5552 36020 5580 36051
rect 5626 36048 5632 36100
rect 5684 36088 5690 36100
rect 5721 36091 5779 36097
rect 5721 36088 5733 36091
rect 5684 36060 5733 36088
rect 5684 36048 5690 36060
rect 5721 36057 5733 36060
rect 5767 36057 5779 36091
rect 5721 36051 5779 36057
rect 6178 36048 6184 36100
rect 6236 36088 6242 36100
rect 6236 36060 7144 36088
rect 6236 36048 6242 36060
rect 7009 36023 7067 36029
rect 7009 36020 7021 36023
rect 5552 35992 7021 36020
rect 3053 35983 3111 35989
rect 7009 35989 7021 35992
rect 7055 35989 7067 36023
rect 7116 36020 7144 36060
rect 7466 36048 7472 36100
rect 7524 36048 7530 36100
rect 9508 36088 9536 36119
rect 7576 36060 9536 36088
rect 7576 36020 7604 36060
rect 7116 35992 7604 36020
rect 8573 36023 8631 36029
rect 7009 35983 7067 35989
rect 8573 35989 8585 36023
rect 8619 36020 8631 36023
rect 8846 36020 8852 36032
rect 8619 35992 8852 36020
rect 8619 35989 8631 35992
rect 8573 35983 8631 35989
rect 8846 35980 8852 35992
rect 8904 35980 8910 36032
rect 9309 36023 9367 36029
rect 9309 35989 9321 36023
rect 9355 36020 9367 36023
rect 9582 36020 9588 36032
rect 9355 35992 9588 36020
rect 9355 35989 9367 35992
rect 9309 35983 9367 35989
rect 9582 35980 9588 35992
rect 9640 35980 9646 36032
rect 9677 36023 9735 36029
rect 9677 35989 9689 36023
rect 9723 36020 9735 36023
rect 10134 36020 10140 36032
rect 9723 35992 10140 36020
rect 9723 35989 9735 35992
rect 9677 35983 9735 35989
rect 10134 35980 10140 35992
rect 10192 35980 10198 36032
rect 1104 35930 10120 35952
rect 1104 35878 3010 35930
rect 3062 35878 3074 35930
rect 3126 35878 3138 35930
rect 3190 35878 3202 35930
rect 3254 35878 3266 35930
rect 3318 35878 9010 35930
rect 9062 35878 9074 35930
rect 9126 35878 9138 35930
rect 9190 35878 9202 35930
rect 9254 35878 9266 35930
rect 9318 35878 10120 35930
rect 1104 35856 10120 35878
rect 1949 35819 2007 35825
rect 1949 35785 1961 35819
rect 1995 35816 2007 35819
rect 4154 35816 4160 35828
rect 1995 35788 4160 35816
rect 1995 35785 2007 35788
rect 1949 35779 2007 35785
rect 4154 35776 4160 35788
rect 4212 35776 4218 35828
rect 4338 35776 4344 35828
rect 4396 35776 4402 35828
rect 6549 35819 6607 35825
rect 6549 35785 6561 35819
rect 6595 35816 6607 35819
rect 7006 35816 7012 35828
rect 6595 35788 7012 35816
rect 6595 35785 6607 35788
rect 6549 35779 6607 35785
rect 7006 35776 7012 35788
rect 7064 35776 7070 35828
rect 7653 35819 7711 35825
rect 7653 35785 7665 35819
rect 7699 35816 7711 35819
rect 8386 35816 8392 35828
rect 7699 35788 8392 35816
rect 7699 35785 7711 35788
rect 7653 35779 7711 35785
rect 8386 35776 8392 35788
rect 8444 35776 8450 35828
rect 7742 35748 7748 35760
rect 6932 35720 7748 35748
rect 6932 35692 6960 35720
rect 7742 35708 7748 35720
rect 7800 35708 7806 35760
rect 1486 35640 1492 35692
rect 1544 35640 1550 35692
rect 1762 35640 1768 35692
rect 1820 35640 1826 35692
rect 2225 35683 2283 35689
rect 2225 35649 2237 35683
rect 2271 35680 2283 35683
rect 2314 35680 2320 35692
rect 2271 35652 2320 35680
rect 2271 35649 2283 35652
rect 2225 35643 2283 35649
rect 2314 35640 2320 35652
rect 2372 35640 2378 35692
rect 2498 35640 2504 35692
rect 2556 35680 2562 35692
rect 2556 35652 2820 35680
rect 2556 35640 2562 35652
rect 2792 35624 2820 35652
rect 3694 35640 3700 35692
rect 3752 35640 3758 35692
rect 6365 35683 6423 35689
rect 6365 35649 6377 35683
rect 6411 35680 6423 35683
rect 6914 35680 6920 35692
rect 6411 35652 6920 35680
rect 6411 35649 6423 35652
rect 6365 35643 6423 35649
rect 6914 35640 6920 35652
rect 6972 35640 6978 35692
rect 8294 35640 8300 35692
rect 8352 35640 8358 35692
rect 8570 35640 8576 35692
rect 8628 35640 8634 35692
rect 2682 35572 2688 35624
rect 2740 35572 2746 35624
rect 2774 35572 2780 35624
rect 2832 35572 2838 35624
rect 2866 35572 2872 35624
rect 2924 35612 2930 35624
rect 3145 35615 3203 35621
rect 3145 35612 3157 35615
rect 2924 35584 3157 35612
rect 2924 35572 2930 35584
rect 3145 35581 3157 35584
rect 3191 35581 3203 35615
rect 3145 35575 3203 35581
rect 3418 35572 3424 35624
rect 3476 35572 3482 35624
rect 3510 35572 3516 35624
rect 3568 35621 3574 35624
rect 3568 35615 3617 35621
rect 3568 35581 3571 35615
rect 3605 35612 3617 35615
rect 3878 35612 3884 35624
rect 3605 35584 3884 35612
rect 3605 35581 3617 35584
rect 3568 35575 3617 35581
rect 3568 35572 3574 35575
rect 3878 35572 3884 35584
rect 3936 35572 3942 35624
rect 8478 35621 8484 35624
rect 8456 35615 8484 35621
rect 8456 35581 8468 35615
rect 8456 35575 8484 35581
rect 8478 35572 8484 35575
rect 8536 35572 8542 35624
rect 8846 35572 8852 35624
rect 8904 35572 8910 35624
rect 9306 35572 9312 35624
rect 9364 35572 9370 35624
rect 9398 35572 9404 35624
rect 9456 35612 9462 35624
rect 9493 35615 9551 35621
rect 9493 35612 9505 35615
rect 9456 35584 9505 35612
rect 9456 35572 9462 35584
rect 9493 35581 9505 35584
rect 9539 35581 9551 35615
rect 9493 35575 9551 35581
rect 1673 35547 1731 35553
rect 1673 35513 1685 35547
rect 1719 35544 1731 35547
rect 3234 35544 3240 35556
rect 1719 35516 3240 35544
rect 1719 35513 1731 35516
rect 1673 35507 1731 35513
rect 3234 35504 3240 35516
rect 3292 35504 3298 35556
rect 5074 35504 5080 35556
rect 5132 35544 5138 35556
rect 7006 35544 7012 35556
rect 5132 35516 7012 35544
rect 5132 35504 5138 35516
rect 7006 35504 7012 35516
rect 7064 35504 7070 35556
rect 7466 35504 7472 35556
rect 7524 35544 7530 35556
rect 7834 35544 7840 35556
rect 7524 35516 7840 35544
rect 7524 35504 7530 35516
rect 7834 35504 7840 35516
rect 7892 35504 7898 35556
rect 2409 35479 2467 35485
rect 2409 35445 2421 35479
rect 2455 35476 2467 35479
rect 5902 35476 5908 35488
rect 2455 35448 5908 35476
rect 2455 35445 2467 35448
rect 2409 35439 2467 35445
rect 5902 35436 5908 35448
rect 5960 35436 5966 35488
rect 8202 35436 8208 35488
rect 8260 35476 8266 35488
rect 8478 35476 8484 35488
rect 8260 35448 8484 35476
rect 8260 35436 8266 35448
rect 8478 35436 8484 35448
rect 8536 35436 8542 35488
rect 1104 35386 10120 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 7950 35386
rect 8002 35334 8014 35386
rect 8066 35334 8078 35386
rect 8130 35334 8142 35386
rect 8194 35334 8206 35386
rect 8258 35334 10120 35386
rect 1104 35312 10120 35334
rect 1949 35275 2007 35281
rect 1949 35241 1961 35275
rect 1995 35272 2007 35275
rect 2406 35272 2412 35284
rect 1995 35244 2412 35272
rect 1995 35241 2007 35244
rect 1949 35235 2007 35241
rect 2406 35232 2412 35244
rect 2464 35232 2470 35284
rect 6454 35232 6460 35284
rect 6512 35272 6518 35284
rect 8205 35275 8263 35281
rect 6512 35244 7880 35272
rect 6512 35232 6518 35244
rect 6730 35164 6736 35216
rect 6788 35204 6794 35216
rect 7190 35204 7196 35216
rect 6788 35176 7196 35204
rect 6788 35164 6794 35176
rect 7190 35164 7196 35176
rect 7248 35164 7254 35216
rect 7852 35204 7880 35244
rect 8205 35241 8217 35275
rect 8251 35272 8263 35275
rect 8294 35272 8300 35284
rect 8251 35244 8300 35272
rect 8251 35241 8263 35244
rect 8205 35235 8263 35241
rect 8294 35232 8300 35244
rect 8352 35232 8358 35284
rect 9306 35272 9312 35284
rect 8404 35244 9312 35272
rect 8404 35204 8432 35244
rect 9306 35232 9312 35244
rect 9364 35232 9370 35284
rect 7852 35176 8432 35204
rect 8665 35207 8723 35213
rect 8665 35173 8677 35207
rect 8711 35204 8723 35207
rect 9950 35204 9956 35216
rect 8711 35176 9956 35204
rect 8711 35173 8723 35176
rect 8665 35167 8723 35173
rect 9950 35164 9956 35176
rect 10008 35164 10014 35216
rect 1118 35096 1124 35148
rect 1176 35096 1182 35148
rect 1670 35096 1676 35148
rect 1728 35136 1734 35148
rect 4522 35136 4528 35148
rect 1728 35108 4528 35136
rect 1728 35096 1734 35108
rect 4522 35096 4528 35108
rect 4580 35096 4586 35148
rect 1136 35068 1164 35096
rect 1765 35071 1823 35077
rect 1765 35068 1777 35071
rect 1136 35040 1777 35068
rect 1765 35037 1777 35040
rect 1811 35037 1823 35071
rect 1765 35031 1823 35037
rect 1780 35000 1808 35031
rect 5350 35028 5356 35080
rect 5408 35028 5414 35080
rect 5629 35071 5687 35077
rect 5629 35037 5641 35071
rect 5675 35037 5687 35071
rect 5629 35031 5687 35037
rect 5721 35071 5779 35077
rect 5721 35037 5733 35071
rect 5767 35068 5779 35071
rect 6730 35068 6736 35080
rect 5767 35040 6736 35068
rect 5767 35037 5779 35040
rect 5721 35031 5779 35037
rect 1946 35000 1952 35012
rect 1780 34972 1952 35000
rect 1946 34960 1952 34972
rect 2004 34960 2010 35012
rect 5644 35000 5672 35031
rect 6730 35028 6736 35040
rect 6788 35028 6794 35080
rect 7098 35028 7104 35080
rect 7156 35068 7162 35080
rect 7193 35071 7251 35077
rect 7193 35068 7205 35071
rect 7156 35040 7205 35068
rect 7156 35028 7162 35040
rect 7193 35037 7205 35040
rect 7239 35037 7251 35071
rect 7193 35031 7251 35037
rect 7469 35071 7527 35077
rect 7469 35037 7481 35071
rect 7515 35068 7527 35071
rect 7558 35068 7564 35080
rect 7515 35040 7564 35068
rect 7515 35037 7527 35040
rect 7469 35031 7527 35037
rect 7558 35028 7564 35040
rect 7616 35028 7622 35080
rect 8481 35071 8539 35077
rect 8481 35037 8493 35071
rect 8527 35037 8539 35071
rect 8481 35031 8539 35037
rect 5810 35000 5816 35012
rect 5644 34972 5816 35000
rect 5810 34960 5816 34972
rect 5868 34960 5874 35012
rect 5988 35003 6046 35009
rect 5988 34969 6000 35003
rect 6034 35000 6046 35003
rect 6086 35000 6092 35012
rect 6034 34972 6092 35000
rect 6034 34969 6046 34972
rect 5988 34963 6046 34969
rect 6086 34960 6092 34972
rect 6144 34960 6150 35012
rect 6638 34960 6644 35012
rect 6696 35000 6702 35012
rect 8496 35000 8524 35031
rect 8938 35028 8944 35080
rect 8996 35028 9002 35080
rect 9309 35071 9367 35077
rect 9309 35068 9321 35071
rect 9048 35040 9321 35068
rect 6696 34972 8524 35000
rect 6696 34960 6702 34972
rect 4430 34892 4436 34944
rect 4488 34932 4494 34944
rect 4617 34935 4675 34941
rect 4617 34932 4629 34935
rect 4488 34904 4629 34932
rect 4488 34892 4494 34904
rect 4617 34901 4629 34904
rect 4663 34901 4675 34935
rect 4617 34895 4675 34901
rect 4798 34892 4804 34944
rect 4856 34932 4862 34944
rect 6914 34932 6920 34944
rect 4856 34904 6920 34932
rect 4856 34892 4862 34904
rect 6914 34892 6920 34904
rect 6972 34892 6978 34944
rect 7101 34935 7159 34941
rect 7101 34901 7113 34935
rect 7147 34932 7159 34935
rect 7466 34932 7472 34944
rect 7147 34904 7472 34932
rect 7147 34901 7159 34904
rect 7101 34895 7159 34901
rect 7466 34892 7472 34904
rect 7524 34892 7530 34944
rect 7558 34892 7564 34944
rect 7616 34932 7622 34944
rect 9048 34932 9076 35040
rect 9309 35037 9321 35040
rect 9355 35037 9367 35071
rect 9309 35031 9367 35037
rect 10226 35000 10232 35012
rect 9140 34972 10232 35000
rect 9140 34941 9168 34972
rect 10226 34960 10232 34972
rect 10284 34960 10290 35012
rect 7616 34904 9076 34932
rect 9125 34935 9183 34941
rect 7616 34892 7622 34904
rect 9125 34901 9137 34935
rect 9171 34901 9183 34935
rect 9125 34895 9183 34901
rect 9493 34935 9551 34941
rect 9493 34901 9505 34935
rect 9539 34932 9551 34935
rect 10594 34932 10600 34944
rect 9539 34904 10600 34932
rect 9539 34901 9551 34904
rect 9493 34895 9551 34901
rect 10594 34892 10600 34904
rect 10652 34892 10658 34944
rect 1104 34842 10120 34864
rect 1104 34790 3010 34842
rect 3062 34790 3074 34842
rect 3126 34790 3138 34842
rect 3190 34790 3202 34842
rect 3254 34790 3266 34842
rect 3318 34790 9010 34842
rect 9062 34790 9074 34842
rect 9126 34790 9138 34842
rect 9190 34790 9202 34842
rect 9254 34790 9266 34842
rect 9318 34790 10120 34842
rect 1104 34768 10120 34790
rect 1026 34688 1032 34740
rect 1084 34728 1090 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 1084 34700 1593 34728
rect 1084 34688 1090 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 1581 34691 1639 34697
rect 5166 34688 5172 34740
rect 5224 34688 5230 34740
rect 6546 34688 6552 34740
rect 6604 34688 6610 34740
rect 7742 34688 7748 34740
rect 7800 34728 7806 34740
rect 8662 34728 8668 34740
rect 7800 34700 8668 34728
rect 7800 34688 7806 34700
rect 8662 34688 8668 34700
rect 8720 34688 8726 34740
rect 934 34620 940 34672
rect 992 34660 998 34672
rect 1857 34663 1915 34669
rect 1857 34660 1869 34663
rect 992 34632 1869 34660
rect 992 34620 998 34632
rect 1857 34629 1869 34632
rect 1903 34629 1915 34663
rect 1857 34623 1915 34629
rect 5442 34620 5448 34672
rect 5500 34660 5506 34672
rect 6270 34660 6276 34672
rect 5500 34632 6276 34660
rect 5500 34620 5506 34632
rect 6270 34620 6276 34632
rect 6328 34620 6334 34672
rect 6914 34620 6920 34672
rect 6972 34620 6978 34672
rect 7834 34620 7840 34672
rect 7892 34660 7898 34672
rect 8021 34663 8079 34669
rect 8021 34660 8033 34663
rect 7892 34632 8033 34660
rect 7892 34620 7898 34632
rect 8021 34629 8033 34632
rect 8067 34629 8079 34663
rect 8021 34623 8079 34629
rect 382 34552 388 34604
rect 440 34592 446 34604
rect 1489 34595 1547 34601
rect 1489 34592 1501 34595
rect 440 34564 1501 34592
rect 440 34552 446 34564
rect 1489 34561 1501 34564
rect 1535 34561 1547 34595
rect 1489 34555 1547 34561
rect 2774 34552 2780 34604
rect 2832 34592 2838 34604
rect 3237 34595 3295 34601
rect 3237 34592 3249 34595
rect 2832 34564 3249 34592
rect 2832 34552 2838 34564
rect 3237 34561 3249 34564
rect 3283 34592 3295 34595
rect 4798 34592 4804 34604
rect 3283 34564 4804 34592
rect 3283 34561 3295 34564
rect 3237 34555 3295 34561
rect 4798 34552 4804 34564
rect 4856 34552 4862 34604
rect 5350 34552 5356 34604
rect 5408 34592 5414 34604
rect 5905 34595 5963 34601
rect 5905 34592 5917 34595
rect 5408 34564 5917 34592
rect 5408 34552 5414 34564
rect 5905 34561 5917 34564
rect 5951 34592 5963 34595
rect 6365 34595 6423 34601
rect 6365 34592 6377 34595
rect 5951 34564 6377 34592
rect 5951 34561 5963 34564
rect 5905 34555 5963 34561
rect 6365 34561 6377 34564
rect 6411 34592 6423 34595
rect 6638 34592 6644 34604
rect 6411 34564 6644 34592
rect 6411 34561 6423 34564
rect 6365 34555 6423 34561
rect 6638 34552 6644 34564
rect 6696 34552 6702 34604
rect 6932 34592 6960 34620
rect 7193 34595 7251 34601
rect 7193 34592 7205 34595
rect 6932 34564 7205 34592
rect 7193 34561 7205 34564
rect 7239 34561 7251 34595
rect 7193 34555 7251 34561
rect 2041 34527 2099 34533
rect 2041 34524 2053 34527
rect 1320 34496 2053 34524
rect 1320 34400 1348 34496
rect 2041 34493 2053 34496
rect 2087 34493 2099 34527
rect 2041 34487 2099 34493
rect 2961 34527 3019 34533
rect 2961 34493 2973 34527
rect 3007 34493 3019 34527
rect 2961 34487 3019 34493
rect 5077 34527 5135 34533
rect 5077 34493 5089 34527
rect 5123 34524 5135 34527
rect 5442 34524 5448 34536
rect 5123 34496 5448 34524
rect 5123 34493 5135 34496
rect 5077 34487 5135 34493
rect 1762 34416 1768 34468
rect 1820 34456 1826 34468
rect 1946 34456 1952 34468
rect 1820 34428 1952 34456
rect 1820 34416 1826 34428
rect 1946 34416 1952 34428
rect 2004 34456 2010 34468
rect 2976 34456 3004 34487
rect 5442 34484 5448 34496
rect 5500 34484 5506 34536
rect 6181 34527 6239 34533
rect 6181 34493 6193 34527
rect 6227 34524 6239 34527
rect 6270 34524 6276 34536
rect 6227 34496 6276 34524
rect 6227 34493 6239 34496
rect 6181 34487 6239 34493
rect 6270 34484 6276 34496
rect 6328 34484 6334 34536
rect 6914 34484 6920 34536
rect 6972 34484 6978 34536
rect 9309 34459 9367 34465
rect 9309 34456 9321 34459
rect 2004 34428 3004 34456
rect 7576 34428 9321 34456
rect 2004 34416 2010 34428
rect 1302 34348 1308 34400
rect 1360 34348 1366 34400
rect 3970 34348 3976 34400
rect 4028 34348 4034 34400
rect 4062 34348 4068 34400
rect 4120 34348 4126 34400
rect 4706 34348 4712 34400
rect 4764 34388 4770 34400
rect 6086 34388 6092 34400
rect 4764 34360 6092 34388
rect 4764 34348 4770 34360
rect 6086 34348 6092 34360
rect 6144 34348 6150 34400
rect 6730 34348 6736 34400
rect 6788 34388 6794 34400
rect 7576 34388 7604 34428
rect 9309 34425 9321 34428
rect 9355 34425 9367 34459
rect 9309 34419 9367 34425
rect 6788 34360 7604 34388
rect 6788 34348 6794 34360
rect 7834 34348 7840 34400
rect 7892 34388 7898 34400
rect 7929 34391 7987 34397
rect 7929 34388 7941 34391
rect 7892 34360 7941 34388
rect 7892 34348 7898 34360
rect 7929 34357 7941 34360
rect 7975 34357 7987 34391
rect 7929 34351 7987 34357
rect 1104 34298 10120 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 7950 34298
rect 8002 34246 8014 34298
rect 8066 34246 8078 34298
rect 8130 34246 8142 34298
rect 8194 34246 8206 34298
rect 8258 34246 10120 34298
rect 1104 34224 10120 34246
rect 14 34144 20 34196
rect 72 34184 78 34196
rect 3418 34184 3424 34196
rect 72 34156 3424 34184
rect 72 34144 78 34156
rect 3418 34144 3424 34156
rect 3476 34144 3482 34196
rect 6730 34144 6736 34196
rect 6788 34184 6794 34196
rect 9398 34184 9404 34196
rect 6788 34156 9404 34184
rect 6788 34144 6794 34156
rect 9398 34144 9404 34156
rect 9456 34144 9462 34196
rect 1118 34076 1124 34128
rect 1176 34116 1182 34128
rect 1581 34119 1639 34125
rect 1581 34116 1593 34119
rect 1176 34088 1593 34116
rect 1176 34076 1182 34088
rect 1581 34085 1593 34088
rect 1627 34085 1639 34119
rect 1581 34079 1639 34085
rect 3970 34076 3976 34128
rect 4028 34076 4034 34128
rect 4430 34076 4436 34128
rect 4488 34076 4494 34128
rect 6822 34076 6828 34128
rect 6880 34116 6886 34128
rect 8665 34119 8723 34125
rect 6880 34088 7144 34116
rect 6880 34076 6886 34088
rect 1673 34051 1731 34057
rect 1673 34048 1685 34051
rect 1320 34020 1685 34048
rect 1320 33844 1348 34020
rect 1673 34017 1685 34020
rect 1719 34017 1731 34051
rect 3988 34048 4016 34076
rect 7116 34057 7144 34088
rect 8665 34085 8677 34119
rect 8711 34116 8723 34119
rect 9950 34116 9956 34128
rect 8711 34088 9956 34116
rect 8711 34085 8723 34088
rect 8665 34079 8723 34085
rect 9950 34076 9956 34088
rect 10008 34076 10014 34128
rect 4985 34051 5043 34057
rect 4985 34048 4997 34051
rect 3988 34020 4997 34048
rect 1673 34011 1731 34017
rect 4985 34017 4997 34020
rect 5031 34017 5043 34051
rect 4985 34011 5043 34017
rect 7101 34051 7159 34057
rect 7101 34017 7113 34051
rect 7147 34017 7159 34051
rect 10778 34048 10784 34060
rect 7101 34011 7159 34017
rect 8036 34020 10784 34048
rect 1397 33983 1455 33989
rect 1397 33949 1409 33983
rect 1443 33949 1455 33983
rect 1397 33943 1455 33949
rect 1949 33983 2007 33989
rect 1949 33949 1961 33983
rect 1995 33980 2007 33983
rect 2314 33980 2320 33992
rect 1995 33952 2320 33980
rect 1995 33949 2007 33952
rect 1949 33943 2007 33949
rect 1412 33912 1440 33943
rect 1964 33912 1992 33943
rect 2314 33940 2320 33952
rect 2372 33940 2378 33992
rect 2406 33940 2412 33992
rect 2464 33980 2470 33992
rect 3421 33983 3479 33989
rect 3421 33980 3433 33983
rect 2464 33952 3433 33980
rect 2464 33940 2470 33952
rect 3421 33949 3433 33952
rect 3467 33949 3479 33983
rect 3421 33943 3479 33949
rect 3510 33940 3516 33992
rect 3568 33980 3574 33992
rect 3789 33983 3847 33989
rect 3789 33980 3801 33983
rect 3568 33952 3801 33980
rect 3568 33940 3574 33952
rect 3789 33949 3801 33952
rect 3835 33949 3847 33983
rect 3789 33943 3847 33949
rect 3970 33940 3976 33992
rect 4028 33940 4034 33992
rect 4706 33940 4712 33992
rect 4764 33940 4770 33992
rect 4798 33940 4804 33992
rect 4856 33989 4862 33992
rect 4856 33983 4884 33989
rect 4872 33949 4884 33983
rect 4856 33943 4884 33949
rect 5629 33983 5687 33989
rect 5629 33949 5641 33983
rect 5675 33980 5687 33983
rect 5721 33983 5779 33989
rect 5721 33980 5733 33983
rect 5675 33952 5733 33980
rect 5675 33949 5687 33952
rect 5629 33943 5687 33949
rect 5721 33949 5733 33952
rect 5767 33949 5779 33983
rect 5721 33943 5779 33949
rect 4856 33940 4862 33943
rect 6638 33940 6644 33992
rect 6696 33980 6702 33992
rect 7377 33983 7435 33989
rect 7377 33980 7389 33983
rect 6696 33952 7389 33980
rect 6696 33940 6702 33952
rect 7377 33949 7389 33952
rect 7423 33980 7435 33983
rect 7650 33980 7656 33992
rect 7423 33952 7656 33980
rect 7423 33949 7435 33952
rect 7377 33943 7435 33949
rect 7650 33940 7656 33952
rect 7708 33940 7714 33992
rect 8036 33912 8064 34020
rect 10778 34008 10784 34020
rect 10836 34008 10842 34060
rect 8202 33940 8208 33992
rect 8260 33940 8266 33992
rect 8294 33940 8300 33992
rect 8352 33980 8358 33992
rect 8481 33983 8539 33989
rect 8481 33980 8493 33983
rect 8352 33952 8493 33980
rect 8352 33940 8358 33952
rect 8481 33949 8493 33952
rect 8527 33949 8539 33983
rect 8481 33943 8539 33949
rect 9122 33940 9128 33992
rect 9180 33940 9186 33992
rect 9490 33940 9496 33992
rect 9548 33940 9554 33992
rect 8754 33912 8760 33924
rect 1412 33884 1992 33912
rect 5920 33884 8064 33912
rect 8128 33884 8760 33912
rect 1762 33844 1768 33856
rect 1320 33816 1768 33844
rect 1762 33804 1768 33816
rect 1820 33804 1826 33856
rect 2685 33847 2743 33853
rect 2685 33813 2697 33847
rect 2731 33844 2743 33847
rect 3510 33844 3516 33856
rect 2731 33816 3516 33844
rect 2731 33813 2743 33816
rect 2685 33807 2743 33813
rect 3510 33804 3516 33816
rect 3568 33804 3574 33856
rect 3605 33847 3663 33853
rect 3605 33813 3617 33847
rect 3651 33844 3663 33847
rect 3694 33844 3700 33856
rect 3651 33816 3700 33844
rect 3651 33813 3663 33816
rect 3605 33807 3663 33813
rect 3694 33804 3700 33816
rect 3752 33804 3758 33856
rect 5920 33853 5948 33884
rect 8128 33853 8156 33884
rect 8754 33872 8760 33884
rect 8812 33872 8818 33924
rect 10686 33912 10692 33924
rect 9324 33884 10692 33912
rect 5905 33847 5963 33853
rect 5905 33813 5917 33847
rect 5951 33813 5963 33847
rect 5905 33807 5963 33813
rect 8113 33847 8171 33853
rect 8113 33813 8125 33847
rect 8159 33813 8171 33847
rect 8113 33807 8171 33813
rect 8389 33847 8447 33853
rect 8389 33813 8401 33847
rect 8435 33844 8447 33847
rect 8662 33844 8668 33856
rect 8435 33816 8668 33844
rect 8435 33813 8447 33816
rect 8389 33807 8447 33813
rect 8662 33804 8668 33816
rect 8720 33804 8726 33856
rect 9324 33853 9352 33884
rect 10686 33872 10692 33884
rect 10744 33872 10750 33924
rect 9309 33847 9367 33853
rect 9309 33813 9321 33847
rect 9355 33813 9367 33847
rect 9309 33807 9367 33813
rect 9674 33804 9680 33856
rect 9732 33804 9738 33856
rect 1104 33754 10120 33776
rect 1104 33702 3010 33754
rect 3062 33702 3074 33754
rect 3126 33702 3138 33754
rect 3190 33702 3202 33754
rect 3254 33702 3266 33754
rect 3318 33702 9010 33754
rect 9062 33702 9074 33754
rect 9126 33702 9138 33754
rect 9190 33702 9202 33754
rect 9254 33702 9266 33754
rect 9318 33702 10120 33754
rect 1104 33680 10120 33702
rect 1581 33643 1639 33649
rect 1581 33609 1593 33643
rect 1627 33640 1639 33643
rect 6914 33640 6920 33652
rect 1627 33612 6920 33640
rect 1627 33609 1639 33612
rect 1581 33603 1639 33609
rect 6914 33600 6920 33612
rect 6972 33600 6978 33652
rect 8202 33600 8208 33652
rect 8260 33640 8266 33652
rect 9401 33643 9459 33649
rect 9401 33640 9413 33643
rect 8260 33612 9413 33640
rect 8260 33600 8266 33612
rect 9401 33609 9413 33612
rect 9447 33609 9459 33643
rect 9401 33603 9459 33609
rect 1210 33532 1216 33584
rect 1268 33572 1274 33584
rect 1268 33544 1900 33572
rect 1268 33532 1274 33544
rect 750 33464 756 33516
rect 808 33504 814 33516
rect 1872 33513 1900 33544
rect 2406 33532 2412 33584
rect 2464 33532 2470 33584
rect 1489 33507 1547 33513
rect 1489 33504 1501 33507
rect 808 33476 1501 33504
rect 808 33464 814 33476
rect 1489 33473 1501 33476
rect 1535 33473 1547 33507
rect 1489 33467 1547 33473
rect 1857 33507 1915 33513
rect 1857 33473 1869 33507
rect 1903 33473 1915 33507
rect 1857 33467 1915 33473
rect 8754 33464 8760 33516
rect 8812 33464 8818 33516
rect 1578 33396 1584 33448
rect 1636 33436 1642 33448
rect 2406 33436 2412 33448
rect 1636 33408 2412 33436
rect 1636 33396 1642 33408
rect 2406 33396 2412 33408
rect 2464 33396 2470 33448
rect 3050 33396 3056 33448
rect 3108 33396 3114 33448
rect 3234 33445 3240 33448
rect 3212 33439 3240 33445
rect 3212 33405 3224 33439
rect 3212 33399 3240 33405
rect 3234 33396 3240 33399
rect 3292 33396 3298 33448
rect 3326 33396 3332 33448
rect 3384 33396 3390 33448
rect 3510 33396 3516 33448
rect 3568 33436 3574 33448
rect 3605 33439 3663 33445
rect 3605 33436 3617 33439
rect 3568 33408 3617 33436
rect 3568 33396 3574 33408
rect 3605 33405 3617 33408
rect 3651 33405 3663 33439
rect 3605 33399 3663 33405
rect 4065 33439 4123 33445
rect 4065 33405 4077 33439
rect 4111 33436 4123 33439
rect 4154 33436 4160 33448
rect 4111 33408 4160 33436
rect 4111 33405 4123 33408
rect 4065 33399 4123 33405
rect 4154 33396 4160 33408
rect 4212 33396 4218 33448
rect 4246 33396 4252 33448
rect 4304 33436 4310 33448
rect 4798 33436 4804 33448
rect 4304 33408 4804 33436
rect 4304 33396 4310 33408
rect 4798 33396 4804 33408
rect 4856 33396 4862 33448
rect 7282 33396 7288 33448
rect 7340 33436 7346 33448
rect 7561 33439 7619 33445
rect 7561 33436 7573 33439
rect 7340 33408 7573 33436
rect 7340 33396 7346 33408
rect 7561 33405 7573 33408
rect 7607 33405 7619 33439
rect 7561 33399 7619 33405
rect 7742 33396 7748 33448
rect 7800 33396 7806 33448
rect 7834 33396 7840 33448
rect 7892 33436 7898 33448
rect 8205 33439 8263 33445
rect 8205 33436 8217 33439
rect 7892 33408 8217 33436
rect 7892 33396 7898 33408
rect 8205 33405 8217 33408
rect 8251 33405 8263 33439
rect 8481 33439 8539 33445
rect 8481 33436 8493 33439
rect 8205 33399 8263 33405
rect 8312 33408 8493 33436
rect 1118 33328 1124 33380
rect 1176 33368 1182 33380
rect 1670 33368 1676 33380
rect 1176 33340 1676 33368
rect 1176 33328 1182 33340
rect 1670 33328 1676 33340
rect 1728 33328 1734 33380
rect 2041 33371 2099 33377
rect 2041 33337 2053 33371
rect 2087 33368 2099 33371
rect 4172 33368 4200 33396
rect 6546 33368 6552 33380
rect 2087 33340 2544 33368
rect 4172 33340 6552 33368
rect 2087 33337 2099 33340
rect 2041 33331 2099 33337
rect 2516 33300 2544 33340
rect 6546 33328 6552 33340
rect 6604 33328 6610 33380
rect 7466 33328 7472 33380
rect 7524 33368 7530 33380
rect 8312 33368 8340 33408
rect 8481 33405 8493 33408
rect 8527 33405 8539 33439
rect 8481 33399 8539 33405
rect 8619 33439 8677 33445
rect 8619 33405 8631 33439
rect 8665 33436 8677 33439
rect 9950 33436 9956 33448
rect 8665 33408 9956 33436
rect 8665 33405 8677 33408
rect 8619 33399 8677 33405
rect 9950 33396 9956 33408
rect 10008 33396 10014 33448
rect 7524 33340 8340 33368
rect 7524 33328 7530 33340
rect 2958 33300 2964 33312
rect 2516 33272 2964 33300
rect 2958 33260 2964 33272
rect 3016 33260 3022 33312
rect 3786 33260 3792 33312
rect 3844 33300 3850 33312
rect 4154 33300 4160 33312
rect 3844 33272 4160 33300
rect 3844 33260 3850 33272
rect 4154 33260 4160 33272
rect 4212 33260 4218 33312
rect 8312 33300 8340 33340
rect 9490 33328 9496 33380
rect 9548 33328 9554 33380
rect 10042 33300 10048 33312
rect 8312 33272 10048 33300
rect 10042 33260 10048 33272
rect 10100 33260 10106 33312
rect 1104 33210 10120 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 7950 33210
rect 8002 33158 8014 33210
rect 8066 33158 8078 33210
rect 8130 33158 8142 33210
rect 8194 33158 8206 33210
rect 8258 33158 10120 33210
rect 1104 33136 10120 33158
rect 1581 33099 1639 33105
rect 1581 33065 1593 33099
rect 1627 33096 1639 33099
rect 2685 33099 2743 33105
rect 1627 33068 2360 33096
rect 1627 33065 1639 33068
rect 1581 33059 1639 33065
rect 2332 33028 2360 33068
rect 2685 33065 2697 33099
rect 2731 33096 2743 33099
rect 3050 33096 3056 33108
rect 2731 33068 3056 33096
rect 2731 33065 2743 33068
rect 2685 33059 2743 33065
rect 3050 33056 3056 33068
rect 3108 33056 3114 33108
rect 3234 33056 3240 33108
rect 3292 33096 3298 33108
rect 3970 33096 3976 33108
rect 3292 33068 3976 33096
rect 3292 33056 3298 33068
rect 3970 33056 3976 33068
rect 4028 33096 4034 33108
rect 4430 33096 4436 33108
rect 4028 33068 4436 33096
rect 4028 33056 4034 33068
rect 4430 33056 4436 33068
rect 4488 33056 4494 33108
rect 7098 33096 7104 33108
rect 5920 33068 7104 33096
rect 3602 33028 3608 33040
rect 2332 33000 3608 33028
rect 3602 32988 3608 33000
rect 3660 32988 3666 33040
rect 3786 32988 3792 33040
rect 3844 33028 3850 33040
rect 4338 33028 4344 33040
rect 3844 33000 4344 33028
rect 3844 32988 3850 33000
rect 4338 32988 4344 33000
rect 4396 32988 4402 33040
rect 5920 33028 5948 33068
rect 7098 33056 7104 33068
rect 7156 33056 7162 33108
rect 7466 33056 7472 33108
rect 7524 33096 7530 33108
rect 7524 33068 8800 33096
rect 7524 33056 7530 33068
rect 5828 33000 5948 33028
rect 6825 33031 6883 33037
rect 1302 32920 1308 32972
rect 1360 32960 1366 32972
rect 1578 32960 1584 32972
rect 1360 32932 1584 32960
rect 1360 32920 1366 32932
rect 1578 32920 1584 32932
rect 1636 32920 1642 32972
rect 2958 32920 2964 32972
rect 3016 32960 3022 32972
rect 4798 32960 4804 32972
rect 3016 32932 4804 32960
rect 3016 32920 3022 32932
rect 4798 32920 4804 32932
rect 4856 32960 4862 32972
rect 5828 32969 5856 33000
rect 6825 32997 6837 33031
rect 6871 33028 6883 33031
rect 7561 33031 7619 33037
rect 7561 33028 7573 33031
rect 6871 33000 7573 33028
rect 6871 32997 6883 33000
rect 6825 32991 6883 32997
rect 7561 32997 7573 33000
rect 7607 32997 7619 33031
rect 7561 32991 7619 32997
rect 5813 32963 5871 32969
rect 5813 32960 5825 32963
rect 4856 32932 5825 32960
rect 4856 32920 4862 32932
rect 5813 32929 5825 32932
rect 5859 32929 5871 32963
rect 5813 32923 5871 32929
rect 6546 32920 6552 32972
rect 6604 32960 6610 32972
rect 7650 32960 7656 32972
rect 6604 32932 7656 32960
rect 6604 32920 6610 32932
rect 7650 32920 7656 32932
rect 7708 32960 7714 32972
rect 7837 32963 7895 32969
rect 7837 32960 7849 32963
rect 7708 32932 7849 32960
rect 7708 32920 7714 32932
rect 7837 32929 7849 32932
rect 7883 32929 7895 32963
rect 7837 32923 7895 32929
rect 7975 32963 8033 32969
rect 7975 32929 7987 32963
rect 8021 32960 8033 32963
rect 8772 32960 8800 33068
rect 9309 33031 9367 33037
rect 9309 32997 9321 33031
rect 9355 33028 9367 33031
rect 10226 33028 10232 33040
rect 9355 33000 10232 33028
rect 9355 32997 9367 33000
rect 9309 32991 9367 32997
rect 10226 32988 10232 33000
rect 10284 32988 10290 33040
rect 8021 32932 8733 32960
rect 8772 32932 9536 32960
rect 8021 32929 8033 32932
rect 7975 32923 8033 32929
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1412 32824 1440 32855
rect 1670 32852 1676 32904
rect 1728 32852 1734 32904
rect 1946 32892 1952 32904
rect 1780 32864 1952 32892
rect 1780 32824 1808 32864
rect 1946 32852 1952 32864
rect 2004 32852 2010 32904
rect 6089 32895 6147 32901
rect 6089 32861 6101 32895
rect 6135 32861 6147 32895
rect 6089 32855 6147 32861
rect 1412 32796 1808 32824
rect 6104 32824 6132 32855
rect 6730 32852 6736 32904
rect 6788 32892 6794 32904
rect 6917 32895 6975 32901
rect 6917 32892 6929 32895
rect 6788 32864 6929 32892
rect 6788 32852 6794 32864
rect 6917 32861 6929 32864
rect 6963 32861 6975 32895
rect 6917 32855 6975 32861
rect 7098 32852 7104 32904
rect 7156 32852 7162 32904
rect 8110 32852 8116 32904
rect 8168 32852 8174 32904
rect 8705 32892 8733 32932
rect 8846 32892 8852 32904
rect 8705 32864 8852 32892
rect 6270 32824 6276 32836
rect 6104 32796 6276 32824
rect 6270 32784 6276 32796
rect 6328 32784 6334 32836
rect 8772 32824 8800 32864
rect 8846 32852 8852 32864
rect 8904 32852 8910 32904
rect 9508 32901 9536 32932
rect 9033 32895 9091 32901
rect 9033 32861 9045 32895
rect 9079 32892 9091 32895
rect 9125 32895 9183 32901
rect 9125 32892 9137 32895
rect 9079 32864 9137 32892
rect 9079 32861 9091 32864
rect 9033 32855 9091 32861
rect 9125 32861 9137 32864
rect 9171 32861 9183 32895
rect 9125 32855 9183 32861
rect 9493 32895 9551 32901
rect 9493 32861 9505 32895
rect 9539 32861 9551 32895
rect 9493 32855 9551 32861
rect 11146 32824 11152 32836
rect 8772 32796 11152 32824
rect 11146 32784 11152 32796
rect 11204 32784 11210 32836
rect 658 32716 664 32768
rect 716 32756 722 32768
rect 2774 32756 2780 32768
rect 716 32728 2780 32756
rect 716 32716 722 32728
rect 2774 32716 2780 32728
rect 2832 32716 2838 32768
rect 8202 32716 8208 32768
rect 8260 32756 8266 32768
rect 8757 32759 8815 32765
rect 8757 32756 8769 32759
rect 8260 32728 8769 32756
rect 8260 32716 8266 32728
rect 8757 32725 8769 32728
rect 8803 32725 8815 32759
rect 8757 32719 8815 32725
rect 8846 32716 8852 32768
rect 8904 32756 8910 32768
rect 8941 32759 8999 32765
rect 8941 32756 8953 32759
rect 8904 32728 8953 32756
rect 8904 32716 8910 32728
rect 8941 32725 8953 32728
rect 8987 32725 8999 32759
rect 8941 32719 8999 32725
rect 9677 32759 9735 32765
rect 9677 32725 9689 32759
rect 9723 32756 9735 32759
rect 10410 32756 10416 32768
rect 9723 32728 10416 32756
rect 9723 32725 9735 32728
rect 9677 32719 9735 32725
rect 10410 32716 10416 32728
rect 10468 32716 10474 32768
rect 1104 32666 10120 32688
rect 1104 32614 3010 32666
rect 3062 32614 3074 32666
rect 3126 32614 3138 32666
rect 3190 32614 3202 32666
rect 3254 32614 3266 32666
rect 3318 32614 9010 32666
rect 9062 32614 9074 32666
rect 9126 32614 9138 32666
rect 9190 32614 9202 32666
rect 9254 32614 9266 32666
rect 9318 32614 10120 32666
rect 1104 32592 10120 32614
rect 1670 32512 1676 32564
rect 1728 32552 1734 32564
rect 1946 32552 1952 32564
rect 1728 32524 1952 32552
rect 1728 32512 1734 32524
rect 1946 32512 1952 32524
rect 2004 32512 2010 32564
rect 2866 32512 2872 32564
rect 2924 32552 2930 32564
rect 3418 32552 3424 32564
rect 2924 32524 3424 32552
rect 2924 32512 2930 32524
rect 3418 32512 3424 32524
rect 3476 32512 3482 32564
rect 3602 32512 3608 32564
rect 3660 32552 3666 32564
rect 6181 32555 6239 32561
rect 3660 32524 5396 32552
rect 3660 32512 3666 32524
rect 5368 32484 5396 32524
rect 6181 32521 6193 32555
rect 6227 32552 6239 32555
rect 8110 32552 8116 32564
rect 6227 32524 8116 32552
rect 6227 32521 6239 32524
rect 6181 32515 6239 32521
rect 8110 32512 8116 32524
rect 8168 32512 8174 32564
rect 8665 32555 8723 32561
rect 8220 32524 8524 32552
rect 8220 32484 8248 32524
rect 5368 32456 8248 32484
rect 8386 32444 8392 32496
rect 8444 32444 8450 32496
rect 8496 32484 8524 32524
rect 8665 32521 8677 32555
rect 8711 32552 8723 32555
rect 9858 32552 9864 32564
rect 8711 32524 9864 32552
rect 8711 32521 8723 32524
rect 8665 32515 8723 32521
rect 9858 32512 9864 32524
rect 9916 32512 9922 32564
rect 8496 32456 9536 32484
rect 1486 32376 1492 32428
rect 1544 32376 1550 32428
rect 3421 32419 3479 32425
rect 3421 32416 3433 32419
rect 2746 32388 3433 32416
rect 1762 32240 1768 32292
rect 1820 32280 1826 32292
rect 2746 32280 2774 32388
rect 3421 32385 3433 32388
rect 3467 32385 3479 32419
rect 3421 32379 3479 32385
rect 4338 32376 4344 32428
rect 4396 32416 4402 32428
rect 4893 32419 4951 32425
rect 4893 32416 4905 32419
rect 4396 32388 4905 32416
rect 4396 32376 4402 32388
rect 4893 32385 4905 32388
rect 4939 32385 4951 32419
rect 5445 32419 5503 32425
rect 5445 32416 5457 32419
rect 4893 32379 4951 32385
rect 5000 32388 5457 32416
rect 3234 32308 3240 32360
rect 3292 32348 3298 32360
rect 5000 32348 5028 32388
rect 5445 32385 5457 32388
rect 5491 32385 5503 32419
rect 5445 32379 5503 32385
rect 6546 32376 6552 32428
rect 6604 32416 6610 32428
rect 7101 32419 7159 32425
rect 7101 32416 7113 32419
rect 6604 32388 7113 32416
rect 6604 32376 6610 32388
rect 7101 32385 7113 32388
rect 7147 32385 7159 32419
rect 7101 32379 7159 32385
rect 8202 32376 8208 32428
rect 8260 32376 8266 32428
rect 8404 32416 8432 32444
rect 8481 32419 8539 32425
rect 8481 32416 8493 32419
rect 8404 32388 8493 32416
rect 8481 32385 8493 32388
rect 8527 32385 8539 32419
rect 8481 32379 8539 32385
rect 8757 32419 8815 32425
rect 8757 32385 8769 32419
rect 8803 32385 8815 32419
rect 8757 32379 8815 32385
rect 3292 32320 5028 32348
rect 5169 32351 5227 32357
rect 3292 32308 3298 32320
rect 5169 32317 5181 32351
rect 5215 32317 5227 32351
rect 5169 32311 5227 32317
rect 1820 32252 2774 32280
rect 1820 32240 1826 32252
rect 4798 32240 4804 32292
rect 4856 32280 4862 32292
rect 5184 32280 5212 32311
rect 6822 32308 6828 32360
rect 6880 32308 6886 32360
rect 8386 32308 8392 32360
rect 8444 32348 8450 32360
rect 8772 32348 8800 32379
rect 8938 32376 8944 32428
rect 8996 32416 9002 32428
rect 9508 32425 9536 32456
rect 9125 32419 9183 32425
rect 9125 32416 9137 32419
rect 8996 32388 9137 32416
rect 8996 32376 9002 32388
rect 9125 32385 9137 32388
rect 9171 32385 9183 32419
rect 9125 32379 9183 32385
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32385 9551 32419
rect 9493 32379 9551 32385
rect 8444 32320 8800 32348
rect 8444 32308 8450 32320
rect 4856 32252 5212 32280
rect 7837 32283 7895 32289
rect 4856 32240 4862 32252
rect 7837 32249 7849 32283
rect 7883 32280 7895 32283
rect 8846 32280 8852 32292
rect 7883 32252 8852 32280
rect 7883 32249 7895 32252
rect 7837 32243 7895 32249
rect 8846 32240 8852 32252
rect 8904 32240 8910 32292
rect 8941 32283 8999 32289
rect 8941 32249 8953 32283
rect 8987 32280 8999 32283
rect 10226 32280 10232 32292
rect 8987 32252 10232 32280
rect 8987 32249 8999 32252
rect 8941 32243 8999 32249
rect 10226 32240 10232 32252
rect 10284 32240 10290 32292
rect 1210 32172 1216 32224
rect 1268 32212 1274 32224
rect 1581 32215 1639 32221
rect 1581 32212 1593 32215
rect 1268 32184 1593 32212
rect 1268 32172 1274 32184
rect 1581 32181 1593 32184
rect 1627 32181 1639 32215
rect 1581 32175 1639 32181
rect 2774 32172 2780 32224
rect 2832 32212 2838 32224
rect 3605 32215 3663 32221
rect 3605 32212 3617 32215
rect 2832 32184 3617 32212
rect 2832 32172 2838 32184
rect 3605 32181 3617 32184
rect 3651 32181 3663 32215
rect 3605 32175 3663 32181
rect 3878 32172 3884 32224
rect 3936 32212 3942 32224
rect 4706 32212 4712 32224
rect 3936 32184 4712 32212
rect 3936 32172 3942 32184
rect 4706 32172 4712 32184
rect 4764 32172 4770 32224
rect 5077 32215 5135 32221
rect 5077 32181 5089 32215
rect 5123 32212 5135 32215
rect 6086 32212 6092 32224
rect 5123 32184 6092 32212
rect 5123 32181 5135 32184
rect 5077 32175 5135 32181
rect 6086 32172 6092 32184
rect 6144 32172 6150 32224
rect 6733 32215 6791 32221
rect 6733 32181 6745 32215
rect 6779 32212 6791 32215
rect 8294 32212 8300 32224
rect 6779 32184 8300 32212
rect 6779 32181 6791 32184
rect 6733 32175 6791 32181
rect 8294 32172 8300 32184
rect 8352 32172 8358 32224
rect 8389 32215 8447 32221
rect 8389 32181 8401 32215
rect 8435 32212 8447 32215
rect 9214 32212 9220 32224
rect 8435 32184 9220 32212
rect 8435 32181 8447 32184
rect 8389 32175 8447 32181
rect 9214 32172 9220 32184
rect 9272 32172 9278 32224
rect 9309 32215 9367 32221
rect 9309 32181 9321 32215
rect 9355 32212 9367 32215
rect 9398 32212 9404 32224
rect 9355 32184 9404 32212
rect 9355 32181 9367 32184
rect 9309 32175 9367 32181
rect 9398 32172 9404 32184
rect 9456 32172 9462 32224
rect 9674 32172 9680 32224
rect 9732 32172 9738 32224
rect 1104 32122 10120 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 7950 32122
rect 8002 32070 8014 32122
rect 8066 32070 8078 32122
rect 8130 32070 8142 32122
rect 8194 32070 8206 32122
rect 8258 32070 10120 32122
rect 1104 32048 10120 32070
rect 1762 31968 1768 32020
rect 1820 31968 1826 32020
rect 2498 32008 2504 32020
rect 2056 31980 2504 32008
rect 2056 31940 2084 31980
rect 2498 31968 2504 31980
rect 2556 31968 2562 32020
rect 4338 31968 4344 32020
rect 4396 31968 4402 32020
rect 5626 31968 5632 32020
rect 5684 32008 5690 32020
rect 5684 31980 7972 32008
rect 5684 31968 5690 31980
rect 3878 31940 3884 31952
rect 1688 31912 2084 31940
rect 2884 31912 3884 31940
rect 934 31832 940 31884
rect 992 31872 998 31884
rect 1688 31881 1716 31912
rect 1673 31875 1731 31881
rect 1673 31872 1685 31875
rect 992 31844 1685 31872
rect 992 31832 998 31844
rect 1673 31841 1685 31844
rect 1719 31841 1731 31875
rect 1673 31835 1731 31841
rect 2222 31832 2228 31884
rect 2280 31872 2286 31884
rect 2547 31875 2605 31881
rect 2547 31872 2559 31875
rect 2280 31844 2559 31872
rect 2280 31832 2286 31844
rect 2547 31841 2559 31844
rect 2593 31841 2605 31875
rect 2547 31835 2605 31841
rect 2685 31875 2743 31881
rect 2685 31841 2697 31875
rect 2731 31872 2743 31875
rect 2884 31872 2912 31912
rect 3878 31900 3884 31912
rect 3936 31900 3942 31952
rect 5534 31900 5540 31952
rect 5592 31900 5598 31952
rect 7944 31940 7972 31980
rect 9214 31968 9220 32020
rect 9272 32008 9278 32020
rect 10226 32008 10232 32020
rect 9272 31980 10232 32008
rect 9272 31968 9278 31980
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 9122 31940 9128 31952
rect 7944 31912 9128 31940
rect 9122 31900 9128 31912
rect 9180 31900 9186 31952
rect 9309 31943 9367 31949
rect 9309 31909 9321 31943
rect 9355 31940 9367 31943
rect 9490 31940 9496 31952
rect 9355 31912 9496 31940
rect 9355 31909 9367 31912
rect 9309 31903 9367 31909
rect 9490 31900 9496 31912
rect 9548 31900 9554 31952
rect 9582 31900 9588 31952
rect 9640 31940 9646 31952
rect 9677 31943 9735 31949
rect 9677 31940 9689 31943
rect 9640 31912 9689 31940
rect 9640 31900 9646 31912
rect 9677 31909 9689 31912
rect 9723 31909 9735 31943
rect 9677 31903 9735 31909
rect 2731 31844 2912 31872
rect 2961 31875 3019 31881
rect 2731 31841 2743 31844
rect 2685 31835 2743 31841
rect 2961 31841 2973 31875
rect 3007 31872 3019 31875
rect 3050 31872 3056 31884
rect 3007 31844 3056 31872
rect 3007 31841 3019 31844
rect 2961 31835 3019 31841
rect 3050 31832 3056 31844
rect 3108 31832 3114 31884
rect 4430 31832 4436 31884
rect 4488 31832 4494 31884
rect 4982 31832 4988 31884
rect 5040 31832 5046 31884
rect 5810 31832 5816 31884
rect 5868 31872 5874 31884
rect 6822 31872 6828 31884
rect 5868 31844 6828 31872
rect 5868 31832 5874 31844
rect 6822 31832 6828 31844
rect 6880 31872 6886 31884
rect 7285 31875 7343 31881
rect 7285 31872 7297 31875
rect 6880 31844 7297 31872
rect 6880 31832 6886 31844
rect 7285 31841 7297 31844
rect 7331 31841 7343 31875
rect 7285 31835 7343 31841
rect 842 31764 848 31816
rect 900 31804 906 31816
rect 1489 31807 1547 31813
rect 1489 31804 1501 31807
rect 900 31776 1501 31804
rect 900 31764 906 31776
rect 1489 31773 1501 31776
rect 1535 31773 1547 31807
rect 1489 31767 1547 31773
rect 2406 31764 2412 31816
rect 2464 31764 2470 31816
rect 3421 31807 3479 31813
rect 3421 31773 3433 31807
rect 3467 31773 3479 31807
rect 3421 31767 3479 31773
rect 3436 31736 3464 31767
rect 3510 31764 3516 31816
rect 3568 31804 3574 31816
rect 3605 31807 3663 31813
rect 3605 31804 3617 31807
rect 3568 31776 3617 31804
rect 3568 31764 3574 31776
rect 3605 31773 3617 31776
rect 3651 31804 3663 31807
rect 3878 31804 3884 31816
rect 3651 31776 3884 31804
rect 3651 31773 3663 31776
rect 3605 31767 3663 31773
rect 3878 31764 3884 31776
rect 3936 31764 3942 31816
rect 4448 31736 4476 31832
rect 5074 31764 5080 31816
rect 5132 31813 5138 31816
rect 5132 31807 5181 31813
rect 5132 31773 5135 31807
rect 5169 31773 5181 31807
rect 5132 31767 5181 31773
rect 5132 31764 5138 31767
rect 5258 31764 5264 31816
rect 5316 31764 5322 31816
rect 5994 31764 6000 31816
rect 6052 31764 6058 31816
rect 6181 31807 6239 31813
rect 6181 31804 6193 31807
rect 6104 31776 6193 31804
rect 3436 31708 4568 31736
rect 4540 31680 4568 31708
rect 1670 31628 1676 31680
rect 1728 31668 1734 31680
rect 1946 31668 1952 31680
rect 1728 31640 1952 31668
rect 1728 31628 1734 31640
rect 1946 31628 1952 31640
rect 2004 31628 2010 31680
rect 3234 31628 3240 31680
rect 3292 31668 3298 31680
rect 3510 31668 3516 31680
rect 3292 31640 3516 31668
rect 3292 31628 3298 31640
rect 3510 31628 3516 31640
rect 3568 31628 3574 31680
rect 4522 31628 4528 31680
rect 4580 31668 4586 31680
rect 5258 31668 5264 31680
rect 4580 31640 5264 31668
rect 4580 31628 4586 31640
rect 5258 31628 5264 31640
rect 5316 31628 5322 31680
rect 5442 31628 5448 31680
rect 5500 31668 5506 31680
rect 6104 31668 6132 31776
rect 6181 31773 6193 31776
rect 6227 31773 6239 31807
rect 7561 31807 7619 31813
rect 7561 31804 7573 31807
rect 7539 31776 7573 31804
rect 6181 31767 6239 31773
rect 7561 31773 7573 31776
rect 7607 31773 7619 31807
rect 7561 31767 7619 31773
rect 5500 31640 6132 31668
rect 5500 31628 5506 31640
rect 7190 31628 7196 31680
rect 7248 31668 7254 31680
rect 7576 31668 7604 31767
rect 8570 31764 8576 31816
rect 8628 31764 8634 31816
rect 8662 31764 8668 31816
rect 8720 31804 8726 31816
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 8720 31776 9137 31804
rect 8720 31764 8726 31776
rect 9125 31773 9137 31776
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 9306 31764 9312 31816
rect 9364 31804 9370 31816
rect 9493 31807 9551 31813
rect 9493 31804 9505 31807
rect 9364 31776 9505 31804
rect 9364 31764 9370 31776
rect 9493 31773 9505 31776
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 8110 31696 8116 31748
rect 8168 31736 8174 31748
rect 8938 31736 8944 31748
rect 8168 31708 8944 31736
rect 8168 31696 8174 31708
rect 8938 31696 8944 31708
rect 8996 31696 9002 31748
rect 7248 31640 7604 31668
rect 7248 31628 7254 31640
rect 8294 31628 8300 31680
rect 8352 31628 8358 31680
rect 8754 31628 8760 31680
rect 8812 31628 8818 31680
rect 1104 31578 10120 31600
rect 1104 31526 3010 31578
rect 3062 31526 3074 31578
rect 3126 31526 3138 31578
rect 3190 31526 3202 31578
rect 3254 31526 3266 31578
rect 3318 31526 9010 31578
rect 9062 31526 9074 31578
rect 9126 31526 9138 31578
rect 9190 31526 9202 31578
rect 9254 31526 9266 31578
rect 9318 31526 10120 31578
rect 1104 31504 10120 31526
rect 1486 31424 1492 31476
rect 1544 31424 1550 31476
rect 2501 31467 2559 31473
rect 2501 31433 2513 31467
rect 2547 31464 2559 31467
rect 2866 31464 2872 31476
rect 2547 31436 2872 31464
rect 2547 31433 2559 31436
rect 2501 31427 2559 31433
rect 2866 31424 2872 31436
rect 2924 31424 2930 31476
rect 3513 31467 3571 31473
rect 3513 31433 3525 31467
rect 3559 31464 3571 31467
rect 3602 31464 3608 31476
rect 3559 31436 3608 31464
rect 3559 31433 3571 31436
rect 3513 31427 3571 31433
rect 3602 31424 3608 31436
rect 3660 31424 3666 31476
rect 3697 31467 3755 31473
rect 3697 31433 3709 31467
rect 3743 31464 3755 31467
rect 3743 31436 5396 31464
rect 3743 31433 3755 31436
rect 3697 31427 3755 31433
rect 1504 31396 1532 31424
rect 2038 31396 2044 31408
rect 1504 31368 2044 31396
rect 1302 31288 1308 31340
rect 1360 31328 1366 31340
rect 1489 31331 1547 31337
rect 1489 31328 1501 31331
rect 1360 31300 1501 31328
rect 1360 31288 1366 31300
rect 1489 31297 1501 31300
rect 1535 31328 1547 31331
rect 1670 31328 1676 31340
rect 1535 31300 1676 31328
rect 1535 31297 1547 31300
rect 1489 31291 1547 31297
rect 1670 31288 1676 31300
rect 1728 31288 1734 31340
rect 1780 31337 1808 31368
rect 2038 31356 2044 31368
rect 2096 31356 2102 31408
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31297 1823 31331
rect 1765 31291 1823 31297
rect 3326 31288 3332 31340
rect 3384 31288 3390 31340
rect 4522 31337 4528 31340
rect 4500 31331 4528 31337
rect 4500 31297 4512 31331
rect 4500 31291 4528 31297
rect 4522 31288 4528 31291
rect 4580 31288 4586 31340
rect 5368 31328 5396 31436
rect 5994 31424 6000 31476
rect 6052 31464 6058 31476
rect 8110 31464 8116 31476
rect 6052 31436 8116 31464
rect 6052 31424 6058 31436
rect 8110 31424 8116 31436
rect 8168 31424 8174 31476
rect 8570 31424 8576 31476
rect 8628 31464 8634 31476
rect 9493 31467 9551 31473
rect 9493 31464 9505 31467
rect 8628 31436 9505 31464
rect 8628 31424 8634 31436
rect 9493 31433 9505 31436
rect 9539 31433 9551 31467
rect 9493 31427 9551 31433
rect 6454 31356 6460 31408
rect 6512 31396 6518 31408
rect 6914 31396 6920 31408
rect 6512 31368 6920 31396
rect 6512 31356 6518 31368
rect 6914 31356 6920 31368
rect 6972 31356 6978 31408
rect 5629 31331 5687 31337
rect 5629 31328 5641 31331
rect 5368 31300 5641 31328
rect 5629 31297 5641 31300
rect 5675 31297 5687 31331
rect 5629 31291 5687 31297
rect 7742 31288 7748 31340
rect 7800 31328 7806 31340
rect 7837 31331 7895 31337
rect 7837 31328 7849 31331
rect 7800 31300 7849 31328
rect 7800 31288 7806 31300
rect 7837 31297 7849 31300
rect 7883 31297 7895 31331
rect 7837 31291 7895 31297
rect 8570 31288 8576 31340
rect 8628 31288 8634 31340
rect 8846 31288 8852 31340
rect 8904 31288 8910 31340
rect 9766 31288 9772 31340
rect 9824 31288 9830 31340
rect 3602 31220 3608 31272
rect 3660 31260 3666 31272
rect 4341 31263 4399 31269
rect 4341 31260 4353 31263
rect 3660 31232 4353 31260
rect 3660 31220 3666 31232
rect 4341 31229 4353 31232
rect 4387 31229 4399 31263
rect 4341 31223 4399 31229
rect 4617 31263 4675 31269
rect 4617 31229 4629 31263
rect 4663 31260 4675 31263
rect 4798 31260 4804 31272
rect 4663 31232 4804 31260
rect 4663 31229 4675 31232
rect 4617 31223 4675 31229
rect 4798 31220 4804 31232
rect 4856 31220 4862 31272
rect 5353 31263 5411 31269
rect 5353 31229 5365 31263
rect 5399 31260 5411 31263
rect 5442 31260 5448 31272
rect 5399 31232 5448 31260
rect 5399 31229 5411 31232
rect 5353 31223 5411 31229
rect 5442 31220 5448 31232
rect 5500 31220 5506 31272
rect 5537 31263 5595 31269
rect 5537 31229 5549 31263
rect 5583 31229 5595 31263
rect 5537 31223 5595 31229
rect 4246 31084 4252 31136
rect 4304 31124 4310 31136
rect 4816 31124 4844 31220
rect 4890 31152 4896 31204
rect 4948 31152 4954 31204
rect 5166 31152 5172 31204
rect 5224 31192 5230 31204
rect 5552 31192 5580 31223
rect 7650 31220 7656 31272
rect 7708 31220 7714 31272
rect 8294 31220 8300 31272
rect 8352 31220 8358 31272
rect 8386 31220 8392 31272
rect 8444 31260 8450 31272
rect 8588 31260 8616 31288
rect 8444 31232 8616 31260
rect 8444 31220 8450 31232
rect 8662 31220 8668 31272
rect 8720 31269 8726 31272
rect 8720 31263 8748 31269
rect 8736 31229 8748 31263
rect 8720 31223 8748 31229
rect 8720 31220 8726 31223
rect 9030 31220 9036 31272
rect 9088 31260 9094 31272
rect 9398 31260 9404 31272
rect 9088 31232 9404 31260
rect 9088 31220 9094 31232
rect 9398 31220 9404 31232
rect 9456 31260 9462 31272
rect 10134 31260 10140 31272
rect 9456 31232 10140 31260
rect 9456 31220 9462 31232
rect 10134 31220 10140 31232
rect 10192 31220 10198 31272
rect 5626 31192 5632 31204
rect 5224 31164 5632 31192
rect 5224 31152 5230 31164
rect 5626 31152 5632 31164
rect 5684 31152 5690 31204
rect 4304 31096 4844 31124
rect 4304 31084 4310 31096
rect 5074 31084 5080 31136
rect 5132 31124 5138 31136
rect 5534 31124 5540 31136
rect 5132 31096 5540 31124
rect 5132 31084 5138 31096
rect 5534 31084 5540 31096
rect 5592 31084 5598 31136
rect 5813 31127 5871 31133
rect 5813 31093 5825 31127
rect 5859 31124 5871 31127
rect 8570 31124 8576 31136
rect 5859 31096 8576 31124
rect 5859 31093 5871 31096
rect 5813 31087 5871 31093
rect 8570 31084 8576 31096
rect 8628 31084 8634 31136
rect 8846 31084 8852 31136
rect 8904 31124 8910 31136
rect 9585 31127 9643 31133
rect 9585 31124 9597 31127
rect 8904 31096 9597 31124
rect 8904 31084 8910 31096
rect 9585 31093 9597 31096
rect 9631 31093 9643 31127
rect 9585 31087 9643 31093
rect 1104 31034 10120 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 7950 31034
rect 8002 30982 8014 31034
rect 8066 30982 8078 31034
rect 8130 30982 8142 31034
rect 8194 30982 8206 31034
rect 8258 30982 10120 31034
rect 1104 30960 10120 30982
rect 2406 30880 2412 30932
rect 2464 30920 2470 30932
rect 2501 30923 2559 30929
rect 2501 30920 2513 30923
rect 2464 30892 2513 30920
rect 2464 30880 2470 30892
rect 2501 30889 2513 30892
rect 2547 30889 2559 30923
rect 2501 30883 2559 30889
rect 3602 30880 3608 30932
rect 3660 30880 3666 30932
rect 3973 30923 4031 30929
rect 3973 30889 3985 30923
rect 4019 30920 4031 30923
rect 5994 30920 6000 30932
rect 4019 30892 6000 30920
rect 4019 30889 4031 30892
rect 3973 30883 4031 30889
rect 5994 30880 6000 30892
rect 6052 30880 6058 30932
rect 7558 30880 7564 30932
rect 7616 30920 7622 30932
rect 7653 30923 7711 30929
rect 7653 30920 7665 30923
rect 7616 30892 7665 30920
rect 7616 30880 7622 30892
rect 7653 30889 7665 30892
rect 7699 30889 7711 30923
rect 7653 30883 7711 30889
rect 9309 30923 9367 30929
rect 9309 30889 9321 30923
rect 9355 30920 9367 30923
rect 10226 30920 10232 30932
rect 9355 30892 10232 30920
rect 9355 30889 9367 30892
rect 9309 30883 9367 30889
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 2590 30852 2596 30864
rect 2424 30824 2596 30852
rect 2424 30728 2452 30824
rect 2590 30812 2596 30824
rect 2648 30812 2654 30864
rect 4522 30812 4528 30864
rect 4580 30852 4586 30864
rect 5534 30852 5540 30864
rect 4580 30824 5540 30852
rect 4580 30812 4586 30824
rect 5534 30812 5540 30824
rect 5592 30812 5598 30864
rect 8205 30855 8263 30861
rect 8205 30821 8217 30855
rect 8251 30852 8263 30855
rect 9674 30852 9680 30864
rect 8251 30824 9680 30852
rect 8251 30821 8263 30824
rect 8205 30815 8263 30821
rect 9674 30812 9680 30824
rect 9732 30812 9738 30864
rect 3326 30744 3332 30796
rect 3384 30784 3390 30796
rect 3384 30756 4016 30784
rect 3384 30744 3390 30756
rect 1489 30719 1547 30725
rect 1489 30685 1501 30719
rect 1535 30716 1547 30719
rect 1670 30716 1676 30728
rect 1535 30688 1676 30716
rect 1535 30685 1547 30688
rect 1489 30679 1547 30685
rect 1670 30676 1676 30688
rect 1728 30676 1734 30728
rect 1765 30719 1823 30725
rect 1765 30685 1777 30719
rect 1811 30716 1823 30719
rect 2406 30716 2412 30728
rect 1811 30688 2412 30716
rect 1811 30685 1823 30688
rect 1765 30679 1823 30685
rect 2406 30676 2412 30688
rect 2464 30676 2470 30728
rect 2590 30676 2596 30728
rect 2648 30676 2654 30728
rect 2869 30719 2927 30725
rect 2869 30685 2881 30719
rect 2915 30716 2927 30719
rect 3510 30716 3516 30728
rect 2915 30688 3516 30716
rect 2915 30685 2927 30688
rect 2869 30679 2927 30685
rect 3510 30676 3516 30688
rect 3568 30716 3574 30728
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3568 30688 3801 30716
rect 3568 30676 3574 30688
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3988 30716 4016 30756
rect 6178 30744 6184 30796
rect 6236 30784 6242 30796
rect 6273 30787 6331 30793
rect 6273 30784 6285 30787
rect 6236 30756 6285 30784
rect 6236 30744 6242 30756
rect 6273 30753 6285 30756
rect 6319 30753 6331 30787
rect 6273 30747 6331 30753
rect 8662 30744 8668 30796
rect 8720 30784 8726 30796
rect 8720 30756 9536 30784
rect 8720 30744 8726 30756
rect 4706 30716 4712 30728
rect 3988 30688 4712 30716
rect 3789 30679 3847 30685
rect 4706 30676 4712 30688
rect 4764 30716 4770 30728
rect 6454 30716 6460 30728
rect 4764 30688 6460 30716
rect 4764 30676 4770 30688
rect 6454 30676 6460 30688
rect 6512 30716 6518 30728
rect 6549 30719 6607 30725
rect 6549 30716 6561 30719
rect 6512 30688 6561 30716
rect 6512 30676 6518 30688
rect 6549 30685 6561 30688
rect 6595 30685 6607 30719
rect 6549 30679 6607 30685
rect 7190 30676 7196 30728
rect 7248 30716 7254 30728
rect 7469 30719 7527 30725
rect 7469 30716 7481 30719
rect 7248 30688 7481 30716
rect 7248 30676 7254 30688
rect 7469 30685 7481 30688
rect 7515 30685 7527 30719
rect 7469 30679 7527 30685
rect 8386 30676 8392 30728
rect 8444 30676 8450 30728
rect 8481 30719 8539 30725
rect 8481 30685 8493 30719
rect 8527 30685 8539 30719
rect 8481 30679 8539 30685
rect 6270 30608 6276 30660
rect 6328 30648 6334 30660
rect 8496 30648 8524 30679
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9508 30725 9536 30756
rect 9950 30744 9956 30796
rect 10008 30784 10014 30796
rect 10008 30756 10456 30784
rect 10008 30744 10014 30756
rect 9125 30719 9183 30725
rect 9125 30716 9137 30719
rect 8812 30688 9137 30716
rect 8812 30676 8818 30688
rect 9125 30685 9137 30688
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 9493 30719 9551 30725
rect 9493 30685 9505 30719
rect 9539 30685 9551 30719
rect 9493 30679 9551 30685
rect 9950 30648 9956 30660
rect 6328 30620 8524 30648
rect 8680 30620 9956 30648
rect 6328 30608 6334 30620
rect 2866 30540 2872 30592
rect 2924 30580 2930 30592
rect 5810 30580 5816 30592
rect 2924 30552 5816 30580
rect 2924 30540 2930 30552
rect 5810 30540 5816 30552
rect 5868 30540 5874 30592
rect 7285 30583 7343 30589
rect 7285 30549 7297 30583
rect 7331 30580 7343 30583
rect 8386 30580 8392 30592
rect 7331 30552 8392 30580
rect 7331 30549 7343 30552
rect 7285 30543 7343 30549
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 8680 30589 8708 30620
rect 9950 30608 9956 30620
rect 10008 30608 10014 30660
rect 10042 30608 10048 30660
rect 10100 30648 10106 30660
rect 10318 30648 10324 30660
rect 10100 30620 10324 30648
rect 10100 30608 10106 30620
rect 10318 30608 10324 30620
rect 10376 30608 10382 30660
rect 8665 30583 8723 30589
rect 8665 30549 8677 30583
rect 8711 30549 8723 30583
rect 8665 30543 8723 30549
rect 9306 30540 9312 30592
rect 9364 30580 9370 30592
rect 9490 30580 9496 30592
rect 9364 30552 9496 30580
rect 9364 30540 9370 30552
rect 9490 30540 9496 30552
rect 9548 30540 9554 30592
rect 9582 30540 9588 30592
rect 9640 30580 9646 30592
rect 9677 30583 9735 30589
rect 9677 30580 9689 30583
rect 9640 30552 9689 30580
rect 9640 30540 9646 30552
rect 9677 30549 9689 30552
rect 9723 30549 9735 30583
rect 9677 30543 9735 30549
rect 10134 30540 10140 30592
rect 10192 30580 10198 30592
rect 10428 30580 10456 30756
rect 10192 30552 10456 30580
rect 10192 30540 10198 30552
rect 1104 30490 10120 30512
rect 1104 30438 3010 30490
rect 3062 30438 3074 30490
rect 3126 30438 3138 30490
rect 3190 30438 3202 30490
rect 3254 30438 3266 30490
rect 3318 30438 9010 30490
rect 9062 30438 9074 30490
rect 9126 30438 9138 30490
rect 9190 30438 9202 30490
rect 9254 30438 9266 30490
rect 9318 30438 10120 30490
rect 1104 30416 10120 30438
rect 1486 30336 1492 30388
rect 1544 30376 1550 30388
rect 1544 30348 1624 30376
rect 1544 30336 1550 30348
rect 1486 30200 1492 30252
rect 1544 30200 1550 30252
rect 1596 30172 1624 30348
rect 4522 30336 4528 30388
rect 4580 30376 4586 30388
rect 5074 30376 5080 30388
rect 4580 30348 5080 30376
rect 4580 30336 4586 30348
rect 5074 30336 5080 30348
rect 5132 30336 5138 30388
rect 7742 30336 7748 30388
rect 7800 30376 7806 30388
rect 9214 30376 9220 30388
rect 7800 30348 9220 30376
rect 7800 30336 7806 30348
rect 9214 30336 9220 30348
rect 9272 30336 9278 30388
rect 1673 30311 1731 30317
rect 1673 30277 1685 30311
rect 1719 30308 1731 30311
rect 1762 30308 1768 30320
rect 1719 30280 1768 30308
rect 1719 30277 1731 30280
rect 1673 30271 1731 30277
rect 1762 30268 1768 30280
rect 1820 30268 1826 30320
rect 3326 30268 3332 30320
rect 3384 30268 3390 30320
rect 9033 30311 9091 30317
rect 9033 30277 9045 30311
rect 9079 30308 9091 30311
rect 9766 30308 9772 30320
rect 9079 30280 9772 30308
rect 9079 30277 9091 30280
rect 9033 30271 9091 30277
rect 9766 30268 9772 30280
rect 9824 30268 9830 30320
rect 3145 30243 3203 30249
rect 3145 30209 3157 30243
rect 3191 30240 3203 30243
rect 3344 30240 3372 30268
rect 4706 30240 4712 30252
rect 3191 30212 4712 30240
rect 3191 30209 3203 30212
rect 3145 30203 3203 30209
rect 4706 30200 4712 30212
rect 4764 30200 4770 30252
rect 6365 30243 6423 30249
rect 6365 30209 6377 30243
rect 6411 30240 6423 30243
rect 6454 30240 6460 30252
rect 6411 30212 6460 30240
rect 6411 30209 6423 30212
rect 6365 30203 6423 30209
rect 6454 30200 6460 30212
rect 6512 30200 6518 30252
rect 7098 30200 7104 30252
rect 7156 30240 7162 30252
rect 7377 30243 7435 30249
rect 7377 30240 7389 30243
rect 7156 30212 7389 30240
rect 7156 30200 7162 30212
rect 7377 30209 7389 30212
rect 7423 30209 7435 30243
rect 7377 30203 7435 30209
rect 8110 30200 8116 30252
rect 8168 30200 8174 30252
rect 8386 30200 8392 30252
rect 8444 30200 8450 30252
rect 9125 30243 9183 30249
rect 9125 30209 9137 30243
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 1762 30172 1768 30184
rect 1596 30144 1768 30172
rect 1762 30132 1768 30144
rect 1820 30132 1826 30184
rect 2590 30132 2596 30184
rect 2648 30172 2654 30184
rect 2869 30175 2927 30181
rect 2869 30172 2881 30175
rect 2648 30144 2881 30172
rect 2648 30132 2654 30144
rect 2869 30141 2881 30144
rect 2915 30141 2927 30175
rect 2869 30135 2927 30141
rect 3510 30132 3516 30184
rect 3568 30172 3574 30184
rect 6822 30172 6828 30184
rect 3568 30144 6828 30172
rect 3568 30132 3574 30144
rect 6822 30132 6828 30144
rect 6880 30132 6886 30184
rect 7193 30175 7251 30181
rect 7193 30141 7205 30175
rect 7239 30172 7251 30175
rect 7742 30172 7748 30184
rect 7239 30144 7748 30172
rect 7239 30141 7251 30144
rect 7193 30135 7251 30141
rect 7742 30132 7748 30144
rect 7800 30132 7806 30184
rect 8294 30181 8300 30184
rect 8251 30175 8300 30181
rect 8251 30141 8263 30175
rect 8297 30141 8300 30175
rect 8251 30135 8300 30141
rect 8294 30132 8300 30135
rect 8352 30132 8358 30184
rect 8570 30132 8576 30184
rect 8628 30172 8634 30184
rect 9140 30172 9168 30203
rect 9306 30200 9312 30252
rect 9364 30240 9370 30252
rect 9493 30243 9551 30249
rect 9493 30240 9505 30243
rect 9364 30212 9505 30240
rect 9364 30200 9370 30212
rect 9493 30209 9505 30212
rect 9539 30209 9551 30243
rect 9493 30203 9551 30209
rect 9674 30172 9680 30184
rect 8628 30144 9168 30172
rect 9232 30144 9680 30172
rect 8628 30132 8634 30144
rect 3881 30107 3939 30113
rect 3881 30073 3893 30107
rect 3927 30104 3939 30107
rect 4890 30104 4896 30116
rect 3927 30076 4896 30104
rect 3927 30073 3939 30076
rect 3881 30067 3939 30073
rect 4890 30064 4896 30076
rect 4948 30064 4954 30116
rect 7558 30064 7564 30116
rect 7616 30104 7622 30116
rect 7837 30107 7895 30113
rect 7837 30104 7849 30107
rect 7616 30076 7849 30104
rect 7616 30064 7622 30076
rect 7837 30073 7849 30076
rect 7883 30073 7895 30107
rect 7837 30067 7895 30073
rect 106 29996 112 30048
rect 164 30036 170 30048
rect 1581 30039 1639 30045
rect 1581 30036 1593 30039
rect 164 30008 1593 30036
rect 164 29996 170 30008
rect 1581 30005 1593 30008
rect 1627 30005 1639 30039
rect 1581 29999 1639 30005
rect 1670 29996 1676 30048
rect 1728 30036 1734 30048
rect 3694 30036 3700 30048
rect 1728 30008 3700 30036
rect 1728 29996 1734 30008
rect 3694 29996 3700 30008
rect 3752 29996 3758 30048
rect 6549 30039 6607 30045
rect 6549 30005 6561 30039
rect 6595 30036 6607 30039
rect 9232 30036 9260 30144
rect 9674 30132 9680 30144
rect 9732 30132 9738 30184
rect 9309 30107 9367 30113
rect 9309 30073 9321 30107
rect 9355 30104 9367 30107
rect 10318 30104 10324 30116
rect 9355 30076 10324 30104
rect 9355 30073 9367 30076
rect 9309 30067 9367 30073
rect 10318 30064 10324 30076
rect 10376 30064 10382 30116
rect 6595 30008 9260 30036
rect 9677 30039 9735 30045
rect 6595 30005 6607 30008
rect 6549 29999 6607 30005
rect 9677 30005 9689 30039
rect 9723 30036 9735 30039
rect 10594 30036 10600 30048
rect 9723 30008 10600 30036
rect 9723 30005 9735 30008
rect 9677 29999 9735 30005
rect 10594 29996 10600 30008
rect 10652 29996 10658 30048
rect 1104 29946 10120 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 7950 29946
rect 8002 29894 8014 29946
rect 8066 29894 8078 29946
rect 8130 29894 8142 29946
rect 8194 29894 8206 29946
rect 8258 29894 10120 29946
rect 1104 29872 10120 29894
rect 1581 29835 1639 29841
rect 1581 29801 1593 29835
rect 1627 29832 1639 29835
rect 5350 29832 5356 29844
rect 1627 29804 5356 29832
rect 1627 29801 1639 29804
rect 1581 29795 1639 29801
rect 5350 29792 5356 29804
rect 5408 29792 5414 29844
rect 6454 29792 6460 29844
rect 6512 29792 6518 29844
rect 7190 29792 7196 29844
rect 7248 29832 7254 29844
rect 7466 29832 7472 29844
rect 7248 29804 7472 29832
rect 7248 29792 7254 29804
rect 7466 29792 7472 29804
rect 7524 29792 7530 29844
rect 7558 29792 7564 29844
rect 7616 29792 7622 29844
rect 8941 29835 8999 29841
rect 8941 29832 8953 29835
rect 7852 29804 8953 29832
rect 1394 29724 1400 29776
rect 1452 29764 1458 29776
rect 1765 29767 1823 29773
rect 1765 29764 1777 29767
rect 1452 29736 1777 29764
rect 1452 29724 1458 29736
rect 1765 29733 1777 29736
rect 1811 29733 1823 29767
rect 1765 29727 1823 29733
rect 2222 29724 2228 29776
rect 2280 29764 2286 29776
rect 2406 29764 2412 29776
rect 2280 29736 2412 29764
rect 2280 29724 2286 29736
rect 2406 29724 2412 29736
rect 2464 29724 2470 29776
rect 2682 29724 2688 29776
rect 2740 29764 2746 29776
rect 3418 29764 3424 29776
rect 2740 29736 3424 29764
rect 2740 29724 2746 29736
rect 3418 29724 3424 29736
rect 3476 29724 3482 29776
rect 5166 29656 5172 29708
rect 5224 29696 5230 29708
rect 5261 29699 5319 29705
rect 5261 29696 5273 29699
rect 5224 29668 5273 29696
rect 5224 29656 5230 29668
rect 5261 29665 5273 29668
rect 5307 29665 5319 29699
rect 5261 29659 5319 29665
rect 5350 29656 5356 29708
rect 5408 29696 5414 29708
rect 5813 29699 5871 29705
rect 5813 29696 5825 29699
rect 5408 29668 5825 29696
rect 5408 29656 5414 29668
rect 5813 29665 5825 29668
rect 5859 29665 5871 29699
rect 5813 29659 5871 29665
rect 6178 29656 6184 29708
rect 6236 29696 6242 29708
rect 6549 29699 6607 29705
rect 6549 29696 6561 29699
rect 6236 29668 6561 29696
rect 6236 29656 6242 29668
rect 6549 29665 6561 29668
rect 6595 29665 6607 29699
rect 6549 29659 6607 29665
rect 1394 29588 1400 29640
rect 1452 29588 1458 29640
rect 1949 29631 2007 29637
rect 1949 29597 1961 29631
rect 1995 29628 2007 29631
rect 2590 29628 2596 29640
rect 1995 29600 2596 29628
rect 1995 29597 2007 29600
rect 1949 29591 2007 29597
rect 2590 29588 2596 29600
rect 2648 29588 2654 29640
rect 4617 29631 4675 29637
rect 4617 29597 4629 29631
rect 4663 29628 4675 29631
rect 4706 29628 4712 29640
rect 4663 29600 4712 29628
rect 4663 29597 4675 29600
rect 4617 29591 4675 29597
rect 4706 29588 4712 29600
rect 4764 29588 4770 29640
rect 4801 29631 4859 29637
rect 4801 29597 4813 29631
rect 4847 29597 4859 29631
rect 4801 29591 4859 29597
rect 1578 29452 1584 29504
rect 1636 29492 1642 29504
rect 2314 29492 2320 29504
rect 1636 29464 2320 29492
rect 1636 29452 1642 29464
rect 2314 29452 2320 29464
rect 2372 29452 2378 29504
rect 3602 29452 3608 29504
rect 3660 29492 3666 29504
rect 4062 29492 4068 29504
rect 3660 29464 4068 29492
rect 3660 29452 3666 29464
rect 4062 29452 4068 29464
rect 4120 29452 4126 29504
rect 4816 29492 4844 29591
rect 5534 29588 5540 29640
rect 5592 29588 5598 29640
rect 5626 29588 5632 29640
rect 5684 29637 5690 29640
rect 5684 29631 5712 29637
rect 5700 29597 5712 29631
rect 5684 29591 5712 29597
rect 5684 29588 5690 29591
rect 6822 29588 6828 29640
rect 6880 29588 6886 29640
rect 7852 29637 7880 29804
rect 8941 29801 8953 29804
rect 8987 29801 8999 29835
rect 8941 29795 8999 29801
rect 8018 29724 8024 29776
rect 8076 29724 8082 29776
rect 8297 29767 8355 29773
rect 8297 29733 8309 29767
rect 8343 29764 8355 29767
rect 9766 29764 9772 29776
rect 8343 29736 9772 29764
rect 8343 29733 8355 29736
rect 8297 29727 8355 29733
rect 9766 29724 9772 29736
rect 9824 29724 9830 29776
rect 9398 29696 9404 29708
rect 8036 29668 9404 29696
rect 8036 29640 8064 29668
rect 9398 29656 9404 29668
rect 9456 29656 9462 29708
rect 9490 29656 9496 29708
rect 9548 29656 9554 29708
rect 7837 29631 7895 29637
rect 7837 29597 7849 29631
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 8018 29588 8024 29640
rect 8076 29588 8082 29640
rect 8110 29588 8116 29640
rect 8168 29588 8174 29640
rect 8478 29588 8484 29640
rect 8536 29588 8542 29640
rect 9030 29588 9036 29640
rect 9088 29628 9094 29640
rect 10686 29628 10692 29640
rect 9088 29600 10692 29628
rect 9088 29588 9094 29600
rect 10686 29588 10692 29600
rect 10744 29588 10750 29640
rect 9950 29560 9956 29572
rect 8680 29532 9956 29560
rect 5442 29492 5448 29504
rect 4816 29464 5448 29492
rect 5442 29452 5448 29464
rect 5500 29452 5506 29504
rect 5534 29452 5540 29504
rect 5592 29492 5598 29504
rect 5810 29492 5816 29504
rect 5592 29464 5816 29492
rect 5592 29452 5598 29464
rect 5810 29452 5816 29464
rect 5868 29452 5874 29504
rect 8680 29501 8708 29532
rect 9950 29520 9956 29532
rect 10008 29520 10014 29572
rect 8665 29495 8723 29501
rect 8665 29461 8677 29495
rect 8711 29461 8723 29495
rect 8665 29455 8723 29461
rect 9214 29452 9220 29504
rect 9272 29492 9278 29504
rect 9309 29495 9367 29501
rect 9309 29492 9321 29495
rect 9272 29464 9321 29492
rect 9272 29452 9278 29464
rect 9309 29461 9321 29464
rect 9355 29492 9367 29495
rect 9582 29492 9588 29504
rect 9355 29464 9588 29492
rect 9355 29461 9367 29464
rect 9309 29455 9367 29461
rect 9582 29452 9588 29464
rect 9640 29452 9646 29504
rect 1104 29402 10120 29424
rect 1104 29350 3010 29402
rect 3062 29350 3074 29402
rect 3126 29350 3138 29402
rect 3190 29350 3202 29402
rect 3254 29350 3266 29402
rect 3318 29350 9010 29402
rect 9062 29350 9074 29402
rect 9126 29350 9138 29402
rect 9190 29350 9202 29402
rect 9254 29350 9266 29402
rect 9318 29350 10120 29402
rect 1104 29328 10120 29350
rect 658 29248 664 29300
rect 716 29288 722 29300
rect 1581 29291 1639 29297
rect 1581 29288 1593 29291
rect 716 29260 1593 29288
rect 716 29248 722 29260
rect 1581 29257 1593 29260
rect 1627 29257 1639 29291
rect 1581 29251 1639 29257
rect 2314 29248 2320 29300
rect 2372 29288 2378 29300
rect 2372 29260 2912 29288
rect 2372 29248 2378 29260
rect 1762 29180 1768 29232
rect 1820 29180 1826 29232
rect 382 29112 388 29164
rect 440 29152 446 29164
rect 1397 29155 1455 29161
rect 1397 29152 1409 29155
rect 440 29124 1409 29152
rect 440 29112 446 29124
rect 1397 29121 1409 29124
rect 1443 29121 1455 29155
rect 1780 29152 1808 29180
rect 2041 29155 2099 29161
rect 2041 29152 2053 29155
rect 1780 29124 2053 29152
rect 1397 29115 1455 29121
rect 2041 29121 2053 29124
rect 2087 29152 2099 29155
rect 2884 29152 2912 29260
rect 5166 29248 5172 29300
rect 5224 29248 5230 29300
rect 5276 29260 9168 29288
rect 2958 29180 2964 29232
rect 3016 29220 3022 29232
rect 3510 29220 3516 29232
rect 3016 29192 3516 29220
rect 3016 29180 3022 29192
rect 3510 29180 3516 29192
rect 3568 29180 3574 29232
rect 3602 29180 3608 29232
rect 3660 29220 3666 29232
rect 5276 29220 5304 29260
rect 7190 29220 7196 29232
rect 3660 29192 5304 29220
rect 7024 29192 7196 29220
rect 3660 29180 3666 29192
rect 4433 29155 4491 29161
rect 4433 29152 4445 29155
rect 2087 29124 2820 29152
rect 2884 29124 4445 29152
rect 2087 29121 2099 29124
rect 2041 29115 2099 29121
rect 1762 29044 1768 29096
rect 1820 29044 1826 29096
rect 2792 29084 2820 29124
rect 4433 29121 4445 29124
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 2792 29056 2912 29084
rect 2682 28908 2688 28960
rect 2740 28948 2746 28960
rect 2777 28951 2835 28957
rect 2777 28948 2789 28951
rect 2740 28920 2789 28948
rect 2740 28908 2746 28920
rect 2777 28917 2789 28920
rect 2823 28917 2835 28951
rect 2884 28948 2912 29056
rect 4154 29044 4160 29096
rect 4212 29044 4218 29096
rect 7024 29016 7052 29192
rect 7190 29180 7196 29192
rect 7248 29180 7254 29232
rect 7098 29112 7104 29164
rect 7156 29152 7162 29164
rect 7377 29155 7435 29161
rect 7377 29152 7389 29155
rect 7156 29124 7389 29152
rect 7156 29112 7162 29124
rect 7377 29121 7389 29124
rect 7423 29152 7435 29155
rect 7558 29152 7564 29164
rect 7423 29124 7564 29152
rect 7423 29121 7435 29124
rect 7377 29115 7435 29121
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 8110 29112 8116 29164
rect 8168 29112 8174 29164
rect 9140 29161 9168 29260
rect 9125 29155 9183 29161
rect 9125 29121 9137 29155
rect 9171 29121 9183 29155
rect 9125 29115 9183 29121
rect 9214 29112 9220 29164
rect 9272 29152 9278 29164
rect 9493 29155 9551 29161
rect 9493 29152 9505 29155
rect 9272 29124 9505 29152
rect 9272 29112 9278 29124
rect 9493 29121 9505 29124
rect 9539 29121 9551 29155
rect 9493 29115 9551 29121
rect 9674 29112 9680 29164
rect 9732 29152 9738 29164
rect 9732 29124 9996 29152
rect 9732 29112 9738 29124
rect 9968 29096 9996 29124
rect 7193 29087 7251 29093
rect 7193 29053 7205 29087
rect 7239 29053 7251 29087
rect 7193 29047 7251 29053
rect 7098 29016 7104 29028
rect 7024 28988 7104 29016
rect 7098 28976 7104 28988
rect 7156 28976 7162 29028
rect 7208 29016 7236 29047
rect 7466 29044 7472 29096
rect 7524 29084 7530 29096
rect 8202 29084 8208 29096
rect 8260 29093 8266 29096
rect 8260 29087 8288 29093
rect 7524 29056 8208 29084
rect 7524 29044 7530 29056
rect 8202 29044 8208 29056
rect 8276 29053 8288 29087
rect 8260 29047 8288 29053
rect 8260 29044 8266 29047
rect 8386 29044 8392 29096
rect 8444 29044 8450 29096
rect 8754 29044 8760 29096
rect 8812 29084 8818 29096
rect 9858 29084 9864 29096
rect 8812 29056 9864 29084
rect 8812 29044 8818 29056
rect 9858 29044 9864 29056
rect 9916 29044 9922 29096
rect 9950 29044 9956 29096
rect 10008 29044 10014 29096
rect 7742 29016 7748 29028
rect 7208 28988 7748 29016
rect 7742 28976 7748 28988
rect 7800 28976 7806 29028
rect 7834 28976 7840 29028
rect 7892 28976 7898 29028
rect 9309 29019 9367 29025
rect 9309 28985 9321 29019
rect 9355 29016 9367 29019
rect 9582 29016 9588 29028
rect 9355 28988 9588 29016
rect 9355 28985 9367 28988
rect 9309 28979 9367 28985
rect 9582 28976 9588 28988
rect 9640 28976 9646 29028
rect 9674 28976 9680 29028
rect 9732 28976 9738 29028
rect 4246 28948 4252 28960
rect 2884 28920 4252 28948
rect 2777 28911 2835 28917
rect 4246 28908 4252 28920
rect 4304 28908 4310 28960
rect 4430 28908 4436 28960
rect 4488 28948 4494 28960
rect 5166 28948 5172 28960
rect 4488 28920 5172 28948
rect 4488 28908 4494 28920
rect 5166 28908 5172 28920
rect 5224 28908 5230 28960
rect 7374 28908 7380 28960
rect 7432 28948 7438 28960
rect 7926 28948 7932 28960
rect 7432 28920 7932 28948
rect 7432 28908 7438 28920
rect 7926 28908 7932 28920
rect 7984 28908 7990 28960
rect 8570 28908 8576 28960
rect 8628 28948 8634 28960
rect 9033 28951 9091 28957
rect 9033 28948 9045 28951
rect 8628 28920 9045 28948
rect 8628 28908 8634 28920
rect 9033 28917 9045 28920
rect 9079 28917 9091 28951
rect 9033 28911 9091 28917
rect 1104 28858 10120 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 7950 28858
rect 8002 28806 8014 28858
rect 8066 28806 8078 28858
rect 8130 28806 8142 28858
rect 8194 28806 8206 28858
rect 8258 28806 10120 28858
rect 1104 28784 10120 28806
rect 1394 28704 1400 28756
rect 1452 28744 1458 28756
rect 1581 28747 1639 28753
rect 1581 28744 1593 28747
rect 1452 28716 1593 28744
rect 1452 28704 1458 28716
rect 1581 28713 1593 28716
rect 1627 28713 1639 28747
rect 3234 28744 3240 28756
rect 1581 28707 1639 28713
rect 1872 28716 3240 28744
rect 1210 28636 1216 28688
rect 1268 28676 1274 28688
rect 1872 28676 1900 28716
rect 3234 28704 3240 28716
rect 3292 28704 3298 28756
rect 3602 28704 3608 28756
rect 3660 28704 3666 28756
rect 4798 28744 4804 28756
rect 3712 28716 4804 28744
rect 3712 28676 3740 28716
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 4985 28747 5043 28753
rect 4985 28713 4997 28747
rect 5031 28744 5043 28747
rect 5350 28744 5356 28756
rect 5031 28716 5356 28744
rect 5031 28713 5043 28716
rect 4985 28707 5043 28713
rect 5350 28704 5356 28716
rect 5408 28704 5414 28756
rect 7469 28747 7527 28753
rect 7469 28713 7481 28747
rect 7515 28744 7527 28747
rect 8386 28744 8392 28756
rect 7515 28716 8392 28744
rect 7515 28713 7527 28716
rect 7469 28707 7527 28713
rect 8386 28704 8392 28716
rect 8444 28704 8450 28756
rect 9398 28744 9404 28756
rect 8496 28716 9404 28744
rect 1268 28648 1900 28676
rect 2746 28648 3740 28676
rect 1268 28636 1274 28648
rect 2746 28608 2774 28648
rect 7926 28636 7932 28688
rect 7984 28676 7990 28688
rect 8496 28676 8524 28716
rect 9398 28704 9404 28716
rect 9456 28704 9462 28756
rect 7984 28648 8524 28676
rect 9309 28679 9367 28685
rect 7984 28636 7990 28648
rect 9309 28645 9321 28679
rect 9355 28676 9367 28679
rect 10226 28676 10232 28688
rect 9355 28648 10232 28676
rect 9355 28645 9367 28648
rect 9309 28639 9367 28645
rect 10226 28636 10232 28648
rect 10284 28636 10290 28688
rect 2332 28580 2774 28608
rect 1489 28543 1547 28549
rect 1489 28509 1501 28543
rect 1535 28540 1547 28543
rect 1762 28540 1768 28552
rect 1535 28512 1768 28540
rect 1535 28509 1547 28512
rect 1489 28503 1547 28509
rect 1762 28500 1768 28512
rect 1820 28500 1826 28552
rect 2041 28543 2099 28549
rect 2041 28509 2053 28543
rect 2087 28540 2099 28543
rect 2130 28540 2136 28552
rect 2087 28512 2136 28540
rect 2087 28509 2099 28512
rect 2041 28503 2099 28509
rect 2130 28500 2136 28512
rect 2188 28500 2194 28552
rect 382 28432 388 28484
rect 440 28472 446 28484
rect 2332 28472 2360 28580
rect 3326 28568 3332 28620
rect 3384 28608 3390 28620
rect 3602 28608 3608 28620
rect 3384 28580 3608 28608
rect 3384 28568 3390 28580
rect 3602 28568 3608 28580
rect 3660 28568 3666 28620
rect 5442 28568 5448 28620
rect 5500 28608 5506 28620
rect 5500 28580 6132 28608
rect 5500 28568 5506 28580
rect 3421 28543 3479 28549
rect 3421 28540 3433 28543
rect 440 28444 2360 28472
rect 2562 28512 3433 28540
rect 440 28432 446 28444
rect 2406 28364 2412 28416
rect 2464 28404 2470 28416
rect 2562 28404 2590 28512
rect 3421 28509 3433 28512
rect 3467 28509 3479 28543
rect 3421 28503 3479 28509
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28540 4031 28543
rect 4154 28540 4160 28552
rect 4019 28512 4160 28540
rect 4019 28509 4031 28512
rect 3973 28503 4031 28509
rect 4154 28500 4160 28512
rect 4212 28500 4218 28552
rect 4246 28500 4252 28552
rect 4304 28500 4310 28552
rect 4982 28500 4988 28552
rect 5040 28540 5046 28552
rect 5537 28543 5595 28549
rect 5537 28540 5549 28543
rect 5040 28512 5549 28540
rect 5040 28500 5046 28512
rect 5537 28509 5549 28512
rect 5583 28509 5595 28543
rect 6104 28540 6132 28580
rect 6178 28568 6184 28620
rect 6236 28608 6242 28620
rect 6457 28611 6515 28617
rect 6457 28608 6469 28611
rect 6236 28580 6469 28608
rect 6236 28568 6242 28580
rect 6457 28577 6469 28580
rect 6503 28577 6515 28611
rect 10318 28608 10324 28620
rect 6457 28571 6515 28577
rect 7116 28580 10324 28608
rect 7116 28552 7144 28580
rect 10318 28568 10324 28580
rect 10376 28568 10382 28620
rect 6733 28543 6791 28549
rect 6104 28512 6684 28540
rect 5537 28503 5595 28509
rect 3234 28432 3240 28484
rect 3292 28472 3298 28484
rect 4798 28472 4804 28484
rect 3292 28444 4804 28472
rect 3292 28432 3298 28444
rect 4798 28432 4804 28444
rect 4856 28432 4862 28484
rect 5721 28475 5779 28481
rect 5721 28441 5733 28475
rect 5767 28472 5779 28475
rect 5902 28472 5908 28484
rect 5767 28444 5908 28472
rect 5767 28441 5779 28444
rect 5721 28435 5779 28441
rect 5902 28432 5908 28444
rect 5960 28472 5966 28484
rect 6546 28472 6552 28484
rect 5960 28444 6552 28472
rect 5960 28432 5966 28444
rect 6546 28432 6552 28444
rect 6604 28432 6610 28484
rect 6656 28472 6684 28512
rect 6733 28509 6745 28543
rect 6779 28540 6791 28543
rect 7098 28540 7104 28552
rect 6779 28512 7104 28540
rect 6779 28509 6791 28512
rect 6733 28503 6791 28509
rect 7098 28500 7104 28512
rect 7156 28500 7162 28552
rect 8570 28500 8576 28552
rect 8628 28500 8634 28552
rect 8662 28500 8668 28552
rect 8720 28540 8726 28552
rect 9125 28543 9183 28549
rect 9125 28540 9137 28543
rect 8720 28512 9137 28540
rect 8720 28500 8726 28512
rect 9125 28509 9137 28512
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 9398 28500 9404 28552
rect 9456 28540 9462 28552
rect 9493 28543 9551 28549
rect 9493 28540 9505 28543
rect 9456 28512 9505 28540
rect 9456 28500 9462 28512
rect 9493 28509 9505 28512
rect 9539 28509 9551 28543
rect 9493 28503 9551 28509
rect 11054 28472 11060 28484
rect 6656 28444 11060 28472
rect 11054 28432 11060 28444
rect 11112 28432 11118 28484
rect 2464 28376 2590 28404
rect 2777 28407 2835 28413
rect 2464 28364 2470 28376
rect 2777 28373 2789 28407
rect 2823 28404 2835 28407
rect 3510 28404 3516 28416
rect 2823 28376 3516 28404
rect 2823 28373 2835 28376
rect 2777 28367 2835 28373
rect 3510 28364 3516 28376
rect 3568 28364 3574 28416
rect 4430 28364 4436 28416
rect 4488 28404 4494 28416
rect 5074 28404 5080 28416
rect 4488 28376 5080 28404
rect 4488 28364 4494 28376
rect 5074 28364 5080 28376
rect 5132 28404 5138 28416
rect 5353 28407 5411 28413
rect 5353 28404 5365 28407
rect 5132 28376 5365 28404
rect 5132 28364 5138 28376
rect 5353 28373 5365 28376
rect 5399 28373 5411 28407
rect 5353 28367 5411 28373
rect 5442 28364 5448 28416
rect 5500 28404 5506 28416
rect 5813 28407 5871 28413
rect 5813 28404 5825 28407
rect 5500 28376 5825 28404
rect 5500 28364 5506 28376
rect 5813 28373 5825 28376
rect 5859 28404 5871 28407
rect 6730 28404 6736 28416
rect 5859 28376 6736 28404
rect 5859 28373 5871 28376
rect 5813 28367 5871 28373
rect 6730 28364 6736 28376
rect 6788 28364 6794 28416
rect 8754 28364 8760 28416
rect 8812 28364 8818 28416
rect 9677 28407 9735 28413
rect 9677 28373 9689 28407
rect 9723 28404 9735 28407
rect 10410 28404 10416 28416
rect 9723 28376 10416 28404
rect 9723 28373 9735 28376
rect 9677 28367 9735 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 1104 28314 10120 28336
rect 1104 28262 3010 28314
rect 3062 28262 3074 28314
rect 3126 28262 3138 28314
rect 3190 28262 3202 28314
rect 3254 28262 3266 28314
rect 3318 28262 9010 28314
rect 9062 28262 9074 28314
rect 9126 28262 9138 28314
rect 9190 28262 9202 28314
rect 9254 28262 9266 28314
rect 9318 28262 10120 28314
rect 1104 28240 10120 28262
rect 2406 28160 2412 28212
rect 2464 28160 2470 28212
rect 2608 28172 4108 28200
rect 1762 28092 1768 28144
rect 1820 28132 1826 28144
rect 2608 28132 2636 28172
rect 1820 28104 2636 28132
rect 1820 28092 1826 28104
rect 1394 28024 1400 28076
rect 1452 28024 1458 28076
rect 4080 28064 4108 28172
rect 4154 28160 4160 28212
rect 4212 28160 4218 28212
rect 5810 28160 5816 28212
rect 5868 28200 5874 28212
rect 6822 28200 6828 28212
rect 5868 28172 6828 28200
rect 5868 28160 5874 28172
rect 4172 28132 4200 28160
rect 4798 28132 4804 28144
rect 4172 28104 4804 28132
rect 4798 28092 4804 28104
rect 4856 28132 4862 28144
rect 4856 28104 6040 28132
rect 4856 28092 4862 28104
rect 5442 28064 5448 28076
rect 4080 28036 5448 28064
rect 5442 28024 5448 28036
rect 5500 28024 5506 28076
rect 5721 28067 5779 28073
rect 5721 28033 5733 28067
rect 5767 28064 5779 28067
rect 5810 28064 5816 28076
rect 5767 28036 5816 28064
rect 5767 28033 5779 28036
rect 5721 28027 5779 28033
rect 5810 28024 5816 28036
rect 5868 28024 5874 28076
rect 6012 28073 6040 28104
rect 5997 28067 6055 28073
rect 5997 28033 6009 28067
rect 6043 28033 6055 28067
rect 5997 28027 6055 28033
rect 6178 28024 6184 28076
rect 6236 28064 6242 28076
rect 6748 28073 6776 28172
rect 6822 28160 6828 28172
rect 6880 28160 6886 28212
rect 7469 28203 7527 28209
rect 7469 28169 7481 28203
rect 7515 28200 7527 28203
rect 7834 28200 7840 28212
rect 7515 28172 7840 28200
rect 7515 28169 7527 28172
rect 7469 28163 7527 28169
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 8110 28160 8116 28212
rect 8168 28160 8174 28212
rect 9401 28203 9459 28209
rect 9401 28169 9413 28203
rect 9447 28200 9459 28203
rect 9490 28200 9496 28212
rect 9447 28172 9496 28200
rect 9447 28169 9459 28172
rect 9401 28163 9459 28169
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 6914 28092 6920 28144
rect 6972 28132 6978 28144
rect 6972 28104 8616 28132
rect 6972 28092 6978 28104
rect 8588 28076 8616 28104
rect 6457 28067 6515 28073
rect 6457 28064 6469 28067
rect 6236 28036 6469 28064
rect 6236 28024 6242 28036
rect 6457 28033 6469 28036
rect 6503 28033 6515 28067
rect 6457 28027 6515 28033
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28033 6791 28067
rect 6733 28027 6791 28033
rect 7834 28024 7840 28076
rect 7892 28064 7898 28076
rect 8297 28067 8355 28073
rect 8297 28064 8309 28067
rect 7892 28036 8309 28064
rect 7892 28024 7898 28036
rect 8297 28033 8309 28036
rect 8343 28064 8355 28067
rect 8389 28067 8447 28073
rect 8389 28064 8401 28067
rect 8343 28036 8401 28064
rect 8343 28033 8355 28036
rect 8297 28027 8355 28033
rect 8389 28033 8401 28036
rect 8435 28033 8447 28067
rect 8389 28027 8447 28033
rect 8570 28024 8576 28076
rect 8628 28064 8634 28076
rect 8665 28067 8723 28073
rect 8665 28064 8677 28067
rect 8628 28036 8677 28064
rect 8628 28024 8634 28036
rect 8665 28033 8677 28036
rect 8711 28033 8723 28067
rect 8665 28027 8723 28033
rect 8754 28024 8760 28076
rect 8812 28064 8818 28076
rect 9493 28067 9551 28073
rect 9493 28064 9505 28067
rect 8812 28036 9505 28064
rect 8812 28024 8818 28036
rect 9493 28033 9505 28036
rect 9539 28033 9551 28067
rect 9493 28027 9551 28033
rect 2682 27956 2688 28008
rect 2740 27996 2746 28008
rect 3234 28005 3240 28008
rect 3053 27999 3111 28005
rect 3053 27996 3065 27999
rect 2740 27968 3065 27996
rect 2740 27956 2746 27968
rect 3053 27965 3065 27968
rect 3099 27965 3111 27999
rect 3053 27959 3111 27965
rect 3212 27999 3240 28005
rect 3212 27965 3224 27999
rect 3212 27959 3240 27965
rect 3234 27956 3240 27959
rect 3292 27956 3298 28008
rect 3329 27999 3387 28005
rect 3329 27965 3341 27999
rect 3375 27996 3387 27999
rect 3375 27968 3740 27996
rect 3375 27965 3387 27968
rect 3329 27959 3387 27965
rect 3510 27888 3516 27940
rect 3568 27928 3574 27940
rect 3605 27931 3663 27937
rect 3605 27928 3617 27931
rect 3568 27900 3617 27928
rect 3568 27888 3574 27900
rect 3605 27897 3617 27900
rect 3651 27897 3663 27931
rect 3605 27891 3663 27897
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 1670 27860 1676 27872
rect 1627 27832 1676 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 1670 27820 1676 27832
rect 1728 27820 1734 27872
rect 3050 27820 3056 27872
rect 3108 27860 3114 27872
rect 3712 27860 3740 27968
rect 4062 27956 4068 28008
rect 4120 27956 4126 28008
rect 4246 27956 4252 28008
rect 4304 27956 4310 28008
rect 3108 27832 3740 27860
rect 3108 27820 3114 27832
rect 3878 27820 3884 27872
rect 3936 27860 3942 27872
rect 4985 27863 5043 27869
rect 4985 27860 4997 27863
rect 3936 27832 4997 27860
rect 3936 27820 3942 27832
rect 4985 27829 4997 27832
rect 5031 27829 5043 27863
rect 4985 27823 5043 27829
rect 6822 27820 6828 27872
rect 6880 27860 6886 27872
rect 7926 27860 7932 27872
rect 6880 27832 7932 27860
rect 6880 27820 6886 27832
rect 7926 27820 7932 27832
rect 7984 27820 7990 27872
rect 9674 27820 9680 27872
rect 9732 27820 9738 27872
rect 1104 27770 10120 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 7950 27770
rect 8002 27718 8014 27770
rect 8066 27718 8078 27770
rect 8130 27718 8142 27770
rect 8194 27718 8206 27770
rect 8258 27718 10120 27770
rect 1104 27696 10120 27718
rect 1210 27616 1216 27668
rect 1268 27656 1274 27668
rect 2866 27656 2872 27668
rect 1268 27628 2872 27656
rect 1268 27616 1274 27628
rect 2866 27616 2872 27628
rect 2924 27616 2930 27668
rect 3234 27616 3240 27668
rect 3292 27656 3298 27668
rect 3786 27656 3792 27668
rect 3292 27628 3792 27656
rect 3292 27616 3298 27628
rect 3786 27616 3792 27628
rect 3844 27616 3850 27668
rect 4433 27659 4491 27665
rect 4433 27625 4445 27659
rect 4479 27656 4491 27659
rect 4479 27628 5488 27656
rect 4479 27625 4491 27628
rect 4433 27619 4491 27625
rect 4430 27520 4436 27532
rect 2700 27492 4436 27520
rect 2222 27412 2228 27464
rect 2280 27452 2286 27464
rect 2317 27455 2375 27461
rect 2317 27452 2329 27455
rect 2280 27424 2329 27452
rect 2280 27412 2286 27424
rect 2317 27421 2329 27424
rect 2363 27421 2375 27455
rect 2317 27415 2375 27421
rect 2590 27412 2596 27464
rect 2648 27452 2654 27464
rect 2700 27452 2728 27492
rect 4430 27480 4436 27492
rect 4488 27480 4494 27532
rect 5460 27520 5488 27628
rect 5534 27616 5540 27668
rect 5592 27656 5598 27668
rect 5810 27656 5816 27668
rect 5592 27628 5816 27656
rect 5592 27616 5598 27628
rect 5810 27616 5816 27628
rect 5868 27616 5874 27668
rect 5994 27616 6000 27668
rect 6052 27656 6058 27668
rect 8386 27656 8392 27668
rect 6052 27628 8392 27656
rect 6052 27616 6058 27628
rect 8386 27616 8392 27628
rect 8444 27616 8450 27668
rect 8754 27548 8760 27600
rect 8812 27548 8818 27600
rect 9309 27591 9367 27597
rect 9309 27557 9321 27591
rect 9355 27588 9367 27591
rect 10226 27588 10232 27600
rect 9355 27560 10232 27588
rect 9355 27557 9367 27560
rect 9309 27551 9367 27557
rect 10226 27548 10232 27560
rect 10284 27548 10290 27600
rect 5460 27492 9536 27520
rect 2648 27424 2728 27452
rect 2648 27412 2654 27424
rect 3510 27412 3516 27464
rect 3568 27452 3574 27464
rect 4249 27455 4307 27461
rect 4249 27452 4261 27455
rect 3568 27424 4261 27452
rect 3568 27412 3574 27424
rect 4249 27421 4261 27424
rect 4295 27421 4307 27455
rect 4249 27415 4307 27421
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27421 4583 27455
rect 4525 27415 4583 27421
rect 4801 27455 4859 27461
rect 4801 27421 4813 27455
rect 4847 27452 4859 27455
rect 4890 27452 4896 27464
rect 4847 27424 4896 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 4540 27328 4568 27415
rect 4890 27412 4896 27424
rect 4948 27412 4954 27464
rect 5074 27412 5080 27464
rect 5132 27452 5138 27464
rect 7006 27452 7012 27464
rect 5132 27424 7012 27452
rect 5132 27412 5138 27424
rect 7006 27412 7012 27424
rect 7064 27452 7070 27464
rect 7834 27452 7840 27464
rect 7064 27424 7840 27452
rect 7064 27412 7070 27424
rect 7834 27412 7840 27424
rect 7892 27452 7898 27464
rect 8297 27455 8355 27461
rect 8297 27452 8309 27455
rect 7892 27424 8309 27452
rect 7892 27412 7898 27424
rect 8297 27421 8309 27424
rect 8343 27421 8355 27455
rect 8297 27415 8355 27421
rect 8570 27412 8576 27464
rect 8628 27412 8634 27464
rect 9122 27412 9128 27464
rect 9180 27412 9186 27464
rect 9508 27461 9536 27492
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 10134 27412 10140 27464
rect 10192 27452 10198 27464
rect 10594 27452 10600 27464
rect 10192 27424 10600 27452
rect 10192 27412 10198 27424
rect 10594 27412 10600 27424
rect 10652 27412 10658 27464
rect 7098 27344 7104 27396
rect 7156 27384 7162 27396
rect 8113 27387 8171 27393
rect 8113 27384 8125 27387
rect 7156 27356 8125 27384
rect 7156 27344 7162 27356
rect 8113 27353 8125 27356
rect 8159 27353 8171 27387
rect 8113 27347 8171 27353
rect 8662 27344 8668 27396
rect 8720 27384 8726 27396
rect 10962 27384 10968 27396
rect 8720 27356 10968 27384
rect 8720 27344 8726 27356
rect 10962 27344 10968 27356
rect 11020 27344 11026 27396
rect 842 27276 848 27328
rect 900 27316 906 27328
rect 1581 27319 1639 27325
rect 1581 27316 1593 27319
rect 900 27288 1593 27316
rect 900 27276 906 27288
rect 1581 27285 1593 27288
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 2038 27276 2044 27328
rect 2096 27316 2102 27328
rect 4338 27316 4344 27328
rect 2096 27288 4344 27316
rect 2096 27276 2102 27288
rect 4338 27276 4344 27288
rect 4396 27276 4402 27328
rect 4522 27276 4528 27328
rect 4580 27276 4586 27328
rect 4890 27276 4896 27328
rect 4948 27316 4954 27328
rect 5442 27316 5448 27328
rect 4948 27288 5448 27316
rect 4948 27276 4954 27288
rect 5442 27276 5448 27288
rect 5500 27276 5506 27328
rect 5537 27319 5595 27325
rect 5537 27285 5549 27319
rect 5583 27316 5595 27319
rect 6270 27316 6276 27328
rect 5583 27288 6276 27316
rect 5583 27285 5595 27288
rect 5537 27279 5595 27285
rect 6270 27276 6276 27288
rect 6328 27276 6334 27328
rect 6914 27276 6920 27328
rect 6972 27316 6978 27328
rect 9490 27316 9496 27328
rect 6972 27288 9496 27316
rect 6972 27276 6978 27288
rect 9490 27276 9496 27288
rect 9548 27276 9554 27328
rect 9677 27319 9735 27325
rect 9677 27285 9689 27319
rect 9723 27316 9735 27319
rect 10778 27316 10784 27328
rect 9723 27288 10784 27316
rect 9723 27285 9735 27288
rect 9677 27279 9735 27285
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 1104 27226 10120 27248
rect 1104 27174 3010 27226
rect 3062 27174 3074 27226
rect 3126 27174 3138 27226
rect 3190 27174 3202 27226
rect 3254 27174 3266 27226
rect 3318 27174 9010 27226
rect 9062 27174 9074 27226
rect 9126 27174 9138 27226
rect 9190 27174 9202 27226
rect 9254 27174 9266 27226
rect 9318 27174 10120 27226
rect 1104 27152 10120 27174
rect 2038 27112 2044 27124
rect 1412 27084 2044 27112
rect 1412 27044 1440 27084
rect 2038 27072 2044 27084
rect 2096 27072 2102 27124
rect 2961 27115 3019 27121
rect 2961 27081 2973 27115
rect 3007 27112 3019 27115
rect 3510 27112 3516 27124
rect 3007 27084 3516 27112
rect 3007 27081 3019 27084
rect 2961 27075 3019 27081
rect 3510 27072 3516 27084
rect 3568 27072 3574 27124
rect 3786 27072 3792 27124
rect 3844 27112 3850 27124
rect 4062 27112 4068 27124
rect 3844 27084 4068 27112
rect 3844 27072 3850 27084
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4614 27072 4620 27124
rect 4672 27112 4678 27124
rect 4672 27084 5396 27112
rect 4672 27072 4678 27084
rect 1320 27016 1440 27044
rect 1320 26772 1348 27016
rect 1486 27004 1492 27056
rect 1544 27044 1550 27056
rect 1946 27044 1952 27056
rect 1544 27016 1952 27044
rect 1544 27004 1550 27016
rect 1946 27004 1952 27016
rect 2004 27004 2010 27056
rect 2314 27004 2320 27056
rect 2372 27044 2378 27056
rect 2498 27044 2504 27056
rect 2372 27016 2504 27044
rect 2372 27004 2378 27016
rect 2498 27004 2504 27016
rect 2556 27004 2562 27056
rect 5258 27044 5264 27056
rect 4816 27016 5264 27044
rect 1394 26936 1400 26988
rect 1452 26936 1458 26988
rect 1670 26936 1676 26988
rect 1728 26976 1734 26988
rect 2133 26979 2191 26985
rect 2133 26976 2145 26979
rect 1728 26948 2145 26976
rect 1728 26936 1734 26948
rect 2133 26945 2145 26948
rect 2179 26976 2191 26979
rect 2222 26976 2228 26988
rect 2179 26948 2228 26976
rect 2179 26945 2191 26948
rect 2133 26939 2191 26945
rect 2222 26936 2228 26948
rect 2280 26936 2286 26988
rect 4816 26985 4844 27016
rect 5258 27004 5264 27016
rect 5316 27004 5322 27056
rect 4801 26979 4859 26985
rect 4801 26945 4813 26979
rect 4847 26945 4859 26979
rect 4801 26939 4859 26945
rect 5166 26936 5172 26988
rect 5224 26976 5230 26988
rect 5368 26976 5396 27084
rect 6454 27072 6460 27124
rect 6512 27112 6518 27124
rect 7834 27112 7840 27124
rect 6512 27084 7840 27112
rect 6512 27072 6518 27084
rect 7834 27072 7840 27084
rect 7892 27072 7898 27124
rect 9309 27115 9367 27121
rect 9309 27081 9321 27115
rect 9355 27112 9367 27115
rect 10318 27112 10324 27124
rect 9355 27084 10324 27112
rect 9355 27081 9367 27084
rect 9309 27075 9367 27081
rect 10318 27072 10324 27084
rect 10376 27072 10382 27124
rect 10502 27044 10508 27056
rect 8772 27016 10508 27044
rect 5224 26948 5396 26976
rect 6733 26979 6791 26985
rect 5224 26936 5230 26948
rect 6733 26945 6745 26979
rect 6779 26976 6791 26979
rect 6914 26976 6920 26988
rect 6779 26948 6920 26976
rect 6779 26945 6791 26948
rect 6733 26939 6791 26945
rect 6914 26936 6920 26948
rect 6972 26936 6978 26988
rect 8772 26985 8800 27016
rect 10502 27004 10508 27016
rect 10560 27004 10566 27056
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26945 8539 26979
rect 8481 26939 8539 26945
rect 8757 26979 8815 26985
rect 8757 26945 8769 26979
rect 8803 26945 8815 26979
rect 8757 26939 8815 26945
rect 9125 26979 9183 26985
rect 9125 26945 9137 26979
rect 9171 26976 9183 26979
rect 9398 26976 9404 26988
rect 9171 26948 9404 26976
rect 9171 26945 9183 26948
rect 9125 26939 9183 26945
rect 1762 26868 1768 26920
rect 1820 26908 1826 26920
rect 1857 26911 1915 26917
rect 1857 26908 1869 26911
rect 1820 26880 1869 26908
rect 1820 26868 1826 26880
rect 1857 26877 1869 26880
rect 1903 26877 1915 26911
rect 1857 26871 1915 26877
rect 3234 26868 3240 26920
rect 3292 26908 3298 26920
rect 3786 26917 3792 26920
rect 3605 26911 3663 26917
rect 3605 26908 3617 26911
rect 3292 26880 3617 26908
rect 3292 26868 3298 26880
rect 3605 26877 3617 26880
rect 3651 26877 3663 26911
rect 3605 26871 3663 26877
rect 3764 26911 3792 26917
rect 3764 26877 3776 26911
rect 3764 26871 3792 26877
rect 3786 26868 3792 26871
rect 3844 26868 3850 26920
rect 3881 26911 3939 26917
rect 3881 26877 3893 26911
rect 3927 26908 3939 26911
rect 4430 26908 4436 26920
rect 3927 26880 4436 26908
rect 3927 26877 3939 26880
rect 3881 26871 3939 26877
rect 4430 26868 4436 26880
rect 4488 26868 4494 26920
rect 4614 26868 4620 26920
rect 4672 26868 4678 26920
rect 4890 26868 4896 26920
rect 4948 26868 4954 26920
rect 2869 26843 2927 26849
rect 2869 26809 2881 26843
rect 2915 26840 2927 26843
rect 4157 26843 4215 26849
rect 2915 26812 3280 26840
rect 2915 26809 2927 26812
rect 2869 26803 2927 26809
rect 1044 26744 1348 26772
rect 1581 26775 1639 26781
rect 1044 26568 1072 26744
rect 1581 26741 1593 26775
rect 1627 26772 1639 26775
rect 2774 26772 2780 26784
rect 1627 26744 2780 26772
rect 1627 26741 1639 26744
rect 1581 26735 1639 26741
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 3252 26772 3280 26812
rect 4157 26809 4169 26843
rect 4203 26809 4215 26843
rect 4157 26803 4215 26809
rect 4172 26772 4200 26803
rect 6454 26800 6460 26852
rect 6512 26840 6518 26852
rect 8496 26840 8524 26939
rect 9398 26936 9404 26948
rect 9456 26936 9462 26988
rect 9490 26936 9496 26988
rect 9548 26936 9554 26988
rect 9766 26908 9772 26920
rect 8680 26880 9772 26908
rect 8680 26849 8708 26880
rect 9766 26868 9772 26880
rect 9824 26868 9830 26920
rect 10042 26868 10048 26920
rect 10100 26908 10106 26920
rect 10502 26908 10508 26920
rect 10100 26880 10508 26908
rect 10100 26868 10106 26880
rect 10502 26868 10508 26880
rect 10560 26868 10566 26920
rect 6512 26812 8524 26840
rect 8665 26843 8723 26849
rect 6512 26800 6518 26812
rect 8665 26809 8677 26843
rect 8711 26809 8723 26843
rect 8665 26803 8723 26809
rect 8941 26843 8999 26849
rect 8941 26809 8953 26843
rect 8987 26840 8999 26843
rect 9306 26840 9312 26852
rect 8987 26812 9312 26840
rect 8987 26809 8999 26812
rect 8941 26803 8999 26809
rect 9306 26800 9312 26812
rect 9364 26800 9370 26852
rect 3252 26744 4200 26772
rect 5350 26732 5356 26784
rect 5408 26772 5414 26784
rect 5718 26772 5724 26784
rect 5408 26744 5724 26772
rect 5408 26732 5414 26744
rect 5718 26732 5724 26744
rect 5776 26732 5782 26784
rect 5810 26732 5816 26784
rect 5868 26772 5874 26784
rect 5905 26775 5963 26781
rect 5905 26772 5917 26775
rect 5868 26744 5917 26772
rect 5868 26732 5874 26744
rect 5905 26741 5917 26744
rect 5951 26741 5963 26775
rect 5905 26735 5963 26741
rect 6917 26775 6975 26781
rect 6917 26741 6929 26775
rect 6963 26772 6975 26775
rect 8754 26772 8760 26784
rect 6963 26744 8760 26772
rect 6963 26741 6975 26744
rect 6917 26735 6975 26741
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 9674 26732 9680 26784
rect 9732 26732 9738 26784
rect 1104 26682 10120 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 7950 26682
rect 8002 26630 8014 26682
rect 8066 26630 8078 26682
rect 8130 26630 8142 26682
rect 8194 26630 8206 26682
rect 8258 26630 10120 26682
rect 1104 26608 10120 26630
rect 1581 26571 1639 26577
rect 1581 26568 1593 26571
rect 1044 26540 1593 26568
rect 1581 26537 1593 26540
rect 1627 26537 1639 26571
rect 1581 26531 1639 26537
rect 3234 26528 3240 26580
rect 3292 26528 3298 26580
rect 3694 26528 3700 26580
rect 3752 26568 3758 26580
rect 4617 26571 4675 26577
rect 4617 26568 4629 26571
rect 3752 26540 4629 26568
rect 3752 26528 3758 26540
rect 4617 26537 4629 26540
rect 4663 26568 4675 26571
rect 4890 26568 4896 26580
rect 4663 26540 4896 26568
rect 4663 26537 4675 26540
rect 4617 26531 4675 26537
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 5074 26528 5080 26580
rect 5132 26568 5138 26580
rect 5132 26540 6684 26568
rect 5132 26528 5138 26540
rect 5626 26460 5632 26512
rect 5684 26500 5690 26512
rect 5721 26503 5779 26509
rect 5721 26500 5733 26503
rect 5684 26472 5733 26500
rect 5684 26460 5690 26472
rect 5721 26469 5733 26472
rect 5767 26469 5779 26503
rect 6656 26500 6684 26540
rect 6914 26528 6920 26580
rect 6972 26528 6978 26580
rect 9582 26528 9588 26580
rect 9640 26568 9646 26580
rect 9677 26571 9735 26577
rect 9677 26568 9689 26571
rect 9640 26540 9689 26568
rect 9640 26528 9646 26540
rect 9677 26537 9689 26540
rect 9723 26537 9735 26571
rect 9677 26531 9735 26537
rect 8205 26503 8263 26509
rect 6656 26472 6960 26500
rect 5721 26463 5779 26469
rect 4890 26392 4896 26444
rect 4948 26432 4954 26444
rect 5077 26435 5135 26441
rect 5077 26432 5089 26435
rect 4948 26404 5089 26432
rect 4948 26392 4954 26404
rect 5077 26401 5089 26404
rect 5123 26401 5135 26435
rect 5077 26395 5135 26401
rect 6270 26392 6276 26444
rect 6328 26392 6334 26444
rect 658 26324 664 26376
rect 716 26364 722 26376
rect 1397 26367 1455 26373
rect 1397 26364 1409 26367
rect 716 26336 1409 26364
rect 716 26324 722 26336
rect 1397 26333 1409 26336
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 1670 26324 1676 26376
rect 1728 26364 1734 26376
rect 1765 26367 1823 26373
rect 1765 26364 1777 26367
rect 1728 26336 1777 26364
rect 1728 26324 1734 26336
rect 1765 26333 1777 26336
rect 1811 26333 1823 26367
rect 1765 26327 1823 26333
rect 1854 26324 1860 26376
rect 1912 26364 1918 26376
rect 2225 26367 2283 26373
rect 2225 26364 2237 26367
rect 1912 26336 2237 26364
rect 1912 26324 1918 26336
rect 2225 26333 2237 26336
rect 2271 26333 2283 26367
rect 2225 26327 2283 26333
rect 2406 26324 2412 26376
rect 2464 26364 2470 26376
rect 2501 26367 2559 26373
rect 2501 26364 2513 26367
rect 2464 26336 2513 26364
rect 2464 26324 2470 26336
rect 2501 26333 2513 26336
rect 2547 26364 2559 26367
rect 2774 26364 2780 26376
rect 2547 26336 2780 26364
rect 2547 26333 2559 26336
rect 2501 26327 2559 26333
rect 2774 26324 2780 26336
rect 2832 26324 2838 26376
rect 3786 26324 3792 26376
rect 3844 26364 3850 26376
rect 3844 26336 3924 26364
rect 3844 26324 3850 26336
rect 3896 26240 3924 26336
rect 4982 26324 4988 26376
rect 5040 26324 5046 26376
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26333 5319 26367
rect 5994 26340 6000 26392
rect 6052 26340 6058 26392
rect 6086 26340 6092 26392
rect 6144 26380 6150 26392
rect 6144 26373 6157 26380
rect 6932 26376 6960 26472
rect 8205 26469 8217 26503
rect 8251 26500 8263 26503
rect 8478 26500 8484 26512
rect 8251 26472 8484 26500
rect 8251 26469 8263 26472
rect 8205 26463 8263 26469
rect 8478 26460 8484 26472
rect 8536 26460 8542 26512
rect 9309 26503 9367 26509
rect 9309 26469 9321 26503
rect 9355 26500 9367 26503
rect 10226 26500 10232 26512
rect 9355 26472 10232 26500
rect 9355 26469 9367 26472
rect 9309 26463 9367 26469
rect 10226 26460 10232 26472
rect 10284 26460 10290 26512
rect 6144 26367 6193 26373
rect 6144 26340 6147 26367
rect 5261 26327 5319 26333
rect 5997 26333 6009 26340
rect 6043 26333 6055 26340
rect 6129 26336 6147 26340
rect 5997 26327 6055 26333
rect 6135 26333 6147 26336
rect 6181 26333 6193 26367
rect 6135 26327 6193 26333
rect 4522 26256 4528 26308
rect 4580 26256 4586 26308
rect 4614 26256 4620 26308
rect 4672 26296 4678 26308
rect 5276 26296 5304 26327
rect 6914 26324 6920 26376
rect 6972 26364 6978 26376
rect 7193 26367 7251 26373
rect 7193 26364 7205 26367
rect 6972 26336 7205 26364
rect 6972 26324 6978 26336
rect 7193 26333 7205 26336
rect 7239 26333 7251 26367
rect 7193 26327 7251 26333
rect 7469 26367 7527 26373
rect 7469 26333 7481 26367
rect 7515 26364 7527 26367
rect 7926 26364 7932 26376
rect 7515 26336 7932 26364
rect 7515 26333 7527 26336
rect 7469 26327 7527 26333
rect 7926 26324 7932 26336
rect 7984 26324 7990 26376
rect 8202 26324 8208 26376
rect 8260 26364 8266 26376
rect 8846 26364 8852 26376
rect 8260 26336 8852 26364
rect 8260 26324 8266 26336
rect 8846 26324 8852 26336
rect 8904 26324 8910 26376
rect 8938 26324 8944 26376
rect 8996 26364 9002 26376
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8996 26336 9137 26364
rect 8996 26324 9002 26336
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9490 26324 9496 26376
rect 9548 26324 9554 26376
rect 8294 26296 8300 26308
rect 4672 26268 5304 26296
rect 4672 26256 4678 26268
rect 1946 26188 1952 26240
rect 2004 26188 2010 26240
rect 2958 26188 2964 26240
rect 3016 26228 3022 26240
rect 3786 26228 3792 26240
rect 3016 26200 3792 26228
rect 3016 26188 3022 26200
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 3878 26188 3884 26240
rect 3936 26188 3942 26240
rect 4798 26188 4804 26240
rect 4856 26188 4862 26240
rect 5276 26228 5304 26268
rect 6748 26268 8300 26296
rect 6748 26228 6776 26268
rect 8294 26256 8300 26268
rect 8352 26296 8358 26308
rect 10594 26296 10600 26308
rect 8352 26268 10600 26296
rect 8352 26256 8358 26268
rect 10594 26256 10600 26268
rect 10652 26256 10658 26308
rect 5276 26200 6776 26228
rect 7834 26188 7840 26240
rect 7892 26228 7898 26240
rect 7892 26200 10640 26228
rect 7892 26188 7898 26200
rect 10612 26172 10640 26200
rect 1104 26138 10120 26160
rect 1104 26086 3010 26138
rect 3062 26086 3074 26138
rect 3126 26086 3138 26138
rect 3190 26086 3202 26138
rect 3254 26086 3266 26138
rect 3318 26086 9010 26138
rect 9062 26086 9074 26138
rect 9126 26086 9138 26138
rect 9190 26086 9202 26138
rect 9254 26086 9266 26138
rect 9318 26086 10120 26138
rect 10594 26120 10600 26172
rect 10652 26120 10658 26172
rect 1104 26064 10120 26086
rect 198 25984 204 26036
rect 256 26024 262 26036
rect 3418 26024 3424 26036
rect 256 25996 3424 26024
rect 256 25984 262 25996
rect 3418 25984 3424 25996
rect 3476 25984 3482 26036
rect 3878 25984 3884 26036
rect 3936 26024 3942 26036
rect 6086 26024 6092 26036
rect 3936 25996 6092 26024
rect 3936 25984 3942 25996
rect 6086 25984 6092 25996
rect 6144 25984 6150 26036
rect 7558 25984 7564 26036
rect 7616 26024 7622 26036
rect 7834 26024 7840 26036
rect 7616 25996 7840 26024
rect 7616 25984 7622 25996
rect 7834 25984 7840 25996
rect 7892 25984 7898 26036
rect 8478 26024 8484 26036
rect 8036 25996 8484 26024
rect 1762 25916 1768 25968
rect 1820 25956 1826 25968
rect 1820 25928 2544 25956
rect 1820 25916 1826 25928
rect 2317 25891 2375 25897
rect 2317 25857 2329 25891
rect 2363 25888 2375 25891
rect 2406 25888 2412 25900
rect 2363 25860 2412 25888
rect 2363 25857 2375 25860
rect 2317 25851 2375 25857
rect 2406 25848 2412 25860
rect 2464 25848 2470 25900
rect 2516 25888 2544 25928
rect 2958 25916 2964 25968
rect 3016 25956 3022 25968
rect 6270 25956 6276 25968
rect 3016 25928 6276 25956
rect 3016 25916 3022 25928
rect 6270 25916 6276 25928
rect 6328 25956 6334 25968
rect 6328 25928 6868 25956
rect 6328 25916 6334 25928
rect 2590 25888 2596 25900
rect 2516 25860 2596 25888
rect 2590 25848 2596 25860
rect 2648 25848 2654 25900
rect 3237 25891 3295 25897
rect 3237 25857 3249 25891
rect 3283 25888 3295 25891
rect 3602 25888 3608 25900
rect 3283 25860 3608 25888
rect 3283 25857 3295 25860
rect 3237 25851 3295 25857
rect 3602 25848 3608 25860
rect 3660 25848 3666 25900
rect 6549 25891 6607 25897
rect 6549 25857 6561 25891
rect 6595 25888 6607 25891
rect 6730 25888 6736 25900
rect 6595 25860 6736 25888
rect 6595 25857 6607 25860
rect 6549 25851 6607 25857
rect 6730 25848 6736 25860
rect 6788 25848 6794 25900
rect 6840 25897 6868 25928
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25857 6883 25891
rect 6825 25851 6883 25857
rect 7282 25848 7288 25900
rect 7340 25888 7346 25900
rect 7837 25891 7895 25897
rect 7837 25888 7849 25891
rect 7340 25860 7849 25888
rect 7340 25848 7346 25860
rect 7837 25857 7849 25860
rect 7883 25857 7895 25891
rect 8036 25888 8064 25996
rect 8478 25984 8484 25996
rect 8536 25984 8542 26036
rect 8036 25860 8248 25888
rect 7837 25851 7895 25857
rect 3513 25823 3571 25829
rect 3513 25789 3525 25823
rect 3559 25820 3571 25823
rect 3694 25820 3700 25832
rect 3559 25792 3700 25820
rect 3559 25789 3571 25792
rect 3513 25783 3571 25789
rect 3694 25780 3700 25792
rect 3752 25780 3758 25832
rect 7650 25780 7656 25832
rect 7708 25820 7714 25832
rect 8021 25823 8079 25829
rect 8021 25820 8033 25823
rect 7708 25792 8033 25820
rect 7708 25780 7714 25792
rect 8021 25789 8033 25792
rect 8067 25789 8079 25823
rect 8220 25820 8248 25860
rect 8938 25829 8944 25832
rect 8481 25823 8539 25829
rect 8481 25820 8493 25823
rect 8220 25792 8493 25820
rect 8021 25783 8079 25789
rect 8481 25789 8493 25792
rect 8527 25789 8539 25823
rect 8757 25823 8815 25829
rect 8757 25820 8769 25823
rect 8481 25783 8539 25789
rect 8588 25792 8769 25820
rect 8294 25712 8300 25764
rect 8352 25752 8358 25764
rect 8588 25752 8616 25792
rect 8757 25789 8769 25792
rect 8803 25789 8815 25823
rect 8757 25783 8815 25789
rect 8895 25823 8944 25829
rect 8895 25789 8907 25823
rect 8941 25789 8944 25823
rect 8895 25783 8944 25789
rect 8938 25780 8944 25783
rect 8996 25780 9002 25832
rect 9033 25823 9091 25829
rect 9033 25789 9045 25823
rect 9079 25820 9091 25823
rect 9079 25792 9536 25820
rect 9079 25789 9091 25792
rect 9033 25783 9091 25789
rect 9508 25764 9536 25792
rect 8352 25724 8616 25752
rect 8352 25712 8358 25724
rect 9490 25712 9496 25764
rect 9548 25712 9554 25764
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 2498 25684 2504 25696
rect 1627 25656 2504 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 2498 25644 2504 25656
rect 2556 25644 2562 25696
rect 6822 25644 6828 25696
rect 6880 25684 6886 25696
rect 7561 25687 7619 25693
rect 7561 25684 7573 25687
rect 6880 25656 7573 25684
rect 6880 25644 6886 25656
rect 7561 25653 7573 25656
rect 7607 25653 7619 25687
rect 7561 25647 7619 25653
rect 8570 25644 8576 25696
rect 8628 25684 8634 25696
rect 9677 25687 9735 25693
rect 9677 25684 9689 25687
rect 8628 25656 9689 25684
rect 8628 25644 8634 25656
rect 9677 25653 9689 25656
rect 9723 25653 9735 25687
rect 9677 25647 9735 25653
rect 1104 25594 10120 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 7950 25594
rect 8002 25542 8014 25594
rect 8066 25542 8078 25594
rect 8130 25542 8142 25594
rect 8194 25542 8206 25594
rect 8258 25542 10120 25594
rect 1104 25520 10120 25542
rect 290 25440 296 25492
rect 348 25480 354 25492
rect 1949 25483 2007 25489
rect 1949 25480 1961 25483
rect 348 25452 1961 25480
rect 348 25440 354 25452
rect 1949 25449 1961 25452
rect 1995 25449 2007 25483
rect 1949 25443 2007 25449
rect 2866 25440 2872 25492
rect 2924 25480 2930 25492
rect 3050 25480 3056 25492
rect 2924 25452 3056 25480
rect 2924 25440 2930 25452
rect 3050 25440 3056 25452
rect 3108 25440 3114 25492
rect 4816 25452 6408 25480
rect 4816 25424 4844 25452
rect 4798 25372 4804 25424
rect 4856 25372 4862 25424
rect 4614 25344 4620 25356
rect 2746 25316 4620 25344
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 1765 25279 1823 25285
rect 1765 25245 1777 25279
rect 1811 25276 1823 25279
rect 2498 25276 2504 25288
rect 1811 25248 2504 25276
rect 1811 25245 1823 25248
rect 1765 25239 1823 25245
rect 2498 25236 2504 25248
rect 2556 25236 2562 25288
rect 2746 25208 2774 25316
rect 4614 25304 4620 25316
rect 4672 25304 4678 25356
rect 4816 25285 4844 25372
rect 6380 25353 6408 25452
rect 7558 25440 7564 25492
rect 7616 25480 7622 25492
rect 7926 25480 7932 25492
rect 7616 25452 7932 25480
rect 7616 25440 7622 25452
rect 7926 25440 7932 25452
rect 7984 25440 7990 25492
rect 8481 25483 8539 25489
rect 8481 25449 8493 25483
rect 8527 25480 8539 25483
rect 9490 25480 9496 25492
rect 8527 25452 9496 25480
rect 8527 25449 8539 25452
rect 8481 25443 8539 25449
rect 9490 25440 9496 25452
rect 9548 25440 9554 25492
rect 8938 25412 8944 25424
rect 8312 25384 8944 25412
rect 6365 25347 6423 25353
rect 6365 25313 6377 25347
rect 6411 25313 6423 25347
rect 7469 25347 7527 25353
rect 7469 25344 7481 25347
rect 6365 25307 6423 25313
rect 6932 25316 7144 25344
rect 6932 25288 6960 25316
rect 7116 25288 7144 25316
rect 7392 25316 7481 25344
rect 4801 25279 4859 25285
rect 4801 25245 4813 25279
rect 4847 25245 4859 25279
rect 4801 25239 4859 25245
rect 4982 25236 4988 25288
rect 5040 25276 5046 25288
rect 5077 25279 5135 25285
rect 5077 25276 5089 25279
rect 5040 25248 5089 25276
rect 5040 25236 5046 25248
rect 5077 25245 5089 25248
rect 5123 25276 5135 25279
rect 5166 25276 5172 25288
rect 5123 25248 5172 25276
rect 5123 25245 5135 25248
rect 5077 25239 5135 25245
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 5442 25236 5448 25288
rect 5500 25276 5506 25288
rect 6641 25279 6699 25285
rect 6641 25276 6653 25279
rect 5500 25248 6653 25276
rect 5500 25236 5506 25248
rect 6641 25245 6653 25248
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6914 25236 6920 25288
rect 6972 25236 6978 25288
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 7392 25276 7420 25316
rect 7469 25313 7481 25316
rect 7515 25313 7527 25347
rect 7469 25307 7527 25313
rect 7156 25248 7420 25276
rect 7745 25279 7803 25285
rect 7156 25236 7162 25248
rect 7745 25245 7757 25279
rect 7791 25276 7803 25279
rect 8018 25276 8024 25288
rect 7791 25248 8024 25276
rect 7791 25245 7803 25248
rect 7745 25239 7803 25245
rect 8018 25236 8024 25248
rect 8076 25236 8082 25288
rect 8202 25236 8208 25288
rect 8260 25276 8266 25288
rect 8312 25276 8340 25384
rect 8938 25372 8944 25384
rect 8996 25372 9002 25424
rect 9309 25415 9367 25421
rect 9309 25381 9321 25415
rect 9355 25412 9367 25415
rect 10226 25412 10232 25424
rect 9355 25384 10232 25412
rect 9355 25381 9367 25384
rect 9309 25375 9367 25381
rect 10226 25372 10232 25384
rect 10284 25372 10290 25424
rect 10318 25372 10324 25424
rect 10376 25412 10382 25424
rect 11146 25412 11152 25424
rect 10376 25384 11152 25412
rect 10376 25372 10382 25384
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 8260 25248 8340 25276
rect 8404 25316 9536 25344
rect 8260 25236 8266 25248
rect 3050 25208 3056 25220
rect 1596 25180 2774 25208
rect 2884 25180 3056 25208
rect 1596 25149 1624 25180
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25109 1639 25143
rect 1581 25103 1639 25109
rect 2222 25100 2228 25152
rect 2280 25140 2286 25152
rect 2884 25140 2912 25180
rect 3050 25168 3056 25180
rect 3108 25168 3114 25220
rect 7558 25168 7564 25220
rect 7616 25208 7622 25220
rect 8404 25208 8432 25316
rect 8570 25236 8576 25288
rect 8628 25236 8634 25288
rect 9030 25276 9036 25288
rect 8680 25248 9036 25276
rect 7616 25180 8432 25208
rect 7616 25168 7622 25180
rect 2280 25112 2912 25140
rect 2280 25100 2286 25112
rect 5810 25100 5816 25152
rect 5868 25100 5874 25152
rect 6914 25100 6920 25152
rect 6972 25140 6978 25152
rect 7377 25143 7435 25149
rect 7377 25140 7389 25143
rect 6972 25112 7389 25140
rect 6972 25100 6978 25112
rect 7377 25109 7389 25112
rect 7423 25109 7435 25143
rect 7377 25103 7435 25109
rect 7926 25100 7932 25152
rect 7984 25140 7990 25152
rect 8202 25140 8208 25152
rect 7984 25112 8208 25140
rect 7984 25100 7990 25112
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 8680 25140 8708 25248
rect 9030 25236 9036 25248
rect 9088 25236 9094 25288
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9398 25276 9404 25288
rect 9171 25248 9404 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9398 25236 9404 25248
rect 9456 25236 9462 25288
rect 9508 25285 9536 25316
rect 10134 25304 10140 25356
rect 10192 25344 10198 25356
rect 10870 25344 10876 25356
rect 10192 25316 10876 25344
rect 10192 25304 10198 25316
rect 10870 25304 10876 25316
rect 10928 25304 10934 25356
rect 9493 25279 9551 25285
rect 9493 25245 9505 25279
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 10042 25208 10048 25220
rect 8772 25180 10048 25208
rect 8772 25149 8800 25180
rect 10042 25168 10048 25180
rect 10100 25168 10106 25220
rect 8352 25112 8708 25140
rect 8757 25143 8815 25149
rect 8352 25100 8358 25112
rect 8757 25109 8769 25143
rect 8803 25109 8815 25143
rect 8757 25103 8815 25109
rect 9674 25100 9680 25152
rect 9732 25100 9738 25152
rect 1104 25050 10120 25072
rect 1104 24998 3010 25050
rect 3062 24998 3074 25050
rect 3126 24998 3138 25050
rect 3190 24998 3202 25050
rect 3254 24998 3266 25050
rect 3318 24998 9010 25050
rect 9062 24998 9074 25050
rect 9126 24998 9138 25050
rect 9190 24998 9202 25050
rect 9254 24998 9266 25050
rect 9318 24998 10120 25050
rect 1104 24976 10120 24998
rect 2958 24896 2964 24948
rect 3016 24936 3022 24948
rect 3878 24936 3884 24948
rect 3016 24908 3884 24936
rect 3016 24896 3022 24908
rect 3878 24896 3884 24908
rect 3936 24896 3942 24948
rect 4982 24896 4988 24948
rect 5040 24936 5046 24948
rect 5442 24936 5448 24948
rect 5040 24908 5448 24936
rect 5040 24896 5046 24908
rect 5442 24896 5448 24908
rect 5500 24896 5506 24948
rect 5629 24939 5687 24945
rect 5629 24905 5641 24939
rect 5675 24936 5687 24939
rect 6730 24936 6736 24948
rect 5675 24908 6736 24936
rect 5675 24905 5687 24908
rect 5629 24899 5687 24905
rect 6730 24896 6736 24908
rect 6788 24896 6794 24948
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 7248 24908 8984 24936
rect 7248 24896 7254 24908
rect 1394 24760 1400 24812
rect 1452 24760 1458 24812
rect 2130 24760 2136 24812
rect 2188 24800 2194 24812
rect 2685 24803 2743 24809
rect 2685 24800 2697 24803
rect 2188 24772 2697 24800
rect 2188 24760 2194 24772
rect 2685 24769 2697 24772
rect 2731 24769 2743 24803
rect 2685 24763 2743 24769
rect 5442 24760 5448 24812
rect 5500 24760 5506 24812
rect 7098 24760 7104 24812
rect 7156 24800 7162 24812
rect 7377 24803 7435 24809
rect 7377 24800 7389 24803
rect 7156 24772 7389 24800
rect 7156 24760 7162 24772
rect 7377 24769 7389 24772
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 8110 24760 8116 24812
rect 8168 24760 8174 24812
rect 8202 24760 8208 24812
rect 8260 24809 8266 24812
rect 8260 24803 8288 24809
rect 8276 24769 8288 24803
rect 8956 24800 8984 24908
rect 9217 24871 9275 24877
rect 9217 24837 9229 24871
rect 9263 24868 9275 24871
rect 9398 24868 9404 24880
rect 9263 24840 9404 24868
rect 9263 24837 9275 24840
rect 9217 24831 9275 24837
rect 9398 24828 9404 24840
rect 9456 24868 9462 24880
rect 9456 24840 9628 24868
rect 9456 24828 9462 24840
rect 9493 24803 9551 24809
rect 9493 24800 9505 24803
rect 8956 24772 9505 24800
rect 8260 24763 8288 24769
rect 9493 24769 9505 24772
rect 9539 24769 9551 24803
rect 9600 24800 9628 24840
rect 10778 24800 10784 24812
rect 9600 24772 10784 24800
rect 9493 24763 9551 24769
rect 8260 24760 8266 24763
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 658 24692 664 24744
rect 716 24732 722 24744
rect 2222 24732 2228 24744
rect 716 24704 2228 24732
rect 716 24692 722 24704
rect 2222 24692 2228 24704
rect 2280 24692 2286 24744
rect 2406 24692 2412 24744
rect 2464 24692 2470 24744
rect 3142 24692 3148 24744
rect 3200 24732 3206 24744
rect 3513 24735 3571 24741
rect 3513 24732 3525 24735
rect 3200 24704 3525 24732
rect 3200 24692 3206 24704
rect 3513 24701 3525 24704
rect 3559 24701 3571 24735
rect 3513 24695 3571 24701
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24732 3755 24735
rect 3786 24732 3792 24744
rect 3743 24704 3792 24732
rect 3743 24701 3755 24704
rect 3697 24695 3755 24701
rect 3786 24692 3792 24704
rect 3844 24692 3850 24744
rect 4614 24741 4620 24744
rect 4433 24735 4491 24741
rect 4433 24732 4445 24735
rect 4264 24704 4445 24732
rect 1578 24624 1584 24676
rect 1636 24624 1642 24676
rect 4154 24624 4160 24676
rect 4212 24624 4218 24676
rect 3421 24599 3479 24605
rect 3421 24565 3433 24599
rect 3467 24596 3479 24599
rect 3878 24596 3884 24608
rect 3467 24568 3884 24596
rect 3467 24565 3479 24568
rect 3421 24559 3479 24565
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 4264 24596 4292 24704
rect 4433 24701 4445 24704
rect 4479 24701 4491 24735
rect 4433 24695 4491 24701
rect 4571 24735 4620 24741
rect 4571 24701 4583 24735
rect 4617 24701 4620 24735
rect 4571 24695 4620 24701
rect 4614 24692 4620 24695
rect 4672 24692 4678 24744
rect 4706 24692 4712 24744
rect 4764 24692 4770 24744
rect 7190 24692 7196 24744
rect 7248 24692 7254 24744
rect 7926 24732 7932 24744
rect 7760 24704 7932 24732
rect 6270 24664 6276 24676
rect 5092 24636 6276 24664
rect 5092 24596 5120 24636
rect 6270 24624 6276 24636
rect 6328 24664 6334 24676
rect 7760 24664 7788 24704
rect 7926 24692 7932 24704
rect 7984 24692 7990 24744
rect 8386 24692 8392 24744
rect 8444 24692 8450 24744
rect 8570 24692 8576 24744
rect 8628 24732 8634 24744
rect 8938 24732 8944 24744
rect 8628 24704 8944 24732
rect 8628 24692 8634 24704
rect 8938 24692 8944 24704
rect 8996 24692 9002 24744
rect 6328 24636 7788 24664
rect 6328 24624 6334 24636
rect 7834 24624 7840 24676
rect 7892 24624 7898 24676
rect 9490 24624 9496 24676
rect 9548 24664 9554 24676
rect 9766 24664 9772 24676
rect 9548 24636 9772 24664
rect 9548 24624 9554 24636
rect 9766 24624 9772 24636
rect 9824 24624 9830 24676
rect 4264 24568 5120 24596
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5353 24599 5411 24605
rect 5353 24596 5365 24599
rect 5224 24568 5365 24596
rect 5224 24556 5230 24568
rect 5353 24565 5365 24568
rect 5399 24565 5411 24599
rect 5353 24559 5411 24565
rect 6638 24556 6644 24608
rect 6696 24596 6702 24608
rect 7190 24596 7196 24608
rect 6696 24568 7196 24596
rect 6696 24556 6702 24568
rect 7190 24556 7196 24568
rect 7248 24556 7254 24608
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 8110 24596 8116 24608
rect 7340 24568 8116 24596
rect 7340 24556 7346 24568
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 8570 24556 8576 24608
rect 8628 24596 8634 24608
rect 9033 24599 9091 24605
rect 9033 24596 9045 24599
rect 8628 24568 9045 24596
rect 8628 24556 8634 24568
rect 9033 24565 9045 24568
rect 9079 24565 9091 24599
rect 9033 24559 9091 24565
rect 9674 24556 9680 24608
rect 9732 24556 9738 24608
rect 1104 24506 10120 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 7950 24506
rect 8002 24454 8014 24506
rect 8066 24454 8078 24506
rect 8130 24454 8142 24506
rect 8194 24454 8206 24506
rect 8258 24454 10120 24506
rect 1104 24432 10120 24454
rect 1486 24352 1492 24404
rect 1544 24392 1550 24404
rect 1581 24395 1639 24401
rect 1581 24392 1593 24395
rect 1544 24364 1593 24392
rect 1544 24352 1550 24364
rect 1581 24361 1593 24364
rect 1627 24361 1639 24395
rect 1581 24355 1639 24361
rect 5169 24395 5227 24401
rect 5169 24361 5181 24395
rect 5215 24392 5227 24395
rect 6454 24392 6460 24404
rect 5215 24364 6460 24392
rect 5215 24361 5227 24364
rect 5169 24355 5227 24361
rect 6454 24352 6460 24364
rect 6512 24352 6518 24404
rect 8113 24395 8171 24401
rect 8113 24361 8125 24395
rect 8159 24392 8171 24395
rect 8386 24392 8392 24404
rect 8159 24364 8392 24392
rect 8159 24361 8171 24364
rect 8113 24355 8171 24361
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 9677 24395 9735 24401
rect 9677 24361 9689 24395
rect 9723 24392 9735 24395
rect 9766 24392 9772 24404
rect 9723 24364 9772 24392
rect 9723 24361 9735 24364
rect 9677 24355 9735 24361
rect 9766 24352 9772 24364
rect 9824 24352 9830 24404
rect 4890 24284 4896 24336
rect 4948 24324 4954 24336
rect 5350 24324 5356 24336
rect 4948 24296 5356 24324
rect 4948 24284 4954 24296
rect 5350 24284 5356 24296
rect 5408 24284 5414 24336
rect 6270 24284 6276 24336
rect 6328 24284 6334 24336
rect 6365 24327 6423 24333
rect 6365 24293 6377 24327
rect 6411 24324 6423 24327
rect 6914 24324 6920 24336
rect 6411 24296 6920 24324
rect 6411 24293 6423 24296
rect 6365 24287 6423 24293
rect 6914 24284 6920 24296
rect 6972 24284 6978 24336
rect 8938 24324 8944 24336
rect 8036 24296 8944 24324
rect 1854 24216 1860 24268
rect 1912 24256 1918 24268
rect 2130 24256 2136 24268
rect 1912 24228 2136 24256
rect 1912 24216 1918 24228
rect 2130 24216 2136 24228
rect 2188 24256 2194 24268
rect 2406 24256 2412 24268
rect 2188 24228 2412 24256
rect 2188 24216 2194 24228
rect 2406 24216 2412 24228
rect 2464 24216 2470 24268
rect 5951 24259 6009 24265
rect 5951 24256 5963 24259
rect 5276 24228 5963 24256
rect 1394 24148 1400 24200
rect 1452 24148 1458 24200
rect 2314 24148 2320 24200
rect 2372 24188 2378 24200
rect 2685 24191 2743 24197
rect 2685 24188 2697 24191
rect 2372 24160 2697 24188
rect 2372 24148 2378 24160
rect 2685 24157 2697 24160
rect 2731 24157 2743 24191
rect 2685 24151 2743 24157
rect 2222 24080 2228 24132
rect 2280 24120 2286 24132
rect 4154 24120 4160 24132
rect 2280 24092 4160 24120
rect 2280 24080 2286 24092
rect 4154 24080 4160 24092
rect 4212 24080 4218 24132
rect 2314 24012 2320 24064
rect 2372 24052 2378 24064
rect 2590 24052 2596 24064
rect 2372 24024 2596 24052
rect 2372 24012 2378 24024
rect 2590 24012 2596 24024
rect 2648 24012 2654 24064
rect 3421 24055 3479 24061
rect 3421 24021 3433 24055
rect 3467 24052 3479 24055
rect 4430 24052 4436 24064
rect 3467 24024 4436 24052
rect 3467 24021 3479 24024
rect 3421 24015 3479 24021
rect 4430 24012 4436 24024
rect 4488 24012 4494 24064
rect 4614 24012 4620 24064
rect 4672 24052 4678 24064
rect 5276 24052 5304 24228
rect 5951 24225 5963 24228
rect 5997 24225 6009 24259
rect 6288 24256 6316 24284
rect 5951 24219 6009 24225
rect 6104 24228 6316 24256
rect 5810 24148 5816 24200
rect 5868 24148 5874 24200
rect 6104 24197 6132 24228
rect 8036 24200 8064 24296
rect 8938 24284 8944 24296
rect 8996 24284 9002 24336
rect 9309 24327 9367 24333
rect 9309 24293 9321 24327
rect 9355 24324 9367 24327
rect 10226 24324 10232 24336
rect 9355 24296 10232 24324
rect 9355 24293 9367 24296
rect 9309 24287 9367 24293
rect 10226 24284 10232 24296
rect 10284 24284 10290 24336
rect 8846 24216 8852 24268
rect 8904 24256 8910 24268
rect 8904 24228 9536 24256
rect 8904 24216 8910 24228
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24157 6147 24191
rect 6089 24151 6147 24157
rect 6638 24148 6644 24200
rect 6696 24188 6702 24200
rect 6825 24191 6883 24197
rect 6825 24188 6837 24191
rect 6696 24160 6837 24188
rect 6696 24148 6702 24160
rect 6825 24157 6837 24160
rect 6871 24157 6883 24191
rect 6825 24151 6883 24157
rect 7009 24191 7067 24197
rect 7009 24157 7021 24191
rect 7055 24157 7067 24191
rect 7009 24151 7067 24157
rect 7101 24191 7159 24197
rect 7101 24157 7113 24191
rect 7147 24188 7159 24191
rect 7282 24188 7288 24200
rect 7147 24160 7288 24188
rect 7147 24157 7159 24160
rect 7101 24151 7159 24157
rect 7024 24120 7052 24151
rect 7282 24148 7288 24160
rect 7340 24148 7346 24200
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 8018 24188 8024 24200
rect 7423 24160 8024 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 8018 24148 8024 24160
rect 8076 24148 8082 24200
rect 8570 24148 8576 24200
rect 8628 24148 8634 24200
rect 9122 24148 9128 24200
rect 9180 24148 9186 24200
rect 9508 24197 9536 24228
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24157 9551 24191
rect 9493 24151 9551 24157
rect 7926 24120 7932 24132
rect 7024 24092 7932 24120
rect 7926 24080 7932 24092
rect 7984 24080 7990 24132
rect 6454 24052 6460 24064
rect 4672 24024 6460 24052
rect 4672 24012 4678 24024
rect 6454 24012 6460 24024
rect 6512 24012 6518 24064
rect 8754 24012 8760 24064
rect 8812 24012 8818 24064
rect 1104 23962 10120 23984
rect 1104 23910 3010 23962
rect 3062 23910 3074 23962
rect 3126 23910 3138 23962
rect 3190 23910 3202 23962
rect 3254 23910 3266 23962
rect 3318 23910 9010 23962
rect 9062 23910 9074 23962
rect 9126 23910 9138 23962
rect 9190 23910 9202 23962
rect 9254 23910 9266 23962
rect 9318 23910 10120 23962
rect 1104 23888 10120 23910
rect 2222 23808 2228 23860
rect 2280 23848 2286 23860
rect 3053 23851 3111 23857
rect 3053 23848 3065 23851
rect 2280 23820 3065 23848
rect 2280 23808 2286 23820
rect 3053 23817 3065 23820
rect 3099 23817 3111 23851
rect 3053 23811 3111 23817
rect 5077 23851 5135 23857
rect 5077 23817 5089 23851
rect 5123 23848 5135 23851
rect 5442 23848 5448 23860
rect 5123 23820 5448 23848
rect 5123 23817 5135 23820
rect 5077 23811 5135 23817
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 7742 23848 7748 23860
rect 5592 23820 7748 23848
rect 5592 23808 5598 23820
rect 7742 23808 7748 23820
rect 7800 23808 7806 23860
rect 7834 23808 7840 23860
rect 7892 23848 7898 23860
rect 8297 23851 8355 23857
rect 8297 23848 8309 23851
rect 7892 23820 8309 23848
rect 7892 23808 7898 23820
rect 8297 23817 8309 23820
rect 8343 23817 8355 23851
rect 8297 23811 8355 23817
rect 8662 23808 8668 23860
rect 8720 23848 8726 23860
rect 9306 23848 9312 23860
rect 8720 23820 9312 23848
rect 8720 23808 8726 23820
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 9674 23808 9680 23860
rect 9732 23808 9738 23860
rect 2130 23740 2136 23792
rect 2188 23780 2194 23792
rect 2590 23780 2596 23792
rect 2188 23752 2596 23780
rect 2188 23740 2194 23752
rect 2590 23740 2596 23752
rect 2648 23740 2654 23792
rect 3234 23740 3240 23792
rect 3292 23780 3298 23792
rect 3292 23752 3464 23780
rect 3292 23740 3298 23752
rect 1486 23672 1492 23724
rect 1544 23712 1550 23724
rect 3436 23721 3464 23752
rect 6362 23740 6368 23792
rect 6420 23780 6426 23792
rect 6730 23780 6736 23792
rect 6420 23752 6736 23780
rect 6420 23740 6426 23752
rect 6730 23740 6736 23752
rect 6788 23740 6794 23792
rect 7374 23740 7380 23792
rect 7432 23780 7438 23792
rect 7432 23752 8524 23780
rect 7432 23740 7438 23752
rect 2317 23715 2375 23721
rect 2317 23712 2329 23715
rect 1544 23684 2329 23712
rect 1544 23672 1550 23684
rect 2317 23681 2329 23684
rect 2363 23681 2375 23715
rect 2317 23675 2375 23681
rect 3421 23715 3479 23721
rect 3421 23681 3433 23715
rect 3467 23681 3479 23715
rect 3421 23675 3479 23681
rect 4154 23672 4160 23724
rect 4212 23672 4218 23724
rect 4430 23672 4436 23724
rect 4488 23672 4494 23724
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5902 23672 5908 23724
rect 5960 23712 5966 23724
rect 7561 23715 7619 23721
rect 7561 23712 7573 23715
rect 5960 23684 7573 23712
rect 5960 23672 5966 23684
rect 7561 23681 7573 23684
rect 7607 23712 7619 23715
rect 8202 23712 8208 23724
rect 7607 23684 8208 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 8202 23672 8208 23684
rect 8260 23712 8266 23724
rect 8389 23715 8447 23721
rect 8389 23712 8401 23715
rect 8260 23684 8401 23712
rect 8260 23672 8266 23684
rect 8389 23681 8401 23684
rect 8435 23681 8447 23715
rect 8389 23675 8447 23681
rect 1854 23604 1860 23656
rect 1912 23644 1918 23656
rect 2041 23647 2099 23653
rect 2041 23644 2053 23647
rect 1912 23616 2053 23644
rect 1912 23604 1918 23616
rect 2041 23613 2053 23616
rect 2087 23613 2099 23647
rect 2041 23607 2099 23613
rect 3237 23647 3295 23653
rect 3237 23613 3249 23647
rect 3283 23613 3295 23647
rect 3237 23607 3295 23613
rect 3252 23508 3280 23607
rect 3878 23604 3884 23656
rect 3936 23604 3942 23656
rect 4295 23647 4353 23653
rect 4295 23613 4307 23647
rect 4341 23644 4353 23647
rect 6270 23644 6276 23656
rect 4341 23616 6276 23644
rect 4341 23613 4353 23616
rect 4295 23607 4353 23613
rect 6270 23604 6276 23616
rect 6328 23604 6334 23656
rect 7282 23604 7288 23656
rect 7340 23604 7346 23656
rect 8496 23644 8524 23752
rect 8846 23740 8852 23792
rect 8904 23780 8910 23792
rect 8904 23752 9536 23780
rect 8904 23740 8910 23752
rect 8754 23672 8760 23724
rect 8812 23712 8818 23724
rect 9508 23721 9536 23752
rect 9125 23715 9183 23721
rect 9125 23712 9137 23715
rect 8812 23684 9137 23712
rect 8812 23672 8818 23684
rect 9125 23681 9137 23684
rect 9171 23681 9183 23715
rect 9125 23675 9183 23681
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23681 9551 23715
rect 9493 23675 9551 23681
rect 10962 23644 10968 23656
rect 8496 23616 10968 23644
rect 10962 23604 10968 23616
rect 11020 23604 11026 23656
rect 5442 23536 5448 23588
rect 5500 23576 5506 23588
rect 7300 23576 7328 23604
rect 5500 23548 7328 23576
rect 8573 23579 8631 23585
rect 5500 23536 5506 23548
rect 8573 23545 8585 23579
rect 8619 23576 8631 23579
rect 9858 23576 9864 23588
rect 8619 23548 9864 23576
rect 8619 23545 8631 23548
rect 8573 23539 8631 23545
rect 9858 23536 9864 23548
rect 9916 23536 9922 23588
rect 4614 23508 4620 23520
rect 3252 23480 4620 23508
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 5353 23511 5411 23517
rect 5353 23477 5365 23511
rect 5399 23508 5411 23511
rect 8478 23508 8484 23520
rect 5399 23480 8484 23508
rect 5399 23477 5411 23480
rect 5353 23471 5411 23477
rect 8478 23468 8484 23480
rect 8536 23468 8542 23520
rect 9309 23511 9367 23517
rect 9309 23477 9321 23511
rect 9355 23508 9367 23511
rect 10226 23508 10232 23520
rect 9355 23480 10232 23508
rect 9355 23477 9367 23480
rect 9309 23471 9367 23477
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 106 23400 112 23452
rect 164 23400 170 23452
rect 1104 23418 10120 23440
rect 124 22964 152 23400
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 7950 23418
rect 8002 23366 8014 23418
rect 8066 23366 8078 23418
rect 8130 23366 8142 23418
rect 8194 23366 8206 23418
rect 8258 23366 10120 23418
rect 1104 23344 10120 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 2866 23304 2872 23316
rect 1627 23276 2872 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 2866 23264 2872 23276
rect 2924 23264 2930 23316
rect 2961 23307 3019 23313
rect 2961 23273 2973 23307
rect 3007 23304 3019 23307
rect 4706 23304 4712 23316
rect 3007 23276 4712 23304
rect 3007 23273 3019 23276
rect 2961 23267 3019 23273
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 6822 23264 6828 23316
rect 6880 23304 6886 23316
rect 7374 23304 7380 23316
rect 6880 23276 7380 23304
rect 6880 23264 6886 23276
rect 7374 23264 7380 23276
rect 7432 23264 7438 23316
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 7742 23304 7748 23316
rect 7616 23276 7748 23304
rect 7616 23264 7622 23276
rect 7742 23264 7748 23276
rect 7800 23264 7806 23316
rect 8754 23264 8760 23316
rect 8812 23304 8818 23316
rect 9582 23304 9588 23316
rect 8812 23276 9588 23304
rect 8812 23264 8818 23276
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 474 23196 480 23248
rect 532 23236 538 23248
rect 1857 23239 1915 23245
rect 1857 23236 1869 23239
rect 532 23208 1869 23236
rect 532 23196 538 23208
rect 1857 23205 1869 23208
rect 1903 23205 1915 23239
rect 1857 23199 1915 23205
rect 1946 23196 1952 23248
rect 2004 23196 2010 23248
rect 9674 23196 9680 23248
rect 9732 23196 9738 23248
rect 1964 23168 1992 23196
rect 1688 23140 1992 23168
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 1688 23109 1716 23140
rect 2590 23128 2596 23180
rect 2648 23168 2654 23180
rect 4614 23168 4620 23180
rect 2648 23140 4620 23168
rect 2648 23128 2654 23140
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 6362 23128 6368 23180
rect 6420 23168 6426 23180
rect 6733 23171 6791 23177
rect 6733 23168 6745 23171
rect 6420 23140 6745 23168
rect 6420 23128 6426 23140
rect 6733 23137 6745 23140
rect 6779 23137 6791 23171
rect 6733 23131 6791 23137
rect 7006 23128 7012 23180
rect 7064 23168 7070 23180
rect 7745 23171 7803 23177
rect 7745 23168 7757 23171
rect 7064 23140 7757 23168
rect 7064 23128 7070 23140
rect 7745 23137 7757 23140
rect 7791 23137 7803 23171
rect 7745 23131 7803 23137
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23069 1731 23103
rect 1673 23063 1731 23069
rect 1854 23060 1860 23112
rect 1912 23100 1918 23112
rect 1949 23103 2007 23109
rect 1949 23100 1961 23103
rect 1912 23072 1961 23100
rect 1912 23060 1918 23072
rect 1949 23069 1961 23072
rect 1995 23069 2007 23103
rect 1949 23063 2007 23069
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23069 2283 23103
rect 2225 23063 2283 23069
rect 1578 22992 1584 23044
rect 1636 23032 1642 23044
rect 2038 23032 2044 23044
rect 1636 23004 2044 23032
rect 1636 22992 1642 23004
rect 2038 22992 2044 23004
rect 2096 23032 2102 23044
rect 2240 23032 2268 23063
rect 5718 23060 5724 23112
rect 5776 23100 5782 23112
rect 7760 23100 7788 23131
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 9582 23168 9588 23180
rect 9456 23140 9588 23168
rect 9456 23128 9462 23140
rect 9582 23128 9588 23140
rect 9640 23128 9646 23180
rect 7926 23100 7932 23112
rect 5776 23072 6684 23100
rect 7760 23072 7932 23100
rect 5776 23060 5782 23072
rect 2096 23004 2268 23032
rect 2096 22992 2102 23004
rect 4798 22992 4804 23044
rect 4856 23032 4862 23044
rect 6549 23035 6607 23041
rect 6549 23032 6561 23035
rect 4856 23004 6561 23032
rect 4856 22992 4862 23004
rect 6549 23001 6561 23004
rect 6595 23001 6607 23035
rect 6656 23032 6684 23072
rect 7926 23060 7932 23072
rect 7984 23060 7990 23112
rect 8018 23060 8024 23112
rect 8076 23060 8082 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 8128 23072 9137 23100
rect 8128 23032 8156 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9125 23063 9183 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 6656 23004 8156 23032
rect 6549 22995 6607 23001
rect 8570 22992 8576 23044
rect 8628 23032 8634 23044
rect 9508 23032 9536 23063
rect 8628 23004 9536 23032
rect 8628 22992 8634 23004
rect 2682 22964 2688 22976
rect 124 22936 2688 22964
rect 2682 22924 2688 22936
rect 2740 22924 2746 22976
rect 3786 22924 3792 22976
rect 3844 22964 3850 22976
rect 5350 22964 5356 22976
rect 3844 22936 5356 22964
rect 3844 22924 3850 22936
rect 5350 22924 5356 22936
rect 5408 22924 5414 22976
rect 5994 22924 6000 22976
rect 6052 22964 6058 22976
rect 6181 22967 6239 22973
rect 6181 22964 6193 22967
rect 6052 22936 6193 22964
rect 6052 22924 6058 22936
rect 6181 22933 6193 22936
rect 6227 22933 6239 22967
rect 6181 22927 6239 22933
rect 6270 22924 6276 22976
rect 6328 22964 6334 22976
rect 6641 22967 6699 22973
rect 6641 22964 6653 22967
rect 6328 22936 6653 22964
rect 6328 22924 6334 22936
rect 6641 22933 6653 22936
rect 6687 22933 6699 22967
rect 6641 22927 6699 22933
rect 8757 22967 8815 22973
rect 8757 22933 8769 22967
rect 8803 22964 8815 22967
rect 8846 22964 8852 22976
rect 8803 22936 8852 22964
rect 8803 22933 8815 22936
rect 8757 22927 8815 22933
rect 8846 22924 8852 22936
rect 8904 22924 8910 22976
rect 9309 22967 9367 22973
rect 9309 22933 9321 22967
rect 9355 22964 9367 22967
rect 10226 22964 10232 22976
rect 9355 22936 10232 22964
rect 9355 22933 9367 22936
rect 9309 22927 9367 22933
rect 10226 22924 10232 22936
rect 10284 22924 10290 22976
rect 1104 22874 10120 22896
rect 1104 22822 3010 22874
rect 3062 22822 3074 22874
rect 3126 22822 3138 22874
rect 3190 22822 3202 22874
rect 3254 22822 3266 22874
rect 3318 22822 9010 22874
rect 9062 22822 9074 22874
rect 9126 22822 9138 22874
rect 9190 22822 9202 22874
rect 9254 22822 9266 22874
rect 9318 22822 10120 22874
rect 1104 22800 10120 22822
rect 10226 22788 10232 22840
rect 10284 22828 10290 22840
rect 10594 22828 10600 22840
rect 10284 22800 10600 22828
rect 10284 22788 10290 22800
rect 10594 22788 10600 22800
rect 10652 22788 10658 22840
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 1627 22732 6224 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 2774 22692 2780 22704
rect 1688 22664 2780 22692
rect 1394 22584 1400 22636
rect 1452 22584 1458 22636
rect 1486 22584 1492 22636
rect 1544 22624 1550 22636
rect 1688 22633 1716 22664
rect 2774 22652 2780 22664
rect 2832 22652 2838 22704
rect 4614 22692 4620 22704
rect 4264 22664 4620 22692
rect 1673 22627 1731 22633
rect 1673 22624 1685 22627
rect 1544 22596 1685 22624
rect 1544 22584 1550 22596
rect 1673 22593 1685 22596
rect 1719 22593 1731 22627
rect 1673 22587 1731 22593
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22624 2007 22627
rect 2038 22624 2044 22636
rect 1995 22596 2044 22624
rect 1995 22593 2007 22596
rect 1949 22587 2007 22593
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 4264 22633 4292 22664
rect 4614 22652 4620 22664
rect 4672 22652 4678 22704
rect 4249 22627 4307 22633
rect 4249 22593 4261 22627
rect 4295 22593 4307 22627
rect 4249 22587 4307 22593
rect 4525 22627 4583 22633
rect 4525 22593 4537 22627
rect 4571 22624 4583 22627
rect 4982 22624 4988 22636
rect 4571 22596 4988 22624
rect 4571 22593 4583 22596
rect 4525 22587 4583 22593
rect 4982 22584 4988 22596
rect 5040 22624 5046 22636
rect 5166 22624 5172 22636
rect 5040 22596 5172 22624
rect 5040 22584 5046 22596
rect 5166 22584 5172 22596
rect 5224 22584 5230 22636
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6196 22624 6224 22732
rect 6362 22720 6368 22772
rect 6420 22720 6426 22772
rect 7006 22720 7012 22772
rect 7064 22760 7070 22772
rect 9033 22763 9091 22769
rect 9033 22760 9045 22763
rect 7064 22732 9045 22760
rect 7064 22720 7070 22732
rect 9033 22729 9045 22732
rect 9079 22729 9091 22763
rect 9033 22723 9091 22729
rect 9493 22763 9551 22769
rect 9493 22729 9505 22763
rect 9539 22729 9551 22763
rect 9493 22723 9551 22729
rect 6270 22652 6276 22704
rect 6328 22692 6334 22704
rect 6328 22664 7236 22692
rect 6328 22652 6334 22664
rect 6730 22624 6736 22636
rect 6196 22596 6736 22624
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 7006 22584 7012 22636
rect 7064 22624 7070 22636
rect 7101 22627 7159 22633
rect 7101 22624 7113 22627
rect 7064 22596 7113 22624
rect 7064 22584 7070 22596
rect 7101 22593 7113 22596
rect 7147 22593 7159 22627
rect 7208 22624 7236 22664
rect 7558 22652 7564 22704
rect 7616 22692 7622 22704
rect 9125 22695 9183 22701
rect 9125 22692 9137 22695
rect 7616 22664 9137 22692
rect 7616 22652 7622 22664
rect 9125 22661 9137 22664
rect 9171 22661 9183 22695
rect 9125 22655 9183 22661
rect 8389 22627 8447 22633
rect 8389 22624 8401 22627
rect 7208 22596 8401 22624
rect 7101 22587 7159 22593
rect 8389 22593 8401 22596
rect 8435 22593 8447 22627
rect 9508 22624 9536 22723
rect 9769 22627 9827 22633
rect 9769 22624 9781 22627
rect 9508 22596 9781 22624
rect 8389 22587 8447 22593
rect 9769 22593 9781 22596
rect 9815 22593 9827 22627
rect 9769 22587 9827 22593
rect 5258 22516 5264 22568
rect 5316 22516 5322 22568
rect 5626 22516 5632 22568
rect 5684 22556 5690 22568
rect 6362 22556 6368 22568
rect 5684 22528 6368 22556
rect 5684 22516 5690 22528
rect 6362 22516 6368 22528
rect 6420 22516 6426 22568
rect 7377 22559 7435 22565
rect 7377 22525 7389 22559
rect 7423 22556 7435 22559
rect 7926 22556 7932 22568
rect 7423 22528 7932 22556
rect 7423 22525 7435 22528
rect 7377 22519 7435 22525
rect 7926 22516 7932 22528
rect 7984 22516 7990 22568
rect 8846 22516 8852 22568
rect 8904 22516 8910 22568
rect 4982 22448 4988 22500
rect 5040 22488 5046 22500
rect 5276 22488 5304 22516
rect 5040 22460 5304 22488
rect 8573 22491 8631 22497
rect 5040 22448 5046 22460
rect 8573 22457 8585 22491
rect 8619 22488 8631 22491
rect 9858 22488 9864 22500
rect 8619 22460 9864 22488
rect 8619 22457 8631 22460
rect 8573 22451 8631 22457
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 2590 22380 2596 22432
rect 2648 22420 2654 22432
rect 2685 22423 2743 22429
rect 2685 22420 2697 22423
rect 2648 22392 2697 22420
rect 2648 22380 2654 22392
rect 2685 22389 2697 22392
rect 2731 22389 2743 22423
rect 2685 22383 2743 22389
rect 3418 22380 3424 22432
rect 3476 22420 3482 22432
rect 4338 22420 4344 22432
rect 3476 22392 4344 22420
rect 3476 22380 3482 22392
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 5258 22380 5264 22432
rect 5316 22380 5322 22432
rect 6178 22380 6184 22432
rect 6236 22380 6242 22432
rect 6730 22380 6736 22432
rect 6788 22420 6794 22432
rect 9585 22423 9643 22429
rect 9585 22420 9597 22423
rect 6788 22392 9597 22420
rect 6788 22380 6794 22392
rect 9585 22389 9597 22392
rect 9631 22389 9643 22423
rect 9585 22383 9643 22389
rect 1104 22330 10120 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 7950 22330
rect 8002 22278 8014 22330
rect 8066 22278 8078 22330
rect 8130 22278 8142 22330
rect 8194 22278 8206 22330
rect 8258 22278 10120 22330
rect 1104 22256 10120 22278
rect 3878 22176 3884 22228
rect 3936 22176 3942 22228
rect 6730 22176 6736 22228
rect 6788 22216 6794 22228
rect 6788 22188 6914 22216
rect 6788 22176 6794 22188
rect 1486 22040 1492 22092
rect 1544 22080 1550 22092
rect 1765 22083 1823 22089
rect 1765 22080 1777 22083
rect 1544 22052 1777 22080
rect 1544 22040 1550 22052
rect 1765 22049 1777 22052
rect 1811 22049 1823 22083
rect 1765 22043 1823 22049
rect 198 21972 204 22024
rect 256 22012 262 22024
rect 566 22012 572 22024
rect 256 21984 572 22012
rect 256 21972 262 21984
rect 566 21972 572 21984
rect 624 21972 630 22024
rect 1394 21972 1400 22024
rect 1452 22012 1458 22024
rect 1504 22012 1532 22040
rect 3896 22024 3924 22176
rect 4062 22108 4068 22160
rect 4120 22148 4126 22160
rect 4522 22148 4528 22160
rect 4120 22120 4528 22148
rect 4120 22108 4126 22120
rect 4522 22108 4528 22120
rect 4580 22108 4586 22160
rect 5258 22108 5264 22160
rect 5316 22108 5322 22160
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 5534 22080 5540 22092
rect 4212 22052 5540 22080
rect 4212 22040 4218 22052
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 5626 22040 5632 22092
rect 5684 22089 5690 22092
rect 5684 22083 5712 22089
rect 5700 22049 5712 22083
rect 5684 22043 5712 22049
rect 5684 22040 5690 22043
rect 6886 22024 6914 22188
rect 7006 22176 7012 22228
rect 7064 22176 7070 22228
rect 7466 22176 7472 22228
rect 7524 22176 7530 22228
rect 8294 22176 8300 22228
rect 8352 22216 8358 22228
rect 8389 22219 8447 22225
rect 8389 22216 8401 22219
rect 8352 22188 8401 22216
rect 8352 22176 8358 22188
rect 8389 22185 8401 22188
rect 8435 22185 8447 22219
rect 8389 22179 8447 22185
rect 7024 22080 7052 22176
rect 7190 22108 7196 22160
rect 7248 22148 7254 22160
rect 7484 22148 7512 22176
rect 7248 22120 7512 22148
rect 7248 22108 7254 22120
rect 9582 22108 9588 22160
rect 9640 22148 9646 22160
rect 10594 22148 10600 22160
rect 9640 22120 10600 22148
rect 9640 22108 9646 22120
rect 10594 22108 10600 22120
rect 10652 22108 10658 22160
rect 7926 22080 7932 22092
rect 7024 22052 7932 22080
rect 7926 22040 7932 22052
rect 7984 22040 7990 22092
rect 9398 22040 9404 22092
rect 9456 22080 9462 22092
rect 11146 22080 11152 22092
rect 9456 22052 11152 22080
rect 9456 22040 9462 22052
rect 11146 22040 11152 22052
rect 11204 22040 11210 22092
rect 1452 21984 1532 22012
rect 2041 22015 2099 22021
rect 1452 21972 1458 21984
rect 2041 21981 2053 22015
rect 2087 21981 2099 22015
rect 2041 21975 2099 21981
rect 1578 21904 1584 21956
rect 1636 21944 1642 21956
rect 2056 21944 2084 21975
rect 3234 21972 3240 22024
rect 3292 22012 3298 22024
rect 3510 22012 3516 22024
rect 3292 21984 3516 22012
rect 3292 21972 3298 21984
rect 3510 21972 3516 21984
rect 3568 21972 3574 22024
rect 3878 21972 3884 22024
rect 3936 21972 3942 22024
rect 4522 21972 4528 22024
rect 4580 22012 4586 22024
rect 4617 22015 4675 22021
rect 4617 22012 4629 22015
rect 4580 21984 4629 22012
rect 4580 21972 4586 21984
rect 4617 21981 4629 21984
rect 4663 21981 4675 22015
rect 4617 21975 4675 21981
rect 4798 21972 4804 22024
rect 4856 21972 4862 22024
rect 5810 21972 5816 22024
rect 5868 21972 5874 22024
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 22012 6515 22015
rect 6549 22015 6607 22021
rect 6549 22012 6561 22015
rect 6503 21984 6561 22012
rect 6503 21981 6515 21984
rect 6457 21975 6515 21981
rect 6549 21981 6561 21984
rect 6595 21981 6607 22015
rect 6549 21975 6607 21981
rect 6822 21972 6828 22024
rect 6880 21984 6914 22024
rect 6880 21972 6886 21984
rect 8202 21972 8208 22024
rect 8260 21972 8266 22024
rect 8478 21972 8484 22024
rect 8536 21972 8542 22024
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8812 21984 9137 22012
rect 8812 21972 8818 21984
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 9125 21975 9183 21981
rect 9214 21972 9220 22024
rect 9272 22012 9278 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 9272 21984 9505 22012
rect 9272 21972 9278 21984
rect 9493 21981 9505 21984
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 1636 21916 2084 21944
rect 1636 21904 1642 21916
rect 2222 21904 2228 21956
rect 2280 21944 2286 21956
rect 9858 21944 9864 21956
rect 2280 21916 3832 21944
rect 2280 21904 2286 21916
rect 2777 21879 2835 21885
rect 2777 21845 2789 21879
rect 2823 21876 2835 21879
rect 3694 21876 3700 21888
rect 2823 21848 3700 21876
rect 2823 21845 2835 21848
rect 2777 21839 2835 21845
rect 3694 21836 3700 21848
rect 3752 21836 3758 21888
rect 3804 21876 3832 21916
rect 8680 21916 9864 21944
rect 5442 21876 5448 21888
rect 3804 21848 5448 21876
rect 5442 21836 5448 21848
rect 5500 21836 5506 21888
rect 6733 21879 6791 21885
rect 6733 21845 6745 21879
rect 6779 21876 6791 21879
rect 7006 21876 7012 21888
rect 6779 21848 7012 21876
rect 6779 21845 6791 21848
rect 6733 21839 6791 21845
rect 7006 21836 7012 21848
rect 7064 21836 7070 21888
rect 8680 21885 8708 21916
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 8665 21879 8723 21885
rect 8665 21845 8677 21879
rect 8711 21845 8723 21879
rect 8665 21839 8723 21845
rect 8754 21836 8760 21888
rect 8812 21876 8818 21888
rect 9214 21876 9220 21888
rect 8812 21848 9220 21876
rect 8812 21836 8818 21848
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 9582 21876 9588 21888
rect 9355 21848 9588 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 9766 21876 9772 21888
rect 9723 21848 9772 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 1104 21786 10120 21808
rect 1104 21734 3010 21786
rect 3062 21734 3074 21786
rect 3126 21734 3138 21786
rect 3190 21734 3202 21786
rect 3254 21734 3266 21786
rect 3318 21734 9010 21786
rect 9062 21734 9074 21786
rect 9126 21734 9138 21786
rect 9190 21734 9202 21786
rect 9254 21734 9266 21786
rect 9318 21734 10120 21786
rect 1104 21712 10120 21734
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21672 2467 21675
rect 2455 21644 5396 21672
rect 2455 21641 2467 21644
rect 2409 21635 2467 21641
rect 1578 21564 1584 21616
rect 1636 21604 1642 21616
rect 1762 21604 1768 21616
rect 1636 21576 1768 21604
rect 1636 21564 1642 21576
rect 1762 21564 1768 21576
rect 1820 21564 1826 21616
rect 4356 21576 5304 21604
rect 1394 21536 1400 21548
rect 952 21508 1400 21536
rect 952 20992 980 21508
rect 1394 21496 1400 21508
rect 1452 21496 1458 21548
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 4356 21545 4384 21576
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21536 4491 21539
rect 4614 21536 4620 21548
rect 4479 21508 4620 21536
rect 4479 21505 4491 21508
rect 4433 21499 4491 21505
rect 4614 21496 4620 21508
rect 4672 21496 4678 21548
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21536 4767 21539
rect 4798 21536 4804 21548
rect 4755 21508 4804 21536
rect 4755 21505 4767 21508
rect 4709 21499 4767 21505
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 4982 21496 4988 21548
rect 5040 21536 5046 21548
rect 5040 21508 5120 21536
rect 5040 21496 5046 21508
rect 2590 21428 2596 21480
rect 2648 21468 2654 21480
rect 3326 21477 3332 21480
rect 3145 21471 3203 21477
rect 3145 21468 3157 21471
rect 2648 21440 3157 21468
rect 2648 21428 2654 21440
rect 3145 21437 3157 21440
rect 3191 21437 3203 21471
rect 3145 21431 3203 21437
rect 3304 21471 3332 21477
rect 3304 21437 3316 21471
rect 3304 21431 3332 21437
rect 3326 21428 3332 21431
rect 3384 21428 3390 21480
rect 3421 21471 3479 21477
rect 3421 21437 3433 21471
rect 3467 21468 3479 21471
rect 3467 21440 3648 21468
rect 3467 21437 3479 21440
rect 3421 21431 3479 21437
rect 3620 21400 3648 21440
rect 3694 21428 3700 21480
rect 3752 21428 3758 21480
rect 4154 21428 4160 21480
rect 4212 21428 4218 21480
rect 4338 21400 4344 21412
rect 3620 21372 4344 21400
rect 4338 21360 4344 21372
rect 4396 21360 4402 21412
rect 5092 21400 5120 21508
rect 5276 21468 5304 21576
rect 5368 21536 5396 21644
rect 5442 21632 5448 21684
rect 5500 21632 5506 21684
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 9309 21675 9367 21681
rect 9309 21672 9321 21675
rect 8260 21644 9321 21672
rect 8260 21632 8266 21644
rect 9309 21641 9321 21644
rect 9355 21641 9367 21675
rect 9309 21635 9367 21641
rect 9674 21632 9680 21684
rect 9732 21632 9738 21684
rect 7466 21564 7472 21616
rect 7524 21564 7530 21616
rect 5810 21536 5816 21548
rect 5368 21508 5816 21536
rect 5810 21496 5816 21508
rect 5868 21496 5874 21548
rect 7006 21496 7012 21548
rect 7064 21536 7070 21548
rect 7484 21536 7512 21564
rect 7064 21508 7512 21536
rect 7064 21496 7070 21508
rect 9398 21496 9404 21548
rect 9456 21536 9462 21548
rect 9493 21539 9551 21545
rect 9493 21536 9505 21539
rect 9456 21508 9505 21536
rect 9456 21496 9462 21508
rect 9493 21505 9505 21508
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 5350 21468 5356 21480
rect 5276 21440 5356 21468
rect 5350 21428 5356 21440
rect 5408 21428 5414 21480
rect 7466 21428 7472 21480
rect 7524 21428 7530 21480
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7616 21440 7665 21468
rect 7616 21428 7622 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 8389 21471 8447 21477
rect 8389 21468 8401 21471
rect 7653 21431 7711 21437
rect 8220 21440 8401 21468
rect 5534 21400 5540 21412
rect 5092 21372 5540 21400
rect 5534 21360 5540 21372
rect 5592 21360 5598 21412
rect 7668 21400 7696 21431
rect 8220 21412 8248 21440
rect 8389 21437 8401 21440
rect 8435 21437 8447 21471
rect 8389 21431 8447 21437
rect 8478 21428 8484 21480
rect 8536 21477 8542 21480
rect 8536 21471 8564 21477
rect 8552 21437 8564 21471
rect 8536 21431 8564 21437
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21468 8723 21471
rect 9030 21468 9036 21480
rect 8711 21440 9036 21468
rect 8711 21437 8723 21440
rect 8665 21431 8723 21437
rect 8536 21428 8542 21431
rect 9030 21428 9036 21440
rect 9088 21428 9094 21480
rect 7742 21400 7748 21412
rect 7668 21372 7748 21400
rect 7742 21360 7748 21372
rect 7800 21360 7806 21412
rect 8113 21403 8171 21409
rect 8113 21369 8125 21403
rect 8159 21369 8171 21403
rect 8113 21363 8171 21369
rect 1026 21292 1032 21344
rect 1084 21332 1090 21344
rect 1762 21332 1768 21344
rect 1084 21304 1768 21332
rect 1084 21292 1090 21304
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 2501 21335 2559 21341
rect 2501 21301 2513 21335
rect 2547 21332 2559 21335
rect 4062 21332 4068 21344
rect 2547 21304 4068 21332
rect 2547 21301 2559 21304
rect 2501 21295 2559 21301
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 4154 21292 4160 21344
rect 4212 21332 4218 21344
rect 8128 21332 8156 21363
rect 8202 21360 8208 21412
rect 8260 21360 8266 21412
rect 4212 21304 8156 21332
rect 4212 21292 4218 21304
rect 1104 21242 10120 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 7950 21242
rect 8002 21190 8014 21242
rect 8066 21190 8078 21242
rect 8130 21190 8142 21242
rect 8194 21190 8206 21242
rect 8258 21190 10120 21242
rect 1104 21168 10120 21190
rect 10226 21156 10232 21208
rect 10284 21196 10290 21208
rect 10686 21196 10692 21208
rect 10284 21168 10692 21196
rect 10284 21156 10290 21168
rect 10686 21156 10692 21168
rect 10744 21156 10750 21208
rect 3237 21131 3295 21137
rect 3237 21097 3249 21131
rect 3283 21128 3295 21131
rect 4154 21128 4160 21140
rect 3283 21100 4160 21128
rect 3283 21097 3295 21100
rect 3237 21091 3295 21097
rect 4154 21088 4160 21100
rect 4212 21088 4218 21140
rect 4246 21088 4252 21140
rect 4304 21088 4310 21140
rect 5074 21088 5080 21140
rect 5132 21088 5138 21140
rect 6454 21088 6460 21140
rect 6512 21128 6518 21140
rect 6638 21128 6644 21140
rect 6512 21100 6644 21128
rect 6512 21088 6518 21100
rect 6638 21088 6644 21100
rect 6696 21088 6702 21140
rect 8294 21128 8300 21140
rect 7116 21100 8300 21128
rect 3326 21020 3332 21072
rect 3384 21060 3390 21072
rect 3694 21060 3700 21072
rect 3384 21032 3700 21060
rect 3384 21020 3390 21032
rect 3694 21020 3700 21032
rect 3752 21020 3758 21072
rect 4338 21020 4344 21072
rect 4396 21060 4402 21072
rect 7116 21060 7144 21100
rect 4396 21032 7144 21060
rect 4396 21020 4402 21032
rect 2222 20992 2228 21004
rect 952 20964 2228 20992
rect 2222 20952 2228 20964
rect 2280 20952 2286 21004
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 4246 20992 4252 21004
rect 4028 20964 4252 20992
rect 4028 20952 4034 20964
rect 4246 20952 4252 20964
rect 4304 20952 4310 21004
rect 6454 20992 6460 21004
rect 4448 20964 6460 20992
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 1673 20927 1731 20933
rect 1673 20924 1685 20927
rect 1504 20896 1685 20924
rect 842 20816 848 20868
rect 900 20856 906 20868
rect 1504 20856 1532 20896
rect 1673 20893 1685 20896
rect 1719 20893 1731 20927
rect 1673 20887 1731 20893
rect 2498 20884 2504 20936
rect 2556 20884 2562 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 4448 20856 4476 20964
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 7558 20952 7564 21004
rect 7616 20952 7622 21004
rect 7668 20992 7696 21100
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 8754 21088 8760 21140
rect 8812 21128 8818 21140
rect 9398 21128 9404 21140
rect 8812 21100 9404 21128
rect 8812 21088 8818 21100
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 9674 21088 9680 21140
rect 9732 21088 9738 21140
rect 9309 21063 9367 21069
rect 9309 21029 9321 21063
rect 9355 21060 9367 21063
rect 10226 21060 10232 21072
rect 9355 21032 10232 21060
rect 9355 21029 9367 21032
rect 9309 21023 9367 21029
rect 10226 21020 10232 21032
rect 10284 21020 10290 21072
rect 7668 20964 7880 20992
rect 4798 20884 4804 20936
rect 4856 20924 4862 20936
rect 4893 20927 4951 20933
rect 4893 20924 4905 20927
rect 4856 20896 4905 20924
rect 4856 20884 4862 20896
rect 4893 20893 4905 20896
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 6917 20927 6975 20933
rect 6917 20893 6929 20927
rect 6963 20893 6975 20927
rect 6917 20887 6975 20893
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7190 20924 7196 20952
rect 7147 20900 7196 20924
rect 7248 20900 7254 20952
rect 7852 20933 7880 20964
rect 7926 20952 7932 21004
rect 7984 21001 7990 21004
rect 7984 20995 8012 21001
rect 8000 20961 8012 20995
rect 7984 20955 8012 20961
rect 7984 20952 7990 20955
rect 7837 20927 7895 20933
rect 7147 20896 7236 20900
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7837 20893 7849 20927
rect 7883 20893 7895 20927
rect 7837 20887 7895 20893
rect 900 20828 1532 20856
rect 1596 20828 4476 20856
rect 900 20816 906 20828
rect 1596 20797 1624 20828
rect 4522 20816 4528 20868
rect 4580 20856 4586 20868
rect 6270 20856 6276 20868
rect 4580 20828 6276 20856
rect 4580 20816 4586 20828
rect 6270 20816 6276 20828
rect 6328 20816 6334 20868
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20757 1639 20791
rect 1581 20751 1639 20757
rect 1854 20748 1860 20800
rect 1912 20748 1918 20800
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 4154 20788 4160 20800
rect 3936 20760 4160 20788
rect 3936 20748 3942 20760
rect 4154 20748 4160 20760
rect 4212 20748 4218 20800
rect 5166 20748 5172 20800
rect 5224 20788 5230 20800
rect 5810 20788 5816 20800
rect 5224 20760 5816 20788
rect 5224 20748 5230 20760
rect 5810 20748 5816 20760
rect 5868 20748 5874 20800
rect 6932 20788 6960 20887
rect 8110 20884 8116 20936
rect 8168 20884 8174 20936
rect 8754 20884 8760 20936
rect 8812 20924 8818 20936
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8812 20896 9137 20924
rect 8812 20884 8818 20896
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 9493 20927 9551 20933
rect 9493 20893 9505 20927
rect 9539 20924 9551 20927
rect 10042 20924 10048 20936
rect 9539 20896 10048 20924
rect 9539 20893 9551 20896
rect 9493 20887 9551 20893
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 8202 20788 8208 20800
rect 6932 20760 8208 20788
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 8570 20748 8576 20800
rect 8628 20788 8634 20800
rect 8757 20791 8815 20797
rect 8757 20788 8769 20791
rect 8628 20760 8769 20788
rect 8628 20748 8634 20760
rect 8757 20757 8769 20760
rect 8803 20757 8815 20791
rect 8757 20751 8815 20757
rect 1104 20698 10120 20720
rect 1104 20646 3010 20698
rect 3062 20646 3074 20698
rect 3126 20646 3138 20698
rect 3190 20646 3202 20698
rect 3254 20646 3266 20698
rect 3318 20646 9010 20698
rect 9062 20646 9074 20698
rect 9126 20646 9138 20698
rect 9190 20646 9202 20698
rect 9254 20646 9266 20698
rect 9318 20646 10120 20698
rect 1104 20624 10120 20646
rect 1762 20544 1768 20596
rect 1820 20584 1826 20596
rect 3786 20584 3792 20596
rect 1820 20556 3792 20584
rect 1820 20544 1826 20556
rect 3786 20544 3792 20556
rect 3844 20544 3850 20596
rect 7653 20587 7711 20593
rect 7653 20553 7665 20587
rect 7699 20584 7711 20587
rect 8110 20584 8116 20596
rect 7699 20556 8116 20584
rect 7699 20553 7711 20556
rect 7653 20547 7711 20553
rect 8110 20544 8116 20556
rect 8168 20544 8174 20596
rect 8662 20544 8668 20596
rect 8720 20544 8726 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 3602 20476 3608 20528
rect 3660 20516 3666 20528
rect 6270 20516 6276 20528
rect 3660 20488 6276 20516
rect 3660 20476 3666 20488
rect 6270 20476 6276 20488
rect 6328 20476 6334 20528
rect 7282 20476 7288 20528
rect 7340 20516 7346 20528
rect 9582 20516 9588 20528
rect 7340 20488 9588 20516
rect 7340 20476 7346 20488
rect 9582 20476 9588 20488
rect 9640 20476 9646 20528
rect 1946 20408 1952 20460
rect 2004 20448 2010 20460
rect 2133 20451 2191 20457
rect 2133 20448 2145 20451
rect 2004 20420 2145 20448
rect 2004 20408 2010 20420
rect 2133 20417 2145 20420
rect 2179 20448 2191 20451
rect 3878 20448 3884 20460
rect 2179 20420 3884 20448
rect 2179 20417 2191 20420
rect 2133 20411 2191 20417
rect 3878 20408 3884 20420
rect 3936 20408 3942 20460
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 6917 20451 6975 20457
rect 6917 20448 6929 20451
rect 6512 20420 6929 20448
rect 6512 20408 6518 20420
rect 6917 20417 6929 20420
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 7190 20408 7196 20460
rect 7248 20448 7254 20460
rect 7742 20448 7748 20460
rect 7248 20420 7748 20448
rect 7248 20408 7254 20420
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20448 8539 20451
rect 8570 20448 8576 20460
rect 8527 20420 8576 20448
rect 8527 20417 8539 20420
rect 8481 20411 8539 20417
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 8757 20451 8815 20457
rect 8757 20417 8769 20451
rect 8803 20417 8815 20451
rect 8757 20411 8815 20417
rect 6362 20340 6368 20392
rect 6420 20380 6426 20392
rect 6641 20383 6699 20389
rect 6641 20380 6653 20383
rect 6420 20352 6653 20380
rect 6420 20340 6426 20352
rect 6641 20349 6653 20352
rect 6687 20349 6699 20383
rect 6641 20343 6699 20349
rect 7282 20340 7288 20392
rect 7340 20380 7346 20392
rect 8772 20380 8800 20411
rect 9030 20408 9036 20460
rect 9088 20448 9094 20460
rect 9125 20451 9183 20457
rect 9125 20448 9137 20451
rect 9088 20420 9137 20448
rect 9088 20408 9094 20420
rect 9125 20417 9137 20420
rect 9171 20417 9183 20451
rect 9125 20411 9183 20417
rect 9214 20408 9220 20460
rect 9272 20448 9278 20460
rect 9493 20451 9551 20457
rect 9493 20448 9505 20451
rect 9272 20420 9505 20448
rect 9272 20408 9278 20420
rect 9493 20417 9505 20420
rect 9539 20417 9551 20451
rect 9493 20411 9551 20417
rect 7340 20352 8800 20380
rect 7340 20340 7346 20352
rect 8938 20340 8944 20392
rect 8996 20380 9002 20392
rect 9766 20380 9772 20392
rect 8996 20352 9772 20380
rect 8996 20340 9002 20352
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 1854 20272 1860 20324
rect 1912 20312 1918 20324
rect 5166 20312 5172 20324
rect 1912 20284 5172 20312
rect 1912 20272 1918 20284
rect 5166 20272 5172 20284
rect 5224 20272 5230 20324
rect 7650 20272 7656 20324
rect 7708 20312 7714 20324
rect 7926 20312 7932 20324
rect 7708 20284 7932 20312
rect 7708 20272 7714 20284
rect 7926 20272 7932 20284
rect 7984 20272 7990 20324
rect 9309 20315 9367 20321
rect 9309 20281 9321 20315
rect 9355 20312 9367 20315
rect 10226 20312 10232 20324
rect 9355 20284 10232 20312
rect 9355 20281 9367 20284
rect 9309 20275 9367 20281
rect 10226 20272 10232 20284
rect 10284 20272 10290 20324
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 1949 20247 2007 20253
rect 1949 20244 1961 20247
rect 1820 20216 1961 20244
rect 1820 20204 1826 20216
rect 1949 20213 1961 20216
rect 1995 20244 2007 20247
rect 2038 20244 2044 20256
rect 1995 20216 2044 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 8941 20247 8999 20253
rect 8941 20213 8953 20247
rect 8987 20244 8999 20247
rect 10042 20244 10048 20256
rect 8987 20216 10048 20244
rect 8987 20213 8999 20216
rect 8941 20207 8999 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 1104 20154 10120 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 7950 20154
rect 8002 20102 8014 20154
rect 8066 20102 8078 20154
rect 8130 20102 8142 20154
rect 8194 20102 8206 20154
rect 8258 20102 10120 20154
rect 1104 20080 10120 20102
rect 1394 20000 1400 20052
rect 1452 20040 1458 20052
rect 2590 20040 2596 20052
rect 1452 20012 2596 20040
rect 1452 20000 1458 20012
rect 2590 20000 2596 20012
rect 2648 20040 2654 20052
rect 2648 20012 2774 20040
rect 2648 20000 2654 20012
rect 1762 19864 1768 19916
rect 1820 19864 1826 19916
rect 2746 19904 2774 20012
rect 4522 20000 4528 20052
rect 4580 20000 4586 20052
rect 7377 20043 7435 20049
rect 7377 20009 7389 20043
rect 7423 20040 7435 20043
rect 7558 20040 7564 20052
rect 7423 20012 7564 20040
rect 7423 20009 7435 20012
rect 7377 20003 7435 20009
rect 7558 20000 7564 20012
rect 7616 20000 7622 20052
rect 8754 20000 8760 20052
rect 8812 20000 8818 20052
rect 9674 20000 9680 20052
rect 9732 20000 9738 20052
rect 9309 19975 9367 19981
rect 9309 19941 9321 19975
rect 9355 19972 9367 19975
rect 10226 19972 10232 19984
rect 9355 19944 10232 19972
rect 9355 19941 9367 19944
rect 9309 19935 9367 19941
rect 10226 19932 10232 19944
rect 10284 19932 10290 19984
rect 6362 19904 6368 19916
rect 2746 19876 6368 19904
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 1394 19796 1400 19848
rect 1452 19796 1458 19848
rect 1780 19768 1808 19864
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19836 2099 19839
rect 2498 19836 2504 19848
rect 2087 19808 2504 19836
rect 2087 19805 2099 19808
rect 2041 19799 2099 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 2866 19796 2872 19848
rect 2924 19836 2930 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 2924 19808 4353 19836
rect 2924 19796 2930 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 5166 19796 5172 19848
rect 5224 19836 5230 19848
rect 5994 19836 6000 19848
rect 5224 19808 6000 19836
rect 5224 19796 5230 19808
rect 5994 19796 6000 19808
rect 6052 19836 6058 19848
rect 6638 19836 6644 19848
rect 6052 19808 6644 19836
rect 6052 19796 6058 19808
rect 6638 19796 6644 19808
rect 6696 19796 6702 19848
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19805 7527 19839
rect 7469 19799 7527 19805
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19805 7803 19839
rect 7745 19799 7803 19805
rect 7484 19768 7512 19799
rect 7558 19768 7564 19780
rect 1780 19740 2544 19768
rect 7484 19740 7564 19768
rect 2516 19712 2544 19740
rect 7558 19728 7564 19740
rect 7616 19728 7622 19780
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 1762 19700 1768 19712
rect 1627 19672 1768 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 2498 19660 2504 19712
rect 2556 19660 2562 19712
rect 2777 19703 2835 19709
rect 2777 19669 2789 19703
rect 2823 19700 2835 19703
rect 4062 19700 4068 19712
rect 2823 19672 4068 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 6454 19660 6460 19712
rect 6512 19700 6518 19712
rect 7760 19700 7788 19799
rect 8570 19796 8576 19848
rect 8628 19796 8634 19848
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 10502 19836 10508 19848
rect 9539 19808 10508 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 7926 19728 7932 19780
rect 7984 19768 7990 19780
rect 9214 19768 9220 19780
rect 7984 19740 9220 19768
rect 7984 19728 7990 19740
rect 9214 19728 9220 19740
rect 9272 19728 9278 19780
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10410 19768 10416 19780
rect 9916 19740 10416 19768
rect 9916 19728 9922 19740
rect 10410 19728 10416 19740
rect 10468 19728 10474 19780
rect 6512 19672 7788 19700
rect 8481 19703 8539 19709
rect 6512 19660 6518 19672
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8754 19700 8760 19712
rect 8527 19672 8760 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 1104 19610 10120 19632
rect 1104 19558 3010 19610
rect 3062 19558 3074 19610
rect 3126 19558 3138 19610
rect 3190 19558 3202 19610
rect 3254 19558 3266 19610
rect 3318 19558 9010 19610
rect 9062 19558 9074 19610
rect 9126 19558 9138 19610
rect 9190 19558 9202 19610
rect 9254 19558 9266 19610
rect 9318 19558 10120 19610
rect 1104 19536 10120 19558
rect 2866 19456 2872 19508
rect 2924 19456 2930 19508
rect 4985 19499 5043 19505
rect 4985 19465 4997 19499
rect 5031 19496 5043 19499
rect 7282 19496 7288 19508
rect 5031 19468 7288 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 7926 19496 7932 19508
rect 7392 19468 7932 19496
rect 2498 19428 2504 19440
rect 1596 19400 2504 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 1596 19292 1624 19400
rect 2498 19388 2504 19400
rect 2556 19388 2562 19440
rect 7392 19428 7420 19468
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 8628 19468 9413 19496
rect 8628 19456 8634 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9401 19459 9459 19465
rect 9674 19456 9680 19508
rect 9732 19456 9738 19508
rect 4908 19400 7420 19428
rect 1670 19320 1676 19372
rect 1728 19360 1734 19372
rect 2041 19363 2099 19369
rect 2041 19360 2053 19363
rect 1728 19332 2053 19360
rect 1728 19320 1734 19332
rect 2041 19329 2053 19332
rect 2087 19329 2099 19363
rect 2041 19323 2099 19329
rect 3602 19320 3608 19372
rect 3660 19369 3666 19372
rect 3660 19363 3709 19369
rect 3660 19329 3663 19363
rect 3697 19329 3709 19363
rect 3660 19323 3709 19329
rect 3660 19320 3666 19323
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 4801 19363 4859 19369
rect 4801 19360 4813 19363
rect 4396 19332 4813 19360
rect 4396 19320 4402 19332
rect 4801 19329 4813 19332
rect 4847 19329 4859 19363
rect 4801 19323 4859 19329
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1596 19264 1777 19292
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 3513 19295 3571 19301
rect 3513 19292 3525 19295
rect 1765 19255 1823 19261
rect 2792 19264 3525 19292
rect 2792 19233 2820 19264
rect 3513 19261 3525 19264
rect 3559 19261 3571 19295
rect 3513 19255 3571 19261
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 3835 19264 4016 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 2777 19227 2835 19233
rect 2777 19193 2789 19227
rect 2823 19193 2835 19227
rect 2777 19187 2835 19193
rect 3988 19224 4016 19264
rect 4062 19252 4068 19304
rect 4120 19252 4126 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 4614 19292 4620 19304
rect 4571 19264 4620 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 4614 19252 4620 19264
rect 4672 19252 4678 19304
rect 4706 19252 4712 19304
rect 4764 19252 4770 19304
rect 4798 19224 4804 19236
rect 3988 19196 4804 19224
rect 1578 19116 1584 19168
rect 1636 19116 1642 19168
rect 3694 19116 3700 19168
rect 3752 19156 3758 19168
rect 3988 19156 4016 19196
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 3752 19128 4016 19156
rect 3752 19116 3758 19128
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4908 19156 4936 19400
rect 7742 19388 7748 19440
rect 7800 19388 7806 19440
rect 6270 19320 6276 19372
rect 6328 19360 6334 19372
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 6328 19332 6377 19360
rect 6328 19320 6334 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6638 19320 6644 19372
rect 6696 19320 6702 19372
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7561 19363 7619 19369
rect 7561 19360 7573 19363
rect 7524 19332 7573 19360
rect 7524 19320 7530 19332
rect 7561 19329 7573 19332
rect 7607 19329 7619 19363
rect 7760 19360 7788 19388
rect 8481 19363 8539 19369
rect 7760 19332 7880 19360
rect 7561 19323 7619 19329
rect 7742 19252 7748 19304
rect 7800 19252 7806 19304
rect 7852 19292 7880 19332
rect 8481 19329 8493 19363
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 7926 19292 7932 19304
rect 7852 19264 7932 19292
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8496 19292 8524 19323
rect 9490 19320 9496 19372
rect 9548 19320 9554 19372
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 10686 19360 10692 19372
rect 10376 19332 10692 19360
rect 10376 19320 10382 19332
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 8312 19264 8524 19292
rect 7377 19227 7435 19233
rect 7377 19193 7389 19227
rect 7423 19224 7435 19227
rect 8205 19227 8263 19233
rect 8205 19224 8217 19227
rect 7423 19196 8217 19224
rect 7423 19193 7435 19196
rect 7377 19187 7435 19193
rect 8205 19193 8217 19196
rect 8251 19193 8263 19227
rect 8205 19187 8263 19193
rect 4120 19128 4936 19156
rect 4120 19116 4126 19128
rect 5902 19116 5908 19168
rect 5960 19156 5966 19168
rect 7190 19156 7196 19168
rect 5960 19128 7196 19156
rect 5960 19116 5966 19128
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 8312 19156 8340 19264
rect 8570 19252 8576 19304
rect 8628 19301 8634 19304
rect 8628 19295 8656 19301
rect 8644 19261 8656 19295
rect 8628 19255 8656 19261
rect 8757 19295 8815 19301
rect 8757 19261 8769 19295
rect 8803 19292 8815 19295
rect 9122 19292 9128 19304
rect 8803 19264 9128 19292
rect 8803 19261 8815 19264
rect 8757 19255 8815 19261
rect 8628 19252 8634 19255
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 9398 19252 9404 19304
rect 9456 19292 9462 19304
rect 10870 19292 10876 19304
rect 9456 19264 10876 19292
rect 9456 19252 9462 19264
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 10042 19224 10048 19236
rect 9140 19196 10048 19224
rect 8662 19156 8668 19168
rect 8312 19128 8668 19156
rect 8662 19116 8668 19128
rect 8720 19156 8726 19168
rect 9140 19156 9168 19196
rect 10042 19184 10048 19196
rect 10100 19184 10106 19236
rect 8720 19128 9168 19156
rect 8720 19116 8726 19128
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 9858 19156 9864 19168
rect 9640 19128 9864 19156
rect 9640 19116 9646 19128
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 1104 19066 10120 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 7950 19066
rect 8002 19014 8014 19066
rect 8066 19014 8078 19066
rect 8130 19014 8142 19066
rect 8194 19014 8206 19066
rect 8258 19014 10120 19066
rect 1104 18992 10120 19014
rect 3789 18955 3847 18961
rect 3789 18921 3801 18955
rect 3835 18952 3847 18955
rect 4338 18952 4344 18964
rect 3835 18924 4344 18952
rect 3835 18921 3847 18924
rect 3789 18915 3847 18921
rect 4338 18912 4344 18924
rect 4396 18912 4402 18964
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 4764 18924 5672 18952
rect 4764 18912 4770 18924
rect 2961 18887 3019 18893
rect 2961 18853 2973 18887
rect 3007 18884 3019 18887
rect 3878 18884 3884 18896
rect 3007 18856 3884 18884
rect 3007 18853 3019 18856
rect 2961 18847 3019 18853
rect 3878 18844 3884 18856
rect 3936 18844 3942 18896
rect 5074 18884 5080 18896
rect 4908 18856 5080 18884
rect 1670 18776 1676 18828
rect 1728 18816 1734 18828
rect 1946 18816 1952 18828
rect 1728 18788 1952 18816
rect 1728 18776 1734 18788
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 3694 18776 3700 18828
rect 3752 18816 3758 18828
rect 4571 18819 4629 18825
rect 4571 18816 4583 18819
rect 3752 18788 4583 18816
rect 3752 18776 3758 18788
rect 4571 18785 4583 18788
rect 4617 18785 4629 18819
rect 4571 18779 4629 18785
rect 4706 18776 4712 18828
rect 4764 18816 4770 18828
rect 4908 18816 4936 18856
rect 5074 18844 5080 18856
rect 5132 18844 5138 18896
rect 5166 18844 5172 18896
rect 5224 18844 5230 18896
rect 4764 18788 4936 18816
rect 4985 18819 5043 18825
rect 4764 18776 4770 18788
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5184 18816 5212 18844
rect 5644 18825 5672 18924
rect 5902 18912 5908 18964
rect 5960 18912 5966 18964
rect 6822 18912 6828 18964
rect 6880 18952 6886 18964
rect 6880 18924 7604 18952
rect 6880 18912 6886 18924
rect 7576 18884 7604 18924
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 8205 18955 8263 18961
rect 8205 18952 8217 18955
rect 7892 18924 8217 18952
rect 7892 18912 7898 18924
rect 8205 18921 8217 18924
rect 8251 18921 8263 18955
rect 8205 18915 8263 18921
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 8570 18952 8576 18964
rect 8352 18924 8576 18952
rect 8352 18912 8358 18924
rect 8570 18912 8576 18924
rect 8628 18912 8634 18964
rect 9674 18912 9680 18964
rect 9732 18912 9738 18964
rect 9030 18884 9036 18896
rect 7576 18856 9036 18884
rect 9030 18844 9036 18856
rect 9088 18844 9094 18896
rect 9217 18887 9275 18893
rect 9217 18853 9229 18887
rect 9263 18884 9275 18887
rect 10226 18884 10232 18896
rect 9263 18856 10232 18884
rect 9263 18853 9275 18856
rect 9217 18847 9275 18853
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 5031 18788 5212 18816
rect 5629 18819 5687 18825
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5629 18785 5641 18819
rect 5675 18816 5687 18819
rect 5902 18816 5908 18828
rect 5675 18788 5908 18816
rect 5675 18785 5687 18788
rect 5629 18779 5687 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 9858 18816 9864 18828
rect 8404 18788 9864 18816
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18748 2283 18751
rect 3602 18748 3608 18760
rect 2271 18720 3608 18748
rect 2271 18717 2283 18720
rect 2225 18711 2283 18717
rect 1486 18640 1492 18692
rect 1544 18680 1550 18692
rect 2240 18680 2268 18711
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 4430 18708 4436 18760
rect 4488 18708 4494 18760
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 5810 18748 5816 18760
rect 5767 18720 5816 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 1544 18652 2268 18680
rect 5460 18680 5488 18711
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 6362 18708 6368 18760
rect 6420 18748 6426 18760
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6420 18720 6929 18748
rect 6420 18708 6426 18720
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7098 18708 7104 18760
rect 7156 18748 7162 18760
rect 8404 18757 8432 18788
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 7193 18751 7251 18757
rect 7193 18748 7205 18751
rect 7156 18720 7205 18748
rect 7156 18708 7162 18720
rect 7193 18717 7205 18720
rect 7239 18717 7251 18751
rect 7193 18711 7251 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 8487 18751 8545 18757
rect 8487 18717 8499 18751
rect 8533 18717 8545 18751
rect 8487 18711 8545 18717
rect 7558 18680 7564 18692
rect 5460 18652 7564 18680
rect 1544 18640 1550 18652
rect 7558 18640 7564 18652
rect 7616 18640 7622 18692
rect 8502 18680 8530 18711
rect 9030 18708 9036 18760
rect 9088 18748 9094 18760
rect 9401 18751 9459 18757
rect 9401 18748 9413 18751
rect 9088 18720 9413 18748
rect 9088 18708 9094 18720
rect 9401 18717 9413 18720
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9674 18748 9680 18760
rect 9539 18720 9680 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10226 18748 10232 18760
rect 10008 18720 10232 18748
rect 10008 18708 10014 18720
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 8754 18680 8760 18692
rect 7668 18652 8530 18680
rect 8588 18652 8760 18680
rect 2958 18572 2964 18624
rect 3016 18612 3022 18624
rect 3694 18612 3700 18624
rect 3016 18584 3700 18612
rect 3016 18572 3022 18584
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 7668 18612 7696 18652
rect 4764 18584 7696 18612
rect 7929 18615 7987 18621
rect 4764 18572 4770 18584
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8588 18612 8616 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 7975 18584 8616 18612
rect 8665 18615 8723 18621
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8665 18581 8677 18615
rect 8711 18612 8723 18615
rect 9950 18612 9956 18624
rect 8711 18584 9956 18612
rect 8711 18581 8723 18584
rect 8665 18575 8723 18581
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 1104 18522 10120 18544
rect 1104 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 3202 18522
rect 3254 18470 3266 18522
rect 3318 18470 9010 18522
rect 9062 18470 9074 18522
rect 9126 18470 9138 18522
rect 9190 18470 9202 18522
rect 9254 18470 9266 18522
rect 9318 18470 10120 18522
rect 1104 18448 10120 18470
rect 1302 18368 1308 18420
rect 1360 18408 1366 18420
rect 4709 18411 4767 18417
rect 4709 18408 4721 18411
rect 1360 18380 4721 18408
rect 1360 18368 1366 18380
rect 4709 18377 4721 18380
rect 4755 18377 4767 18411
rect 4709 18371 4767 18377
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6236 18380 9536 18408
rect 6236 18368 6242 18380
rect 382 18300 388 18352
rect 440 18340 446 18352
rect 658 18340 664 18352
rect 440 18312 664 18340
rect 440 18300 446 18312
rect 658 18300 664 18312
rect 716 18300 722 18352
rect 2774 18340 2780 18352
rect 1320 18312 2780 18340
rect 1320 18284 1348 18312
rect 2774 18300 2780 18312
rect 2832 18340 2838 18352
rect 3421 18343 3479 18349
rect 3421 18340 3433 18343
rect 2832 18312 3433 18340
rect 2832 18300 2838 18312
rect 3421 18309 3433 18312
rect 3467 18309 3479 18343
rect 3421 18303 3479 18309
rect 198 18232 204 18284
rect 256 18232 262 18284
rect 1302 18232 1308 18284
rect 1360 18232 1366 18284
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1673 18235 1731 18241
rect 216 18080 244 18232
rect 658 18164 664 18216
rect 716 18204 722 18216
rect 1688 18204 1716 18235
rect 1946 18232 1952 18284
rect 2004 18272 2010 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 2004 18244 2053 18272
rect 2004 18232 2010 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2406 18272 2412 18284
rect 2363 18244 2412 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 716 18176 1716 18204
rect 716 18164 722 18176
rect 1762 18164 1768 18216
rect 1820 18204 1826 18216
rect 1820 18176 1900 18204
rect 1820 18164 1826 18176
rect 1486 18096 1492 18148
rect 1544 18136 1550 18148
rect 1670 18136 1676 18148
rect 1544 18108 1676 18136
rect 1544 18096 1550 18108
rect 1670 18096 1676 18108
rect 1728 18096 1734 18148
rect 1872 18145 1900 18176
rect 1857 18139 1915 18145
rect 1857 18105 1869 18139
rect 1903 18105 1915 18139
rect 1857 18099 1915 18105
rect 198 18028 204 18080
rect 256 18028 262 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 1044 18040 1593 18068
rect 1044 17796 1072 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 2056 18068 2084 18235
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 5399 18244 6377 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 6365 18241 6377 18244
rect 6411 18272 6423 18275
rect 6546 18272 6552 18284
rect 6411 18244 6552 18272
rect 6411 18241 6423 18244
rect 6365 18235 6423 18241
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 7006 18272 7012 18284
rect 6696 18244 7012 18272
rect 6696 18232 6702 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 7432 18244 7880 18272
rect 7432 18232 7438 18244
rect 7558 18164 7564 18216
rect 7616 18164 7622 18216
rect 7742 18164 7748 18216
rect 7800 18164 7806 18216
rect 7852 18204 7880 18244
rect 8754 18232 8760 18284
rect 8812 18232 8818 18284
rect 9508 18281 9536 18380
rect 9674 18368 9680 18420
rect 9732 18368 9738 18420
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 8205 18207 8263 18213
rect 8205 18204 8217 18207
rect 7852 18176 8217 18204
rect 8205 18173 8217 18176
rect 8251 18173 8263 18207
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8205 18167 8263 18173
rect 8312 18176 8493 18204
rect 3053 18139 3111 18145
rect 3053 18105 3065 18139
rect 3099 18136 3111 18139
rect 4430 18136 4436 18148
rect 3099 18108 4436 18136
rect 3099 18105 3111 18108
rect 3053 18099 3111 18105
rect 4430 18096 4436 18108
rect 4488 18096 4494 18148
rect 5537 18139 5595 18145
rect 5537 18105 5549 18139
rect 5583 18136 5595 18139
rect 6362 18136 6368 18148
rect 5583 18108 6368 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 6362 18096 6368 18108
rect 6420 18096 6426 18148
rect 7576 18136 7604 18164
rect 7300 18108 7604 18136
rect 7300 18080 7328 18108
rect 8110 18096 8116 18148
rect 8168 18136 8174 18148
rect 8312 18136 8340 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 8570 18164 8576 18216
rect 8628 18213 8634 18216
rect 8628 18207 8656 18213
rect 8644 18173 8656 18207
rect 8628 18167 8656 18173
rect 8628 18164 8634 18167
rect 8168 18108 8340 18136
rect 8168 18096 8174 18108
rect 2682 18068 2688 18080
rect 2056 18040 2688 18068
rect 1581 18031 1639 18037
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 5350 18068 5356 18080
rect 4856 18040 5356 18068
rect 4856 18028 4862 18040
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 7282 18028 7288 18080
rect 7340 18028 7346 18080
rect 7377 18071 7435 18077
rect 7377 18037 7389 18071
rect 7423 18068 7435 18071
rect 7834 18068 7840 18080
rect 7423 18040 7840 18068
rect 7423 18037 7435 18040
rect 7377 18031 7435 18037
rect 7834 18028 7840 18040
rect 7892 18028 7898 18080
rect 8846 18028 8852 18080
rect 8904 18068 8910 18080
rect 9401 18071 9459 18077
rect 9401 18068 9413 18071
rect 8904 18040 9413 18068
rect 8904 18028 8910 18040
rect 9401 18037 9413 18040
rect 9447 18037 9459 18071
rect 9401 18031 9459 18037
rect 1104 17978 10120 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 7950 17978
rect 8002 17926 8014 17978
rect 8066 17926 8078 17978
rect 8130 17926 8142 17978
rect 8194 17926 8206 17978
rect 8258 17926 10120 17978
rect 1104 17904 10120 17926
rect 1210 17824 1216 17876
rect 1268 17864 1274 17876
rect 1670 17864 1676 17876
rect 1268 17836 1676 17864
rect 1268 17824 1274 17836
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 2501 17867 2559 17873
rect 2501 17833 2513 17867
rect 2547 17864 2559 17867
rect 2774 17864 2780 17876
rect 2547 17836 2780 17864
rect 2547 17833 2559 17836
rect 2501 17827 2559 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 6270 17824 6276 17876
rect 6328 17824 6334 17876
rect 6730 17824 6736 17876
rect 6788 17824 6794 17876
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7558 17864 7564 17876
rect 7055 17836 7564 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 8481 17867 8539 17873
rect 8481 17833 8493 17867
rect 8527 17864 8539 17867
rect 9398 17864 9404 17876
rect 8527 17836 9404 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 8113 17799 8171 17805
rect 1044 17768 1624 17796
rect 1210 17620 1216 17672
rect 1268 17660 1274 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 1268 17632 1409 17660
rect 1268 17620 1274 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1596 17660 1624 17768
rect 8113 17765 8125 17799
rect 8159 17796 8171 17799
rect 8754 17796 8760 17808
rect 8159 17768 8760 17796
rect 8159 17765 8171 17768
rect 8113 17759 8171 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 3418 17728 3424 17740
rect 1719 17700 3424 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 3418 17688 3424 17700
rect 3476 17688 3482 17740
rect 6362 17688 6368 17740
rect 6420 17728 6426 17740
rect 7101 17731 7159 17737
rect 7101 17728 7113 17731
rect 6420 17700 7113 17728
rect 6420 17688 6426 17700
rect 7101 17697 7113 17700
rect 7147 17697 7159 17731
rect 7101 17691 7159 17697
rect 8220 17700 8984 17728
rect 1762 17660 1768 17672
rect 1596 17632 1768 17660
rect 1397 17623 1455 17629
rect 1762 17620 1768 17632
rect 1820 17620 1826 17672
rect 1946 17620 1952 17672
rect 2004 17660 2010 17672
rect 2222 17660 2228 17672
rect 2004 17632 2228 17660
rect 2004 17620 2010 17632
rect 2222 17620 2228 17632
rect 2280 17660 2286 17672
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 2280 17632 2329 17660
rect 2280 17620 2286 17632
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 5994 17620 6000 17672
rect 6052 17660 6058 17672
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 6052 17632 6101 17660
rect 6052 17620 6058 17632
rect 6089 17629 6101 17632
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 6454 17620 6460 17672
rect 6512 17660 6518 17672
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 6512 17632 6561 17660
rect 6512 17620 6518 17632
rect 6549 17629 6561 17632
rect 6595 17629 6607 17663
rect 6549 17623 6607 17629
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17629 6883 17663
rect 6825 17623 6883 17629
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17660 7435 17663
rect 7650 17660 7656 17672
rect 7423 17632 7656 17660
rect 7423 17629 7435 17632
rect 7377 17623 7435 17629
rect 3326 17552 3332 17604
rect 3384 17592 3390 17604
rect 5166 17592 5172 17604
rect 3384 17564 5172 17592
rect 3384 17552 3390 17564
rect 5166 17552 5172 17564
rect 5224 17552 5230 17604
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 2501 17527 2559 17533
rect 2501 17524 2513 17527
rect 1452 17496 2513 17524
rect 1452 17484 1458 17496
rect 2501 17493 2513 17496
rect 2547 17493 2559 17527
rect 6564 17524 6592 17623
rect 6840 17592 6868 17623
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 8220 17592 8248 17700
rect 8294 17620 8300 17672
rect 8352 17620 8358 17672
rect 8386 17620 8392 17672
rect 8444 17620 8450 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 8846 17660 8852 17672
rect 8619 17632 8852 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8846 17620 8852 17632
rect 8904 17620 8910 17672
rect 8956 17660 8984 17700
rect 9030 17688 9036 17740
rect 9088 17728 9094 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 9088 17700 9505 17728
rect 9088 17688 9094 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 9766 17688 9772 17740
rect 9824 17688 9830 17740
rect 9674 17660 9680 17672
rect 8956 17632 9680 17660
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 6840 17564 8248 17592
rect 8404 17592 8432 17620
rect 8404 17564 8800 17592
rect 7006 17524 7012 17536
rect 6564 17496 7012 17524
rect 2501 17487 2559 17493
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 7190 17484 7196 17536
rect 7248 17524 7254 17536
rect 8386 17524 8392 17536
rect 7248 17496 8392 17524
rect 7248 17484 7254 17496
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 8772 17533 8800 17564
rect 8757 17527 8815 17533
rect 8757 17493 8769 17527
rect 8803 17493 8815 17527
rect 8757 17487 8815 17493
rect 934 17416 940 17468
rect 992 17416 998 17468
rect 1104 17434 10120 17456
rect 952 17128 980 17416
rect 1104 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 3202 17434
rect 3254 17382 3266 17434
rect 3318 17382 9010 17434
rect 9062 17382 9074 17434
rect 9126 17382 9138 17434
rect 9190 17382 9202 17434
rect 9254 17382 9266 17434
rect 9318 17382 10120 17434
rect 1104 17360 10120 17382
rect 2958 17320 2964 17332
rect 2700 17292 2964 17320
rect 1486 17212 1492 17264
rect 1544 17212 1550 17264
rect 1394 17144 1400 17196
rect 1452 17144 1458 17196
rect 1504 17184 1532 17212
rect 2700 17193 2728 17292
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 3694 17280 3700 17332
rect 3752 17320 3758 17332
rect 4338 17320 4344 17332
rect 3752 17292 4344 17320
rect 3752 17280 3758 17292
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 5074 17280 5080 17332
rect 5132 17320 5138 17332
rect 7558 17320 7564 17332
rect 5132 17292 7564 17320
rect 5132 17280 5138 17292
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 8352 17292 9413 17320
rect 8352 17280 8358 17292
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 9490 17212 9496 17264
rect 9548 17212 9554 17264
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 10962 17252 10968 17264
rect 9640 17224 10968 17252
rect 9640 17212 9646 17224
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 1504 17156 1685 17184
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2685 17187 2743 17193
rect 2685 17153 2697 17187
rect 2731 17153 2743 17187
rect 2685 17147 2743 17153
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4433 17187 4491 17193
rect 4433 17184 4445 17187
rect 4387 17156 4445 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4433 17153 4445 17156
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 934 17076 940 17128
rect 992 17076 998 17128
rect 2498 17076 2504 17128
rect 2556 17076 2562 17128
rect 3436 17116 3464 17147
rect 7098 17144 7104 17196
rect 7156 17184 7162 17196
rect 7742 17184 7748 17196
rect 7156 17156 7748 17184
rect 7156 17144 7162 17156
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 3602 17125 3608 17128
rect 3252 17088 3464 17116
rect 3559 17119 3608 17125
rect 3252 17060 3280 17088
rect 3559 17085 3571 17119
rect 3605 17085 3608 17119
rect 3559 17079 3608 17085
rect 3602 17076 3608 17079
rect 3660 17076 3666 17128
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 3743 17088 4108 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 2774 17008 2780 17060
rect 2832 17048 2838 17060
rect 3145 17051 3203 17057
rect 3145 17048 3157 17051
rect 2832 17020 3157 17048
rect 2832 17008 2838 17020
rect 3145 17017 3157 17020
rect 3191 17017 3203 17051
rect 3145 17011 3203 17017
rect 3234 17008 3240 17060
rect 3292 17008 3298 17060
rect 2409 16983 2467 16989
rect 2409 16949 2421 16983
rect 2455 16980 2467 16983
rect 4080 16980 4108 17088
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7340 17088 7573 17116
rect 7340 17076 7346 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 8205 17119 8263 17125
rect 8205 17116 8217 17119
rect 7892 17088 8217 17116
rect 7892 17076 7898 17088
rect 8205 17085 8217 17088
rect 8251 17085 8263 17119
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 8205 17079 8263 17085
rect 8312 17088 8493 17116
rect 4617 17051 4675 17057
rect 4617 17017 4629 17051
rect 4663 17048 4675 17051
rect 5074 17048 5080 17060
rect 4663 17020 5080 17048
rect 4663 17017 4675 17020
rect 4617 17011 4675 17017
rect 5074 17008 5080 17020
rect 5132 17008 5138 17060
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 8312 17048 8340 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 8570 17076 8576 17128
rect 8628 17125 8634 17128
rect 8628 17119 8656 17125
rect 8644 17085 8656 17119
rect 8628 17079 8656 17085
rect 8628 17076 8634 17079
rect 8168 17020 8340 17048
rect 8168 17008 8174 17020
rect 2455 16952 4108 16980
rect 2455 16949 2467 16952
rect 2409 16943 2467 16949
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 8570 16980 8576 16992
rect 7892 16952 8576 16980
rect 7892 16940 7898 16952
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 1104 16890 10120 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 7950 16890
rect 8002 16838 8014 16890
rect 8066 16838 8078 16890
rect 8130 16838 8142 16890
rect 8194 16838 8206 16890
rect 8258 16838 10120 16890
rect 1104 16816 10120 16838
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 2406 16776 2412 16788
rect 2188 16748 2412 16776
rect 2188 16736 2194 16748
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 2774 16736 2780 16788
rect 2832 16736 2838 16788
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 5132 16748 8217 16776
rect 5132 16736 5138 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 9539 16779 9597 16785
rect 9539 16745 9551 16779
rect 9585 16776 9597 16779
rect 10594 16776 10600 16788
rect 9585 16748 10600 16776
rect 9585 16745 9597 16748
rect 9539 16739 9597 16745
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 5718 16668 5724 16720
rect 5776 16708 5782 16720
rect 6730 16708 6736 16720
rect 5776 16680 6736 16708
rect 5776 16668 5782 16680
rect 6730 16668 6736 16680
rect 6788 16668 6794 16720
rect 7558 16668 7564 16720
rect 7616 16708 7622 16720
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 7616 16680 8493 16708
rect 7616 16668 7622 16680
rect 8481 16677 8493 16680
rect 8527 16677 8539 16711
rect 8481 16671 8539 16677
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 11054 16708 11060 16720
rect 8628 16680 11060 16708
rect 8628 16668 8634 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 1394 16600 1400 16652
rect 1452 16640 1458 16652
rect 1765 16643 1823 16649
rect 1765 16640 1777 16643
rect 1452 16612 1777 16640
rect 1452 16600 1458 16612
rect 1765 16609 1777 16612
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 6178 16640 6184 16652
rect 5592 16612 6184 16640
rect 5592 16600 5598 16612
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 9416 16612 9628 16640
rect 290 16532 296 16584
rect 348 16572 354 16584
rect 1118 16572 1124 16584
rect 348 16544 1124 16572
rect 348 16532 354 16544
rect 1118 16532 1124 16544
rect 1176 16532 1182 16584
rect 1578 16532 1584 16584
rect 1636 16572 1642 16584
rect 2038 16572 2044 16584
rect 1636 16544 2044 16572
rect 1636 16532 1642 16544
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16572 5319 16575
rect 5307 16544 6316 16572
rect 5307 16541 5319 16544
rect 5261 16535 5319 16541
rect 6288 16504 6316 16544
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 6733 16575 6791 16581
rect 6733 16572 6745 16575
rect 6420 16544 6745 16572
rect 6420 16532 6426 16544
rect 6733 16541 6745 16544
rect 6779 16541 6791 16575
rect 6733 16535 6791 16541
rect 7006 16532 7012 16584
rect 7064 16532 7070 16584
rect 8297 16575 8355 16581
rect 8297 16541 8309 16575
rect 8343 16572 8355 16575
rect 9416 16572 9444 16612
rect 8343 16544 9444 16572
rect 9600 16572 9628 16612
rect 9766 16600 9772 16652
rect 9824 16600 9830 16652
rect 9858 16572 9864 16584
rect 9600 16544 9864 16572
rect 8343 16541 8355 16544
rect 8297 16535 8355 16541
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 8665 16507 8723 16513
rect 6288 16476 8248 16504
rect 290 16396 296 16448
rect 348 16436 354 16448
rect 4154 16436 4160 16448
rect 348 16408 4160 16436
rect 348 16396 354 16408
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 4982 16436 4988 16448
rect 4571 16408 4988 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 4982 16396 4988 16408
rect 5040 16396 5046 16448
rect 6086 16396 6092 16448
rect 6144 16436 6150 16448
rect 6288 16436 6316 16476
rect 6144 16408 6316 16436
rect 7745 16439 7803 16445
rect 6144 16396 6150 16408
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 8110 16436 8116 16448
rect 7791 16408 8116 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 8220 16436 8248 16476
rect 8665 16473 8677 16507
rect 8711 16504 8723 16507
rect 9766 16504 9772 16516
rect 8711 16476 9772 16504
rect 8711 16473 8723 16476
rect 8665 16467 8723 16473
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 9306 16436 9312 16448
rect 8220 16408 9312 16436
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 1104 16346 10120 16368
rect 1104 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 3202 16346
rect 3254 16294 3266 16346
rect 3318 16294 9010 16346
rect 9062 16294 9074 16346
rect 9126 16294 9138 16346
rect 9190 16294 9202 16346
rect 9254 16294 9266 16346
rect 9318 16294 10120 16346
rect 1104 16272 10120 16294
rect 2498 16192 2504 16244
rect 2556 16232 2562 16244
rect 2556 16204 4384 16232
rect 2556 16192 2562 16204
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 1670 16056 1676 16108
rect 1728 16056 1734 16108
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2498 16096 2504 16108
rect 2455 16068 2504 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 3602 16056 3608 16108
rect 3660 16056 3666 16108
rect 2593 16031 2651 16037
rect 2593 15997 2605 16031
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 1670 15920 1676 15972
rect 1728 15960 1734 15972
rect 2130 15960 2136 15972
rect 1728 15932 2136 15960
rect 1728 15920 1734 15932
rect 2130 15920 2136 15932
rect 2188 15920 2194 15972
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2314 15892 2320 15904
rect 2096 15864 2320 15892
rect 2096 15852 2102 15864
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 2608 15892 2636 15991
rect 3326 15988 3332 16040
rect 3384 15988 3390 16040
rect 3467 16031 3525 16037
rect 3467 15997 3479 16031
rect 3513 16028 3525 16031
rect 4246 16028 4252 16040
rect 3513 16000 4252 16028
rect 3513 15997 3525 16000
rect 3467 15991 3525 15997
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 4356 16037 4384 16204
rect 5994 16192 6000 16244
rect 6052 16192 6058 16244
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 9585 16235 9643 16241
rect 9585 16232 9597 16235
rect 8444 16204 9597 16232
rect 8444 16192 8450 16204
rect 9585 16201 9597 16204
rect 9631 16201 9643 16235
rect 9585 16195 9643 16201
rect 6012 16164 6040 16192
rect 6012 16136 6684 16164
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 16028 4399 16031
rect 4430 16028 4436 16040
rect 4387 16000 4436 16028
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4890 16028 4896 16040
rect 4571 16000 4896 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 4982 15988 4988 16040
rect 5040 15988 5046 16040
rect 5276 16028 5304 16059
rect 5534 16056 5540 16108
rect 5592 16056 5598 16108
rect 6656 16105 6684 16136
rect 9674 16124 9680 16176
rect 9732 16124 9738 16176
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 7558 16056 7564 16108
rect 7616 16056 7622 16108
rect 8662 16105 8668 16108
rect 8619 16099 8668 16105
rect 8619 16065 8631 16099
rect 8665 16065 8668 16099
rect 8619 16059 8668 16065
rect 8662 16056 8668 16059
rect 8720 16056 8726 16108
rect 5092 16000 5304 16028
rect 5399 16031 5457 16037
rect 3050 15920 3056 15972
rect 3108 15920 3114 15972
rect 4154 15892 4160 15904
rect 2608 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 4338 15892 4344 15904
rect 4295 15864 4344 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5092 15892 5120 16000
rect 5399 15997 5411 16031
rect 5445 16028 5457 16031
rect 5718 16028 5724 16040
rect 5445 16000 5724 16028
rect 5445 15997 5457 16000
rect 5399 15991 5457 15997
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 6362 15988 6368 16040
rect 6420 15988 6426 16040
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7374 16028 7380 16040
rect 7248 16000 7380 16028
rect 7248 15988 7254 16000
rect 7374 15988 7380 16000
rect 7432 16028 7438 16040
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 7432 16000 7757 16028
rect 7432 15988 7438 16000
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 8110 15988 8116 16040
rect 8168 16028 8174 16040
rect 8205 16031 8263 16037
rect 8205 16028 8217 16031
rect 8168 16000 8217 16028
rect 8168 15988 8174 16000
rect 8205 15997 8217 16000
rect 8251 15997 8263 16031
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 8205 15991 8263 15997
rect 8312 16000 8493 16028
rect 8018 15920 8024 15972
rect 8076 15960 8082 15972
rect 8312 15960 8340 16000
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 16028 8815 16031
rect 8803 16000 9168 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 8076 15932 8340 15960
rect 8076 15920 8082 15932
rect 5534 15892 5540 15904
rect 5040 15864 5540 15892
rect 5040 15852 5046 15864
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6178 15852 6184 15904
rect 6236 15852 6242 15904
rect 7377 15895 7435 15901
rect 7377 15861 7389 15895
rect 7423 15892 7435 15895
rect 9140 15892 9168 16000
rect 7423 15864 9168 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 9398 15852 9404 15904
rect 9456 15852 9462 15904
rect 1104 15802 10120 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 7950 15802
rect 8002 15750 8014 15802
rect 8066 15750 8078 15802
rect 8130 15750 8142 15802
rect 8194 15750 8206 15802
rect 8258 15750 10120 15802
rect 1104 15728 10120 15750
rect 3050 15648 3056 15700
rect 3108 15648 3114 15700
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 4525 15691 4583 15697
rect 4525 15688 4537 15691
rect 4120 15660 4537 15688
rect 4120 15648 4126 15660
rect 4525 15657 4537 15660
rect 4571 15657 4583 15691
rect 5442 15688 5448 15700
rect 4525 15651 4583 15657
rect 4632 15660 5448 15688
rect 1670 15512 1676 15564
rect 1728 15552 1734 15564
rect 1946 15552 1952 15564
rect 1728 15524 1952 15552
rect 1728 15512 1734 15524
rect 1946 15512 1952 15524
rect 2004 15552 2010 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 2004 15524 2053 15552
rect 2004 15512 2010 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 2682 15512 2688 15564
rect 2740 15552 2746 15564
rect 2740 15512 2774 15552
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4632 15561 4660 15660
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5997 15691 6055 15697
rect 5997 15657 6009 15691
rect 6043 15688 6055 15691
rect 6730 15688 6736 15700
rect 6043 15660 6736 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7374 15648 7380 15700
rect 7432 15648 7438 15700
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7708 15660 7849 15688
rect 7708 15648 7714 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 11146 15688 11152 15700
rect 7837 15651 7895 15657
rect 7944 15660 11152 15688
rect 5629 15623 5687 15629
rect 5629 15589 5641 15623
rect 5675 15589 5687 15623
rect 5629 15583 5687 15589
rect 4617 15555 4675 15561
rect 4617 15552 4629 15555
rect 4304 15524 4629 15552
rect 4304 15512 4310 15524
rect 4617 15521 4629 15524
rect 4663 15521 4675 15555
rect 5644 15552 5672 15583
rect 5718 15580 5724 15632
rect 5776 15620 5782 15632
rect 7944 15620 7972 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 8846 15620 8852 15632
rect 5776 15592 7972 15620
rect 8036 15592 8852 15620
rect 5776 15580 5782 15592
rect 5994 15552 6000 15564
rect 5644 15524 6000 15552
rect 4617 15515 4675 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 8036 15552 8064 15592
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 9950 15620 9956 15632
rect 9692 15592 9956 15620
rect 6512 15524 8064 15552
rect 8481 15555 8539 15561
rect 6512 15512 6518 15524
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 9692 15552 9720 15592
rect 9950 15580 9956 15592
rect 10008 15580 10014 15632
rect 8527 15524 9720 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 9766 15512 9772 15564
rect 9824 15512 9830 15564
rect 2314 15444 2320 15496
rect 2372 15444 2378 15496
rect 2746 15416 2774 15512
rect 4338 15444 4344 15496
rect 4396 15444 4402 15496
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15484 4951 15487
rect 4982 15484 4988 15496
rect 4939 15456 4988 15484
rect 4939 15453 4951 15456
rect 4893 15447 4951 15453
rect 4908 15416 4936 15447
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 6178 15484 6184 15496
rect 5859 15456 6184 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 2746 15388 4936 15416
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 7576 15416 7604 15447
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 8754 15444 8760 15496
rect 8812 15444 8818 15496
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 8846 15416 8852 15428
rect 5592 15388 7420 15416
rect 7576 15388 8852 15416
rect 5592 15376 5598 15388
rect 4430 15308 4436 15360
rect 4488 15348 4494 15360
rect 7282 15348 7288 15360
rect 4488 15320 7288 15348
rect 4488 15308 4494 15320
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 7392 15348 7420 15388
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 9508 15348 9536 15447
rect 7392 15320 9536 15348
rect 1104 15258 10120 15280
rect 1104 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 3202 15258
rect 3254 15206 3266 15258
rect 3318 15206 9010 15258
rect 9062 15206 9074 15258
rect 9126 15206 9138 15258
rect 9190 15206 9202 15258
rect 9254 15206 9266 15258
rect 9318 15206 10120 15258
rect 1104 15184 10120 15206
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3602 15144 3608 15156
rect 3007 15116 3608 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 3786 15104 3792 15156
rect 3844 15144 3850 15156
rect 4430 15144 4436 15156
rect 3844 15116 4436 15144
rect 3844 15104 3850 15116
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 7650 15144 7656 15156
rect 7607 15116 7656 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 7800 15116 9260 15144
rect 7800 15104 7806 15116
rect 1486 15036 1492 15088
rect 1544 15076 1550 15088
rect 1544 15048 2268 15076
rect 1544 15036 1550 15048
rect 1026 14968 1032 15020
rect 1084 15008 1090 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1084 14980 1685 15008
rect 1084 14968 1090 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 1946 14968 1952 15020
rect 2004 14968 2010 15020
rect 2240 15017 2268 15048
rect 7006 15036 7012 15088
rect 7064 15076 7070 15088
rect 7760 15076 7788 15104
rect 7064 15048 7788 15076
rect 7064 15036 7070 15048
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 15008 2283 15011
rect 2682 15008 2688 15020
rect 2271 14980 2688 15008
rect 2271 14977 2283 14980
rect 2225 14971 2283 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 5166 14968 5172 15020
rect 5224 15008 5230 15020
rect 6730 15008 6736 15020
rect 5224 14980 6736 15008
rect 5224 14968 5230 14980
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 8386 15017 8392 15020
rect 8364 15011 8392 15017
rect 8364 14977 8376 15011
rect 8364 14971 8392 14977
rect 8386 14968 8392 14971
rect 8444 14968 8450 15020
rect 9232 15008 9260 15116
rect 9674 15036 9680 15088
rect 9732 15036 9738 15088
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 9232 14980 9413 15008
rect 9401 14977 9413 14980
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 6457 14943 6515 14949
rect 6457 14940 6469 14943
rect 6420 14912 6469 14940
rect 6420 14900 6426 14912
rect 6457 14909 6469 14912
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 8205 14943 8263 14949
rect 8205 14940 8217 14943
rect 7616 14912 8217 14940
rect 7616 14900 7622 14912
rect 8205 14909 8217 14912
rect 8251 14909 8263 14943
rect 8205 14903 8263 14909
rect 8481 14943 8539 14949
rect 8481 14909 8493 14943
rect 8527 14940 8539 14943
rect 8662 14940 8668 14952
rect 8527 14912 8668 14940
rect 8527 14909 8539 14912
rect 8481 14903 8539 14909
rect 8662 14900 8668 14912
rect 8720 14900 8726 14952
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 8757 14875 8815 14881
rect 8757 14841 8769 14875
rect 8803 14841 8815 14875
rect 8757 14835 8815 14841
rect 1486 14764 1492 14816
rect 1544 14764 1550 14816
rect 2406 14764 2412 14816
rect 2464 14804 2470 14816
rect 2590 14804 2596 14816
rect 2464 14776 2596 14804
rect 2464 14764 2470 14776
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 8772 14804 8800 14835
rect 9490 14832 9496 14884
rect 9548 14832 9554 14884
rect 7515 14776 8800 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 1104 14714 10120 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 7950 14714
rect 8002 14662 8014 14714
rect 8066 14662 8078 14714
rect 8130 14662 8142 14714
rect 8194 14662 8206 14714
rect 8258 14662 10120 14714
rect 1104 14640 10120 14662
rect 4246 14600 4252 14612
rect 1872 14572 4252 14600
rect 1762 14424 1768 14476
rect 1820 14464 1826 14476
rect 1872 14473 1900 14572
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 6454 14600 6460 14612
rect 4479 14572 6460 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 9306 14560 9312 14612
rect 9364 14560 9370 14612
rect 9585 14603 9643 14609
rect 9585 14569 9597 14603
rect 9631 14600 9643 14603
rect 9950 14600 9956 14612
rect 9631 14572 9956 14600
rect 9631 14569 9643 14572
rect 9585 14563 9643 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 4338 14492 4344 14544
rect 4396 14532 4402 14544
rect 4522 14532 4528 14544
rect 4396 14504 4528 14532
rect 4396 14492 4402 14504
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 6914 14492 6920 14544
rect 6972 14532 6978 14544
rect 7541 14535 7599 14541
rect 7541 14532 7553 14535
rect 6972 14504 7553 14532
rect 6972 14492 6978 14504
rect 7541 14501 7553 14504
rect 7587 14501 7599 14535
rect 10042 14532 10048 14544
rect 7541 14495 7599 14501
rect 9646 14504 10048 14532
rect 1857 14467 1915 14473
rect 1857 14464 1869 14467
rect 1820 14436 1869 14464
rect 1820 14424 1826 14436
rect 1857 14433 1869 14436
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14464 7159 14467
rect 7190 14464 7196 14476
rect 7147 14436 7196 14464
rect 7147 14433 7159 14436
rect 7101 14427 7159 14433
rect 7190 14424 7196 14436
rect 7248 14464 7254 14476
rect 7650 14464 7656 14476
rect 7248 14436 7656 14464
rect 7248 14424 7254 14436
rect 7650 14424 7656 14436
rect 7708 14464 7714 14476
rect 9214 14464 9220 14476
rect 7708 14436 9220 14464
rect 7708 14424 7714 14436
rect 9214 14424 9220 14436
rect 9272 14464 9278 14476
rect 9646 14464 9674 14504
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 9272 14436 9674 14464
rect 9272 14424 9278 14436
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 2133 14399 2191 14405
rect 2133 14396 2145 14399
rect 1673 14359 1731 14365
rect 1872 14368 2145 14396
rect 1486 14220 1492 14272
rect 1544 14220 1550 14272
rect 1688 14260 1716 14359
rect 1872 14340 1900 14368
rect 2133 14365 2145 14368
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4522 14396 4528 14408
rect 4295 14368 4528 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5810 14396 5816 14408
rect 4939 14368 5816 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 1854 14288 1860 14340
rect 1912 14288 1918 14340
rect 3878 14328 3884 14340
rect 2792 14300 3884 14328
rect 2792 14260 2820 14300
rect 3878 14288 3884 14300
rect 3936 14288 3942 14340
rect 4632 14328 4660 14359
rect 5810 14356 5816 14368
rect 5868 14356 5874 14408
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 6546 14396 6552 14408
rect 6503 14368 6552 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 5074 14328 5080 14340
rect 4632 14300 5080 14328
rect 5074 14288 5080 14300
rect 5132 14328 5138 14340
rect 6748 14328 6776 14359
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 6880 14368 6929 14396
rect 6880 14356 6886 14368
rect 6917 14365 6929 14368
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7834 14356 7840 14408
rect 7892 14356 7898 14408
rect 8018 14405 8024 14408
rect 7975 14399 8024 14405
rect 7975 14365 7987 14399
rect 8021 14365 8024 14399
rect 7975 14359 8024 14365
rect 8018 14356 8024 14359
rect 8076 14356 8082 14408
rect 8110 14356 8116 14408
rect 8168 14356 8174 14408
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9398 14396 9404 14408
rect 9171 14368 9404 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 10502 14396 10508 14408
rect 9723 14368 10508 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 5132 14300 6776 14328
rect 5132 14288 5138 14300
rect 1688 14232 2820 14260
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14260 2927 14263
rect 3510 14260 3516 14272
rect 2915 14232 3516 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5629 14263 5687 14269
rect 5629 14260 5641 14263
rect 5592 14232 5641 14260
rect 5592 14220 5598 14232
rect 5629 14229 5641 14232
rect 5675 14229 5687 14263
rect 5629 14223 5687 14229
rect 5721 14263 5779 14269
rect 5721 14229 5733 14263
rect 5767 14260 5779 14263
rect 5810 14260 5816 14272
rect 5767 14232 5816 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 8754 14220 8760 14272
rect 8812 14220 8818 14272
rect 1104 14170 10120 14192
rect 1104 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 3202 14170
rect 3254 14118 3266 14170
rect 3318 14118 9010 14170
rect 9062 14118 9074 14170
rect 9126 14118 9138 14170
rect 9190 14118 9202 14170
rect 9254 14118 9266 14170
rect 9318 14118 10120 14170
rect 1104 14096 10120 14118
rect 2777 14059 2835 14065
rect 2777 14025 2789 14059
rect 2823 14056 2835 14059
rect 4062 14056 4068 14068
rect 2823 14028 4068 14056
rect 2823 14025 2835 14028
rect 2777 14019 2835 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4580 14028 4721 14056
rect 4580 14016 4586 14028
rect 4709 14025 4721 14028
rect 4755 14025 4767 14059
rect 4709 14019 4767 14025
rect 7190 14016 7196 14068
rect 7248 14056 7254 14068
rect 8018 14056 8024 14068
rect 7248 14028 8024 14056
rect 7248 14016 7254 14028
rect 8018 14016 8024 14028
rect 8076 14056 8082 14068
rect 8202 14056 8208 14068
rect 8076 14028 8208 14056
rect 8076 14016 8082 14028
rect 8202 14016 8208 14028
rect 8260 14056 8266 14068
rect 8386 14056 8392 14068
rect 8260 14028 8392 14056
rect 8260 14016 8266 14028
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9585 14059 9643 14065
rect 9585 14056 9597 14059
rect 8720 14028 9597 14056
rect 8720 14016 8726 14028
rect 9585 14025 9597 14028
rect 9631 14025 9643 14059
rect 9585 14019 9643 14025
rect 1670 13948 1676 14000
rect 1728 13988 1734 14000
rect 1728 13960 2084 13988
rect 1728 13948 1734 13960
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 2056 13929 2084 13960
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2590 13920 2596 13932
rect 2087 13892 2596 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3786 13880 3792 13932
rect 3844 13880 3850 13932
rect 4062 13880 4068 13932
rect 4120 13880 4126 13932
rect 5074 13880 5080 13932
rect 5132 13880 5138 13932
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 7650 13880 7656 13932
rect 7708 13880 7714 13932
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 9766 13880 9772 13932
rect 9824 13880 9830 13932
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 2884 13784 2912 13815
rect 3050 13812 3056 13864
rect 3108 13812 3114 13864
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 3927 13855 3985 13861
rect 3927 13821 3939 13855
rect 3973 13852 3985 13855
rect 4246 13852 4252 13864
rect 3973 13824 4252 13852
rect 3973 13821 3985 13824
rect 3927 13815 3985 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 7098 13852 7104 13864
rect 6788 13824 7104 13852
rect 6788 13812 6794 13824
rect 7098 13812 7104 13824
rect 7156 13852 7162 13864
rect 7469 13855 7527 13861
rect 7469 13852 7481 13855
rect 7156 13824 7481 13852
rect 7156 13812 7162 13824
rect 7469 13821 7481 13824
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8506 13855 8564 13861
rect 8506 13852 8518 13855
rect 8260 13824 8518 13852
rect 8260 13812 8266 13824
rect 8506 13821 8518 13824
rect 8552 13821 8564 13855
rect 8506 13815 8564 13821
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 8846 13852 8852 13864
rect 8711 13824 8852 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 2884 13756 3556 13784
rect 3528 13728 3556 13756
rect 7834 13744 7840 13796
rect 7892 13784 7898 13796
rect 8113 13787 8171 13793
rect 8113 13784 8125 13787
rect 7892 13756 8125 13784
rect 7892 13744 7898 13756
rect 8113 13753 8125 13756
rect 8159 13753 8171 13787
rect 8113 13747 8171 13753
rect 3510 13676 3516 13728
rect 3568 13676 3574 13728
rect 6089 13719 6147 13725
rect 6089 13685 6101 13719
rect 6135 13716 6147 13719
rect 6730 13716 6736 13728
rect 6135 13688 6736 13716
rect 6135 13685 6147 13688
rect 6089 13679 6147 13685
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 8386 13716 8392 13728
rect 7708 13688 8392 13716
rect 7708 13676 7714 13688
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 9306 13676 9312 13728
rect 9364 13676 9370 13728
rect 1104 13626 10120 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 7950 13626
rect 8002 13574 8014 13626
rect 8066 13574 8078 13626
rect 8130 13574 8142 13626
rect 8194 13574 8206 13626
rect 8258 13574 10120 13626
rect 1104 13552 10120 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 7650 13512 7656 13524
rect 3108 13484 7656 13512
rect 3108 13472 3114 13484
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 7742 13472 7748 13524
rect 7800 13472 7806 13524
rect 9674 13512 9680 13524
rect 8404 13484 9680 13512
rect 1026 13404 1032 13456
rect 1084 13444 1090 13456
rect 6822 13453 6828 13456
rect 1949 13447 2007 13453
rect 1949 13444 1961 13447
rect 1084 13416 1961 13444
rect 1084 13404 1090 13416
rect 1949 13413 1961 13416
rect 1995 13413 2007 13447
rect 1949 13407 2007 13413
rect 6779 13447 6828 13453
rect 6779 13413 6791 13447
rect 6825 13413 6828 13447
rect 6779 13407 6828 13413
rect 6822 13404 6828 13407
rect 6880 13404 6886 13456
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 7926 13444 7932 13456
rect 7340 13416 7932 13444
rect 7340 13404 7346 13416
rect 7926 13404 7932 13416
rect 7984 13404 7990 13456
rect 8021 13447 8079 13453
rect 8021 13413 8033 13447
rect 8067 13444 8079 13447
rect 8202 13444 8208 13456
rect 8067 13416 8208 13444
rect 8067 13413 8079 13416
rect 8021 13407 8079 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13413 8355 13447
rect 8297 13407 8355 13413
rect 198 13336 204 13388
rect 256 13376 262 13388
rect 4982 13376 4988 13388
rect 256 13348 4988 13376
rect 256 13336 262 13348
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5994 13336 6000 13388
rect 6052 13376 6058 13388
rect 8312 13376 8340 13407
rect 6052 13348 8340 13376
rect 6052 13336 6058 13348
rect 1578 13268 1584 13320
rect 1636 13308 1642 13320
rect 1673 13311 1731 13317
rect 1673 13308 1685 13311
rect 1636 13280 1685 13308
rect 1636 13268 1642 13280
rect 1673 13277 1685 13280
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 1762 13268 1768 13320
rect 1820 13268 1826 13320
rect 6730 13317 6736 13320
rect 6708 13311 6736 13317
rect 6708 13277 6720 13311
rect 6708 13271 6736 13277
rect 6730 13268 6736 13271
rect 6788 13268 6794 13320
rect 7929 13311 7987 13317
rect 7929 13277 7941 13311
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8404 13308 8432 13484
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9214 13404 9220 13456
rect 9272 13444 9278 13456
rect 9950 13444 9956 13456
rect 9272 13416 9956 13444
rect 9272 13404 9278 13416
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 9490 13336 9496 13388
rect 9548 13336 9554 13388
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 10502 13376 10508 13388
rect 9640 13348 10508 13376
rect 9640 13336 9646 13348
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 8251 13280 8432 13308
rect 8481 13311 8539 13317
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 9214 13308 9220 13320
rect 8803 13280 9220 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 566 13200 572 13252
rect 624 13240 630 13252
rect 3602 13240 3608 13252
rect 624 13212 3608 13240
rect 624 13200 630 13212
rect 3602 13200 3608 13212
rect 3660 13200 3666 13252
rect 3878 13200 3884 13252
rect 3936 13240 3942 13252
rect 4338 13240 4344 13252
rect 3936 13212 4344 13240
rect 3936 13200 3942 13212
rect 4338 13200 4344 13212
rect 4396 13200 4402 13252
rect 5902 13200 5908 13252
rect 5960 13240 5966 13252
rect 7650 13240 7656 13252
rect 5960 13212 7656 13240
rect 5960 13200 5966 13212
rect 7650 13200 7656 13212
rect 7708 13200 7714 13252
rect 7944 13240 7972 13271
rect 8386 13240 8392 13252
rect 7944 13212 8392 13240
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 8496 13240 8524 13271
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 9306 13268 9312 13320
rect 9364 13268 9370 13320
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9766 13308 9772 13320
rect 9456 13280 9772 13308
rect 9456 13268 9462 13280
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 10962 13240 10968 13252
rect 8496 13212 10968 13240
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 1486 13132 1492 13184
rect 1544 13132 1550 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 8573 13175 8631 13181
rect 8573 13172 8585 13175
rect 4304 13144 8585 13172
rect 4304 13132 4310 13144
rect 8573 13141 8585 13144
rect 8619 13141 8631 13175
rect 8573 13135 8631 13141
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 8720 13144 8953 13172
rect 8720 13132 8726 13144
rect 8941 13141 8953 13144
rect 8987 13141 8999 13175
rect 8941 13135 8999 13141
rect 9398 13132 9404 13184
rect 9456 13132 9462 13184
rect 1104 13082 10120 13104
rect 1104 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 3202 13082
rect 3254 13030 3266 13082
rect 3318 13030 9010 13082
rect 9062 13030 9074 13082
rect 9126 13030 9138 13082
rect 9190 13030 9202 13082
rect 9254 13030 9266 13082
rect 9318 13030 10120 13082
rect 1104 13008 10120 13030
rect 3510 12968 3516 12980
rect 2976 12940 3516 12968
rect 1486 12860 1492 12912
rect 1544 12900 1550 12912
rect 1670 12900 1676 12912
rect 1544 12872 1676 12900
rect 1544 12860 1550 12872
rect 1670 12860 1676 12872
rect 1728 12860 1734 12912
rect 2498 12900 2504 12912
rect 1780 12872 2504 12900
rect 1780 12832 1808 12872
rect 2498 12860 2504 12872
rect 2556 12860 2562 12912
rect 1688 12804 1808 12832
rect 1688 12776 1716 12804
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1912 12804 1961 12832
rect 1912 12792 1918 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 2976 12832 3004 12940
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 4706 12968 4712 12980
rect 3844 12940 4712 12968
rect 3844 12928 3850 12940
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 4893 12971 4951 12977
rect 4893 12937 4905 12971
rect 4939 12968 4951 12971
rect 5718 12968 5724 12980
rect 4939 12940 5724 12968
rect 4939 12937 4951 12940
rect 4893 12931 4951 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 9217 12971 9275 12977
rect 6788 12940 9076 12968
rect 6788 12928 6794 12940
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 7116 12909 7144 12940
rect 6917 12903 6975 12909
rect 6917 12900 6929 12903
rect 6328 12872 6929 12900
rect 6328 12860 6334 12872
rect 6917 12869 6929 12872
rect 6963 12869 6975 12903
rect 6917 12863 6975 12869
rect 7101 12903 7159 12909
rect 7101 12869 7113 12903
rect 7147 12869 7159 12903
rect 9048 12900 9076 12940
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9398 12968 9404 12980
rect 9263 12940 9404 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10318 12900 10324 12912
rect 9048 12872 9444 12900
rect 7101 12863 7159 12869
rect 9416 12844 9444 12872
rect 9508 12872 10324 12900
rect 3697 12835 3755 12841
rect 2823 12804 3096 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 3068 12776 3096 12804
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4709 12835 4767 12841
rect 4709 12832 4721 12835
rect 4663 12804 4721 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4709 12801 4721 12804
rect 4755 12801 4767 12835
rect 4709 12795 4767 12801
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 2958 12724 2964 12776
rect 3016 12724 3022 12776
rect 3050 12724 3056 12776
rect 3108 12724 3114 12776
rect 3712 12764 3740 12795
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 4856 12804 5764 12832
rect 4856 12792 4862 12804
rect 3878 12773 3884 12776
rect 3553 12736 3740 12764
rect 3835 12767 3884 12773
rect 2685 12699 2743 12705
rect 2685 12665 2697 12699
rect 2731 12696 2743 12699
rect 3421 12699 3479 12705
rect 3421 12696 3433 12699
rect 2731 12668 3433 12696
rect 2731 12665 2743 12668
rect 2685 12659 2743 12665
rect 3421 12665 3433 12668
rect 3467 12665 3479 12699
rect 3421 12659 3479 12665
rect 3553 12628 3581 12736
rect 3835 12733 3847 12767
rect 3881 12733 3884 12767
rect 3835 12727 3884 12733
rect 3878 12724 3884 12727
rect 3936 12724 3942 12776
rect 3973 12767 4031 12773
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 4019 12736 4752 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 4724 12708 4752 12736
rect 5626 12724 5632 12776
rect 5684 12724 5690 12776
rect 5736 12764 5764 12804
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6512 12804 6561 12832
rect 6512 12792 6518 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6822 12792 6828 12844
rect 6880 12792 6886 12844
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7432 12804 7788 12832
rect 7432 12792 7438 12804
rect 5736 12736 6960 12764
rect 4706 12656 4712 12708
rect 4764 12656 4770 12708
rect 5166 12628 5172 12640
rect 3553 12600 5172 12628
rect 5166 12588 5172 12600
rect 5224 12628 5230 12640
rect 5644 12628 5672 12724
rect 6365 12699 6423 12705
rect 6365 12665 6377 12699
rect 6411 12696 6423 12699
rect 6822 12696 6828 12708
rect 6411 12668 6828 12696
rect 6411 12665 6423 12668
rect 6365 12659 6423 12665
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 5224 12600 5672 12628
rect 5224 12588 5230 12600
rect 6730 12588 6736 12640
rect 6788 12588 6794 12640
rect 6932 12628 6960 12736
rect 7006 12724 7012 12776
rect 7064 12764 7070 12776
rect 7561 12767 7619 12773
rect 7561 12764 7573 12767
rect 7064 12736 7573 12764
rect 7064 12724 7070 12736
rect 7561 12733 7573 12736
rect 7607 12733 7619 12767
rect 7760 12764 7788 12804
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 9508 12841 9536 12872
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 10686 12832 10692 12844
rect 9815 12804 10692 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 7926 12764 7932 12776
rect 7760 12736 7932 12764
rect 7561 12727 7619 12733
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 8414 12767 8472 12773
rect 8414 12764 8426 12767
rect 8168 12736 8426 12764
rect 8168 12724 8174 12736
rect 8414 12733 8426 12736
rect 8460 12733 8472 12767
rect 8414 12727 8472 12733
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 8938 12764 8944 12776
rect 8619 12736 8944 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 7374 12656 7380 12708
rect 7432 12696 7438 12708
rect 8021 12699 8079 12705
rect 8021 12696 8033 12699
rect 7432 12668 8033 12696
rect 7432 12656 7438 12668
rect 8021 12665 8033 12668
rect 8067 12665 8079 12699
rect 8021 12659 8079 12665
rect 9309 12699 9367 12705
rect 9309 12665 9321 12699
rect 9355 12696 9367 12699
rect 10594 12696 10600 12708
rect 9355 12668 10600 12696
rect 9355 12665 9367 12668
rect 9309 12659 9367 12665
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 9585 12631 9643 12637
rect 9585 12628 9597 12631
rect 6932 12600 9597 12628
rect 9585 12597 9597 12600
rect 9631 12597 9643 12631
rect 9585 12591 9643 12597
rect 10042 12588 10048 12640
rect 10100 12628 10106 12640
rect 10778 12628 10784 12640
rect 10100 12600 10784 12628
rect 10100 12588 10106 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 1104 12538 10120 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 7950 12538
rect 8002 12486 8014 12538
rect 8066 12486 8078 12538
rect 8130 12486 8142 12538
rect 8194 12486 8206 12538
rect 8258 12486 10120 12538
rect 1104 12464 10120 12486
rect 382 12384 388 12436
rect 440 12424 446 12436
rect 1302 12424 1308 12436
rect 440 12396 1308 12424
rect 440 12384 446 12396
rect 1302 12384 1308 12396
rect 1360 12424 1366 12436
rect 1397 12427 1455 12433
rect 1397 12424 1409 12427
rect 1360 12396 1409 12424
rect 1360 12384 1366 12396
rect 1397 12393 1409 12396
rect 1443 12393 1455 12427
rect 1397 12387 1455 12393
rect 2685 12427 2743 12433
rect 2685 12393 2697 12427
rect 2731 12424 2743 12427
rect 4706 12424 4712 12436
rect 2731 12396 4712 12424
rect 2731 12393 2743 12396
rect 2685 12387 2743 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 6178 12424 6184 12436
rect 5592 12396 6184 12424
rect 5592 12384 5598 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 6788 12396 6837 12424
rect 6788 12384 6794 12396
rect 6825 12393 6837 12396
rect 6871 12393 6883 12427
rect 6825 12387 6883 12393
rect 7116 12396 7604 12424
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2777 12359 2835 12365
rect 2777 12356 2789 12359
rect 2556 12328 2789 12356
rect 2556 12316 2562 12328
rect 2777 12325 2789 12328
rect 2823 12325 2835 12359
rect 2777 12319 2835 12325
rect 5258 12316 5264 12368
rect 5316 12356 5322 12368
rect 5316 12328 5764 12356
rect 5316 12316 5322 12328
rect 5736 12300 5764 12328
rect 6638 12316 6644 12368
rect 6696 12316 6702 12368
rect 1670 12248 1676 12300
rect 1728 12248 1734 12300
rect 2866 12288 2872 12300
rect 2700 12260 2872 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12220 2007 12223
rect 2590 12220 2596 12232
rect 1995 12192 2596 12220
rect 1995 12189 2007 12192
rect 1949 12183 2007 12189
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 1964 12152 1992 12183
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 1728 12124 1992 12152
rect 1728 12112 1734 12124
rect 2222 12112 2228 12164
rect 2280 12152 2286 12164
rect 2700 12152 2728 12260
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 4985 12291 5043 12297
rect 4985 12288 4997 12291
rect 4764 12260 4997 12288
rect 4764 12248 4770 12260
rect 4985 12257 4997 12260
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5776 12260 5917 12288
rect 5776 12248 5782 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6656 12288 6684 12316
rect 7116 12288 7144 12396
rect 7576 12356 7604 12396
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7708 12396 8033 12424
rect 7708 12384 7714 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 8938 12424 8944 12436
rect 8021 12387 8079 12393
rect 8128 12396 8944 12424
rect 8128 12356 8156 12396
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 7576 12328 8156 12356
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 8297 12359 8355 12365
rect 8297 12356 8309 12359
rect 8260 12328 8309 12356
rect 8260 12316 8266 12328
rect 8297 12325 8309 12328
rect 8343 12325 8355 12359
rect 8297 12319 8355 12325
rect 8573 12359 8631 12365
rect 8573 12325 8585 12359
rect 8619 12356 8631 12359
rect 9122 12356 9128 12368
rect 8619 12328 9128 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 9122 12316 9128 12328
rect 9180 12316 9186 12368
rect 9858 12288 9864 12300
rect 6236 12260 7144 12288
rect 8496 12260 9864 12288
rect 6236 12248 6242 12260
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 3881 12223 3939 12229
rect 3881 12220 3893 12223
rect 3752 12192 3893 12220
rect 3752 12180 3758 12192
rect 3881 12189 3893 12192
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 2280 12124 2728 12152
rect 2280 12112 2286 12124
rect 2866 12112 2872 12164
rect 2924 12152 2930 12164
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2924 12124 2973 12152
rect 2924 12112 2930 12124
rect 2961 12121 2973 12124
rect 3007 12121 3019 12155
rect 3896 12152 3924 12183
rect 4154 12180 4160 12232
rect 4212 12180 4218 12232
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12220 5227 12223
rect 5350 12220 5356 12232
rect 5215 12192 5356 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5994 12180 6000 12232
rect 6052 12229 6058 12232
rect 6052 12223 6080 12229
rect 6068 12189 6080 12223
rect 6052 12183 6080 12189
rect 6052 12180 6058 12183
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 6880 12192 7113 12220
rect 6880 12180 6886 12192
rect 7101 12189 7113 12192
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 8496 12229 8524 12260
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 5074 12152 5080 12164
rect 3896 12124 5080 12152
rect 2961 12115 3019 12121
rect 5074 12112 5080 12124
rect 5132 12112 5138 12164
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6788 12124 7205 12152
rect 6788 12112 6794 12124
rect 7193 12121 7205 12124
rect 7239 12121 7251 12155
rect 7193 12115 7251 12121
rect 7285 12155 7343 12161
rect 7285 12121 7297 12155
rect 7331 12121 7343 12155
rect 8772 12152 8800 12183
rect 9490 12180 9496 12232
rect 9548 12180 9554 12232
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 8938 12152 8944 12164
rect 8772 12124 8944 12152
rect 7285 12115 7343 12121
rect 4893 12087 4951 12093
rect 4893 12053 4905 12087
rect 4939 12084 4951 12087
rect 6454 12084 6460 12096
rect 4939 12056 6460 12084
rect 4939 12053 4951 12056
rect 4893 12047 4951 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6880 12056 6929 12084
rect 6880 12044 6886 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 7300 12084 7328 12115
rect 8938 12112 8944 12124
rect 8996 12112 9002 12164
rect 9122 12112 9128 12164
rect 9180 12112 9186 12164
rect 9398 12112 9404 12164
rect 9456 12152 9462 12164
rect 9674 12152 9680 12164
rect 9456 12124 9680 12152
rect 9456 12112 9462 12124
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 8662 12084 8668 12096
rect 7300 12056 8668 12084
rect 6917 12047 6975 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9140 12084 9168 12112
rect 10226 12084 10232 12096
rect 9140 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 1104 11994 10120 12016
rect 1104 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 3202 11994
rect 3254 11942 3266 11994
rect 3318 11942 9010 11994
rect 9062 11942 9074 11994
rect 9126 11942 9138 11994
rect 9190 11942 9202 11994
rect 9254 11942 9266 11994
rect 9318 11942 10120 11994
rect 1104 11920 10120 11942
rect 3510 11880 3516 11892
rect 2746 11852 3516 11880
rect 842 11772 848 11824
rect 900 11812 906 11824
rect 900 11784 2268 11812
rect 900 11772 906 11784
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 2240 11753 2268 11784
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1360 11716 1685 11744
rect 1360 11704 1366 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2271 11716 2544 11744
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1486 11676 1492 11688
rect 992 11648 1492 11676
rect 992 11636 998 11648
rect 1486 11636 1492 11648
rect 1544 11676 1550 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1544 11648 1961 11676
rect 1544 11636 1550 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 2516 11676 2544 11716
rect 2746 11676 2774 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4246 11880 4252 11892
rect 4120 11852 4252 11880
rect 4120 11840 4126 11852
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5169 11883 5227 11889
rect 5169 11849 5181 11883
rect 5215 11880 5227 11883
rect 5258 11880 5264 11892
rect 5215 11852 5264 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 6549 11883 6607 11889
rect 6549 11849 6561 11883
rect 6595 11880 6607 11883
rect 7466 11880 7472 11892
rect 6595 11852 7472 11880
rect 6595 11849 6607 11852
rect 6549 11843 6607 11849
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 9398 11880 9404 11892
rect 8260 11852 9404 11880
rect 8260 11840 8266 11852
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 4062 11704 4068 11756
rect 4120 11753 4126 11756
rect 4120 11747 4148 11753
rect 4136 11713 4148 11747
rect 4120 11707 4148 11713
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 4985 11747 5043 11753
rect 4985 11744 4997 11747
rect 4939 11716 4997 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 4985 11713 4997 11716
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 4120 11704 4126 11707
rect 6454 11704 6460 11756
rect 6512 11704 6518 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7742 11744 7748 11756
rect 7064 11716 7748 11744
rect 7064 11704 7070 11716
rect 7742 11704 7748 11716
rect 7800 11704 7806 11756
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 10778 11744 10784 11756
rect 9723 11716 10784 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 2516 11648 2774 11676
rect 1949 11639 2007 11645
rect 3050 11636 3056 11688
rect 3108 11636 3114 11688
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11676 4307 11679
rect 6270 11676 6276 11688
rect 4295 11648 4660 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 566 11568 572 11620
rect 624 11608 630 11620
rect 1302 11608 1308 11620
rect 624 11580 1308 11608
rect 624 11568 630 11580
rect 1302 11568 1308 11580
rect 1360 11568 1366 11620
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 3697 11611 3755 11617
rect 3697 11608 3709 11611
rect 2924 11580 3709 11608
rect 2924 11568 2930 11580
rect 3697 11577 3709 11580
rect 3743 11577 3755 11611
rect 3697 11571 3755 11577
rect 1486 11500 1492 11552
rect 1544 11500 1550 11552
rect 2222 11500 2228 11552
rect 2280 11540 2286 11552
rect 2406 11540 2412 11552
rect 2280 11512 2412 11540
rect 2280 11500 2286 11512
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 2961 11543 3019 11549
rect 2961 11509 2973 11543
rect 3007 11540 3019 11543
rect 4632 11540 4660 11648
rect 4908 11648 6276 11676
rect 4908 11620 4936 11648
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 7524 11648 7573 11676
rect 7524 11636 7530 11648
rect 7561 11645 7573 11648
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 4890 11568 4896 11620
rect 4948 11568 4954 11620
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 6546 11608 6552 11620
rect 5868 11580 6552 11608
rect 5868 11568 5874 11580
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 7576 11608 7604 11639
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8352 11648 8493 11676
rect 8352 11636 8358 11648
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 8570 11636 8576 11688
rect 8628 11685 8634 11688
rect 8628 11679 8656 11685
rect 8644 11645 8656 11679
rect 8628 11639 8656 11645
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8938 11676 8944 11688
rect 8803 11648 8944 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 8628 11636 8634 11639
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9493 11679 9551 11685
rect 9493 11676 9505 11679
rect 9180 11648 9505 11676
rect 9180 11636 9186 11648
rect 9493 11645 9505 11648
rect 9539 11645 9551 11679
rect 9493 11639 9551 11645
rect 7926 11608 7932 11620
rect 7576 11580 7932 11608
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11577 8263 11611
rect 8205 11571 8263 11577
rect 3007 11512 4660 11540
rect 3007 11509 3019 11512
rect 2961 11503 3019 11509
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 6730 11540 6736 11552
rect 4764 11512 6736 11540
rect 4764 11500 4770 11512
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 8220 11540 8248 11571
rect 6972 11512 8248 11540
rect 8312 11540 8340 11636
rect 8662 11540 8668 11552
rect 8312 11512 8668 11540
rect 6972 11500 6978 11512
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9272 11512 9413 11540
rect 9272 11500 9278 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 1104 11450 10120 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 7950 11450
rect 8002 11398 8014 11450
rect 8066 11398 8078 11450
rect 8130 11398 8142 11450
rect 8194 11398 8206 11450
rect 8258 11398 10120 11450
rect 1104 11376 10120 11398
rect 2866 11296 2872 11348
rect 2924 11296 2930 11348
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 6822 11336 6828 11348
rect 4028 11308 6828 11336
rect 4028 11296 4034 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7282 11296 7288 11348
rect 7340 11296 7346 11348
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7432 11308 8033 11336
rect 7432 11296 7438 11308
rect 8021 11305 8033 11308
rect 8067 11305 8079 11339
rect 8021 11299 8079 11305
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11336 8631 11339
rect 8846 11336 8852 11348
rect 8619 11308 8852 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 10594 11336 10600 11348
rect 9232 11308 10600 11336
rect 842 11228 848 11280
rect 900 11268 906 11280
rect 1489 11271 1547 11277
rect 1489 11268 1501 11271
rect 900 11240 1501 11268
rect 900 11228 906 11240
rect 1489 11237 1501 11240
rect 1535 11237 1547 11271
rect 1489 11231 1547 11237
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 4338 11268 4344 11280
rect 4212 11240 4344 11268
rect 4212 11228 4218 11240
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 5626 11228 5632 11280
rect 5684 11268 5690 11280
rect 6089 11271 6147 11277
rect 6089 11268 6101 11271
rect 5684 11240 6101 11268
rect 5684 11228 5690 11240
rect 6089 11237 6101 11240
rect 6135 11237 6147 11271
rect 6089 11231 6147 11237
rect 7745 11271 7803 11277
rect 7745 11237 7757 11271
rect 7791 11268 7803 11271
rect 9232 11268 9260 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 7791 11240 9260 11268
rect 9677 11271 9735 11277
rect 7791 11237 7803 11240
rect 7745 11231 7803 11237
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 10226 11268 10232 11280
rect 9723 11240 10232 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 10226 11228 10232 11240
rect 10284 11228 10290 11280
rect 934 11160 940 11212
rect 992 11200 998 11212
rect 1857 11203 1915 11209
rect 1857 11200 1869 11203
rect 992 11172 1869 11200
rect 992 11160 998 11172
rect 1857 11169 1869 11172
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1872 11132 1900 11163
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 5534 11200 5540 11212
rect 3292 11172 5540 11200
rect 3292 11160 3298 11172
rect 5534 11160 5540 11172
rect 5592 11200 5598 11212
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 5592 11172 6377 11200
rect 5592 11160 5598 11172
rect 6365 11169 6377 11172
rect 6411 11169 6423 11203
rect 6365 11163 6423 11169
rect 6638 11160 6644 11212
rect 6696 11160 6702 11212
rect 8846 11200 8852 11212
rect 7944 11172 8852 11200
rect 2038 11132 2044 11144
rect 1872 11104 2044 11132
rect 1673 11095 1731 11101
rect 1688 11064 1716 11095
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11132 2191 11135
rect 2406 11132 2412 11144
rect 2179 11104 2412 11132
rect 2179 11101 2191 11104
rect 2133 11095 2191 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 4890 11132 4896 11144
rect 4488 11104 4896 11132
rect 4488 11092 4494 11104
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5074 11092 5080 11144
rect 5132 11132 5138 11144
rect 5445 11135 5503 11141
rect 5445 11132 5457 11135
rect 5132 11104 5457 11132
rect 5132 11092 5138 11104
rect 5445 11101 5457 11104
rect 5491 11101 5503 11135
rect 5445 11095 5503 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 5810 11132 5816 11144
rect 5675 11104 5816 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6454 11092 6460 11144
rect 6512 11141 6518 11144
rect 7944 11141 7972 11172
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 9122 11160 9128 11212
rect 9180 11160 9186 11212
rect 9214 11160 9220 11212
rect 9272 11160 9278 11212
rect 6512 11135 6540 11141
rect 6528 11101 6540 11135
rect 6512 11095 6540 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 6512 11092 6518 11095
rect 1946 11064 1952 11076
rect 1688 11036 1952 11064
rect 1946 11024 1952 11036
rect 2004 11024 2010 11076
rect 8220 11064 8248 11095
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 8757 11135 8815 11141
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9950 11132 9956 11144
rect 8803 11104 9956 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 9858 11064 9864 11076
rect 8220 11036 9864 11064
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 934 10956 940 11008
rect 992 10996 998 11008
rect 1394 10996 1400 11008
rect 992 10968 1400 10996
rect 992 10956 998 10968
rect 1394 10956 1400 10968
rect 1452 10956 1458 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6914 10996 6920 11008
rect 6512 10968 6920 10996
rect 6512 10956 6518 10968
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 8570 10996 8576 11008
rect 7340 10968 8576 10996
rect 7340 10956 7346 10968
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8754 10956 8760 11008
rect 8812 10996 8818 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 8812 10968 9321 10996
rect 8812 10956 8818 10968
rect 9309 10965 9321 10968
rect 9355 10965 9367 10999
rect 9309 10959 9367 10965
rect 1104 10906 10120 10928
rect 1104 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 3202 10906
rect 3254 10854 3266 10906
rect 3318 10854 9010 10906
rect 9062 10854 9074 10906
rect 9126 10854 9138 10906
rect 9190 10854 9202 10906
rect 9254 10854 9266 10906
rect 9318 10854 10120 10906
rect 1104 10832 10120 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 1946 10792 1952 10804
rect 1535 10764 1952 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 5718 10792 5724 10804
rect 3099 10764 5724 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 5718 10752 5724 10764
rect 5776 10792 5782 10804
rect 6822 10792 6828 10804
rect 5776 10764 6828 10792
rect 5776 10752 5782 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 7558 10752 7564 10804
rect 7616 10752 7622 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 8352 10764 9505 10792
rect 8352 10752 8358 10764
rect 9493 10761 9505 10764
rect 9539 10761 9551 10795
rect 9493 10755 9551 10761
rect 2866 10724 2872 10736
rect 1780 10696 2872 10724
rect 1394 10616 1400 10668
rect 1452 10656 1458 10668
rect 1780 10665 1808 10696
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 3694 10684 3700 10736
rect 3752 10724 3758 10736
rect 3789 10727 3847 10733
rect 3789 10724 3801 10727
rect 3752 10696 3801 10724
rect 3752 10684 3758 10696
rect 3789 10693 3801 10696
rect 3835 10693 3847 10727
rect 3789 10687 3847 10693
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 5132 10696 7144 10724
rect 5132 10684 5138 10696
rect 1765 10659 1823 10665
rect 1765 10656 1777 10659
rect 1452 10628 1777 10656
rect 1452 10616 1458 10628
rect 1765 10625 1777 10628
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2406 10656 2412 10668
rect 2363 10628 2412 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 2746 10628 3617 10656
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10557 2099 10591
rect 2041 10551 2099 10557
rect 1949 10523 2007 10529
rect 1949 10489 1961 10523
rect 1995 10520 2007 10523
rect 2056 10520 2084 10551
rect 1995 10492 2084 10520
rect 1995 10489 2007 10492
rect 1949 10483 2007 10489
rect 2056 10452 2084 10492
rect 2498 10452 2504 10464
rect 2056 10424 2504 10452
rect 2498 10412 2504 10424
rect 2556 10452 2562 10464
rect 2746 10452 2774 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 5994 10656 6000 10668
rect 5399 10628 6000 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6788 10628 6837 10656
rect 6788 10616 6794 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4948 10560 5089 10588
rect 4948 10548 4954 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6362 10588 6368 10600
rect 5868 10560 6368 10588
rect 5868 10548 5874 10560
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 7116 10588 7144 10696
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7432 10628 7665 10656
rect 7432 10616 7438 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 8662 10616 8668 10668
rect 8720 10665 8726 10668
rect 8720 10659 8748 10665
rect 8736 10625 8748 10659
rect 8720 10619 8748 10625
rect 8720 10616 8726 10619
rect 9766 10616 9772 10668
rect 9824 10616 9830 10668
rect 7558 10588 7564 10600
rect 7116 10560 7564 10588
rect 7558 10548 7564 10560
rect 7616 10588 7622 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7616 10560 7849 10588
rect 7616 10548 7622 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 7837 10551 7895 10557
rect 8429 10560 8585 10588
rect 5169 10523 5227 10529
rect 5169 10489 5181 10523
rect 5215 10520 5227 10523
rect 5442 10520 5448 10532
rect 5215 10492 5448 10520
rect 5215 10489 5227 10492
rect 5169 10483 5227 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 8294 10480 8300 10532
rect 8352 10480 8358 10532
rect 2556 10424 2774 10452
rect 2556 10412 2562 10424
rect 2866 10412 2872 10464
rect 2924 10452 2930 10464
rect 3697 10455 3755 10461
rect 3697 10452 3709 10455
rect 2924 10424 3709 10452
rect 2924 10412 2930 10424
rect 3697 10421 3709 10424
rect 3743 10421 3755 10455
rect 3697 10415 3755 10421
rect 5258 10412 5264 10464
rect 5316 10412 5322 10464
rect 8429 10452 8457 10560
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8846 10548 8852 10600
rect 8904 10548 8910 10600
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9548 10560 9628 10588
rect 9548 10548 9554 10560
rect 9600 10529 9628 10560
rect 9585 10523 9643 10529
rect 9585 10489 9597 10523
rect 9631 10489 9643 10523
rect 9585 10483 9643 10489
rect 9490 10452 9496 10464
rect 8429 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 1104 10362 10120 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 7950 10362
rect 8002 10310 8014 10362
rect 8066 10310 8078 10362
rect 8130 10310 8142 10362
rect 8194 10310 8206 10362
rect 8258 10310 10120 10362
rect 1104 10288 10120 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1949 10251 2007 10257
rect 1949 10248 1961 10251
rect 1544 10220 1961 10248
rect 1544 10208 1550 10220
rect 1949 10217 1961 10220
rect 1995 10217 2007 10251
rect 4062 10248 4068 10260
rect 1949 10211 2007 10217
rect 2700 10220 4068 10248
rect 2700 10180 2728 10220
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 6178 10248 6184 10260
rect 5040 10220 6184 10248
rect 5040 10208 5046 10220
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8846 10248 8852 10260
rect 7883 10220 8852 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 1964 10152 2728 10180
rect 4801 10183 4859 10189
rect 1964 10056 1992 10152
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 5074 10180 5080 10192
rect 4847 10152 5080 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 5074 10140 5080 10152
rect 5132 10180 5138 10192
rect 5132 10152 5212 10180
rect 5132 10140 5138 10152
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 5184 10121 5212 10152
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 5316 10152 6500 10180
rect 5316 10140 5322 10152
rect 6472 10124 6500 10152
rect 8478 10140 8484 10192
rect 8536 10140 8542 10192
rect 2593 10115 2651 10121
rect 2593 10112 2605 10115
rect 2556 10084 2605 10112
rect 2556 10072 2562 10084
rect 2593 10081 2605 10084
rect 2639 10081 2651 10115
rect 2593 10075 2651 10081
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10081 5227 10115
rect 5169 10075 5227 10081
rect 1026 10004 1032 10056
rect 1084 10044 1090 10056
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1084 10016 1685 10044
rect 1084 10004 1090 10016
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 1946 10044 1952 10056
rect 1903 10016 1952 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2608 9976 2636 10075
rect 6454 10072 6460 10124
rect 6512 10072 6518 10124
rect 6822 10072 6828 10124
rect 6880 10072 6886 10124
rect 7466 10072 7472 10124
rect 7524 10112 7530 10124
rect 8202 10112 8208 10124
rect 7524 10084 8208 10112
rect 7524 10072 7530 10084
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9674 10112 9680 10124
rect 8404 10084 9680 10112
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 2869 10047 2927 10053
rect 2869 10044 2881 10047
rect 2832 10016 2881 10044
rect 2832 10004 2838 10016
rect 2869 10013 2881 10016
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3804 9976 3832 10007
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5261 10047 5319 10053
rect 5261 10044 5273 10047
rect 4764 10016 5273 10044
rect 4764 10004 4770 10016
rect 5261 10013 5273 10016
rect 5307 10013 5319 10047
rect 5261 10007 5319 10013
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 5810 10044 5816 10056
rect 5491 10016 5816 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 8404 10053 8432 10084
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9766 10072 9772 10124
rect 9824 10072 9830 10124
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 7064 10016 7113 10044
rect 7064 10004 7070 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 8389 10047 8447 10053
rect 8389 10013 8401 10047
rect 8435 10013 8447 10047
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 8389 10007 8447 10013
rect 8496 10016 9505 10044
rect 4890 9976 4896 9988
rect 2608 9948 3832 9976
rect 4724 9948 4896 9976
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 4724 9908 4752 9948
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5077 9979 5135 9985
rect 5077 9976 5089 9979
rect 5040 9948 5089 9976
rect 5040 9936 5046 9948
rect 5077 9945 5089 9948
rect 5123 9945 5135 9979
rect 5077 9939 5135 9945
rect 5537 9979 5595 9985
rect 5537 9945 5549 9979
rect 5583 9945 5595 9979
rect 5537 9939 5595 9945
rect 6273 9979 6331 9985
rect 6273 9945 6285 9979
rect 6319 9976 6331 9979
rect 7282 9976 7288 9988
rect 6319 9948 7288 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 3651 9880 4752 9908
rect 5552 9908 5580 9939
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8496 9976 8524 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 8168 9948 8524 9976
rect 8665 9979 8723 9985
rect 8168 9936 8174 9948
rect 8665 9945 8677 9979
rect 8711 9976 8723 9979
rect 10042 9976 10048 9988
rect 8711 9948 10048 9976
rect 8711 9945 8723 9948
rect 8665 9939 8723 9945
rect 10042 9936 10048 9948
rect 10100 9936 10106 9988
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 5552 9880 5917 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 5905 9871 5963 9877
rect 6362 9868 6368 9920
rect 6420 9868 6426 9920
rect 8018 9868 8024 9920
rect 8076 9908 8082 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 8076 9880 8217 9908
rect 8076 9868 8082 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 9490 9908 9496 9920
rect 8619 9880 9496 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 1104 9818 10120 9840
rect 1104 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 3202 9818
rect 3254 9766 3266 9818
rect 3318 9766 9010 9818
rect 9062 9766 9074 9818
rect 9126 9766 9138 9818
rect 9190 9766 9202 9818
rect 9254 9766 9266 9818
rect 9318 9766 10120 9818
rect 1104 9744 10120 9766
rect 474 9664 480 9716
rect 532 9704 538 9716
rect 3878 9704 3884 9716
rect 532 9676 3884 9704
rect 532 9664 538 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4706 9664 4712 9716
rect 4764 9664 4770 9716
rect 5353 9707 5411 9713
rect 5353 9673 5365 9707
rect 5399 9704 5411 9707
rect 5442 9704 5448 9716
rect 5399 9676 5448 9704
rect 5399 9673 5411 9676
rect 5353 9667 5411 9673
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 8110 9704 8116 9716
rect 5684 9676 8116 9704
rect 5684 9664 5690 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8294 9664 8300 9716
rect 8352 9664 8358 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 10870 9704 10876 9716
rect 8628 9676 10876 9704
rect 8628 9664 8634 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 3694 9636 3700 9648
rect 1688 9608 3700 9636
rect 1688 9577 1716 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 4798 9636 4804 9648
rect 4571 9608 4804 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 4798 9596 4804 9608
rect 4856 9596 4862 9648
rect 5810 9596 5816 9648
rect 5868 9645 5874 9648
rect 5868 9639 5917 9645
rect 5868 9605 5871 9639
rect 5905 9605 5917 9639
rect 8754 9636 8760 9648
rect 5868 9599 5917 9605
rect 6932 9608 8760 9636
rect 5868 9596 5874 9599
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2556 9540 2697 9568
rect 2556 9528 2562 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3418 9568 3424 9580
rect 3007 9540 3424 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 4982 9528 4988 9580
rect 5040 9528 5046 9580
rect 5074 9528 5080 9580
rect 5132 9528 5138 9580
rect 5215 9571 5273 9577
rect 5215 9537 5227 9571
rect 5261 9537 5273 9571
rect 5215 9531 5273 9537
rect 5230 9500 5258 9531
rect 5442 9528 5448 9580
rect 5500 9528 5506 9580
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 5962 9570 6020 9576
rect 5962 9536 5974 9570
rect 6008 9536 6020 9570
rect 5092 9472 5258 9500
rect 5092 9444 5120 9472
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5552 9500 5580 9531
rect 5408 9472 5580 9500
rect 5736 9500 5764 9531
rect 5962 9530 6020 9536
rect 5810 9500 5816 9512
rect 5736 9472 5816 9500
rect 5408 9460 5414 9472
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4157 9435 4215 9441
rect 4157 9432 4169 9435
rect 3743 9404 4169 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 4157 9401 4169 9404
rect 4203 9432 4215 9435
rect 4203 9404 4936 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 1486 9324 1492 9376
rect 1544 9324 1550 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4798 9324 4804 9376
rect 4856 9324 4862 9376
rect 4908 9364 4936 9404
rect 5074 9392 5080 9444
rect 5132 9392 5138 9444
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 5629 9435 5687 9441
rect 5629 9432 5641 9435
rect 5500 9404 5641 9432
rect 5500 9392 5506 9404
rect 5629 9401 5641 9404
rect 5675 9401 5687 9435
rect 5977 9432 6005 9530
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6932 9577 6960 9608
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6512 9540 6561 9568
rect 6512 9528 6518 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6917 9571 6975 9577
rect 6917 9537 6929 9571
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7524 9540 7573 9568
rect 7524 9528 7530 9540
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 8386 9528 8392 9580
rect 8444 9568 8450 9580
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 8444 9540 8585 9568
rect 8444 9528 8450 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 6880 9472 7297 9500
rect 6880 9460 6886 9472
rect 7285 9469 7297 9472
rect 7331 9469 7343 9503
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 7285 9463 7343 9469
rect 8588 9472 9505 9500
rect 6086 9432 6092 9444
rect 5977 9404 6092 9432
rect 5629 9395 5687 9401
rect 6086 9392 6092 9404
rect 6144 9432 6150 9444
rect 6144 9404 6592 9432
rect 6144 9392 6150 9404
rect 5258 9364 5264 9376
rect 4908 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 6564 9373 6592 9404
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 6328 9336 6377 9364
rect 6328 9324 6334 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7374 9364 7380 9376
rect 6972 9336 7380 9364
rect 6972 9324 6978 9336
rect 7374 9324 7380 9336
rect 7432 9364 7438 9376
rect 8588 9364 8616 9472
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 9766 9460 9772 9512
rect 9824 9460 9830 9512
rect 7432 9336 8616 9364
rect 8665 9367 8723 9373
rect 7432 9324 7438 9336
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 9490 9364 9496 9376
rect 8711 9336 9496 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 1104 9274 10120 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 7950 9274
rect 8002 9222 8014 9274
rect 8066 9222 8078 9274
rect 8130 9222 8142 9274
rect 8194 9222 8206 9274
rect 8258 9222 10120 9274
rect 1104 9200 10120 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2406 9160 2412 9172
rect 2004 9132 2412 9160
rect 2004 9120 2010 9132
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6454 9160 6460 9172
rect 5868 9132 6460 9160
rect 5868 9120 5874 9132
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 8297 9095 8355 9101
rect 8297 9092 8309 9095
rect 6972 9064 8309 9092
rect 6972 9052 6978 9064
rect 8297 9061 8309 9064
rect 8343 9061 8355 9095
rect 8297 9055 8355 9061
rect 8478 9052 8484 9104
rect 8536 9092 8542 9104
rect 8846 9092 8852 9104
rect 8536 9064 8852 9092
rect 8536 9052 8542 9064
rect 8846 9052 8852 9064
rect 8904 9052 8910 9104
rect 9306 9052 9312 9104
rect 9364 9092 9370 9104
rect 9493 9095 9551 9101
rect 9493 9092 9505 9095
rect 9364 9064 9505 9092
rect 9364 9052 9370 9064
rect 9493 9061 9505 9064
rect 9539 9061 9551 9095
rect 9493 9055 9551 9061
rect 9858 9024 9864 9036
rect 7852 8996 9864 9024
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 4798 8956 4804 8968
rect 1719 8928 4804 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 7852 8965 7880 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8925 7895 8959
rect 7964 8959 8022 8965
rect 7964 8956 7976 8959
rect 7837 8919 7895 8925
rect 7944 8925 7976 8956
rect 8010 8925 8022 8959
rect 7944 8919 8022 8925
rect 8067 8959 8125 8965
rect 8067 8925 8079 8959
rect 8113 8956 8125 8959
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8113 8928 8217 8956
rect 8113 8925 8125 8928
rect 8067 8919 8125 8925
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 7944 8888 7972 8919
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8444 8928 8493 8956
rect 8444 8916 8450 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8481 8919 8539 8925
rect 8588 8928 9137 8956
rect 8588 8888 8616 8928
rect 9125 8925 9137 8928
rect 9171 8956 9183 8959
rect 9398 8956 9404 8968
rect 9171 8928 9404 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 9398 8916 9404 8928
rect 9456 8956 9462 8968
rect 9582 8956 9588 8968
rect 9456 8928 9588 8956
rect 9456 8916 9462 8928
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 7944 8860 8616 8888
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 8904 8860 8953 8888
rect 8904 8848 8910 8860
rect 8941 8857 8953 8860
rect 8987 8857 8999 8891
rect 8941 8851 8999 8857
rect 9674 8848 9680 8900
rect 9732 8848 9738 8900
rect 842 8780 848 8832
rect 900 8820 906 8832
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 900 8792 1501 8820
rect 900 8780 906 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 1489 8783 1547 8789
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2498 8820 2504 8832
rect 2280 8792 2504 8820
rect 2280 8780 2286 8792
rect 2498 8780 2504 8792
rect 2556 8820 2562 8832
rect 6546 8820 6552 8832
rect 2556 8792 6552 8820
rect 2556 8780 2562 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 7558 8820 7564 8832
rect 7064 8792 7564 8820
rect 7064 8780 7070 8792
rect 7558 8780 7564 8792
rect 7616 8820 7622 8832
rect 7653 8823 7711 8829
rect 7653 8820 7665 8823
rect 7616 8792 7665 8820
rect 7616 8780 7622 8792
rect 7653 8789 7665 8792
rect 7699 8820 7711 8823
rect 8202 8820 8208 8832
rect 7699 8792 8208 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8665 8823 8723 8829
rect 8665 8789 8677 8823
rect 8711 8820 8723 8823
rect 8754 8820 8760 8832
rect 8711 8792 8760 8820
rect 8711 8789 8723 8792
rect 8665 8783 8723 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9309 8823 9367 8829
rect 9309 8789 9321 8823
rect 9355 8820 9367 8823
rect 9398 8820 9404 8832
rect 9355 8792 9404 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 1104 8730 10120 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 10120 8730
rect 1104 8656 10120 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1268 8588 1961 8616
rect 1268 8576 1274 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 1949 8579 2007 8585
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 8260 8588 8800 8616
rect 8260 8576 8266 8588
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 1670 8548 1676 8560
rect 1535 8520 1676 8548
rect 1535 8517 1547 8520
rect 1489 8511 1547 8517
rect 1670 8508 1676 8520
rect 1728 8508 1734 8560
rect 1854 8508 1860 8560
rect 1912 8508 1918 8560
rect 8772 8548 8800 8588
rect 8846 8576 8852 8628
rect 8904 8616 8910 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 8904 8588 8953 8616
rect 8904 8576 8910 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 9493 8551 9551 8557
rect 9493 8548 9505 8551
rect 8772 8520 9505 8548
rect 9493 8517 9505 8520
rect 9539 8517 9551 8551
rect 9493 8511 9551 8517
rect 1872 8480 1900 8508
rect 2593 8483 2651 8489
rect 2593 8480 2605 8483
rect 1872 8452 2605 8480
rect 2593 8449 2605 8452
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 4062 8480 4068 8492
rect 3476 8452 4068 8480
rect 3476 8440 3482 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 6362 8480 6368 8492
rect 5868 8452 6368 8480
rect 5868 8440 5874 8452
rect 6362 8440 6368 8452
rect 6420 8480 6426 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6420 8452 7297 8480
rect 6420 8440 6426 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 290 8372 296 8424
rect 348 8412 354 8424
rect 1673 8415 1731 8421
rect 1673 8412 1685 8415
rect 348 8384 1685 8412
rect 348 8372 354 8384
rect 1673 8381 1685 8384
rect 1719 8381 1731 8415
rect 1673 8375 1731 8381
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 2280 8384 2329 8412
rect 2280 8372 2286 8384
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 7006 8412 7012 8424
rect 4764 8384 7012 8412
rect 4764 8372 4770 8384
rect 7006 8372 7012 8384
rect 7064 8412 7070 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 7064 8384 7113 8412
rect 7064 8372 7070 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7300 8412 7328 8443
rect 7374 8412 7380 8424
rect 7300 8384 7380 8412
rect 7101 8375 7159 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 8202 8421 8208 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7852 8384 8033 8412
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8344 3387 8347
rect 4062 8344 4068 8356
rect 3375 8316 4068 8344
rect 3375 8313 3387 8316
rect 3329 8307 3387 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 5718 8304 5724 8356
rect 5776 8344 5782 8356
rect 7745 8347 7803 8353
rect 7745 8344 7757 8347
rect 5776 8316 7757 8344
rect 5776 8304 5782 8316
rect 7745 8313 7757 8316
rect 7791 8313 7803 8347
rect 7745 8307 7803 8313
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 5534 8276 5540 8288
rect 4212 8248 5540 8276
rect 4212 8236 4218 8248
rect 5534 8236 5540 8248
rect 5592 8276 5598 8288
rect 7558 8276 7564 8288
rect 5592 8248 7564 8276
rect 5592 8236 5598 8248
rect 7558 8236 7564 8248
rect 7616 8276 7622 8288
rect 7852 8276 7880 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 8159 8415 8208 8421
rect 8159 8381 8171 8415
rect 8205 8381 8208 8415
rect 8159 8375 8208 8381
rect 8202 8372 8208 8375
rect 8260 8372 8266 8424
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8412 8355 8415
rect 8478 8412 8484 8424
rect 8343 8384 8484 8412
rect 8343 8381 8355 8384
rect 8297 8375 8355 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9416 8412 9444 8443
rect 8720 8384 9444 8412
rect 9585 8415 9643 8421
rect 8720 8372 8726 8384
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 9600 8344 9628 8375
rect 8904 8316 9628 8344
rect 8904 8304 8910 8316
rect 7616 8248 7880 8276
rect 7616 8236 7622 8248
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 9033 8279 9091 8285
rect 9033 8276 9045 8279
rect 8536 8248 9045 8276
rect 8536 8236 8542 8248
rect 9033 8245 9045 8248
rect 9079 8245 9091 8279
rect 9033 8239 9091 8245
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 9398 8276 9404 8288
rect 9272 8248 9404 8276
rect 9272 8236 9278 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 1104 8186 10120 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 10120 8186
rect 1104 8112 10120 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 6362 8072 6368 8084
rect 2547 8044 6368 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 6914 8032 6920 8084
rect 6972 8032 6978 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8662 8072 8668 8084
rect 8619 8044 8668 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 8938 8032 8944 8084
rect 8996 8032 9002 8084
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 10226 8072 10232 8084
rect 9456 8044 10232 8072
rect 9456 8032 9462 8044
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 4798 7964 4804 8016
rect 4856 8004 4862 8016
rect 5258 8004 5264 8016
rect 4856 7976 5264 8004
rect 4856 7964 4862 7976
rect 2222 7896 2228 7948
rect 2280 7936 2286 7948
rect 2498 7936 2504 7948
rect 2280 7908 2504 7936
rect 2280 7896 2286 7908
rect 2498 7896 2504 7908
rect 2556 7936 2562 7948
rect 5092 7945 5120 7976
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 5718 7964 5724 8016
rect 5776 7964 5782 8016
rect 7742 7964 7748 8016
rect 7800 7964 7806 8016
rect 9858 8004 9864 8016
rect 7944 7976 9864 8004
rect 2593 7939 2651 7945
rect 2593 7936 2605 7939
rect 2556 7908 2605 7936
rect 2556 7896 2562 7908
rect 2593 7905 2605 7908
rect 2639 7905 2651 7939
rect 2593 7899 2651 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7905 5135 7939
rect 5350 7936 5356 7948
rect 5077 7899 5135 7905
rect 5276 7908 5356 7936
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 1504 7800 1532 7831
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 5276 7877 5304 7908
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 5997 7939 6055 7945
rect 5997 7936 6009 7939
rect 5684 7908 6009 7936
rect 5684 7896 5690 7908
rect 5997 7905 6009 7908
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 6086 7896 6092 7948
rect 6144 7945 6150 7948
rect 6144 7939 6172 7945
rect 6160 7905 6172 7939
rect 6144 7899 6172 7905
rect 6144 7896 6150 7899
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1728 7840 1777 7868
rect 1728 7828 1734 7840
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 1765 7831 1823 7837
rect 2746 7840 2881 7868
rect 2222 7800 2228 7812
rect 1504 7772 2228 7800
rect 2222 7760 2228 7772
rect 2280 7760 2286 7812
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2746 7800 2774 7840
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 6270 7828 6276 7880
rect 6328 7828 6334 7880
rect 7944 7877 7972 7976
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 9674 7936 9680 7948
rect 8312 7908 9680 7936
rect 8312 7877 8340 7908
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8297 7871 8355 7877
rect 8297 7837 8309 7871
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8812 7840 9137 7868
rect 8812 7828 8818 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 9398 7868 9404 7880
rect 9355 7840 9404 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9490 7828 9496 7880
rect 9548 7828 9554 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 10962 7868 10968 7880
rect 9815 7840 10968 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 2372 7772 2774 7800
rect 2372 7760 2378 7772
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 8113 7803 8171 7809
rect 8113 7800 8125 7803
rect 7340 7772 8125 7800
rect 7340 7760 7346 7772
rect 8113 7769 8125 7772
rect 8159 7769 8171 7803
rect 8113 7763 8171 7769
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 9950 7800 9956 7812
rect 8711 7772 9956 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 9950 7760 9956 7772
rect 10008 7760 10014 7812
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4798 7732 4804 7744
rect 3651 7704 4804 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 6270 7732 6276 7744
rect 5132 7704 6276 7732
rect 5132 7692 5138 7704
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 9585 7735 9643 7741
rect 9585 7732 9597 7735
rect 7616 7704 9597 7732
rect 7616 7692 7622 7704
rect 9585 7701 9597 7704
rect 9631 7701 9643 7735
rect 9585 7695 9643 7701
rect 1104 7642 10120 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 10120 7642
rect 1104 7568 10120 7590
rect 1486 7488 1492 7540
rect 1544 7488 1550 7540
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 2406 7488 2412 7540
rect 2464 7488 2470 7540
rect 3697 7531 3755 7537
rect 3697 7497 3709 7531
rect 3743 7528 3755 7531
rect 3743 7500 5948 7528
rect 3743 7497 3755 7500
rect 3697 7491 3755 7497
rect 2314 7420 2320 7472
rect 2372 7420 2378 7472
rect 2682 7420 2688 7472
rect 2740 7420 2746 7472
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2700 7392 2728 7420
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 1995 7364 2973 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 1688 7256 1716 7355
rect 4154 7352 4160 7404
rect 4212 7352 4218 7404
rect 2222 7284 2228 7336
rect 2280 7324 2286 7336
rect 2685 7327 2743 7333
rect 2685 7324 2697 7327
rect 2280 7296 2697 7324
rect 2280 7284 2286 7296
rect 2685 7293 2697 7296
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 4706 7324 4712 7336
rect 4387 7296 4712 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4798 7284 4804 7336
rect 4856 7284 4862 7336
rect 5258 7333 5264 7336
rect 5077 7327 5135 7333
rect 5077 7324 5089 7327
rect 4908 7296 5089 7324
rect 3970 7256 3976 7268
rect 1688 7228 2820 7256
rect 14 7148 20 7200
rect 72 7188 78 7200
rect 2682 7188 2688 7200
rect 72 7160 2688 7188
rect 72 7148 78 7160
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 2792 7188 2820 7228
rect 3344 7228 3976 7256
rect 3344 7188 3372 7228
rect 3970 7216 3976 7228
rect 4028 7216 4034 7268
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 4908 7256 4936 7296
rect 5077 7293 5089 7296
rect 5123 7293 5135 7327
rect 5077 7287 5135 7293
rect 5215 7327 5264 7333
rect 5215 7293 5227 7327
rect 5261 7293 5264 7327
rect 5215 7287 5264 7293
rect 5258 7284 5264 7287
rect 5316 7284 5322 7336
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7316 5411 7327
rect 5920 7324 5948 7500
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 7190 7528 7196 7540
rect 7147 7500 7196 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7708 7500 7757 7528
rect 7708 7488 7714 7500
rect 7745 7497 7757 7500
rect 7791 7497 7803 7531
rect 9674 7528 9680 7540
rect 7745 7491 7803 7497
rect 7944 7500 9680 7528
rect 7469 7463 7527 7469
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 7515 7432 7880 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 6457 7395 6515 7401
rect 6457 7361 6469 7395
rect 6503 7392 6515 7395
rect 6638 7392 6644 7404
rect 6503 7364 6644 7392
rect 6503 7361 6515 7364
rect 6457 7355 6515 7361
rect 6638 7352 6644 7364
rect 6696 7352 6702 7404
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 5460 7316 5948 7324
rect 5399 7296 5948 7316
rect 5997 7327 6055 7333
rect 5399 7293 5488 7296
rect 5353 7288 5488 7293
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6748 7324 6776 7355
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 7561 7395 7619 7401
rect 7561 7390 7573 7395
rect 7484 7362 7573 7390
rect 7484 7324 7512 7362
rect 7561 7361 7573 7362
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 6043 7296 6776 7324
rect 7208 7296 7512 7324
rect 7852 7324 7880 7432
rect 7944 7401 7972 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 8478 7420 8484 7472
rect 8536 7420 8542 7472
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 9950 7460 9956 7472
rect 8628 7432 9956 7460
rect 8628 7420 8634 7432
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8202 7392 8208 7404
rect 8159 7364 8208 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7392 8447 7395
rect 8662 7392 8668 7404
rect 8435 7364 8668 7392
rect 8435 7361 8447 7364
rect 8389 7355 8447 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8846 7352 8852 7404
rect 8904 7352 8910 7404
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9398 7392 9404 7404
rect 9171 7364 9404 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 8754 7324 8760 7336
rect 7852 7296 8760 7324
rect 6043 7293 6055 7296
rect 5353 7287 5411 7288
rect 5997 7287 6055 7293
rect 4672 7228 4936 7256
rect 6641 7259 6699 7265
rect 4672 7216 4678 7228
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 6822 7256 6828 7268
rect 6687 7228 6828 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 6822 7216 6828 7228
rect 6880 7216 6886 7268
rect 2792 7160 3372 7188
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 7208 7188 7236 7296
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 7466 7256 7472 7268
rect 7340 7228 7472 7256
rect 7340 7216 7346 7228
rect 7466 7216 7472 7228
rect 7524 7216 7530 7268
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 7708 7228 8217 7256
rect 7708 7216 7714 7228
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 8864 7256 8892 7352
rect 9214 7333 9220 7336
rect 9213 7287 9220 7333
rect 9214 7284 9220 7287
rect 9272 7284 9278 7336
rect 9401 7259 9459 7265
rect 9401 7256 9413 7259
rect 8864 7228 9413 7256
rect 8205 7219 8263 7225
rect 9401 7225 9413 7228
rect 9447 7225 9459 7259
rect 9401 7219 9459 7225
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 9585 7259 9643 7265
rect 9585 7256 9597 7259
rect 9548 7228 9597 7256
rect 9548 7216 9554 7228
rect 9585 7225 9597 7228
rect 9631 7225 9643 7259
rect 9585 7219 9643 7225
rect 5408 7160 7236 7188
rect 5408 7148 5414 7160
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7892 7160 8033 7188
rect 7892 7148 7898 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 8570 7148 8576 7200
rect 8628 7148 8634 7200
rect 8846 7148 8852 7200
rect 8904 7188 8910 7200
rect 9033 7191 9091 7197
rect 9033 7188 9045 7191
rect 8904 7160 9045 7188
rect 8904 7148 8910 7160
rect 9033 7157 9045 7160
rect 9079 7188 9091 7191
rect 9214 7188 9220 7200
rect 9079 7160 9220 7188
rect 9079 7157 9091 7160
rect 9033 7151 9091 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9306 7148 9312 7200
rect 9364 7148 9370 7200
rect 1104 7098 10120 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 10120 7098
rect 1104 7024 10120 7046
rect 5350 6984 5356 6996
rect 5000 6956 5356 6984
rect 4430 6808 4436 6860
rect 4488 6848 4494 6860
rect 5000 6857 5028 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5442 6944 5448 6996
rect 5500 6984 5506 6996
rect 5994 6984 6000 6996
rect 5500 6956 6000 6984
rect 5500 6944 5506 6956
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 6825 6987 6883 6993
rect 6825 6984 6837 6987
rect 6696 6956 6837 6984
rect 6696 6944 6702 6956
rect 6825 6953 6837 6956
rect 6871 6953 6883 6987
rect 6825 6947 6883 6953
rect 7837 6987 7895 6993
rect 7837 6953 7849 6987
rect 7883 6984 7895 6987
rect 8846 6984 8852 6996
rect 7883 6956 8852 6984
rect 7883 6953 7895 6956
rect 7837 6947 7895 6953
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 7469 6919 7527 6925
rect 7469 6916 7481 6919
rect 7432 6888 7481 6916
rect 7432 6876 7438 6888
rect 7469 6885 7481 6888
rect 7515 6885 7527 6919
rect 7469 6879 7527 6885
rect 7650 6876 7656 6928
rect 7708 6916 7714 6928
rect 8021 6919 8079 6925
rect 8021 6916 8033 6919
rect 7708 6888 8033 6916
rect 7708 6876 7714 6888
rect 8021 6885 8033 6888
rect 8067 6885 8079 6919
rect 10686 6916 10692 6928
rect 8021 6879 8079 6885
rect 9508 6888 10692 6916
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4488 6820 4997 6848
rect 4488 6808 4494 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6848 5227 6851
rect 5534 6848 5540 6860
rect 5215 6820 5540 6848
rect 5215 6817 5227 6820
rect 5169 6811 5227 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 5905 6851 5963 6857
rect 5905 6848 5917 6851
rect 5776 6820 5917 6848
rect 5776 6808 5782 6820
rect 5905 6817 5917 6820
rect 5951 6817 5963 6851
rect 5905 6811 5963 6817
rect 5994 6808 6000 6860
rect 6052 6857 6058 6860
rect 6052 6851 6080 6857
rect 6068 6817 6080 6851
rect 6052 6811 6080 6817
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 6362 6848 6368 6860
rect 6227 6820 6368 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6052 6808 6058 6811
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6748 6820 7788 6848
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 1912 6752 2145 6780
rect 1912 6740 1918 6752
rect 2133 6749 2145 6752
rect 2179 6749 2191 6783
rect 2133 6743 2191 6749
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6780 2467 6783
rect 2590 6780 2596 6792
rect 2455 6752 2596 6780
rect 2455 6749 2467 6752
rect 2409 6743 2467 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 1397 6647 1455 6653
rect 1397 6613 1409 6647
rect 1443 6644 1455 6647
rect 1670 6644 1676 6656
rect 1443 6616 1676 6644
rect 1443 6613 1455 6616
rect 1397 6607 1455 6613
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 5626 6644 5632 6656
rect 4120 6616 5632 6644
rect 4120 6604 4126 6616
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6748 6644 6776 6820
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7760 6780 7788 6820
rect 7834 6808 7840 6860
rect 7892 6848 7898 6860
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 7892 6820 8309 6848
rect 7892 6808 7898 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 9306 6848 9312 6860
rect 8711 6820 9312 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9508 6857 9536 6888
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7760 6752 8125 6780
rect 7377 6743 7435 6749
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 7392 6712 7420 6743
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8260 6752 8401 6780
rect 8260 6740 8266 6752
rect 8389 6749 8401 6752
rect 8435 6780 8447 6783
rect 8478 6780 8484 6792
rect 8435 6752 8484 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 9674 6712 9680 6724
rect 7392 6684 9680 6712
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 5776 6616 6776 6644
rect 5776 6604 5782 6616
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7193 6647 7251 6653
rect 7193 6644 7205 6647
rect 7156 6616 7205 6644
rect 7156 6604 7162 6616
rect 7193 6613 7205 6616
rect 7239 6613 7251 6647
rect 7193 6607 7251 6613
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7616 6616 7849 6644
rect 7616 6604 7622 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 10318 6644 10324 6656
rect 8812 6616 10324 6644
rect 8812 6604 8818 6616
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 1104 6554 10120 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 10120 6554
rect 1104 6480 10120 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1360 6412 1593 6440
rect 1360 6400 1366 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1728 6412 2145 6440
rect 1728 6400 1734 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 4062 6440 4068 6452
rect 2924 6412 4068 6440
rect 2924 6400 2930 6412
rect 4062 6400 4068 6412
rect 4120 6440 4126 6452
rect 4120 6412 6408 6440
rect 4120 6400 4126 6412
rect 5718 6372 5724 6384
rect 2056 6344 5724 6372
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 2056 6313 2084 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6304 2927 6307
rect 3510 6304 3516 6316
rect 2915 6276 3516 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 3510 6264 3516 6276
rect 3568 6304 3574 6316
rect 6380 6313 6408 6412
rect 7374 6400 7380 6452
rect 7432 6400 7438 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8573 6443 8631 6449
rect 7524 6412 8248 6440
rect 7524 6400 7530 6412
rect 8220 6372 8248 6412
rect 8573 6409 8585 6443
rect 8619 6440 8631 6443
rect 8846 6440 8852 6452
rect 8619 6412 8852 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 10502 6372 10508 6384
rect 7024 6344 7972 6372
rect 8220 6344 10508 6372
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 3568 6276 4353 6304
rect 3568 6264 3574 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6546 6304 6552 6316
rect 6411 6276 6552 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6304 6699 6307
rect 6730 6304 6736 6316
rect 6687 6276 6736 6304
rect 6687 6273 6699 6276
rect 6641 6267 6699 6273
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6205 3203 6239
rect 3145 6199 3203 6205
rect 1854 6060 1860 6112
rect 1912 6060 1918 6112
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 3160 6100 3188 6199
rect 4062 6196 4068 6248
rect 4120 6196 4126 6248
rect 6086 6168 6092 6180
rect 4724 6140 6092 6168
rect 4724 6100 4752 6140
rect 6086 6128 6092 6140
rect 6144 6128 6150 6180
rect 3108 6072 4752 6100
rect 3108 6060 3114 6072
rect 5074 6060 5080 6112
rect 5132 6060 5138 6112
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 7024 6100 7052 6344
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7800 6276 7849 6304
rect 7800 6264 7806 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7944 6304 7972 6344
rect 10502 6332 10508 6344
rect 10560 6332 10566 6384
rect 8846 6313 8852 6316
rect 8814 6307 8852 6313
rect 7944 6276 8156 6304
rect 7837 6267 7895 6273
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6205 7619 6239
rect 8128 6236 8156 6276
rect 8814 6273 8826 6307
rect 8814 6267 8852 6273
rect 8846 6264 8852 6267
rect 8904 6264 8910 6316
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 8128 6208 9505 6236
rect 7561 6199 7619 6205
rect 9493 6205 9505 6208
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 7576 6168 7604 6199
rect 9766 6196 9772 6248
rect 9824 6196 9830 6248
rect 7432 6140 7604 6168
rect 7432 6128 7438 6140
rect 8662 6128 8668 6180
rect 8720 6177 8726 6180
rect 8720 6171 8769 6177
rect 8720 6137 8723 6171
rect 8757 6137 8769 6171
rect 8720 6131 8769 6137
rect 8720 6128 8726 6131
rect 5500 6072 7052 6100
rect 5500 6060 5506 6072
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 10042 6100 10048 6112
rect 7892 6072 10048 6100
rect 7892 6060 7898 6072
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 1104 6010 10120 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 10120 6010
rect 1104 5936 10120 5958
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 3050 5896 3056 5908
rect 2648 5868 3056 5896
rect 2648 5856 2654 5868
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 5442 5896 5448 5908
rect 4212 5868 5448 5896
rect 4212 5856 4218 5868
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7561 5899 7619 5905
rect 6604 5868 7512 5896
rect 6604 5856 6610 5868
rect 2608 5769 2636 5856
rect 3605 5831 3663 5837
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 3651 5800 4384 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 4356 5769 4384 5800
rect 5718 5788 5724 5840
rect 5776 5788 5782 5840
rect 6454 5788 6460 5840
rect 6512 5788 6518 5840
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 6546 5720 6552 5772
rect 6604 5720 6610 5772
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 7484 5760 7512 5868
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 8386 5896 8392 5908
rect 7607 5868 8392 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 9582 5896 9588 5908
rect 8711 5868 9588 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7432 5732 7665 5760
rect 7432 5720 7438 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 9490 5720 9496 5772
rect 9548 5720 9554 5772
rect 2866 5652 2872 5704
rect 2924 5652 2930 5704
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4982 5692 4988 5704
rect 4304 5664 4988 5692
rect 4304 5652 4310 5664
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 5592 5664 6837 5692
rect 5592 5652 5598 5664
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 6825 5655 6883 5661
rect 6932 5664 7941 5692
rect 6273 5627 6331 5633
rect 6273 5593 6285 5627
rect 6319 5624 6331 5627
rect 6730 5624 6736 5636
rect 6319 5596 6736 5624
rect 6319 5593 6331 5596
rect 6273 5587 6331 5593
rect 6730 5584 6736 5596
rect 6788 5584 6794 5636
rect 3786 5516 3792 5568
rect 3844 5516 3850 5568
rect 5902 5516 5908 5568
rect 5960 5556 5966 5568
rect 6932 5556 6960 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 5960 5528 6960 5556
rect 5960 5516 5966 5528
rect 1104 5466 10120 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 10120 5466
rect 1104 5392 10120 5414
rect 3694 5312 3700 5364
rect 3752 5312 3758 5364
rect 4522 5312 4528 5364
rect 4580 5312 4586 5364
rect 8478 5312 8484 5364
rect 8536 5312 8542 5364
rect 9309 5355 9367 5361
rect 9309 5321 9321 5355
rect 9355 5352 9367 5355
rect 9398 5352 9404 5364
rect 9355 5324 9404 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 4433 5287 4491 5293
rect 4433 5284 4445 5287
rect 2924 5256 4445 5284
rect 2924 5244 2930 5256
rect 4433 5253 4445 5256
rect 4479 5284 4491 5287
rect 7282 5284 7288 5296
rect 4479 5256 7288 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 7282 5244 7288 5256
rect 7340 5284 7346 5296
rect 7340 5256 7788 5284
rect 7340 5244 7346 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 2774 5216 2780 5228
rect 1719 5188 2780 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3786 5216 3792 5228
rect 3559 5188 3792 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 5902 5216 5908 5228
rect 5859 5188 5908 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 6086 5176 6092 5228
rect 6144 5176 6150 5228
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7760 5225 7788 5256
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7432 5188 7481 5216
rect 7432 5176 7438 5188
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9674 5216 9680 5228
rect 9539 5188 9680 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 10686 5216 10692 5228
rect 9815 5188 10692 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 4338 5040 4344 5092
rect 4396 5080 4402 5092
rect 5077 5083 5135 5089
rect 5077 5080 5089 5083
rect 4396 5052 5089 5080
rect 4396 5040 4402 5052
rect 5077 5049 5089 5052
rect 5123 5049 5135 5083
rect 5077 5043 5135 5049
rect 1486 4972 1492 5024
rect 1544 4972 1550 5024
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 3476 4984 9597 5012
rect 3476 4972 3482 4984
rect 9585 4981 9597 4984
rect 9631 4981 9643 5015
rect 9585 4975 9643 4981
rect 1104 4922 10120 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 10120 4922
rect 1104 4848 10120 4870
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 4246 4740 4252 4752
rect 1719 4712 4252 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 4246 4700 4252 4712
rect 4304 4700 4310 4752
rect 1026 4632 1032 4684
rect 1084 4672 1090 4684
rect 5721 4675 5779 4681
rect 5721 4672 5733 4675
rect 1084 4644 5733 4672
rect 1084 4632 1090 4644
rect 5721 4641 5733 4644
rect 5767 4641 5779 4675
rect 5721 4635 5779 4641
rect 5537 4607 5595 4613
rect 5537 4573 5549 4607
rect 5583 4604 5595 4607
rect 5902 4604 5908 4616
rect 5583 4576 5908 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 1486 4496 1492 4548
rect 1544 4496 1550 4548
rect 1104 4378 10120 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 10120 4378
rect 1104 4304 10120 4326
rect 750 4224 756 4276
rect 808 4264 814 4276
rect 4154 4264 4160 4276
rect 808 4236 4160 4264
rect 808 4224 814 4236
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 1118 4156 1124 4208
rect 1176 4196 1182 4208
rect 1854 4196 1860 4208
rect 1176 4168 1860 4196
rect 1176 4156 1182 4168
rect 1854 4156 1860 4168
rect 1912 4156 1918 4208
rect 1104 3834 10120 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 10120 3834
rect 1104 3760 10120 3782
rect 1104 3290 10120 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 10120 3290
rect 1104 3216 10120 3238
rect 1104 2746 10120 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 10120 2746
rect 1104 2672 10120 2694
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 3602 2632 3608 2644
rect 2639 2604 3608 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 5534 2632 5540 2644
rect 3936 2604 5540 2632
rect 3936 2592 3942 2604
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 658 2524 664 2576
rect 716 2564 722 2576
rect 2774 2564 2780 2576
rect 716 2536 2780 2564
rect 716 2524 722 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2372 2400 2421 2428
rect 2372 2388 2378 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 1104 2202 10120 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 10120 2202
rect 1104 2128 10120 2150
rect 2682 2048 2688 2100
rect 2740 2088 2746 2100
rect 3234 2088 3240 2100
rect 2740 2060 3240 2088
rect 2740 2048 2746 2060
rect 3234 2048 3240 2060
rect 3292 2048 3298 2100
<< via1 >>
rect 7840 43460 7892 43512
rect 8392 43460 8444 43512
rect 940 43256 992 43308
rect 1400 43256 1452 43308
rect 6736 42508 6788 42560
rect 9220 42508 9272 42560
rect 3010 42406 3062 42458
rect 3074 42406 3126 42458
rect 3138 42406 3190 42458
rect 3202 42406 3254 42458
rect 3266 42406 3318 42458
rect 9010 42406 9062 42458
rect 9074 42406 9126 42458
rect 9138 42406 9190 42458
rect 9202 42406 9254 42458
rect 9266 42406 9318 42458
rect 1492 42304 1544 42356
rect 1860 42304 1912 42356
rect 2320 42304 2372 42356
rect 2780 42304 2832 42356
rect 3424 42347 3476 42356
rect 3424 42313 3433 42347
rect 3433 42313 3467 42347
rect 3467 42313 3476 42347
rect 3424 42304 3476 42313
rect 3700 42304 3752 42356
rect 4160 42304 4212 42356
rect 4620 42304 4672 42356
rect 5080 42304 5132 42356
rect 5540 42304 5592 42356
rect 6000 42347 6052 42356
rect 6000 42313 6009 42347
rect 6009 42313 6043 42347
rect 6043 42313 6052 42347
rect 6000 42304 6052 42313
rect 6460 42304 6512 42356
rect 6920 42304 6972 42356
rect 7380 42304 7432 42356
rect 8392 42347 8444 42356
rect 8392 42313 8401 42347
rect 8401 42313 8435 42347
rect 8435 42313 8444 42347
rect 8392 42304 8444 42313
rect 8760 42304 8812 42356
rect 1124 42168 1176 42220
rect 2320 42168 2372 42220
rect 3976 42236 4028 42288
rect 7196 42236 7248 42288
rect 8484 42236 8536 42288
rect 2412 42032 2464 42084
rect 4988 42211 5040 42220
rect 4988 42177 4997 42211
rect 4997 42177 5031 42211
rect 5031 42177 5040 42211
rect 4988 42168 5040 42177
rect 5448 42211 5500 42220
rect 5448 42177 5457 42211
rect 5457 42177 5491 42211
rect 5491 42177 5500 42211
rect 5448 42168 5500 42177
rect 6184 42211 6236 42220
rect 6184 42177 6193 42211
rect 6193 42177 6227 42211
rect 6227 42177 6236 42211
rect 6184 42168 6236 42177
rect 6552 42211 6604 42220
rect 6552 42177 6561 42211
rect 6561 42177 6595 42211
rect 6595 42177 6604 42211
rect 6552 42168 6604 42177
rect 7472 42211 7524 42220
rect 7472 42177 7481 42211
rect 7481 42177 7515 42211
rect 7515 42177 7524 42211
rect 7472 42168 7524 42177
rect 7840 42211 7892 42220
rect 7840 42177 7849 42211
rect 7849 42177 7883 42211
rect 7883 42177 7892 42211
rect 7840 42168 7892 42177
rect 8576 42211 8628 42220
rect 8576 42177 8585 42211
rect 8585 42177 8619 42211
rect 8619 42177 8628 42211
rect 8576 42168 8628 42177
rect 8760 42100 8812 42152
rect 9496 42100 9548 42152
rect 7380 42032 7432 42084
rect 8300 42032 8352 42084
rect 6920 41964 6972 42016
rect 7012 42007 7064 42016
rect 7012 41973 7021 42007
rect 7021 41973 7055 42007
rect 7055 41973 7064 42007
rect 7012 41964 7064 41973
rect 7288 41964 7340 42016
rect 7748 41964 7800 42016
rect 1950 41862 2002 41914
rect 2014 41862 2066 41914
rect 2078 41862 2130 41914
rect 2142 41862 2194 41914
rect 2206 41862 2258 41914
rect 7950 41862 8002 41914
rect 8014 41862 8066 41914
rect 8078 41862 8130 41914
rect 8142 41862 8194 41914
rect 8206 41862 8258 41914
rect 1400 41803 1452 41812
rect 1400 41769 1409 41803
rect 1409 41769 1443 41803
rect 1443 41769 1452 41803
rect 1400 41760 1452 41769
rect 6552 41803 6604 41812
rect 6552 41769 6561 41803
rect 6561 41769 6595 41803
rect 6595 41769 6604 41803
rect 6552 41760 6604 41769
rect 6736 41803 6788 41812
rect 6736 41769 6745 41803
rect 6745 41769 6779 41803
rect 6779 41769 6788 41803
rect 6736 41760 6788 41769
rect 7472 41803 7524 41812
rect 7472 41769 7481 41803
rect 7481 41769 7515 41803
rect 7515 41769 7524 41803
rect 7472 41760 7524 41769
rect 7840 41760 7892 41812
rect 10140 41760 10192 41812
rect 5448 41692 5500 41744
rect 6000 41624 6052 41676
rect 5448 41556 5500 41608
rect 4988 41488 5040 41540
rect 8392 41624 8444 41676
rect 7012 41556 7064 41608
rect 8024 41599 8076 41608
rect 8024 41565 8033 41599
rect 8033 41565 8067 41599
rect 8067 41565 8076 41599
rect 8024 41556 8076 41565
rect 8116 41556 8168 41608
rect 8852 41556 8904 41608
rect 9404 41556 9456 41608
rect 9588 41556 9640 41608
rect 9680 41556 9732 41608
rect 3792 41420 3844 41472
rect 9680 41463 9732 41472
rect 9680 41429 9689 41463
rect 9689 41429 9723 41463
rect 9723 41429 9732 41463
rect 9680 41420 9732 41429
rect 3010 41318 3062 41370
rect 3074 41318 3126 41370
rect 3138 41318 3190 41370
rect 3202 41318 3254 41370
rect 3266 41318 3318 41370
rect 9010 41318 9062 41370
rect 9074 41318 9126 41370
rect 9138 41318 9190 41370
rect 9202 41318 9254 41370
rect 9266 41318 9318 41370
rect 6184 41216 6236 41268
rect 6920 41216 6972 41268
rect 7380 41259 7432 41268
rect 7380 41225 7389 41259
rect 7389 41225 7423 41259
rect 7423 41225 7432 41259
rect 7380 41216 7432 41225
rect 8024 41216 8076 41268
rect 8852 41216 8904 41268
rect 9404 41216 9456 41268
rect 9496 41259 9548 41268
rect 9496 41225 9505 41259
rect 9505 41225 9539 41259
rect 9539 41225 9548 41259
rect 9496 41216 9548 41225
rect 1492 41123 1544 41132
rect 1492 41089 1501 41123
rect 1501 41089 1535 41123
rect 1535 41089 1544 41123
rect 1492 41080 1544 41089
rect 6828 41080 6880 41132
rect 7012 41123 7064 41132
rect 7012 41089 7021 41123
rect 7021 41089 7055 41123
rect 7055 41089 7064 41123
rect 7012 41080 7064 41089
rect 848 41012 900 41064
rect 7748 41080 7800 41132
rect 7840 41080 7892 41132
rect 8300 41080 8352 41132
rect 9404 41123 9456 41132
rect 9404 41089 9413 41123
rect 9413 41089 9447 41123
rect 9447 41089 9456 41123
rect 9404 41080 9456 41089
rect 9772 41080 9824 41132
rect 1860 40944 1912 40996
rect 3884 40944 3936 40996
rect 8484 40944 8536 40996
rect 8576 40919 8628 40928
rect 8576 40885 8585 40919
rect 8585 40885 8619 40919
rect 8619 40885 8628 40919
rect 8576 40876 8628 40885
rect 10416 40876 10468 40928
rect 1950 40774 2002 40826
rect 2014 40774 2066 40826
rect 2078 40774 2130 40826
rect 2142 40774 2194 40826
rect 2206 40774 2258 40826
rect 7950 40774 8002 40826
rect 8014 40774 8066 40826
rect 8078 40774 8130 40826
rect 8142 40774 8194 40826
rect 8206 40774 8258 40826
rect 7196 40672 7248 40724
rect 8392 40672 8444 40724
rect 8668 40672 8720 40724
rect 7380 40468 7432 40520
rect 8668 40468 8720 40520
rect 9588 40468 9640 40520
rect 1492 40443 1544 40452
rect 1492 40409 1501 40443
rect 1501 40409 1535 40443
rect 1535 40409 1544 40443
rect 1492 40400 1544 40409
rect 1768 40400 1820 40452
rect 7472 40400 7524 40452
rect 7840 40400 7892 40452
rect 6828 40375 6880 40384
rect 6828 40341 6837 40375
rect 6837 40341 6871 40375
rect 6871 40341 6880 40375
rect 6828 40332 6880 40341
rect 7748 40375 7800 40384
rect 7748 40341 7757 40375
rect 7757 40341 7791 40375
rect 7791 40341 7800 40375
rect 7748 40332 7800 40341
rect 8300 40375 8352 40384
rect 8300 40341 8309 40375
rect 8309 40341 8343 40375
rect 8343 40341 8352 40375
rect 8300 40332 8352 40341
rect 9404 40332 9456 40384
rect 9772 40332 9824 40384
rect 3010 40230 3062 40282
rect 3074 40230 3126 40282
rect 3138 40230 3190 40282
rect 3202 40230 3254 40282
rect 3266 40230 3318 40282
rect 9010 40230 9062 40282
rect 9074 40230 9126 40282
rect 9138 40230 9190 40282
rect 9202 40230 9254 40282
rect 9266 40230 9318 40282
rect 4068 40128 4120 40180
rect 572 40060 624 40112
rect 9220 40060 9272 40112
rect 8760 39899 8812 39908
rect 8760 39865 8769 39899
rect 8769 39865 8803 39899
rect 8803 39865 8812 39899
rect 8760 39856 8812 39865
rect 10600 39856 10652 39908
rect 7380 39831 7432 39840
rect 7380 39797 7389 39831
rect 7389 39797 7423 39831
rect 7423 39797 7432 39831
rect 7380 39788 7432 39797
rect 8668 39831 8720 39840
rect 8668 39797 8677 39831
rect 8677 39797 8711 39831
rect 8711 39797 8720 39831
rect 8668 39788 8720 39797
rect 10784 39788 10836 39840
rect 1950 39686 2002 39738
rect 2014 39686 2066 39738
rect 2078 39686 2130 39738
rect 2142 39686 2194 39738
rect 2206 39686 2258 39738
rect 7950 39686 8002 39738
rect 8014 39686 8066 39738
rect 8078 39686 8130 39738
rect 8142 39686 8194 39738
rect 8206 39686 8258 39738
rect 10232 39516 10284 39568
rect 3700 39448 3752 39500
rect 3976 39448 4028 39500
rect 5172 39423 5224 39432
rect 5172 39389 5181 39423
rect 5181 39389 5215 39423
rect 5215 39389 5224 39423
rect 5172 39380 5224 39389
rect 5816 39380 5868 39432
rect 1492 39355 1544 39364
rect 1492 39321 1501 39355
rect 1501 39321 1535 39355
rect 1535 39321 1544 39355
rect 1492 39312 1544 39321
rect 2780 39312 2832 39364
rect 3976 39312 4028 39364
rect 9496 39423 9548 39432
rect 9496 39389 9505 39423
rect 9505 39389 9539 39423
rect 9539 39389 9548 39423
rect 9496 39380 9548 39389
rect 4436 39287 4488 39296
rect 4436 39253 4445 39287
rect 4445 39253 4479 39287
rect 4479 39253 4488 39287
rect 4436 39244 4488 39253
rect 10416 39244 10468 39296
rect 3010 39142 3062 39194
rect 3074 39142 3126 39194
rect 3138 39142 3190 39194
rect 3202 39142 3254 39194
rect 3266 39142 3318 39194
rect 9010 39142 9062 39194
rect 9074 39142 9126 39194
rect 9138 39142 9190 39194
rect 9202 39142 9254 39194
rect 9266 39142 9318 39194
rect 10324 39040 10376 39092
rect 756 38904 808 38956
rect 4344 38904 4396 38956
rect 5816 38972 5868 39024
rect 4988 38904 5040 38956
rect 5724 38947 5776 38956
rect 5724 38913 5733 38947
rect 5733 38913 5767 38947
rect 5767 38913 5776 38947
rect 5724 38904 5776 38913
rect 8760 38947 8812 38956
rect 8760 38913 8769 38947
rect 8769 38913 8803 38947
rect 8803 38913 8812 38947
rect 8760 38904 8812 38913
rect 9128 38947 9180 38956
rect 9128 38913 9137 38947
rect 9137 38913 9171 38947
rect 9171 38913 9180 38947
rect 9128 38904 9180 38913
rect 9496 38947 9548 38956
rect 9496 38913 9505 38947
rect 9505 38913 9539 38947
rect 9539 38913 9548 38947
rect 9496 38904 9548 38913
rect 2596 38768 2648 38820
rect 10140 38768 10192 38820
rect 5264 38700 5316 38752
rect 5356 38700 5408 38752
rect 6276 38700 6328 38752
rect 8852 38700 8904 38752
rect 10508 38700 10560 38752
rect 1950 38598 2002 38650
rect 2014 38598 2066 38650
rect 2078 38598 2130 38650
rect 2142 38598 2194 38650
rect 2206 38598 2258 38650
rect 7950 38598 8002 38650
rect 8014 38598 8066 38650
rect 8078 38598 8130 38650
rect 8142 38598 8194 38650
rect 8206 38598 8258 38650
rect 3424 38496 3476 38548
rect 4712 38496 4764 38548
rect 5724 38496 5776 38548
rect 4436 38428 4488 38480
rect 10048 38428 10100 38480
rect 2688 38360 2740 38412
rect 1584 38292 1636 38344
rect 1492 38267 1544 38276
rect 1492 38233 1501 38267
rect 1501 38233 1535 38267
rect 1535 38233 1544 38267
rect 1492 38224 1544 38233
rect 1860 38224 1912 38276
rect 2504 38292 2556 38344
rect 5356 38403 5408 38412
rect 5356 38369 5365 38403
rect 5365 38369 5399 38403
rect 5399 38369 5408 38403
rect 5356 38360 5408 38369
rect 6460 38403 6512 38412
rect 6460 38369 6469 38403
rect 6469 38369 6503 38403
rect 6503 38369 6512 38403
rect 6460 38360 6512 38369
rect 3424 38224 3476 38276
rect 3516 38224 3568 38276
rect 5080 38335 5132 38344
rect 5080 38301 5089 38335
rect 5089 38301 5123 38335
rect 5123 38301 5132 38335
rect 5080 38292 5132 38301
rect 6184 38335 6236 38344
rect 6184 38301 6193 38335
rect 6193 38301 6227 38335
rect 6227 38301 6236 38335
rect 6184 38292 6236 38301
rect 8484 38335 8536 38344
rect 8484 38301 8493 38335
rect 8493 38301 8527 38335
rect 8527 38301 8536 38335
rect 8484 38292 8536 38301
rect 9128 38335 9180 38344
rect 9128 38301 9137 38335
rect 9137 38301 9171 38335
rect 9171 38301 9180 38335
rect 9128 38292 9180 38301
rect 2872 38156 2924 38208
rect 4160 38156 4212 38208
rect 6644 38156 6696 38208
rect 7840 38156 7892 38208
rect 9956 38224 10008 38276
rect 10968 38156 11020 38208
rect 3010 38054 3062 38106
rect 3074 38054 3126 38106
rect 3138 38054 3190 38106
rect 3202 38054 3254 38106
rect 3266 38054 3318 38106
rect 9010 38054 9062 38106
rect 9074 38054 9126 38106
rect 9138 38054 9190 38106
rect 9202 38054 9254 38106
rect 9266 38054 9318 38106
rect 480 37952 532 38004
rect 3976 37952 4028 38004
rect 4344 37995 4396 38004
rect 4344 37961 4353 37995
rect 4353 37961 4387 37995
rect 4387 37961 4396 37995
rect 4344 37952 4396 37961
rect 1584 37816 1636 37868
rect 1768 37816 1820 37868
rect 4620 37816 4672 37868
rect 5172 37952 5224 38004
rect 6184 37952 6236 38004
rect 10140 37952 10192 38004
rect 5908 37884 5960 37936
rect 5632 37859 5684 37868
rect 5632 37825 5641 37859
rect 5641 37825 5675 37859
rect 5675 37825 5684 37859
rect 5632 37816 5684 37825
rect 6368 37859 6420 37868
rect 6368 37825 6377 37859
rect 6377 37825 6411 37859
rect 6411 37825 6420 37859
rect 6368 37816 6420 37825
rect 8668 37859 8720 37868
rect 8668 37825 8677 37859
rect 8677 37825 8711 37859
rect 8711 37825 8720 37859
rect 8668 37816 8720 37825
rect 8760 37859 8812 37868
rect 8760 37825 8769 37859
rect 8769 37825 8803 37859
rect 8803 37825 8812 37859
rect 8760 37816 8812 37825
rect 2504 37791 2556 37800
rect 2504 37757 2513 37791
rect 2513 37757 2547 37791
rect 2547 37757 2556 37791
rect 2504 37748 2556 37757
rect 2688 37791 2740 37800
rect 2688 37757 2697 37791
rect 2697 37757 2731 37791
rect 2731 37757 2740 37791
rect 2688 37748 2740 37757
rect 2872 37748 2924 37800
rect 3424 37791 3476 37800
rect 3424 37757 3433 37791
rect 3433 37757 3467 37791
rect 3467 37757 3476 37791
rect 3424 37748 3476 37757
rect 3516 37791 3568 37800
rect 3516 37757 3550 37791
rect 3550 37757 3568 37791
rect 3516 37748 3568 37757
rect 4252 37748 4304 37800
rect 7012 37748 7064 37800
rect 5816 37723 5868 37732
rect 5816 37689 5825 37723
rect 5825 37689 5859 37723
rect 5859 37689 5868 37723
rect 5816 37680 5868 37689
rect 10232 37680 10284 37732
rect 4896 37612 4948 37664
rect 6920 37612 6972 37664
rect 8484 37655 8536 37664
rect 8484 37621 8493 37655
rect 8493 37621 8527 37655
rect 8527 37621 8536 37655
rect 8484 37612 8536 37621
rect 10600 37612 10652 37664
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 7950 37510 8002 37562
rect 8014 37510 8066 37562
rect 8078 37510 8130 37562
rect 8142 37510 8194 37562
rect 8206 37510 8258 37562
rect 204 37408 256 37460
rect 5632 37408 5684 37460
rect 6368 37408 6420 37460
rect 6092 37340 6144 37392
rect 7472 37340 7524 37392
rect 5264 37272 5316 37324
rect 7380 37272 7432 37324
rect 7564 37315 7616 37324
rect 7564 37281 7573 37315
rect 7573 37281 7607 37315
rect 7607 37281 7616 37315
rect 7564 37272 7616 37281
rect 1676 37247 1728 37256
rect 1676 37213 1685 37247
rect 1685 37213 1719 37247
rect 1719 37213 1728 37247
rect 1676 37204 1728 37213
rect 1492 37179 1544 37188
rect 1492 37145 1501 37179
rect 1501 37145 1535 37179
rect 1535 37145 1544 37179
rect 1492 37136 1544 37145
rect 1584 37136 1636 37188
rect 1860 37204 1912 37256
rect 2044 37136 2096 37188
rect 4252 37247 4304 37256
rect 4252 37213 4261 37247
rect 4261 37213 4295 37247
rect 4295 37213 4304 37247
rect 4252 37204 4304 37213
rect 4528 37247 4580 37256
rect 4528 37213 4537 37247
rect 4537 37213 4571 37247
rect 4571 37213 4580 37247
rect 4528 37204 4580 37213
rect 4988 37204 5040 37256
rect 2228 37068 2280 37120
rect 4068 37136 4120 37188
rect 3884 37068 3936 37120
rect 5632 37136 5684 37188
rect 5724 37179 5776 37188
rect 5724 37145 5733 37179
rect 5733 37145 5767 37179
rect 5767 37145 5776 37179
rect 5724 37136 5776 37145
rect 6552 37136 6604 37188
rect 9404 37204 9456 37256
rect 8392 37068 8444 37120
rect 10324 37136 10376 37188
rect 9680 37111 9732 37120
rect 9680 37077 9689 37111
rect 9689 37077 9723 37111
rect 9723 37077 9732 37111
rect 9680 37068 9732 37077
rect 3010 36966 3062 37018
rect 3074 36966 3126 37018
rect 3138 36966 3190 37018
rect 3202 36966 3254 37018
rect 3266 36966 3318 37018
rect 9010 36966 9062 37018
rect 9074 36966 9126 37018
rect 9138 36966 9190 37018
rect 9202 36966 9254 37018
rect 9266 36966 9318 37018
rect 1584 36864 1636 36916
rect 4252 36864 4304 36916
rect 5540 36864 5592 36916
rect 8668 36864 8720 36916
rect 1768 36796 1820 36848
rect 3608 36796 3660 36848
rect 4344 36728 4396 36780
rect 4528 36771 4580 36780
rect 4528 36737 4562 36771
rect 4562 36737 4580 36771
rect 4528 36728 4580 36737
rect 1676 36660 1728 36712
rect 3700 36660 3752 36712
rect 3884 36660 3936 36712
rect 4252 36703 4304 36712
rect 4252 36669 4261 36703
rect 4261 36669 4295 36703
rect 4295 36669 4304 36703
rect 4252 36660 4304 36669
rect 3424 36592 3476 36644
rect 1584 36524 1636 36576
rect 2044 36524 2096 36576
rect 3700 36524 3752 36576
rect 4068 36524 4120 36576
rect 6920 36728 6972 36780
rect 7840 36771 7892 36780
rect 7840 36737 7849 36771
rect 7849 36737 7883 36771
rect 7883 36737 7892 36771
rect 7840 36728 7892 36737
rect 9312 36796 9364 36848
rect 9128 36771 9180 36780
rect 9128 36737 9137 36771
rect 9137 36737 9171 36771
rect 9171 36737 9180 36771
rect 9128 36728 9180 36737
rect 7656 36660 7708 36712
rect 8116 36703 8168 36712
rect 8116 36669 8125 36703
rect 8125 36669 8159 36703
rect 8159 36669 8168 36703
rect 8116 36660 8168 36669
rect 8392 36703 8444 36712
rect 8392 36669 8401 36703
rect 8401 36669 8435 36703
rect 8435 36669 8444 36703
rect 8392 36660 8444 36669
rect 8760 36660 8812 36712
rect 10508 36592 10560 36644
rect 10416 36524 10468 36576
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 7950 36422 8002 36474
rect 8014 36422 8066 36474
rect 8078 36422 8130 36474
rect 8142 36422 8194 36474
rect 8206 36422 8258 36474
rect 4252 36363 4304 36372
rect 4252 36329 4261 36363
rect 4261 36329 4295 36363
rect 4295 36329 4304 36363
rect 4252 36320 4304 36329
rect 4068 36252 4120 36304
rect 6736 36252 6788 36304
rect 1216 36184 1268 36236
rect 1492 36184 1544 36236
rect 1676 36184 1728 36236
rect 4436 36184 4488 36236
rect 6000 36184 6052 36236
rect 1124 36116 1176 36168
rect 2320 36159 2372 36168
rect 2320 36125 2329 36159
rect 2329 36125 2363 36159
rect 2363 36125 2372 36159
rect 2320 36116 2372 36125
rect 9404 36320 9456 36372
rect 9496 36252 9548 36304
rect 10232 36252 10284 36304
rect 8300 36184 8352 36236
rect 10876 36184 10928 36236
rect 1492 36091 1544 36100
rect 1492 36057 1501 36091
rect 1501 36057 1535 36091
rect 1535 36057 1544 36091
rect 1492 36048 1544 36057
rect 1676 36091 1728 36100
rect 1676 36057 1685 36091
rect 1685 36057 1719 36091
rect 1719 36057 1728 36091
rect 1676 36048 1728 36057
rect 296 35980 348 36032
rect 7104 36116 7156 36168
rect 7748 36116 7800 36168
rect 8852 36116 8904 36168
rect 2872 35980 2924 36032
rect 5632 36048 5684 36100
rect 6184 36048 6236 36100
rect 7472 36091 7524 36100
rect 7472 36057 7481 36091
rect 7481 36057 7515 36091
rect 7515 36057 7524 36091
rect 7472 36048 7524 36057
rect 8852 35980 8904 36032
rect 9588 35980 9640 36032
rect 10140 35980 10192 36032
rect 3010 35878 3062 35930
rect 3074 35878 3126 35930
rect 3138 35878 3190 35930
rect 3202 35878 3254 35930
rect 3266 35878 3318 35930
rect 9010 35878 9062 35930
rect 9074 35878 9126 35930
rect 9138 35878 9190 35930
rect 9202 35878 9254 35930
rect 9266 35878 9318 35930
rect 4160 35776 4212 35828
rect 4344 35819 4396 35828
rect 4344 35785 4353 35819
rect 4353 35785 4387 35819
rect 4387 35785 4396 35819
rect 4344 35776 4396 35785
rect 7012 35776 7064 35828
rect 8392 35776 8444 35828
rect 7748 35708 7800 35760
rect 1492 35683 1544 35692
rect 1492 35649 1501 35683
rect 1501 35649 1535 35683
rect 1535 35649 1544 35683
rect 1492 35640 1544 35649
rect 1768 35683 1820 35692
rect 1768 35649 1777 35683
rect 1777 35649 1811 35683
rect 1811 35649 1820 35683
rect 1768 35640 1820 35649
rect 2320 35640 2372 35692
rect 2504 35683 2556 35692
rect 2504 35649 2513 35683
rect 2513 35649 2547 35683
rect 2547 35649 2556 35683
rect 2504 35640 2556 35649
rect 3700 35683 3752 35692
rect 3700 35649 3709 35683
rect 3709 35649 3743 35683
rect 3743 35649 3752 35683
rect 3700 35640 3752 35649
rect 6920 35640 6972 35692
rect 8300 35683 8352 35692
rect 8300 35649 8309 35683
rect 8309 35649 8343 35683
rect 8343 35649 8352 35683
rect 8300 35640 8352 35649
rect 8576 35683 8628 35692
rect 8576 35649 8585 35683
rect 8585 35649 8619 35683
rect 8619 35649 8628 35683
rect 8576 35640 8628 35649
rect 2688 35615 2740 35624
rect 2688 35581 2697 35615
rect 2697 35581 2731 35615
rect 2731 35581 2740 35615
rect 2688 35572 2740 35581
rect 2780 35572 2832 35624
rect 2872 35572 2924 35624
rect 3424 35615 3476 35624
rect 3424 35581 3433 35615
rect 3433 35581 3467 35615
rect 3467 35581 3476 35615
rect 3424 35572 3476 35581
rect 3516 35572 3568 35624
rect 3884 35572 3936 35624
rect 8484 35615 8536 35624
rect 8484 35581 8502 35615
rect 8502 35581 8536 35615
rect 8484 35572 8536 35581
rect 8852 35615 8904 35624
rect 8852 35581 8861 35615
rect 8861 35581 8895 35615
rect 8895 35581 8904 35615
rect 8852 35572 8904 35581
rect 9312 35615 9364 35624
rect 9312 35581 9321 35615
rect 9321 35581 9355 35615
rect 9355 35581 9364 35615
rect 9312 35572 9364 35581
rect 9404 35572 9456 35624
rect 3240 35504 3292 35556
rect 5080 35504 5132 35556
rect 7012 35504 7064 35556
rect 7472 35504 7524 35556
rect 7840 35504 7892 35556
rect 5908 35436 5960 35488
rect 8208 35436 8260 35488
rect 8484 35436 8536 35488
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 7950 35334 8002 35386
rect 8014 35334 8066 35386
rect 8078 35334 8130 35386
rect 8142 35334 8194 35386
rect 8206 35334 8258 35386
rect 2412 35232 2464 35284
rect 6460 35232 6512 35284
rect 6736 35164 6788 35216
rect 7196 35164 7248 35216
rect 8300 35232 8352 35284
rect 9312 35232 9364 35284
rect 9956 35164 10008 35216
rect 1124 35096 1176 35148
rect 1676 35096 1728 35148
rect 4528 35096 4580 35148
rect 5356 35071 5408 35080
rect 5356 35037 5365 35071
rect 5365 35037 5399 35071
rect 5399 35037 5408 35071
rect 5356 35028 5408 35037
rect 1952 34960 2004 35012
rect 6736 35028 6788 35080
rect 7104 35028 7156 35080
rect 7564 35028 7616 35080
rect 5816 34960 5868 35012
rect 6092 34960 6144 35012
rect 6644 34960 6696 35012
rect 8944 35071 8996 35080
rect 8944 35037 8953 35071
rect 8953 35037 8987 35071
rect 8987 35037 8996 35071
rect 8944 35028 8996 35037
rect 4436 34892 4488 34944
rect 4804 34892 4856 34944
rect 6920 34892 6972 34944
rect 7472 34892 7524 34944
rect 7564 34892 7616 34944
rect 10232 34960 10284 35012
rect 10600 34892 10652 34944
rect 3010 34790 3062 34842
rect 3074 34790 3126 34842
rect 3138 34790 3190 34842
rect 3202 34790 3254 34842
rect 3266 34790 3318 34842
rect 9010 34790 9062 34842
rect 9074 34790 9126 34842
rect 9138 34790 9190 34842
rect 9202 34790 9254 34842
rect 9266 34790 9318 34842
rect 1032 34688 1084 34740
rect 5172 34731 5224 34740
rect 5172 34697 5181 34731
rect 5181 34697 5215 34731
rect 5215 34697 5224 34731
rect 5172 34688 5224 34697
rect 6552 34731 6604 34740
rect 6552 34697 6561 34731
rect 6561 34697 6595 34731
rect 6595 34697 6604 34731
rect 6552 34688 6604 34697
rect 7748 34688 7800 34740
rect 8668 34688 8720 34740
rect 940 34620 992 34672
rect 5448 34620 5500 34672
rect 6276 34620 6328 34672
rect 6920 34620 6972 34672
rect 7840 34620 7892 34672
rect 388 34552 440 34604
rect 2780 34552 2832 34604
rect 4804 34595 4856 34604
rect 4804 34561 4813 34595
rect 4813 34561 4847 34595
rect 4847 34561 4856 34595
rect 4804 34552 4856 34561
rect 5356 34552 5408 34604
rect 6644 34552 6696 34604
rect 1768 34416 1820 34468
rect 1952 34416 2004 34468
rect 5448 34484 5500 34536
rect 6276 34484 6328 34536
rect 6920 34527 6972 34536
rect 6920 34493 6929 34527
rect 6929 34493 6963 34527
rect 6963 34493 6972 34527
rect 6920 34484 6972 34493
rect 1308 34348 1360 34400
rect 3976 34391 4028 34400
rect 3976 34357 3985 34391
rect 3985 34357 4019 34391
rect 4019 34357 4028 34391
rect 3976 34348 4028 34357
rect 4068 34391 4120 34400
rect 4068 34357 4077 34391
rect 4077 34357 4111 34391
rect 4111 34357 4120 34391
rect 4068 34348 4120 34357
rect 4712 34348 4764 34400
rect 6092 34348 6144 34400
rect 6736 34348 6788 34400
rect 7840 34348 7892 34400
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 7950 34246 8002 34298
rect 8014 34246 8066 34298
rect 8078 34246 8130 34298
rect 8142 34246 8194 34298
rect 8206 34246 8258 34298
rect 20 34144 72 34196
rect 3424 34144 3476 34196
rect 6736 34144 6788 34196
rect 9404 34144 9456 34196
rect 1124 34076 1176 34128
rect 3976 34076 4028 34128
rect 4436 34119 4488 34128
rect 4436 34085 4445 34119
rect 4445 34085 4479 34119
rect 4479 34085 4488 34119
rect 4436 34076 4488 34085
rect 6828 34076 6880 34128
rect 9956 34076 10008 34128
rect 2320 33940 2372 33992
rect 2412 33940 2464 33992
rect 3516 33940 3568 33992
rect 3976 33983 4028 33992
rect 3976 33949 3985 33983
rect 3985 33949 4019 33983
rect 4019 33949 4028 33983
rect 3976 33940 4028 33949
rect 4712 33983 4764 33992
rect 4712 33949 4721 33983
rect 4721 33949 4755 33983
rect 4755 33949 4764 33983
rect 4712 33940 4764 33949
rect 4804 33983 4856 33992
rect 4804 33949 4838 33983
rect 4838 33949 4856 33983
rect 4804 33940 4856 33949
rect 6644 33940 6696 33992
rect 7656 33940 7708 33992
rect 10784 34008 10836 34060
rect 8208 33983 8260 33992
rect 8208 33949 8217 33983
rect 8217 33949 8251 33983
rect 8251 33949 8260 33983
rect 8208 33940 8260 33949
rect 8300 33940 8352 33992
rect 9128 33983 9180 33992
rect 9128 33949 9137 33983
rect 9137 33949 9171 33983
rect 9171 33949 9180 33983
rect 9128 33940 9180 33949
rect 9496 33983 9548 33992
rect 9496 33949 9505 33983
rect 9505 33949 9539 33983
rect 9539 33949 9548 33983
rect 9496 33940 9548 33949
rect 1768 33804 1820 33856
rect 3516 33804 3568 33856
rect 3700 33804 3752 33856
rect 8760 33872 8812 33924
rect 8668 33804 8720 33856
rect 10692 33872 10744 33924
rect 9680 33847 9732 33856
rect 9680 33813 9689 33847
rect 9689 33813 9723 33847
rect 9723 33813 9732 33847
rect 9680 33804 9732 33813
rect 3010 33702 3062 33754
rect 3074 33702 3126 33754
rect 3138 33702 3190 33754
rect 3202 33702 3254 33754
rect 3266 33702 3318 33754
rect 9010 33702 9062 33754
rect 9074 33702 9126 33754
rect 9138 33702 9190 33754
rect 9202 33702 9254 33754
rect 9266 33702 9318 33754
rect 6920 33600 6972 33652
rect 8208 33600 8260 33652
rect 1216 33532 1268 33584
rect 756 33464 808 33516
rect 2412 33575 2464 33584
rect 2412 33541 2421 33575
rect 2421 33541 2455 33575
rect 2455 33541 2464 33575
rect 2412 33532 2464 33541
rect 8760 33507 8812 33516
rect 8760 33473 8769 33507
rect 8769 33473 8803 33507
rect 8803 33473 8812 33507
rect 8760 33464 8812 33473
rect 1584 33396 1636 33448
rect 2412 33396 2464 33448
rect 3056 33439 3108 33448
rect 3056 33405 3065 33439
rect 3065 33405 3099 33439
rect 3099 33405 3108 33439
rect 3056 33396 3108 33405
rect 3240 33439 3292 33448
rect 3240 33405 3258 33439
rect 3258 33405 3292 33439
rect 3240 33396 3292 33405
rect 3332 33439 3384 33448
rect 3332 33405 3341 33439
rect 3341 33405 3375 33439
rect 3375 33405 3384 33439
rect 3332 33396 3384 33405
rect 3516 33396 3568 33448
rect 4160 33396 4212 33448
rect 4252 33439 4304 33448
rect 4252 33405 4261 33439
rect 4261 33405 4295 33439
rect 4295 33405 4304 33439
rect 4252 33396 4304 33405
rect 4804 33396 4856 33448
rect 7288 33396 7340 33448
rect 7748 33439 7800 33448
rect 7748 33405 7757 33439
rect 7757 33405 7791 33439
rect 7791 33405 7800 33439
rect 7748 33396 7800 33405
rect 7840 33396 7892 33448
rect 1124 33328 1176 33380
rect 1676 33328 1728 33380
rect 6552 33328 6604 33380
rect 7472 33328 7524 33380
rect 9956 33396 10008 33448
rect 2964 33260 3016 33312
rect 3792 33260 3844 33312
rect 4160 33260 4212 33312
rect 9496 33371 9548 33380
rect 9496 33337 9505 33371
rect 9505 33337 9539 33371
rect 9539 33337 9548 33371
rect 9496 33328 9548 33337
rect 10048 33260 10100 33312
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 7950 33158 8002 33210
rect 8014 33158 8066 33210
rect 8078 33158 8130 33210
rect 8142 33158 8194 33210
rect 8206 33158 8258 33210
rect 3056 33056 3108 33108
rect 3240 33056 3292 33108
rect 3976 33056 4028 33108
rect 4436 33056 4488 33108
rect 3608 32988 3660 33040
rect 3792 32988 3844 33040
rect 4344 32988 4396 33040
rect 7104 33056 7156 33108
rect 7472 33056 7524 33108
rect 1308 32920 1360 32972
rect 1584 32920 1636 32972
rect 2964 32920 3016 32972
rect 4804 32920 4856 32972
rect 6552 32920 6604 32972
rect 7656 32920 7708 32972
rect 10232 32988 10284 33040
rect 1676 32895 1728 32904
rect 1676 32861 1685 32895
rect 1685 32861 1719 32895
rect 1719 32861 1728 32895
rect 1676 32852 1728 32861
rect 1952 32895 2004 32904
rect 1952 32861 1961 32895
rect 1961 32861 1995 32895
rect 1995 32861 2004 32895
rect 1952 32852 2004 32861
rect 6736 32852 6788 32904
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 8116 32895 8168 32904
rect 8116 32861 8125 32895
rect 8125 32861 8159 32895
rect 8159 32861 8168 32895
rect 8116 32852 8168 32861
rect 6276 32784 6328 32836
rect 8852 32852 8904 32904
rect 11152 32784 11204 32836
rect 664 32716 716 32768
rect 2780 32716 2832 32768
rect 8208 32716 8260 32768
rect 8852 32716 8904 32768
rect 10416 32716 10468 32768
rect 3010 32614 3062 32666
rect 3074 32614 3126 32666
rect 3138 32614 3190 32666
rect 3202 32614 3254 32666
rect 3266 32614 3318 32666
rect 9010 32614 9062 32666
rect 9074 32614 9126 32666
rect 9138 32614 9190 32666
rect 9202 32614 9254 32666
rect 9266 32614 9318 32666
rect 1676 32512 1728 32564
rect 1952 32512 2004 32564
rect 2872 32512 2924 32564
rect 3424 32512 3476 32564
rect 3608 32512 3660 32564
rect 8116 32512 8168 32564
rect 8392 32444 8444 32496
rect 9864 32512 9916 32564
rect 1492 32419 1544 32428
rect 1492 32385 1501 32419
rect 1501 32385 1535 32419
rect 1535 32385 1544 32419
rect 1492 32376 1544 32385
rect 1768 32240 1820 32292
rect 4344 32376 4396 32428
rect 3240 32308 3292 32360
rect 6552 32419 6604 32428
rect 6552 32385 6561 32419
rect 6561 32385 6595 32419
rect 6595 32385 6604 32419
rect 6552 32376 6604 32385
rect 8208 32419 8260 32428
rect 8208 32385 8217 32419
rect 8217 32385 8251 32419
rect 8251 32385 8260 32419
rect 8208 32376 8260 32385
rect 4804 32240 4856 32292
rect 6828 32351 6880 32360
rect 6828 32317 6837 32351
rect 6837 32317 6871 32351
rect 6871 32317 6880 32351
rect 6828 32308 6880 32317
rect 8392 32308 8444 32360
rect 8944 32376 8996 32428
rect 8852 32240 8904 32292
rect 10232 32240 10284 32292
rect 1216 32172 1268 32224
rect 2780 32172 2832 32224
rect 3884 32172 3936 32224
rect 4712 32172 4764 32224
rect 6092 32172 6144 32224
rect 8300 32172 8352 32224
rect 9220 32172 9272 32224
rect 9404 32172 9456 32224
rect 9680 32215 9732 32224
rect 9680 32181 9689 32215
rect 9689 32181 9723 32215
rect 9723 32181 9732 32215
rect 9680 32172 9732 32181
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 7950 32070 8002 32122
rect 8014 32070 8066 32122
rect 8078 32070 8130 32122
rect 8142 32070 8194 32122
rect 8206 32070 8258 32122
rect 1768 32011 1820 32020
rect 1768 31977 1777 32011
rect 1777 31977 1811 32011
rect 1811 31977 1820 32011
rect 1768 31968 1820 31977
rect 2504 31968 2556 32020
rect 4344 32011 4396 32020
rect 4344 31977 4353 32011
rect 4353 31977 4387 32011
rect 4387 31977 4396 32011
rect 4344 31968 4396 31977
rect 5632 31968 5684 32020
rect 940 31832 992 31884
rect 2228 31832 2280 31884
rect 3884 31900 3936 31952
rect 5540 31943 5592 31952
rect 5540 31909 5549 31943
rect 5549 31909 5583 31943
rect 5583 31909 5592 31943
rect 5540 31900 5592 31909
rect 9220 31968 9272 32020
rect 10232 31968 10284 32020
rect 9128 31900 9180 31952
rect 9496 31900 9548 31952
rect 9588 31900 9640 31952
rect 3056 31832 3108 31884
rect 4436 31832 4488 31884
rect 4988 31875 5040 31884
rect 4988 31841 4997 31875
rect 4997 31841 5031 31875
rect 5031 31841 5040 31875
rect 4988 31832 5040 31841
rect 5816 31832 5868 31884
rect 6828 31832 6880 31884
rect 848 31764 900 31816
rect 2412 31807 2464 31816
rect 2412 31773 2421 31807
rect 2421 31773 2455 31807
rect 2455 31773 2464 31807
rect 2412 31764 2464 31773
rect 3516 31764 3568 31816
rect 3884 31764 3936 31816
rect 5080 31764 5132 31816
rect 5264 31807 5316 31816
rect 5264 31773 5273 31807
rect 5273 31773 5307 31807
rect 5307 31773 5316 31807
rect 5264 31764 5316 31773
rect 6000 31807 6052 31816
rect 6000 31773 6009 31807
rect 6009 31773 6043 31807
rect 6043 31773 6052 31807
rect 6000 31764 6052 31773
rect 1676 31628 1728 31680
rect 1952 31628 2004 31680
rect 3240 31628 3292 31680
rect 3516 31628 3568 31680
rect 4528 31628 4580 31680
rect 5264 31628 5316 31680
rect 5448 31628 5500 31680
rect 7196 31628 7248 31680
rect 8576 31807 8628 31816
rect 8576 31773 8585 31807
rect 8585 31773 8619 31807
rect 8619 31773 8628 31807
rect 8576 31764 8628 31773
rect 8668 31764 8720 31816
rect 9312 31764 9364 31816
rect 8116 31696 8168 31748
rect 8944 31696 8996 31748
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 8760 31671 8812 31680
rect 8760 31637 8769 31671
rect 8769 31637 8803 31671
rect 8803 31637 8812 31671
rect 8760 31628 8812 31637
rect 3010 31526 3062 31578
rect 3074 31526 3126 31578
rect 3138 31526 3190 31578
rect 3202 31526 3254 31578
rect 3266 31526 3318 31578
rect 9010 31526 9062 31578
rect 9074 31526 9126 31578
rect 9138 31526 9190 31578
rect 9202 31526 9254 31578
rect 9266 31526 9318 31578
rect 1492 31424 1544 31476
rect 2872 31424 2924 31476
rect 3608 31424 3660 31476
rect 1308 31288 1360 31340
rect 1676 31288 1728 31340
rect 2044 31356 2096 31408
rect 3332 31331 3384 31340
rect 3332 31297 3341 31331
rect 3341 31297 3375 31331
rect 3375 31297 3384 31331
rect 3332 31288 3384 31297
rect 4528 31331 4580 31340
rect 4528 31297 4546 31331
rect 4546 31297 4580 31331
rect 4528 31288 4580 31297
rect 6000 31424 6052 31476
rect 8116 31424 8168 31476
rect 8576 31424 8628 31476
rect 6460 31356 6512 31408
rect 6920 31356 6972 31408
rect 7748 31288 7800 31340
rect 8576 31331 8628 31340
rect 8576 31297 8585 31331
rect 8585 31297 8619 31331
rect 8619 31297 8628 31331
rect 8576 31288 8628 31297
rect 8852 31331 8904 31340
rect 8852 31297 8861 31331
rect 8861 31297 8895 31331
rect 8895 31297 8904 31331
rect 8852 31288 8904 31297
rect 9772 31331 9824 31340
rect 9772 31297 9781 31331
rect 9781 31297 9815 31331
rect 9815 31297 9824 31331
rect 9772 31288 9824 31297
rect 3608 31220 3660 31272
rect 4804 31220 4856 31272
rect 5448 31220 5500 31272
rect 4252 31084 4304 31136
rect 4896 31195 4948 31204
rect 4896 31161 4905 31195
rect 4905 31161 4939 31195
rect 4939 31161 4948 31195
rect 4896 31152 4948 31161
rect 5172 31152 5224 31204
rect 7656 31263 7708 31272
rect 7656 31229 7665 31263
rect 7665 31229 7699 31263
rect 7699 31229 7708 31263
rect 7656 31220 7708 31229
rect 8300 31263 8352 31272
rect 8300 31229 8309 31263
rect 8309 31229 8343 31263
rect 8343 31229 8352 31263
rect 8300 31220 8352 31229
rect 8392 31220 8444 31272
rect 8668 31263 8720 31272
rect 8668 31229 8702 31263
rect 8702 31229 8720 31263
rect 8668 31220 8720 31229
rect 9036 31220 9088 31272
rect 9404 31220 9456 31272
rect 10140 31220 10192 31272
rect 5632 31152 5684 31204
rect 5080 31084 5132 31136
rect 5540 31084 5592 31136
rect 8576 31084 8628 31136
rect 8852 31084 8904 31136
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 7950 30982 8002 31034
rect 8014 30982 8066 31034
rect 8078 30982 8130 31034
rect 8142 30982 8194 31034
rect 8206 30982 8258 31034
rect 2412 30880 2464 30932
rect 3608 30923 3660 30932
rect 3608 30889 3617 30923
rect 3617 30889 3651 30923
rect 3651 30889 3660 30923
rect 3608 30880 3660 30889
rect 6000 30880 6052 30932
rect 7564 30880 7616 30932
rect 10232 30880 10284 30932
rect 2596 30812 2648 30864
rect 4528 30812 4580 30864
rect 5540 30812 5592 30864
rect 9680 30812 9732 30864
rect 3332 30744 3384 30796
rect 1676 30676 1728 30728
rect 2412 30676 2464 30728
rect 2596 30719 2648 30728
rect 2596 30685 2605 30719
rect 2605 30685 2639 30719
rect 2639 30685 2648 30719
rect 2596 30676 2648 30685
rect 3516 30676 3568 30728
rect 6184 30744 6236 30796
rect 8668 30744 8720 30796
rect 4712 30676 4764 30728
rect 6460 30676 6512 30728
rect 7196 30676 7248 30728
rect 8392 30719 8444 30728
rect 8392 30685 8401 30719
rect 8401 30685 8435 30719
rect 8435 30685 8444 30719
rect 8392 30676 8444 30685
rect 6276 30608 6328 30660
rect 8760 30676 8812 30728
rect 9956 30744 10008 30796
rect 2872 30540 2924 30592
rect 5816 30540 5868 30592
rect 8392 30540 8444 30592
rect 9956 30608 10008 30660
rect 10048 30608 10100 30660
rect 10324 30608 10376 30660
rect 9312 30540 9364 30592
rect 9496 30540 9548 30592
rect 9588 30540 9640 30592
rect 10140 30540 10192 30592
rect 3010 30438 3062 30490
rect 3074 30438 3126 30490
rect 3138 30438 3190 30490
rect 3202 30438 3254 30490
rect 3266 30438 3318 30490
rect 9010 30438 9062 30490
rect 9074 30438 9126 30490
rect 9138 30438 9190 30490
rect 9202 30438 9254 30490
rect 9266 30438 9318 30490
rect 1492 30336 1544 30388
rect 1492 30243 1544 30252
rect 1492 30209 1501 30243
rect 1501 30209 1535 30243
rect 1535 30209 1544 30243
rect 1492 30200 1544 30209
rect 4528 30336 4580 30388
rect 5080 30336 5132 30388
rect 7748 30336 7800 30388
rect 9220 30336 9272 30388
rect 1768 30268 1820 30320
rect 3332 30268 3384 30320
rect 9772 30268 9824 30320
rect 4712 30200 4764 30252
rect 6460 30200 6512 30252
rect 7104 30200 7156 30252
rect 8116 30243 8168 30252
rect 8116 30209 8125 30243
rect 8125 30209 8159 30243
rect 8159 30209 8168 30243
rect 8116 30200 8168 30209
rect 8392 30243 8444 30252
rect 8392 30209 8401 30243
rect 8401 30209 8435 30243
rect 8435 30209 8444 30243
rect 8392 30200 8444 30209
rect 1768 30132 1820 30184
rect 2596 30132 2648 30184
rect 3516 30132 3568 30184
rect 6828 30132 6880 30184
rect 7748 30132 7800 30184
rect 8300 30132 8352 30184
rect 8576 30132 8628 30184
rect 9312 30200 9364 30252
rect 4896 30064 4948 30116
rect 7564 30064 7616 30116
rect 112 29996 164 30048
rect 1676 29996 1728 30048
rect 3700 29996 3752 30048
rect 9680 30132 9732 30184
rect 10324 30064 10376 30116
rect 10600 29996 10652 30048
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 7950 29894 8002 29946
rect 8014 29894 8066 29946
rect 8078 29894 8130 29946
rect 8142 29894 8194 29946
rect 8206 29894 8258 29946
rect 5356 29792 5408 29844
rect 6460 29835 6512 29844
rect 6460 29801 6469 29835
rect 6469 29801 6503 29835
rect 6503 29801 6512 29835
rect 6460 29792 6512 29801
rect 7196 29792 7248 29844
rect 7472 29792 7524 29844
rect 7564 29835 7616 29844
rect 7564 29801 7573 29835
rect 7573 29801 7607 29835
rect 7607 29801 7616 29835
rect 7564 29792 7616 29801
rect 1400 29724 1452 29776
rect 2228 29724 2280 29776
rect 2412 29724 2464 29776
rect 2688 29724 2740 29776
rect 3424 29724 3476 29776
rect 5172 29656 5224 29708
rect 5356 29656 5408 29708
rect 6184 29656 6236 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 2596 29588 2648 29640
rect 4712 29588 4764 29640
rect 1584 29452 1636 29504
rect 2320 29452 2372 29504
rect 3608 29452 3660 29504
rect 4068 29452 4120 29504
rect 5540 29631 5592 29640
rect 5540 29597 5549 29631
rect 5549 29597 5583 29631
rect 5583 29597 5592 29631
rect 5540 29588 5592 29597
rect 5632 29631 5684 29640
rect 5632 29597 5666 29631
rect 5666 29597 5684 29631
rect 5632 29588 5684 29597
rect 6828 29631 6880 29640
rect 6828 29597 6837 29631
rect 6837 29597 6871 29631
rect 6871 29597 6880 29631
rect 6828 29588 6880 29597
rect 8024 29767 8076 29776
rect 8024 29733 8033 29767
rect 8033 29733 8067 29767
rect 8067 29733 8076 29767
rect 8024 29724 8076 29733
rect 9772 29724 9824 29776
rect 9404 29699 9456 29708
rect 9404 29665 9413 29699
rect 9413 29665 9447 29699
rect 9447 29665 9456 29699
rect 9404 29656 9456 29665
rect 9496 29699 9548 29708
rect 9496 29665 9505 29699
rect 9505 29665 9539 29699
rect 9539 29665 9548 29699
rect 9496 29656 9548 29665
rect 8024 29588 8076 29640
rect 8116 29631 8168 29640
rect 8116 29597 8125 29631
rect 8125 29597 8159 29631
rect 8159 29597 8168 29631
rect 8116 29588 8168 29597
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 9036 29588 9088 29640
rect 10692 29588 10744 29640
rect 5448 29452 5500 29504
rect 5540 29452 5592 29504
rect 5816 29452 5868 29504
rect 9956 29520 10008 29572
rect 9220 29452 9272 29504
rect 9588 29452 9640 29504
rect 3010 29350 3062 29402
rect 3074 29350 3126 29402
rect 3138 29350 3190 29402
rect 3202 29350 3254 29402
rect 3266 29350 3318 29402
rect 9010 29350 9062 29402
rect 9074 29350 9126 29402
rect 9138 29350 9190 29402
rect 9202 29350 9254 29402
rect 9266 29350 9318 29402
rect 664 29248 716 29300
rect 2320 29248 2372 29300
rect 1768 29180 1820 29232
rect 388 29112 440 29164
rect 5172 29291 5224 29300
rect 5172 29257 5181 29291
rect 5181 29257 5215 29291
rect 5215 29257 5224 29291
rect 5172 29248 5224 29257
rect 2964 29180 3016 29232
rect 3516 29180 3568 29232
rect 3608 29180 3660 29232
rect 1768 29087 1820 29096
rect 1768 29053 1777 29087
rect 1777 29053 1811 29087
rect 1811 29053 1820 29087
rect 1768 29044 1820 29053
rect 2688 28908 2740 28960
rect 4160 29087 4212 29096
rect 4160 29053 4169 29087
rect 4169 29053 4203 29087
rect 4203 29053 4212 29087
rect 4160 29044 4212 29053
rect 7196 29180 7248 29232
rect 7104 29112 7156 29164
rect 7564 29112 7616 29164
rect 8116 29155 8168 29164
rect 8116 29121 8125 29155
rect 8125 29121 8159 29155
rect 8159 29121 8168 29155
rect 8116 29112 8168 29121
rect 9220 29112 9272 29164
rect 9680 29112 9732 29164
rect 7104 28976 7156 29028
rect 7472 29044 7524 29096
rect 8208 29087 8260 29096
rect 8208 29053 8242 29087
rect 8242 29053 8260 29087
rect 8208 29044 8260 29053
rect 8392 29087 8444 29096
rect 8392 29053 8401 29087
rect 8401 29053 8435 29087
rect 8435 29053 8444 29087
rect 8392 29044 8444 29053
rect 8760 29044 8812 29096
rect 9864 29044 9916 29096
rect 9956 29044 10008 29096
rect 7748 28976 7800 29028
rect 7840 29019 7892 29028
rect 7840 28985 7849 29019
rect 7849 28985 7883 29019
rect 7883 28985 7892 29019
rect 7840 28976 7892 28985
rect 9588 28976 9640 29028
rect 9680 29019 9732 29028
rect 9680 28985 9689 29019
rect 9689 28985 9723 29019
rect 9723 28985 9732 29019
rect 9680 28976 9732 28985
rect 4252 28908 4304 28960
rect 4436 28908 4488 28960
rect 5172 28908 5224 28960
rect 7380 28908 7432 28960
rect 7932 28908 7984 28960
rect 8576 28908 8628 28960
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 7950 28806 8002 28858
rect 8014 28806 8066 28858
rect 8078 28806 8130 28858
rect 8142 28806 8194 28858
rect 8206 28806 8258 28858
rect 1400 28704 1452 28756
rect 1216 28636 1268 28688
rect 3240 28704 3292 28756
rect 3608 28747 3660 28756
rect 3608 28713 3617 28747
rect 3617 28713 3651 28747
rect 3651 28713 3660 28747
rect 3608 28704 3660 28713
rect 4804 28704 4856 28756
rect 5356 28704 5408 28756
rect 8392 28704 8444 28756
rect 7932 28636 7984 28688
rect 9404 28704 9456 28756
rect 10232 28636 10284 28688
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 2136 28500 2188 28552
rect 388 28432 440 28484
rect 3332 28568 3384 28620
rect 3608 28568 3660 28620
rect 5448 28568 5500 28620
rect 2412 28364 2464 28416
rect 4160 28500 4212 28552
rect 4252 28543 4304 28552
rect 4252 28509 4261 28543
rect 4261 28509 4295 28543
rect 4295 28509 4304 28543
rect 4252 28500 4304 28509
rect 4988 28500 5040 28552
rect 6184 28568 6236 28620
rect 10324 28568 10376 28620
rect 3240 28432 3292 28484
rect 4804 28432 4856 28484
rect 5908 28432 5960 28484
rect 6552 28432 6604 28484
rect 7104 28500 7156 28552
rect 8576 28543 8628 28552
rect 8576 28509 8585 28543
rect 8585 28509 8619 28543
rect 8619 28509 8628 28543
rect 8576 28500 8628 28509
rect 8668 28500 8720 28552
rect 9404 28500 9456 28552
rect 11060 28432 11112 28484
rect 3516 28364 3568 28416
rect 4436 28364 4488 28416
rect 5080 28364 5132 28416
rect 5448 28364 5500 28416
rect 6736 28364 6788 28416
rect 8760 28407 8812 28416
rect 8760 28373 8769 28407
rect 8769 28373 8803 28407
rect 8803 28373 8812 28407
rect 8760 28364 8812 28373
rect 10416 28364 10468 28416
rect 3010 28262 3062 28314
rect 3074 28262 3126 28314
rect 3138 28262 3190 28314
rect 3202 28262 3254 28314
rect 3266 28262 3318 28314
rect 9010 28262 9062 28314
rect 9074 28262 9126 28314
rect 9138 28262 9190 28314
rect 9202 28262 9254 28314
rect 9266 28262 9318 28314
rect 2412 28203 2464 28212
rect 2412 28169 2421 28203
rect 2421 28169 2455 28203
rect 2455 28169 2464 28203
rect 2412 28160 2464 28169
rect 1768 28092 1820 28144
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 4160 28160 4212 28212
rect 5816 28160 5868 28212
rect 4804 28092 4856 28144
rect 5448 28024 5500 28076
rect 5816 28024 5868 28076
rect 6184 28024 6236 28076
rect 6828 28160 6880 28212
rect 7840 28160 7892 28212
rect 8116 28203 8168 28212
rect 8116 28169 8125 28203
rect 8125 28169 8159 28203
rect 8159 28169 8168 28203
rect 8116 28160 8168 28169
rect 9496 28160 9548 28212
rect 6920 28092 6972 28144
rect 7840 28024 7892 28076
rect 8576 28024 8628 28076
rect 8760 28024 8812 28076
rect 2688 27956 2740 28008
rect 3240 27999 3292 28008
rect 3240 27965 3258 27999
rect 3258 27965 3292 27999
rect 3240 27956 3292 27965
rect 3516 27888 3568 27940
rect 1676 27820 1728 27872
rect 3056 27820 3108 27872
rect 4068 27999 4120 28008
rect 4068 27965 4077 27999
rect 4077 27965 4111 27999
rect 4111 27965 4120 27999
rect 4068 27956 4120 27965
rect 4252 27999 4304 28008
rect 4252 27965 4261 27999
rect 4261 27965 4295 27999
rect 4295 27965 4304 27999
rect 4252 27956 4304 27965
rect 3884 27820 3936 27872
rect 6828 27820 6880 27872
rect 7932 27820 7984 27872
rect 9680 27863 9732 27872
rect 9680 27829 9689 27863
rect 9689 27829 9723 27863
rect 9723 27829 9732 27863
rect 9680 27820 9732 27829
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 7950 27718 8002 27770
rect 8014 27718 8066 27770
rect 8078 27718 8130 27770
rect 8142 27718 8194 27770
rect 8206 27718 8258 27770
rect 1216 27616 1268 27668
rect 2872 27616 2924 27668
rect 3240 27616 3292 27668
rect 3792 27616 3844 27668
rect 2228 27412 2280 27464
rect 2596 27455 2648 27464
rect 2596 27421 2605 27455
rect 2605 27421 2639 27455
rect 2639 27421 2648 27455
rect 4436 27480 4488 27532
rect 5540 27616 5592 27668
rect 5816 27616 5868 27668
rect 6000 27616 6052 27668
rect 8392 27616 8444 27668
rect 8760 27591 8812 27600
rect 8760 27557 8769 27591
rect 8769 27557 8803 27591
rect 8803 27557 8812 27591
rect 8760 27548 8812 27557
rect 10232 27548 10284 27600
rect 2596 27412 2648 27421
rect 3516 27412 3568 27464
rect 4896 27412 4948 27464
rect 5080 27412 5132 27464
rect 7012 27412 7064 27464
rect 7840 27412 7892 27464
rect 8576 27455 8628 27464
rect 8576 27421 8585 27455
rect 8585 27421 8619 27455
rect 8619 27421 8628 27455
rect 8576 27412 8628 27421
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 10140 27412 10192 27464
rect 10600 27412 10652 27464
rect 7104 27344 7156 27396
rect 8668 27344 8720 27396
rect 10968 27344 11020 27396
rect 848 27276 900 27328
rect 2044 27276 2096 27328
rect 4344 27276 4396 27328
rect 4528 27276 4580 27328
rect 4896 27276 4948 27328
rect 5448 27276 5500 27328
rect 6276 27276 6328 27328
rect 6920 27276 6972 27328
rect 9496 27276 9548 27328
rect 10784 27276 10836 27328
rect 3010 27174 3062 27226
rect 3074 27174 3126 27226
rect 3138 27174 3190 27226
rect 3202 27174 3254 27226
rect 3266 27174 3318 27226
rect 9010 27174 9062 27226
rect 9074 27174 9126 27226
rect 9138 27174 9190 27226
rect 9202 27174 9254 27226
rect 9266 27174 9318 27226
rect 2044 27072 2096 27124
rect 3516 27072 3568 27124
rect 3792 27072 3844 27124
rect 4068 27072 4120 27124
rect 4620 27072 4672 27124
rect 1492 27004 1544 27056
rect 1952 27004 2004 27056
rect 2320 27004 2372 27056
rect 2504 27004 2556 27056
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 1676 26936 1728 26988
rect 2228 26936 2280 26988
rect 5264 27004 5316 27056
rect 5172 26979 5224 26988
rect 5172 26945 5181 26979
rect 5181 26945 5215 26979
rect 5215 26945 5224 26979
rect 6460 27072 6512 27124
rect 7840 27072 7892 27124
rect 10324 27072 10376 27124
rect 5172 26936 5224 26945
rect 6920 26936 6972 26988
rect 10508 27004 10560 27056
rect 1768 26868 1820 26920
rect 3240 26868 3292 26920
rect 3792 26911 3844 26920
rect 3792 26877 3810 26911
rect 3810 26877 3844 26911
rect 3792 26868 3844 26877
rect 4436 26868 4488 26920
rect 4620 26911 4672 26920
rect 4620 26877 4629 26911
rect 4629 26877 4663 26911
rect 4663 26877 4672 26911
rect 4620 26868 4672 26877
rect 4896 26911 4948 26920
rect 4896 26877 4905 26911
rect 4905 26877 4939 26911
rect 4939 26877 4948 26911
rect 4896 26868 4948 26877
rect 2780 26732 2832 26784
rect 6460 26800 6512 26852
rect 9404 26936 9456 26988
rect 9496 26979 9548 26988
rect 9496 26945 9505 26979
rect 9505 26945 9539 26979
rect 9539 26945 9548 26979
rect 9496 26936 9548 26945
rect 9772 26868 9824 26920
rect 10048 26868 10100 26920
rect 10508 26868 10560 26920
rect 9312 26800 9364 26852
rect 5356 26732 5408 26784
rect 5724 26732 5776 26784
rect 5816 26732 5868 26784
rect 8760 26732 8812 26784
rect 9680 26775 9732 26784
rect 9680 26741 9689 26775
rect 9689 26741 9723 26775
rect 9723 26741 9732 26775
rect 9680 26732 9732 26741
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 7950 26630 8002 26682
rect 8014 26630 8066 26682
rect 8078 26630 8130 26682
rect 8142 26630 8194 26682
rect 8206 26630 8258 26682
rect 3240 26571 3292 26580
rect 3240 26537 3249 26571
rect 3249 26537 3283 26571
rect 3283 26537 3292 26571
rect 3240 26528 3292 26537
rect 3700 26528 3752 26580
rect 4896 26528 4948 26580
rect 5080 26528 5132 26580
rect 5632 26460 5684 26512
rect 6920 26571 6972 26580
rect 6920 26537 6929 26571
rect 6929 26537 6963 26571
rect 6963 26537 6972 26571
rect 6920 26528 6972 26537
rect 9588 26528 9640 26580
rect 4896 26392 4948 26444
rect 6276 26435 6328 26444
rect 6276 26401 6285 26435
rect 6285 26401 6319 26435
rect 6319 26401 6328 26435
rect 6276 26392 6328 26401
rect 664 26324 716 26376
rect 1676 26324 1728 26376
rect 1860 26324 1912 26376
rect 2412 26324 2464 26376
rect 2780 26324 2832 26376
rect 3792 26324 3844 26376
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 6000 26367 6052 26392
rect 6000 26340 6009 26367
rect 6009 26340 6043 26367
rect 6043 26340 6052 26367
rect 6092 26340 6144 26392
rect 8484 26460 8536 26512
rect 10232 26460 10284 26512
rect 4528 26299 4580 26308
rect 4528 26265 4537 26299
rect 4537 26265 4571 26299
rect 4571 26265 4580 26299
rect 4528 26256 4580 26265
rect 4620 26256 4672 26308
rect 6920 26324 6972 26376
rect 7932 26324 7984 26376
rect 8208 26324 8260 26376
rect 8852 26324 8904 26376
rect 8944 26324 8996 26376
rect 9496 26367 9548 26376
rect 9496 26333 9505 26367
rect 9505 26333 9539 26367
rect 9539 26333 9548 26367
rect 9496 26324 9548 26333
rect 1952 26231 2004 26240
rect 1952 26197 1961 26231
rect 1961 26197 1995 26231
rect 1995 26197 2004 26231
rect 1952 26188 2004 26197
rect 2964 26188 3016 26240
rect 3792 26188 3844 26240
rect 3884 26188 3936 26240
rect 4804 26231 4856 26240
rect 4804 26197 4813 26231
rect 4813 26197 4847 26231
rect 4847 26197 4856 26231
rect 4804 26188 4856 26197
rect 8300 26256 8352 26308
rect 10600 26256 10652 26308
rect 7840 26188 7892 26240
rect 3010 26086 3062 26138
rect 3074 26086 3126 26138
rect 3138 26086 3190 26138
rect 3202 26086 3254 26138
rect 3266 26086 3318 26138
rect 9010 26086 9062 26138
rect 9074 26086 9126 26138
rect 9138 26086 9190 26138
rect 9202 26086 9254 26138
rect 9266 26086 9318 26138
rect 10600 26120 10652 26172
rect 204 25984 256 26036
rect 3424 25984 3476 26036
rect 3884 25984 3936 26036
rect 6092 25984 6144 26036
rect 7564 25984 7616 26036
rect 7840 25984 7892 26036
rect 1768 25916 1820 25968
rect 2412 25848 2464 25900
rect 2964 25916 3016 25968
rect 6276 25916 6328 25968
rect 2596 25891 2648 25900
rect 2596 25857 2605 25891
rect 2605 25857 2639 25891
rect 2639 25857 2648 25891
rect 2596 25848 2648 25857
rect 3608 25848 3660 25900
rect 6736 25848 6788 25900
rect 7288 25848 7340 25900
rect 8484 25984 8536 26036
rect 3700 25780 3752 25832
rect 7656 25780 7708 25832
rect 8300 25712 8352 25764
rect 8944 25780 8996 25832
rect 9496 25712 9548 25764
rect 2504 25644 2556 25696
rect 6828 25644 6880 25696
rect 8576 25644 8628 25696
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 7950 25542 8002 25594
rect 8014 25542 8066 25594
rect 8078 25542 8130 25594
rect 8142 25542 8194 25594
rect 8206 25542 8258 25594
rect 296 25440 348 25492
rect 2872 25440 2924 25492
rect 3056 25440 3108 25492
rect 4804 25372 4856 25424
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 2504 25236 2556 25288
rect 4620 25304 4672 25356
rect 7564 25440 7616 25492
rect 7932 25440 7984 25492
rect 9496 25440 9548 25492
rect 4988 25236 5040 25288
rect 5172 25236 5224 25288
rect 5448 25236 5500 25288
rect 6920 25236 6972 25288
rect 7104 25236 7156 25288
rect 8024 25236 8076 25288
rect 8208 25236 8260 25288
rect 8944 25372 8996 25424
rect 10232 25372 10284 25424
rect 10324 25372 10376 25424
rect 11152 25372 11204 25424
rect 2228 25100 2280 25152
rect 3056 25168 3108 25220
rect 7564 25168 7616 25220
rect 8576 25279 8628 25288
rect 8576 25245 8585 25279
rect 8585 25245 8619 25279
rect 8619 25245 8628 25279
rect 8576 25236 8628 25245
rect 5816 25143 5868 25152
rect 5816 25109 5825 25143
rect 5825 25109 5859 25143
rect 5859 25109 5868 25143
rect 5816 25100 5868 25109
rect 6920 25100 6972 25152
rect 7932 25100 7984 25152
rect 8208 25100 8260 25152
rect 8300 25100 8352 25152
rect 9036 25236 9088 25288
rect 9404 25236 9456 25288
rect 10140 25304 10192 25356
rect 10876 25304 10928 25356
rect 10048 25168 10100 25220
rect 9680 25143 9732 25152
rect 9680 25109 9689 25143
rect 9689 25109 9723 25143
rect 9723 25109 9732 25143
rect 9680 25100 9732 25109
rect 3010 24998 3062 25050
rect 3074 24998 3126 25050
rect 3138 24998 3190 25050
rect 3202 24998 3254 25050
rect 3266 24998 3318 25050
rect 9010 24998 9062 25050
rect 9074 24998 9126 25050
rect 9138 24998 9190 25050
rect 9202 24998 9254 25050
rect 9266 24998 9318 25050
rect 2964 24896 3016 24948
rect 3884 24896 3936 24948
rect 4988 24896 5040 24948
rect 5448 24896 5500 24948
rect 6736 24896 6788 24948
rect 7196 24896 7248 24948
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 2136 24760 2188 24812
rect 5448 24803 5500 24812
rect 5448 24769 5457 24803
rect 5457 24769 5491 24803
rect 5491 24769 5500 24803
rect 5448 24760 5500 24769
rect 7104 24760 7156 24812
rect 8116 24803 8168 24812
rect 8116 24769 8125 24803
rect 8125 24769 8159 24803
rect 8159 24769 8168 24803
rect 8116 24760 8168 24769
rect 8208 24803 8260 24812
rect 8208 24769 8242 24803
rect 8242 24769 8260 24803
rect 9404 24828 9456 24880
rect 8208 24760 8260 24769
rect 10784 24760 10836 24812
rect 664 24692 716 24744
rect 2228 24692 2280 24744
rect 2412 24735 2464 24744
rect 2412 24701 2421 24735
rect 2421 24701 2455 24735
rect 2455 24701 2464 24735
rect 2412 24692 2464 24701
rect 3148 24692 3200 24744
rect 3792 24692 3844 24744
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 4160 24667 4212 24676
rect 4160 24633 4169 24667
rect 4169 24633 4203 24667
rect 4203 24633 4212 24667
rect 4160 24624 4212 24633
rect 3884 24556 3936 24608
rect 4620 24692 4672 24744
rect 4712 24735 4764 24744
rect 4712 24701 4721 24735
rect 4721 24701 4755 24735
rect 4755 24701 4764 24735
rect 4712 24692 4764 24701
rect 7196 24735 7248 24744
rect 7196 24701 7205 24735
rect 7205 24701 7239 24735
rect 7239 24701 7248 24735
rect 7196 24692 7248 24701
rect 6276 24624 6328 24676
rect 7932 24692 7984 24744
rect 8392 24735 8444 24744
rect 8392 24701 8401 24735
rect 8401 24701 8435 24735
rect 8435 24701 8444 24735
rect 8392 24692 8444 24701
rect 8576 24692 8628 24744
rect 8944 24692 8996 24744
rect 7840 24667 7892 24676
rect 7840 24633 7849 24667
rect 7849 24633 7883 24667
rect 7883 24633 7892 24667
rect 7840 24624 7892 24633
rect 9496 24624 9548 24676
rect 9772 24624 9824 24676
rect 5172 24556 5224 24608
rect 6644 24556 6696 24608
rect 7196 24556 7248 24608
rect 7288 24556 7340 24608
rect 8116 24556 8168 24608
rect 8576 24556 8628 24608
rect 9680 24599 9732 24608
rect 9680 24565 9689 24599
rect 9689 24565 9723 24599
rect 9723 24565 9732 24599
rect 9680 24556 9732 24565
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 7950 24454 8002 24506
rect 8014 24454 8066 24506
rect 8078 24454 8130 24506
rect 8142 24454 8194 24506
rect 8206 24454 8258 24506
rect 1492 24352 1544 24404
rect 6460 24352 6512 24404
rect 8392 24352 8444 24404
rect 9772 24352 9824 24404
rect 4896 24284 4948 24336
rect 5356 24284 5408 24336
rect 6276 24284 6328 24336
rect 6920 24284 6972 24336
rect 1860 24216 1912 24268
rect 2136 24216 2188 24268
rect 2412 24259 2464 24268
rect 2412 24225 2421 24259
rect 2421 24225 2455 24259
rect 2455 24225 2464 24259
rect 2412 24216 2464 24225
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 2320 24148 2372 24200
rect 2228 24080 2280 24132
rect 4160 24080 4212 24132
rect 2320 24012 2372 24064
rect 2596 24012 2648 24064
rect 4436 24012 4488 24064
rect 4620 24012 4672 24064
rect 5816 24191 5868 24200
rect 5816 24157 5825 24191
rect 5825 24157 5859 24191
rect 5859 24157 5868 24191
rect 5816 24148 5868 24157
rect 8944 24284 8996 24336
rect 10232 24284 10284 24336
rect 8852 24216 8904 24268
rect 6644 24148 6696 24200
rect 7288 24148 7340 24200
rect 8024 24148 8076 24200
rect 8576 24191 8628 24200
rect 8576 24157 8585 24191
rect 8585 24157 8619 24191
rect 8619 24157 8628 24191
rect 8576 24148 8628 24157
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 7932 24080 7984 24132
rect 6460 24012 6512 24064
rect 8760 24055 8812 24064
rect 8760 24021 8769 24055
rect 8769 24021 8803 24055
rect 8803 24021 8812 24055
rect 8760 24012 8812 24021
rect 3010 23910 3062 23962
rect 3074 23910 3126 23962
rect 3138 23910 3190 23962
rect 3202 23910 3254 23962
rect 3266 23910 3318 23962
rect 9010 23910 9062 23962
rect 9074 23910 9126 23962
rect 9138 23910 9190 23962
rect 9202 23910 9254 23962
rect 9266 23910 9318 23962
rect 2228 23808 2280 23860
rect 5448 23808 5500 23860
rect 5540 23808 5592 23860
rect 7748 23808 7800 23860
rect 7840 23808 7892 23860
rect 8668 23808 8720 23860
rect 9312 23808 9364 23860
rect 9680 23851 9732 23860
rect 9680 23817 9689 23851
rect 9689 23817 9723 23851
rect 9723 23817 9732 23851
rect 9680 23808 9732 23817
rect 2136 23740 2188 23792
rect 2596 23740 2648 23792
rect 3240 23740 3292 23792
rect 1492 23672 1544 23724
rect 6368 23740 6420 23792
rect 6736 23740 6788 23792
rect 7380 23740 7432 23792
rect 4160 23715 4212 23724
rect 4160 23681 4169 23715
rect 4169 23681 4203 23715
rect 4203 23681 4212 23715
rect 4160 23672 4212 23681
rect 4436 23715 4488 23724
rect 4436 23681 4445 23715
rect 4445 23681 4479 23715
rect 4479 23681 4488 23715
rect 4436 23672 4488 23681
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 5908 23672 5960 23724
rect 8208 23672 8260 23724
rect 1860 23604 1912 23656
rect 3884 23647 3936 23656
rect 3884 23613 3893 23647
rect 3893 23613 3927 23647
rect 3927 23613 3936 23647
rect 3884 23604 3936 23613
rect 6276 23604 6328 23656
rect 7288 23647 7340 23656
rect 7288 23613 7297 23647
rect 7297 23613 7331 23647
rect 7331 23613 7340 23647
rect 7288 23604 7340 23613
rect 8852 23740 8904 23792
rect 8760 23672 8812 23724
rect 10968 23604 11020 23656
rect 5448 23536 5500 23588
rect 9864 23536 9916 23588
rect 4620 23468 4672 23520
rect 8484 23468 8536 23520
rect 10232 23468 10284 23520
rect 112 23400 164 23452
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 7950 23366 8002 23418
rect 8014 23366 8066 23418
rect 8078 23366 8130 23418
rect 8142 23366 8194 23418
rect 8206 23366 8258 23418
rect 2872 23264 2924 23316
rect 4712 23264 4764 23316
rect 6828 23264 6880 23316
rect 7380 23264 7432 23316
rect 7564 23264 7616 23316
rect 7748 23264 7800 23316
rect 8760 23264 8812 23316
rect 9588 23264 9640 23316
rect 480 23196 532 23248
rect 1952 23196 2004 23248
rect 9680 23239 9732 23248
rect 9680 23205 9689 23239
rect 9689 23205 9723 23239
rect 9723 23205 9732 23239
rect 9680 23196 9732 23205
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2596 23128 2648 23180
rect 4620 23128 4672 23180
rect 6368 23128 6420 23180
rect 7012 23128 7064 23180
rect 1860 23060 1912 23112
rect 1584 22992 1636 23044
rect 2044 22992 2096 23044
rect 5724 23060 5776 23112
rect 9404 23128 9456 23180
rect 9588 23128 9640 23180
rect 4804 22992 4856 23044
rect 7932 23060 7984 23112
rect 8024 23103 8076 23112
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 8576 22992 8628 23044
rect 2688 22924 2740 22976
rect 3792 22924 3844 22976
rect 5356 22924 5408 22976
rect 6000 22924 6052 22976
rect 6276 22924 6328 22976
rect 8852 22924 8904 22976
rect 10232 22924 10284 22976
rect 3010 22822 3062 22874
rect 3074 22822 3126 22874
rect 3138 22822 3190 22874
rect 3202 22822 3254 22874
rect 3266 22822 3318 22874
rect 9010 22822 9062 22874
rect 9074 22822 9126 22874
rect 9138 22822 9190 22874
rect 9202 22822 9254 22874
rect 9266 22822 9318 22874
rect 10232 22788 10284 22840
rect 10600 22788 10652 22840
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 1492 22584 1544 22636
rect 2780 22652 2832 22704
rect 2044 22584 2096 22636
rect 4620 22652 4672 22704
rect 4988 22584 5040 22636
rect 5172 22584 5224 22636
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 6368 22763 6420 22772
rect 6368 22729 6377 22763
rect 6377 22729 6411 22763
rect 6411 22729 6420 22763
rect 6368 22720 6420 22729
rect 7012 22720 7064 22772
rect 6276 22652 6328 22704
rect 6736 22584 6788 22636
rect 7012 22584 7064 22636
rect 7564 22652 7616 22704
rect 5264 22516 5316 22568
rect 5632 22516 5684 22568
rect 6368 22516 6420 22568
rect 7932 22516 7984 22568
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 4988 22448 5040 22500
rect 9864 22448 9916 22500
rect 2596 22380 2648 22432
rect 3424 22380 3476 22432
rect 4344 22380 4396 22432
rect 5264 22423 5316 22432
rect 5264 22389 5273 22423
rect 5273 22389 5307 22423
rect 5307 22389 5316 22423
rect 5264 22380 5316 22389
rect 6184 22423 6236 22432
rect 6184 22389 6193 22423
rect 6193 22389 6227 22423
rect 6227 22389 6236 22423
rect 6184 22380 6236 22389
rect 6736 22380 6788 22432
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 7950 22278 8002 22330
rect 8014 22278 8066 22330
rect 8078 22278 8130 22330
rect 8142 22278 8194 22330
rect 8206 22278 8258 22330
rect 3884 22176 3936 22228
rect 6736 22176 6788 22228
rect 1492 22040 1544 22092
rect 204 21972 256 22024
rect 572 21972 624 22024
rect 1400 21972 1452 22024
rect 4068 22108 4120 22160
rect 4528 22108 4580 22160
rect 5264 22151 5316 22160
rect 5264 22117 5273 22151
rect 5273 22117 5307 22151
rect 5307 22117 5316 22151
rect 5264 22108 5316 22117
rect 4160 22040 4212 22092
rect 5540 22083 5592 22092
rect 5540 22049 5549 22083
rect 5549 22049 5583 22083
rect 5583 22049 5592 22083
rect 5540 22040 5592 22049
rect 5632 22083 5684 22092
rect 5632 22049 5666 22083
rect 5666 22049 5684 22083
rect 5632 22040 5684 22049
rect 7012 22176 7064 22228
rect 7472 22176 7524 22228
rect 8300 22176 8352 22228
rect 7196 22108 7248 22160
rect 9588 22108 9640 22160
rect 10600 22108 10652 22160
rect 7932 22040 7984 22092
rect 9404 22040 9456 22092
rect 11152 22040 11204 22092
rect 1584 21904 1636 21956
rect 3240 21972 3292 22024
rect 3516 21972 3568 22024
rect 3884 21972 3936 22024
rect 4528 21972 4580 22024
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 5816 22015 5868 22024
rect 5816 21981 5825 22015
rect 5825 21981 5859 22015
rect 5859 21981 5868 22015
rect 5816 21972 5868 21981
rect 6828 21972 6880 22024
rect 8208 22015 8260 22024
rect 8208 21981 8217 22015
rect 8217 21981 8251 22015
rect 8251 21981 8260 22015
rect 8208 21972 8260 21981
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 8760 21972 8812 22024
rect 9220 21972 9272 22024
rect 2228 21904 2280 21956
rect 3700 21836 3752 21888
rect 5448 21836 5500 21888
rect 7012 21836 7064 21888
rect 9864 21904 9916 21956
rect 8760 21836 8812 21888
rect 9220 21836 9272 21888
rect 9588 21836 9640 21888
rect 9772 21836 9824 21888
rect 3010 21734 3062 21786
rect 3074 21734 3126 21786
rect 3138 21734 3190 21786
rect 3202 21734 3254 21786
rect 3266 21734 3318 21786
rect 9010 21734 9062 21786
rect 9074 21734 9126 21786
rect 9138 21734 9190 21786
rect 9202 21734 9254 21786
rect 9266 21734 9318 21786
rect 1584 21564 1636 21616
rect 1768 21564 1820 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 4620 21496 4672 21548
rect 4804 21496 4856 21548
rect 4988 21496 5040 21548
rect 2596 21428 2648 21480
rect 3332 21471 3384 21480
rect 3332 21437 3350 21471
rect 3350 21437 3384 21471
rect 3332 21428 3384 21437
rect 3700 21471 3752 21480
rect 3700 21437 3709 21471
rect 3709 21437 3743 21471
rect 3743 21437 3752 21471
rect 3700 21428 3752 21437
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 4344 21360 4396 21412
rect 5448 21675 5500 21684
rect 5448 21641 5457 21675
rect 5457 21641 5491 21675
rect 5491 21641 5500 21675
rect 5448 21632 5500 21641
rect 8208 21632 8260 21684
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 7472 21564 7524 21616
rect 5816 21496 5868 21548
rect 7012 21496 7064 21548
rect 9404 21496 9456 21548
rect 5356 21428 5408 21480
rect 7472 21471 7524 21480
rect 7472 21437 7481 21471
rect 7481 21437 7515 21471
rect 7515 21437 7524 21471
rect 7472 21428 7524 21437
rect 7564 21428 7616 21480
rect 5540 21360 5592 21412
rect 8484 21471 8536 21480
rect 8484 21437 8518 21471
rect 8518 21437 8536 21471
rect 8484 21428 8536 21437
rect 9036 21428 9088 21480
rect 7748 21360 7800 21412
rect 1032 21292 1084 21344
rect 1768 21292 1820 21344
rect 4068 21292 4120 21344
rect 4160 21292 4212 21344
rect 8208 21360 8260 21412
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 7950 21190 8002 21242
rect 8014 21190 8066 21242
rect 8078 21190 8130 21242
rect 8142 21190 8194 21242
rect 8206 21190 8258 21242
rect 10232 21156 10284 21208
rect 10692 21156 10744 21208
rect 4160 21088 4212 21140
rect 4252 21131 4304 21140
rect 4252 21097 4261 21131
rect 4261 21097 4295 21131
rect 4295 21097 4304 21131
rect 4252 21088 4304 21097
rect 5080 21131 5132 21140
rect 5080 21097 5089 21131
rect 5089 21097 5123 21131
rect 5123 21097 5132 21131
rect 5080 21088 5132 21097
rect 6460 21088 6512 21140
rect 6644 21088 6696 21140
rect 3332 21020 3384 21072
rect 3700 21020 3752 21072
rect 4344 21020 4396 21072
rect 2228 20995 2280 21004
rect 2228 20961 2237 20995
rect 2237 20961 2271 20995
rect 2271 20961 2280 20995
rect 2228 20952 2280 20961
rect 3976 20952 4028 21004
rect 4252 20952 4304 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 848 20816 900 20868
rect 2504 20927 2556 20936
rect 2504 20893 2513 20927
rect 2513 20893 2547 20927
rect 2547 20893 2556 20927
rect 2504 20884 2556 20893
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 6460 20952 6512 21004
rect 7564 20995 7616 21004
rect 7564 20961 7573 20995
rect 7573 20961 7607 20995
rect 7607 20961 7616 20995
rect 7564 20952 7616 20961
rect 8300 21088 8352 21140
rect 8760 21088 8812 21140
rect 9404 21088 9456 21140
rect 9680 21131 9732 21140
rect 9680 21097 9689 21131
rect 9689 21097 9723 21131
rect 9723 21097 9732 21131
rect 9680 21088 9732 21097
rect 10232 21020 10284 21072
rect 4804 20884 4856 20936
rect 7196 20900 7248 20952
rect 7932 20995 7984 21004
rect 7932 20961 7966 20995
rect 7966 20961 7984 20995
rect 7932 20952 7984 20961
rect 4528 20816 4580 20868
rect 6276 20816 6328 20868
rect 1860 20791 1912 20800
rect 1860 20757 1869 20791
rect 1869 20757 1903 20791
rect 1903 20757 1912 20791
rect 1860 20748 1912 20757
rect 3884 20748 3936 20800
rect 4160 20748 4212 20800
rect 5172 20748 5224 20800
rect 5816 20748 5868 20800
rect 8116 20927 8168 20936
rect 8116 20893 8125 20927
rect 8125 20893 8159 20927
rect 8159 20893 8168 20927
rect 8116 20884 8168 20893
rect 8760 20884 8812 20936
rect 10048 20884 10100 20936
rect 8208 20748 8260 20800
rect 8576 20748 8628 20800
rect 3010 20646 3062 20698
rect 3074 20646 3126 20698
rect 3138 20646 3190 20698
rect 3202 20646 3254 20698
rect 3266 20646 3318 20698
rect 9010 20646 9062 20698
rect 9074 20646 9126 20698
rect 9138 20646 9190 20698
rect 9202 20646 9254 20698
rect 9266 20646 9318 20698
rect 1768 20544 1820 20596
rect 3792 20544 3844 20596
rect 8116 20544 8168 20596
rect 8668 20587 8720 20596
rect 8668 20553 8677 20587
rect 8677 20553 8711 20587
rect 8711 20553 8720 20587
rect 8668 20544 8720 20553
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 3608 20476 3660 20528
rect 6276 20476 6328 20528
rect 7288 20476 7340 20528
rect 9588 20476 9640 20528
rect 1952 20408 2004 20460
rect 3884 20408 3936 20460
rect 6460 20408 6512 20460
rect 7196 20408 7248 20460
rect 7748 20408 7800 20460
rect 8576 20408 8628 20460
rect 6368 20340 6420 20392
rect 7288 20340 7340 20392
rect 9036 20408 9088 20460
rect 9220 20408 9272 20460
rect 8944 20340 8996 20392
rect 9772 20340 9824 20392
rect 1860 20272 1912 20324
rect 5172 20272 5224 20324
rect 7656 20272 7708 20324
rect 7932 20272 7984 20324
rect 10232 20272 10284 20324
rect 1768 20204 1820 20256
rect 2044 20204 2096 20256
rect 10048 20204 10100 20256
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 7950 20102 8002 20154
rect 8014 20102 8066 20154
rect 8078 20102 8130 20154
rect 8142 20102 8194 20154
rect 8206 20102 8258 20154
rect 1400 20000 1452 20052
rect 2596 20000 2648 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 4528 20043 4580 20052
rect 4528 20009 4537 20043
rect 4537 20009 4571 20043
rect 4571 20009 4580 20043
rect 4528 20000 4580 20009
rect 7564 20000 7616 20052
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 9680 20043 9732 20052
rect 9680 20009 9689 20043
rect 9689 20009 9723 20043
rect 9723 20009 9732 20043
rect 9680 20000 9732 20009
rect 10232 19932 10284 19984
rect 6368 19907 6420 19916
rect 6368 19873 6377 19907
rect 6377 19873 6411 19907
rect 6411 19873 6420 19907
rect 6368 19864 6420 19873
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 2504 19796 2556 19848
rect 2872 19796 2924 19848
rect 5172 19796 5224 19848
rect 6000 19796 6052 19848
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 7564 19728 7616 19780
rect 1768 19660 1820 19712
rect 2504 19660 2556 19712
rect 4068 19660 4120 19712
rect 6460 19660 6512 19712
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 10508 19796 10560 19848
rect 7932 19728 7984 19780
rect 9220 19728 9272 19780
rect 9864 19728 9916 19780
rect 10416 19728 10468 19780
rect 8760 19660 8812 19712
rect 3010 19558 3062 19610
rect 3074 19558 3126 19610
rect 3138 19558 3190 19610
rect 3202 19558 3254 19610
rect 3266 19558 3318 19610
rect 9010 19558 9062 19610
rect 9074 19558 9126 19610
rect 9138 19558 9190 19610
rect 9202 19558 9254 19610
rect 9266 19558 9318 19610
rect 2872 19499 2924 19508
rect 2872 19465 2881 19499
rect 2881 19465 2915 19499
rect 2915 19465 2924 19499
rect 2872 19456 2924 19465
rect 7288 19456 7340 19508
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2504 19388 2556 19440
rect 7932 19456 7984 19508
rect 8576 19456 8628 19508
rect 9680 19499 9732 19508
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 1676 19320 1728 19372
rect 3608 19320 3660 19372
rect 4344 19320 4396 19372
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 4620 19252 4672 19304
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 3700 19116 3752 19168
rect 4804 19184 4856 19236
rect 4068 19116 4120 19168
rect 7748 19388 7800 19440
rect 6276 19320 6328 19372
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 7472 19320 7524 19372
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 7932 19252 7984 19304
rect 9496 19363 9548 19372
rect 9496 19329 9505 19363
rect 9505 19329 9539 19363
rect 9539 19329 9548 19363
rect 9496 19320 9548 19329
rect 10324 19320 10376 19372
rect 10692 19320 10744 19372
rect 5908 19116 5960 19168
rect 7196 19116 7248 19168
rect 8576 19295 8628 19304
rect 8576 19261 8610 19295
rect 8610 19261 8628 19295
rect 8576 19252 8628 19261
rect 9128 19252 9180 19304
rect 9404 19252 9456 19304
rect 10876 19252 10928 19304
rect 8668 19116 8720 19168
rect 10048 19184 10100 19236
rect 9588 19116 9640 19168
rect 9864 19116 9916 19168
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 7950 19014 8002 19066
rect 8014 19014 8066 19066
rect 8078 19014 8130 19066
rect 8142 19014 8194 19066
rect 8206 19014 8258 19066
rect 4344 18912 4396 18964
rect 4712 18912 4764 18964
rect 3884 18844 3936 18896
rect 1676 18776 1728 18828
rect 1952 18819 2004 18828
rect 1952 18785 1961 18819
rect 1961 18785 1995 18819
rect 1995 18785 2004 18819
rect 1952 18776 2004 18785
rect 3700 18776 3752 18828
rect 4712 18819 4764 18828
rect 4712 18785 4721 18819
rect 4721 18785 4755 18819
rect 4755 18785 4764 18819
rect 5080 18844 5132 18896
rect 5172 18844 5224 18896
rect 4712 18776 4764 18785
rect 5908 18955 5960 18964
rect 5908 18921 5917 18955
rect 5917 18921 5951 18955
rect 5951 18921 5960 18955
rect 5908 18912 5960 18921
rect 6828 18912 6880 18964
rect 7840 18912 7892 18964
rect 8300 18912 8352 18964
rect 8576 18912 8628 18964
rect 9680 18955 9732 18964
rect 9680 18921 9689 18955
rect 9689 18921 9723 18955
rect 9723 18921 9732 18955
rect 9680 18912 9732 18921
rect 9036 18844 9088 18896
rect 10232 18844 10284 18896
rect 5908 18776 5960 18828
rect 1492 18640 1544 18692
rect 3608 18708 3660 18760
rect 4436 18751 4488 18760
rect 4436 18717 4445 18751
rect 4445 18717 4479 18751
rect 4479 18717 4488 18751
rect 4436 18708 4488 18717
rect 5816 18708 5868 18760
rect 6368 18708 6420 18760
rect 7104 18708 7156 18760
rect 9864 18776 9916 18828
rect 7564 18640 7616 18692
rect 9036 18708 9088 18760
rect 9680 18708 9732 18760
rect 9956 18708 10008 18760
rect 10232 18708 10284 18760
rect 2964 18572 3016 18624
rect 3700 18572 3752 18624
rect 4712 18572 4764 18624
rect 8760 18640 8812 18692
rect 9956 18572 10008 18624
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 3202 18470 3254 18522
rect 3266 18470 3318 18522
rect 9010 18470 9062 18522
rect 9074 18470 9126 18522
rect 9138 18470 9190 18522
rect 9202 18470 9254 18522
rect 9266 18470 9318 18522
rect 1308 18368 1360 18420
rect 6184 18368 6236 18420
rect 388 18300 440 18352
rect 664 18300 716 18352
rect 2780 18300 2832 18352
rect 204 18232 256 18284
rect 1308 18232 1360 18284
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 664 18164 716 18216
rect 1952 18232 2004 18284
rect 1768 18164 1820 18216
rect 1492 18096 1544 18148
rect 1676 18096 1728 18148
rect 204 18028 256 18080
rect 2412 18232 2464 18284
rect 6552 18232 6604 18284
rect 6644 18275 6696 18284
rect 6644 18241 6653 18275
rect 6653 18241 6687 18275
rect 6687 18241 6696 18275
rect 6644 18232 6696 18241
rect 7012 18232 7064 18284
rect 7380 18232 7432 18284
rect 7564 18207 7616 18216
rect 7564 18173 7573 18207
rect 7573 18173 7607 18207
rect 7607 18173 7616 18207
rect 7564 18164 7616 18173
rect 7748 18207 7800 18216
rect 7748 18173 7757 18207
rect 7757 18173 7791 18207
rect 7791 18173 7800 18207
rect 7748 18164 7800 18173
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 4436 18096 4488 18148
rect 6368 18096 6420 18148
rect 8116 18096 8168 18148
rect 8576 18207 8628 18216
rect 8576 18173 8610 18207
rect 8610 18173 8628 18207
rect 8576 18164 8628 18173
rect 2688 18028 2740 18080
rect 4804 18028 4856 18080
rect 5356 18028 5408 18080
rect 7288 18028 7340 18080
rect 7840 18028 7892 18080
rect 8852 18028 8904 18080
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 7950 17926 8002 17978
rect 8014 17926 8066 17978
rect 8078 17926 8130 17978
rect 8142 17926 8194 17978
rect 8206 17926 8258 17978
rect 1216 17824 1268 17876
rect 1676 17824 1728 17876
rect 2780 17824 2832 17876
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 6736 17867 6788 17876
rect 6736 17833 6745 17867
rect 6745 17833 6779 17867
rect 6779 17833 6788 17867
rect 6736 17824 6788 17833
rect 7564 17824 7616 17876
rect 9404 17824 9456 17876
rect 1216 17620 1268 17672
rect 8760 17756 8812 17808
rect 3424 17688 3476 17740
rect 6368 17688 6420 17740
rect 1768 17620 1820 17672
rect 1952 17620 2004 17672
rect 2228 17620 2280 17672
rect 6000 17620 6052 17672
rect 6460 17620 6512 17672
rect 3332 17552 3384 17604
rect 5172 17552 5224 17604
rect 1400 17484 1452 17536
rect 7656 17620 7708 17672
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 8300 17620 8352 17629
rect 8392 17620 8444 17672
rect 8852 17620 8904 17672
rect 9036 17688 9088 17740
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 9680 17620 9732 17672
rect 7012 17484 7064 17536
rect 7196 17484 7248 17536
rect 8392 17484 8444 17536
rect 940 17416 992 17468
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 3202 17382 3254 17434
rect 3266 17382 3318 17434
rect 9010 17382 9062 17434
rect 9074 17382 9126 17434
rect 9138 17382 9190 17434
rect 9202 17382 9254 17434
rect 9266 17382 9318 17434
rect 1492 17212 1544 17264
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 2964 17280 3016 17332
rect 3700 17280 3752 17332
rect 4344 17280 4396 17332
rect 5080 17280 5132 17332
rect 7564 17280 7616 17332
rect 8300 17280 8352 17332
rect 9496 17255 9548 17264
rect 9496 17221 9505 17255
rect 9505 17221 9539 17255
rect 9539 17221 9548 17255
rect 9496 17212 9548 17221
rect 9588 17212 9640 17264
rect 10968 17212 11020 17264
rect 940 17076 992 17128
rect 2504 17119 2556 17128
rect 2504 17085 2513 17119
rect 2513 17085 2547 17119
rect 2547 17085 2556 17119
rect 2504 17076 2556 17085
rect 7104 17144 7156 17196
rect 7748 17187 7800 17196
rect 7748 17153 7757 17187
rect 7757 17153 7791 17187
rect 7791 17153 7800 17187
rect 7748 17144 7800 17153
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 3608 17076 3660 17128
rect 2780 17008 2832 17060
rect 3240 17008 3292 17060
rect 7288 17076 7340 17128
rect 7840 17076 7892 17128
rect 5080 17008 5132 17060
rect 8116 17008 8168 17060
rect 8576 17119 8628 17128
rect 8576 17085 8610 17119
rect 8610 17085 8628 17119
rect 8576 17076 8628 17085
rect 7840 16940 7892 16992
rect 8576 16940 8628 16992
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 7950 16838 8002 16890
rect 8014 16838 8066 16890
rect 8078 16838 8130 16890
rect 8142 16838 8194 16890
rect 8206 16838 8258 16890
rect 2136 16736 2188 16788
rect 2412 16736 2464 16788
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 5080 16736 5132 16788
rect 10600 16736 10652 16788
rect 5724 16668 5776 16720
rect 6736 16668 6788 16720
rect 7564 16668 7616 16720
rect 8576 16668 8628 16720
rect 11060 16668 11112 16720
rect 1400 16600 1452 16652
rect 5540 16643 5592 16652
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 6184 16600 6236 16652
rect 296 16532 348 16584
rect 1124 16532 1176 16584
rect 1584 16532 1636 16584
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 6368 16532 6420 16584
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 9864 16532 9916 16584
rect 296 16396 348 16448
rect 4160 16396 4212 16448
rect 4988 16396 5040 16448
rect 6092 16396 6144 16448
rect 8116 16396 8168 16448
rect 9772 16464 9824 16516
rect 9312 16396 9364 16448
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 3202 16294 3254 16346
rect 3266 16294 3318 16346
rect 9010 16294 9062 16346
rect 9074 16294 9126 16346
rect 9138 16294 9190 16346
rect 9202 16294 9254 16346
rect 9266 16294 9318 16346
rect 2504 16192 2556 16244
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2504 16056 2556 16108
rect 3608 16099 3660 16108
rect 3608 16065 3617 16099
rect 3617 16065 3651 16099
rect 3651 16065 3660 16099
rect 3608 16056 3660 16065
rect 1676 15920 1728 15972
rect 2136 15920 2188 15972
rect 2044 15852 2096 15904
rect 2320 15852 2372 15904
rect 3332 16031 3384 16040
rect 3332 15997 3341 16031
rect 3341 15997 3375 16031
rect 3375 15997 3384 16031
rect 3332 15988 3384 15997
rect 4252 15988 4304 16040
rect 6000 16192 6052 16244
rect 8392 16192 8444 16244
rect 4436 15988 4488 16040
rect 4896 15988 4948 16040
rect 4988 16031 5040 16040
rect 4988 15997 4997 16031
rect 4997 15997 5031 16031
rect 5031 15997 5040 16031
rect 4988 15988 5040 15997
rect 5540 16099 5592 16108
rect 5540 16065 5549 16099
rect 5549 16065 5583 16099
rect 5583 16065 5592 16099
rect 5540 16056 5592 16065
rect 9680 16167 9732 16176
rect 9680 16133 9689 16167
rect 9689 16133 9723 16167
rect 9723 16133 9732 16167
rect 9680 16124 9732 16133
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8668 16056 8720 16108
rect 3056 15963 3108 15972
rect 3056 15929 3065 15963
rect 3065 15929 3099 15963
rect 3099 15929 3108 15963
rect 3056 15920 3108 15929
rect 4160 15852 4212 15904
rect 4344 15852 4396 15904
rect 4988 15852 5040 15904
rect 5724 15988 5776 16040
rect 6368 16031 6420 16040
rect 6368 15997 6377 16031
rect 6377 15997 6411 16031
rect 6411 15997 6420 16031
rect 6368 15988 6420 15997
rect 7196 15988 7248 16040
rect 7380 15988 7432 16040
rect 8116 15988 8168 16040
rect 8024 15920 8076 15972
rect 5540 15852 5592 15904
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 7950 15750 8002 15802
rect 8014 15750 8066 15802
rect 8078 15750 8130 15802
rect 8142 15750 8194 15802
rect 8206 15750 8258 15802
rect 3056 15691 3108 15700
rect 3056 15657 3065 15691
rect 3065 15657 3099 15691
rect 3099 15657 3108 15691
rect 3056 15648 3108 15657
rect 4068 15648 4120 15700
rect 1676 15512 1728 15564
rect 1952 15512 2004 15564
rect 2688 15512 2740 15564
rect 4252 15512 4304 15564
rect 5448 15648 5500 15700
rect 6736 15648 6788 15700
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 7380 15648 7432 15657
rect 7656 15648 7708 15700
rect 5724 15580 5776 15632
rect 11152 15648 11204 15700
rect 6000 15512 6052 15564
rect 6460 15512 6512 15564
rect 8852 15580 8904 15632
rect 9956 15580 10008 15632
rect 9772 15555 9824 15564
rect 9772 15521 9781 15555
rect 9781 15521 9815 15555
rect 9815 15521 9824 15555
rect 9772 15512 9824 15521
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 4344 15487 4396 15496
rect 4344 15453 4353 15487
rect 4353 15453 4387 15487
rect 4387 15453 4396 15487
rect 4344 15444 4396 15453
rect 4988 15444 5040 15496
rect 6184 15444 6236 15496
rect 5540 15376 5592 15428
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 8760 15487 8812 15496
rect 8760 15453 8769 15487
rect 8769 15453 8803 15487
rect 8803 15453 8812 15487
rect 8760 15444 8812 15453
rect 4436 15308 4488 15360
rect 7288 15308 7340 15360
rect 8852 15376 8904 15428
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 3202 15206 3254 15258
rect 3266 15206 3318 15258
rect 9010 15206 9062 15258
rect 9074 15206 9126 15258
rect 9138 15206 9190 15258
rect 9202 15206 9254 15258
rect 9266 15206 9318 15258
rect 3608 15104 3660 15156
rect 3792 15104 3844 15156
rect 4436 15104 4488 15156
rect 7656 15104 7708 15156
rect 7748 15104 7800 15156
rect 1492 15036 1544 15088
rect 1032 14968 1084 15020
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 7012 15036 7064 15088
rect 2688 14968 2740 15020
rect 5172 14968 5224 15020
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 8392 15011 8444 15020
rect 8392 14977 8410 15011
rect 8410 14977 8444 15011
rect 8392 14968 8444 14977
rect 9680 15079 9732 15088
rect 9680 15045 9689 15079
rect 9689 15045 9723 15079
rect 9723 15045 9732 15079
rect 9680 15036 9732 15045
rect 6368 14900 6420 14952
rect 7564 14900 7616 14952
rect 8668 14900 8720 14952
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 2412 14764 2464 14816
rect 2596 14764 2648 14816
rect 9496 14875 9548 14884
rect 9496 14841 9505 14875
rect 9505 14841 9539 14875
rect 9539 14841 9548 14875
rect 9496 14832 9548 14841
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 7950 14662 8002 14714
rect 8014 14662 8066 14714
rect 8078 14662 8130 14714
rect 8142 14662 8194 14714
rect 8206 14662 8258 14714
rect 1768 14424 1820 14476
rect 4252 14560 4304 14612
rect 6460 14560 6512 14612
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 9956 14560 10008 14612
rect 4344 14492 4396 14544
rect 4528 14492 4580 14544
rect 6920 14492 6972 14544
rect 7196 14424 7248 14476
rect 7656 14424 7708 14476
rect 9220 14424 9272 14476
rect 10048 14492 10100 14544
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 4528 14356 4580 14408
rect 1860 14288 1912 14340
rect 3884 14288 3936 14340
rect 5816 14356 5868 14408
rect 6552 14356 6604 14408
rect 5080 14288 5132 14340
rect 6828 14356 6880 14408
rect 7840 14399 7892 14408
rect 7840 14365 7849 14399
rect 7849 14365 7883 14399
rect 7883 14365 7892 14399
rect 7840 14356 7892 14365
rect 8024 14356 8076 14408
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 9404 14356 9456 14408
rect 10508 14356 10560 14408
rect 3516 14220 3568 14272
rect 5540 14220 5592 14272
rect 5816 14220 5868 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 3202 14118 3254 14170
rect 3266 14118 3318 14170
rect 9010 14118 9062 14170
rect 9074 14118 9126 14170
rect 9138 14118 9190 14170
rect 9202 14118 9254 14170
rect 9266 14118 9318 14170
rect 4068 14016 4120 14068
rect 4528 14016 4580 14068
rect 7196 14016 7248 14068
rect 8024 14016 8076 14068
rect 8208 14016 8260 14068
rect 8392 14016 8444 14068
rect 8668 14016 8720 14068
rect 1676 13948 1728 14000
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 2596 13880 2648 13932
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 4252 13812 4304 13864
rect 6736 13812 6788 13864
rect 7104 13812 7156 13864
rect 8208 13812 8260 13864
rect 8852 13812 8904 13864
rect 7840 13744 7892 13796
rect 3516 13676 3568 13728
rect 6736 13676 6788 13728
rect 7656 13676 7708 13728
rect 8392 13676 8444 13728
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 7950 13574 8002 13626
rect 8014 13574 8066 13626
rect 8078 13574 8130 13626
rect 8142 13574 8194 13626
rect 8206 13574 8258 13626
rect 3056 13472 3108 13524
rect 7656 13472 7708 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 1032 13404 1084 13456
rect 6828 13404 6880 13456
rect 7288 13404 7340 13456
rect 7932 13404 7984 13456
rect 8208 13404 8260 13456
rect 204 13336 256 13388
rect 4988 13336 5040 13388
rect 6000 13336 6052 13388
rect 1584 13268 1636 13320
rect 1768 13311 1820 13320
rect 1768 13277 1777 13311
rect 1777 13277 1811 13311
rect 1811 13277 1820 13311
rect 1768 13268 1820 13277
rect 6736 13311 6788 13320
rect 6736 13277 6754 13311
rect 6754 13277 6788 13311
rect 6736 13268 6788 13277
rect 9680 13472 9732 13524
rect 9220 13404 9272 13456
rect 9956 13404 10008 13456
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 9588 13336 9640 13388
rect 10508 13336 10560 13388
rect 572 13200 624 13252
rect 3608 13200 3660 13252
rect 3884 13200 3936 13252
rect 4344 13200 4396 13252
rect 5908 13200 5960 13252
rect 7656 13200 7708 13252
rect 8392 13200 8444 13252
rect 9220 13268 9272 13320
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 9404 13268 9456 13320
rect 9772 13268 9824 13320
rect 10968 13200 11020 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 4252 13132 4304 13184
rect 8668 13132 8720 13184
rect 9404 13175 9456 13184
rect 9404 13141 9413 13175
rect 9413 13141 9447 13175
rect 9447 13141 9456 13175
rect 9404 13132 9456 13141
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 3202 13030 3254 13082
rect 3266 13030 3318 13082
rect 9010 13030 9062 13082
rect 9074 13030 9126 13082
rect 9138 13030 9190 13082
rect 9202 13030 9254 13082
rect 9266 13030 9318 13082
rect 1492 12860 1544 12912
rect 1676 12860 1728 12912
rect 2504 12860 2556 12912
rect 1860 12792 1912 12844
rect 3516 12928 3568 12980
rect 3792 12928 3844 12980
rect 4712 12928 4764 12980
rect 5724 12928 5776 12980
rect 6736 12928 6788 12980
rect 6276 12860 6328 12912
rect 9404 12928 9456 12980
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 3056 12724 3108 12776
rect 4804 12792 4856 12844
rect 3884 12724 3936 12776
rect 5632 12724 5684 12776
rect 6460 12792 6512 12844
rect 6828 12835 6880 12844
rect 6828 12801 6837 12835
rect 6837 12801 6871 12835
rect 6871 12801 6880 12835
rect 6828 12792 6880 12801
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 4712 12656 4764 12708
rect 5172 12588 5224 12640
rect 6828 12656 6880 12708
rect 6736 12631 6788 12640
rect 6736 12597 6745 12631
rect 6745 12597 6779 12631
rect 6779 12597 6788 12631
rect 6736 12588 6788 12597
rect 7012 12724 7064 12776
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 9404 12792 9456 12844
rect 10324 12860 10376 12912
rect 10692 12792 10744 12844
rect 7932 12724 7984 12776
rect 8116 12724 8168 12776
rect 8944 12724 8996 12776
rect 7380 12656 7432 12708
rect 10600 12656 10652 12708
rect 10048 12588 10100 12640
rect 10784 12588 10836 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 7950 12486 8002 12538
rect 8014 12486 8066 12538
rect 8078 12486 8130 12538
rect 8142 12486 8194 12538
rect 8206 12486 8258 12538
rect 388 12384 440 12436
rect 1308 12384 1360 12436
rect 4712 12384 4764 12436
rect 5540 12384 5592 12436
rect 6184 12384 6236 12436
rect 6736 12384 6788 12436
rect 2504 12316 2556 12368
rect 5264 12316 5316 12368
rect 6644 12316 6696 12368
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 1676 12112 1728 12164
rect 2596 12180 2648 12232
rect 2228 12112 2280 12164
rect 2872 12248 2924 12300
rect 4712 12248 4764 12300
rect 5632 12291 5684 12300
rect 5632 12257 5641 12291
rect 5641 12257 5675 12291
rect 5675 12257 5684 12291
rect 5632 12248 5684 12257
rect 5724 12248 5776 12300
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 7656 12384 7708 12436
rect 8944 12384 8996 12436
rect 8208 12316 8260 12368
rect 9128 12316 9180 12368
rect 6184 12248 6236 12257
rect 3700 12180 3752 12232
rect 2872 12112 2924 12164
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 5356 12180 5408 12232
rect 6000 12223 6052 12232
rect 6000 12189 6034 12223
rect 6034 12189 6052 12223
rect 6000 12180 6052 12189
rect 6828 12180 6880 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 9864 12248 9916 12300
rect 5080 12112 5132 12164
rect 6736 12112 6788 12164
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 6460 12044 6512 12096
rect 6828 12044 6880 12096
rect 8944 12112 8996 12164
rect 9128 12112 9180 12164
rect 9404 12112 9456 12164
rect 9680 12112 9732 12164
rect 8668 12044 8720 12096
rect 10232 12044 10284 12096
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 3202 11942 3254 11994
rect 3266 11942 3318 11994
rect 9010 11942 9062 11994
rect 9074 11942 9126 11994
rect 9138 11942 9190 11994
rect 9202 11942 9254 11994
rect 9266 11942 9318 11994
rect 848 11772 900 11824
rect 1308 11704 1360 11756
rect 940 11636 992 11688
rect 1492 11636 1544 11688
rect 3516 11840 3568 11892
rect 4068 11840 4120 11892
rect 4252 11840 4304 11892
rect 5264 11840 5316 11892
rect 7472 11840 7524 11892
rect 8208 11840 8260 11892
rect 9404 11840 9456 11892
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 4068 11747 4120 11756
rect 4068 11713 4102 11747
rect 4102 11713 4120 11747
rect 4068 11704 4120 11713
rect 6460 11747 6512 11756
rect 6460 11713 6469 11747
rect 6469 11713 6503 11747
rect 6503 11713 6512 11747
rect 6460 11704 6512 11713
rect 7012 11704 7064 11756
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 10784 11704 10836 11756
rect 3056 11679 3108 11688
rect 3056 11645 3065 11679
rect 3065 11645 3099 11679
rect 3099 11645 3108 11679
rect 3056 11636 3108 11645
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 572 11568 624 11620
rect 1308 11568 1360 11620
rect 2872 11568 2924 11620
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 2228 11500 2280 11552
rect 2412 11500 2464 11552
rect 6276 11636 6328 11688
rect 7472 11636 7524 11688
rect 4896 11568 4948 11620
rect 5816 11568 5868 11620
rect 6552 11568 6604 11620
rect 8300 11636 8352 11688
rect 8576 11679 8628 11688
rect 8576 11645 8610 11679
rect 8610 11645 8628 11679
rect 8576 11636 8628 11645
rect 8944 11636 8996 11688
rect 9128 11636 9180 11688
rect 7932 11568 7984 11620
rect 4712 11500 4764 11552
rect 6736 11500 6788 11552
rect 6920 11500 6972 11552
rect 8668 11500 8720 11552
rect 9220 11500 9272 11552
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 7950 11398 8002 11450
rect 8014 11398 8066 11450
rect 8078 11398 8130 11450
rect 8142 11398 8194 11450
rect 8206 11398 8258 11450
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 3976 11296 4028 11348
rect 6828 11296 6880 11348
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 7380 11296 7432 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8852 11296 8904 11348
rect 848 11228 900 11280
rect 4160 11228 4212 11280
rect 4344 11228 4396 11280
rect 5632 11228 5684 11280
rect 10600 11296 10652 11348
rect 10232 11228 10284 11280
rect 940 11160 992 11212
rect 3240 11160 3292 11212
rect 5540 11160 5592 11212
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 2044 11092 2096 11144
rect 2412 11092 2464 11144
rect 4436 11092 4488 11144
rect 4896 11092 4948 11144
rect 5080 11092 5132 11144
rect 5816 11092 5868 11144
rect 6460 11135 6512 11144
rect 8852 11160 8904 11212
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 6460 11101 6494 11135
rect 6494 11101 6512 11135
rect 6460 11092 6512 11101
rect 1952 11024 2004 11076
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 9956 11092 10008 11144
rect 9864 11024 9916 11076
rect 940 10956 992 11008
rect 1400 10956 1452 11008
rect 6460 10956 6512 11008
rect 6920 10956 6972 11008
rect 7288 10956 7340 11008
rect 8576 10956 8628 11008
rect 8760 10956 8812 11008
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 3202 10854 3254 10906
rect 3266 10854 3318 10906
rect 9010 10854 9062 10906
rect 9074 10854 9126 10906
rect 9138 10854 9190 10906
rect 9202 10854 9254 10906
rect 9266 10854 9318 10906
rect 1952 10752 2004 10804
rect 5724 10752 5776 10804
rect 6828 10752 6880 10804
rect 7564 10795 7616 10804
rect 7564 10761 7573 10795
rect 7573 10761 7607 10795
rect 7607 10761 7616 10795
rect 7564 10752 7616 10761
rect 8300 10752 8352 10804
rect 1400 10616 1452 10668
rect 2872 10684 2924 10736
rect 3700 10684 3752 10736
rect 5080 10684 5132 10736
rect 2412 10616 2464 10668
rect 2504 10412 2556 10464
rect 6000 10616 6052 10668
rect 6736 10616 6788 10668
rect 4896 10548 4948 10600
rect 5816 10548 5868 10600
rect 6368 10548 6420 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 7380 10616 7432 10668
rect 8668 10659 8720 10668
rect 8668 10625 8702 10659
rect 8702 10625 8720 10659
rect 8668 10616 8720 10625
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 7564 10548 7616 10600
rect 5448 10480 5500 10532
rect 8300 10523 8352 10532
rect 8300 10489 8309 10523
rect 8309 10489 8343 10523
rect 8343 10489 8352 10523
rect 8300 10480 8352 10489
rect 2872 10412 2924 10464
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9496 10548 9548 10600
rect 9496 10412 9548 10464
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 7950 10310 8002 10362
rect 8014 10310 8066 10362
rect 8078 10310 8130 10362
rect 8142 10310 8194 10362
rect 8206 10310 8258 10362
rect 1492 10208 1544 10260
rect 4068 10208 4120 10260
rect 4988 10208 5040 10260
rect 6184 10208 6236 10260
rect 8852 10208 8904 10260
rect 5080 10140 5132 10192
rect 2504 10072 2556 10124
rect 5264 10140 5316 10192
rect 8484 10183 8536 10192
rect 8484 10149 8493 10183
rect 8493 10149 8527 10183
rect 8527 10149 8536 10183
rect 8484 10140 8536 10149
rect 1032 10004 1084 10056
rect 1952 10004 2004 10056
rect 6460 10115 6512 10124
rect 6460 10081 6469 10115
rect 6469 10081 6503 10115
rect 6503 10081 6512 10115
rect 6460 10072 6512 10081
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 7472 10072 7524 10124
rect 8208 10072 8260 10124
rect 2780 10004 2832 10056
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4712 10004 4764 10056
rect 5816 10004 5868 10056
rect 7012 10004 7064 10056
rect 9680 10072 9732 10124
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 4896 9936 4948 9988
rect 4988 9936 5040 9988
rect 7288 9936 7340 9988
rect 8116 9936 8168 9988
rect 10048 9936 10100 9988
rect 6368 9911 6420 9920
rect 6368 9877 6377 9911
rect 6377 9877 6411 9911
rect 6411 9877 6420 9911
rect 6368 9868 6420 9877
rect 8024 9868 8076 9920
rect 9496 9868 9548 9920
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 3202 9766 3254 9818
rect 3266 9766 3318 9818
rect 9010 9766 9062 9818
rect 9074 9766 9126 9818
rect 9138 9766 9190 9818
rect 9202 9766 9254 9818
rect 9266 9766 9318 9818
rect 480 9664 532 9716
rect 3884 9664 3936 9716
rect 4712 9707 4764 9716
rect 4712 9673 4721 9707
rect 4721 9673 4755 9707
rect 4755 9673 4764 9707
rect 4712 9664 4764 9673
rect 5448 9664 5500 9716
rect 5632 9664 5684 9716
rect 8116 9664 8168 9716
rect 8300 9707 8352 9716
rect 8300 9673 8309 9707
rect 8309 9673 8343 9707
rect 8343 9673 8352 9707
rect 8300 9664 8352 9673
rect 8576 9664 8628 9716
rect 10876 9664 10928 9716
rect 3700 9596 3752 9648
rect 4804 9596 4856 9648
rect 5816 9596 5868 9648
rect 2504 9528 2556 9580
rect 3424 9528 3476 9580
rect 4988 9571 5040 9580
rect 4988 9537 4997 9571
rect 4997 9537 5031 9571
rect 5031 9537 5040 9571
rect 4988 9528 5040 9537
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 5356 9460 5408 9512
rect 5816 9460 5868 9512
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 4620 9324 4672 9376
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 5080 9392 5132 9444
rect 5448 9392 5500 9444
rect 6460 9528 6512 9580
rect 8760 9596 8812 9648
rect 7472 9528 7524 9580
rect 8392 9528 8444 9580
rect 6828 9460 6880 9512
rect 6092 9392 6144 9444
rect 5264 9324 5316 9376
rect 6276 9324 6328 9376
rect 6920 9324 6972 9376
rect 7380 9324 7432 9376
rect 9772 9503 9824 9512
rect 9772 9469 9781 9503
rect 9781 9469 9815 9503
rect 9815 9469 9824 9503
rect 9772 9460 9824 9469
rect 9496 9324 9548 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 7950 9222 8002 9274
rect 8014 9222 8066 9274
rect 8078 9222 8130 9274
rect 8142 9222 8194 9274
rect 8206 9222 8258 9274
rect 1952 9120 2004 9172
rect 2412 9120 2464 9172
rect 5816 9120 5868 9172
rect 6460 9120 6512 9172
rect 6920 9052 6972 9104
rect 8484 9052 8536 9104
rect 8852 9052 8904 9104
rect 9312 9052 9364 9104
rect 4804 8916 4856 8968
rect 9864 8984 9916 9036
rect 8392 8916 8444 8968
rect 9404 8916 9456 8968
rect 9588 8916 9640 8968
rect 8852 8848 8904 8900
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 848 8780 900 8832
rect 2228 8780 2280 8832
rect 2504 8780 2556 8832
rect 6552 8780 6604 8832
rect 7012 8780 7064 8832
rect 7564 8780 7616 8832
rect 8208 8780 8260 8832
rect 8760 8780 8812 8832
rect 9404 8780 9456 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 1216 8576 1268 8628
rect 8208 8576 8260 8628
rect 1676 8508 1728 8560
rect 1860 8551 1912 8560
rect 1860 8517 1869 8551
rect 1869 8517 1903 8551
rect 1903 8517 1912 8551
rect 1860 8508 1912 8517
rect 8852 8576 8904 8628
rect 3424 8440 3476 8492
rect 4068 8440 4120 8492
rect 5816 8440 5868 8492
rect 6368 8440 6420 8492
rect 296 8372 348 8424
rect 2228 8372 2280 8424
rect 4712 8372 4764 8424
rect 7012 8372 7064 8424
rect 7380 8372 7432 8424
rect 4068 8304 4120 8356
rect 5724 8304 5776 8356
rect 4160 8236 4212 8288
rect 5540 8236 5592 8288
rect 7564 8236 7616 8288
rect 8208 8372 8260 8424
rect 8484 8372 8536 8424
rect 8668 8372 8720 8424
rect 8852 8304 8904 8356
rect 8484 8236 8536 8288
rect 9220 8236 9272 8288
rect 9404 8236 9456 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 6368 8032 6420 8084
rect 6920 8075 6972 8084
rect 6920 8041 6929 8075
rect 6929 8041 6963 8075
rect 6963 8041 6972 8075
rect 6920 8032 6972 8041
rect 8668 8032 8720 8084
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 9404 8032 9456 8084
rect 10232 8032 10284 8084
rect 4804 7964 4856 8016
rect 2228 7896 2280 7948
rect 2504 7896 2556 7948
rect 5264 7964 5316 8016
rect 5724 8007 5776 8016
rect 5724 7973 5733 8007
rect 5733 7973 5767 8007
rect 5767 7973 5776 8007
rect 5724 7964 5776 7973
rect 7748 8007 7800 8016
rect 7748 7973 7757 8007
rect 7757 7973 7791 8007
rect 7791 7973 7800 8007
rect 7748 7964 7800 7973
rect 1676 7828 1728 7880
rect 5356 7896 5408 7948
rect 5632 7896 5684 7948
rect 6092 7939 6144 7948
rect 6092 7905 6126 7939
rect 6126 7905 6144 7939
rect 6092 7896 6144 7905
rect 2228 7760 2280 7812
rect 2320 7760 2372 7812
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 9864 7964 9916 8016
rect 9680 7896 9732 7948
rect 8760 7828 8812 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9404 7828 9456 7880
rect 9496 7871 9548 7880
rect 9496 7837 9505 7871
rect 9505 7837 9539 7871
rect 9539 7837 9548 7871
rect 9496 7828 9548 7837
rect 10968 7828 11020 7880
rect 7288 7760 7340 7812
rect 9956 7760 10008 7812
rect 4804 7692 4856 7744
rect 5080 7692 5132 7744
rect 6276 7692 6328 7744
rect 7564 7692 7616 7744
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 2320 7463 2372 7472
rect 2320 7429 2329 7463
rect 2329 7429 2363 7463
rect 2363 7429 2372 7463
rect 2320 7420 2372 7429
rect 2688 7420 2740 7472
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 2228 7284 2280 7336
rect 4712 7284 4764 7336
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 20 7148 72 7200
rect 2688 7148 2740 7200
rect 3976 7216 4028 7268
rect 4620 7216 4672 7268
rect 5264 7284 5316 7336
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 7196 7488 7248 7540
rect 7656 7488 7708 7540
rect 6644 7352 6696 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 9680 7488 9732 7540
rect 8484 7463 8536 7472
rect 8484 7429 8493 7463
rect 8493 7429 8527 7463
rect 8527 7429 8536 7463
rect 8484 7420 8536 7429
rect 8576 7420 8628 7472
rect 9956 7420 10008 7472
rect 8208 7352 8260 7404
rect 8668 7352 8720 7404
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9404 7352 9456 7404
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 6828 7216 6880 7268
rect 5356 7148 5408 7200
rect 8760 7284 8812 7336
rect 7288 7216 7340 7268
rect 7472 7216 7524 7268
rect 7656 7216 7708 7268
rect 9220 7327 9272 7336
rect 9220 7293 9225 7327
rect 9225 7293 9259 7327
rect 9259 7293 9272 7327
rect 9220 7284 9272 7293
rect 9496 7216 9548 7268
rect 7840 7148 7892 7200
rect 8576 7191 8628 7200
rect 8576 7157 8585 7191
rect 8585 7157 8619 7191
rect 8619 7157 8628 7191
rect 8576 7148 8628 7157
rect 8852 7148 8904 7200
rect 9220 7148 9272 7200
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 4436 6808 4488 6860
rect 5356 6944 5408 6996
rect 5448 6944 5500 6996
rect 6000 6944 6052 6996
rect 6644 6944 6696 6996
rect 8852 6944 8904 6996
rect 7380 6876 7432 6928
rect 7656 6876 7708 6928
rect 5540 6808 5592 6860
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 5724 6808 5776 6860
rect 6000 6851 6052 6860
rect 6000 6817 6034 6851
rect 6034 6817 6052 6851
rect 6000 6808 6052 6817
rect 6368 6808 6420 6860
rect 1860 6740 1912 6792
rect 2596 6740 2648 6792
rect 1676 6604 1728 6656
rect 4068 6604 4120 6656
rect 5632 6604 5684 6656
rect 5724 6604 5776 6656
rect 7840 6808 7892 6860
rect 9312 6808 9364 6860
rect 10692 6876 10744 6928
rect 8208 6740 8260 6792
rect 8484 6740 8536 6792
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 9680 6672 9732 6724
rect 7104 6604 7156 6656
rect 7564 6604 7616 6656
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 8760 6604 8812 6656
rect 10324 6604 10376 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 1308 6400 1360 6452
rect 1676 6400 1728 6452
rect 2872 6400 2924 6452
rect 4068 6400 4120 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 5724 6332 5776 6384
rect 3516 6264 3568 6316
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 7472 6400 7524 6452
rect 8852 6400 8904 6452
rect 6552 6264 6604 6316
rect 6736 6264 6788 6316
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 3056 6060 3108 6112
rect 4068 6239 4120 6248
rect 4068 6205 4077 6239
rect 4077 6205 4111 6239
rect 4111 6205 4120 6239
rect 4068 6196 4120 6205
rect 6092 6128 6144 6180
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 5448 6060 5500 6112
rect 7748 6264 7800 6316
rect 10508 6332 10560 6384
rect 8852 6307 8904 6316
rect 8852 6273 8860 6307
rect 8860 6273 8904 6307
rect 8852 6264 8904 6273
rect 7380 6128 7432 6180
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 8668 6128 8720 6180
rect 7840 6060 7892 6112
rect 10048 6060 10100 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 2596 5856 2648 5908
rect 3056 5856 3108 5908
rect 4160 5856 4212 5908
rect 5448 5856 5500 5908
rect 6552 5856 6604 5908
rect 5724 5831 5776 5840
rect 5724 5797 5733 5831
rect 5733 5797 5767 5831
rect 5767 5797 5776 5831
rect 5724 5788 5776 5797
rect 6460 5831 6512 5840
rect 6460 5797 6469 5831
rect 6469 5797 6503 5831
rect 6503 5797 6512 5831
rect 6460 5788 6512 5797
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 7380 5720 7432 5772
rect 8392 5856 8444 5908
rect 9588 5856 9640 5908
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 4988 5652 5040 5704
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6736 5584 6788 5636
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 5908 5516 5960 5568
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 8484 5355 8536 5364
rect 8484 5321 8493 5355
rect 8493 5321 8527 5355
rect 8527 5321 8536 5355
rect 8484 5312 8536 5321
rect 9404 5312 9456 5364
rect 2872 5244 2924 5296
rect 7288 5244 7340 5296
rect 2780 5176 2832 5228
rect 3792 5176 3844 5228
rect 5908 5176 5960 5228
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6092 5176 6144 5185
rect 7380 5176 7432 5228
rect 9680 5176 9732 5228
rect 10692 5176 10744 5228
rect 4344 5040 4396 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 3424 4972 3476 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 4252 4700 4304 4752
rect 1032 4632 1084 4684
rect 5908 4564 5960 4616
rect 1492 4539 1544 4548
rect 1492 4505 1501 4539
rect 1501 4505 1535 4539
rect 1535 4505 1544 4539
rect 1492 4496 1544 4505
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 756 4224 808 4276
rect 4160 4224 4212 4276
rect 1124 4156 1176 4208
rect 1860 4156 1912 4208
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 3608 2592 3660 2644
rect 3884 2592 3936 2644
rect 5540 2592 5592 2644
rect 664 2524 716 2576
rect 2780 2524 2832 2576
rect 2320 2388 2372 2440
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 2688 2048 2740 2100
rect 3240 2048 3292 2100
<< metal2 >>
rect 938 44944 994 45000
rect 1398 44944 1454 45000
rect 1858 44944 1914 45000
rect 2318 44944 2374 45000
rect 2778 44944 2834 45000
rect 3238 44944 3294 45000
rect 3698 44944 3754 45000
rect 4158 44944 4214 45000
rect 4618 44944 4674 45000
rect 5078 44944 5134 45000
rect 5538 44944 5594 45000
rect 5998 44944 6054 45000
rect 6458 44944 6514 45000
rect 6918 44944 6974 45000
rect 7378 44944 7434 45000
rect 7838 44944 7894 45000
rect 8298 44944 8354 45000
rect 8758 44944 8814 45000
rect 9218 44944 9274 45000
rect 9678 44944 9734 45000
rect 10138 44944 10194 45000
rect 952 43314 980 44944
rect 1412 43466 1440 44944
rect 1412 43438 1532 43466
rect 940 43308 992 43314
rect 940 43250 992 43256
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1124 42220 1176 42226
rect 1124 42162 1176 42168
rect 1136 41414 1164 42162
rect 1412 41818 1440 43250
rect 1504 42362 1532 43438
rect 1872 42362 1900 44944
rect 2332 42362 2360 44944
rect 2792 42362 2820 44944
rect 3252 43466 3280 44944
rect 3252 43438 3464 43466
rect 3010 42460 3318 42469
rect 3010 42458 3016 42460
rect 3072 42458 3096 42460
rect 3152 42458 3176 42460
rect 3232 42458 3256 42460
rect 3312 42458 3318 42460
rect 3072 42406 3074 42458
rect 3254 42406 3256 42458
rect 3010 42404 3016 42406
rect 3072 42404 3096 42406
rect 3152 42404 3176 42406
rect 3232 42404 3256 42406
rect 3312 42404 3318 42406
rect 3010 42395 3318 42404
rect 3436 42362 3464 43438
rect 3712 42362 3740 44944
rect 4172 42362 4200 44944
rect 4632 42362 4660 44944
rect 5092 42362 5120 44944
rect 5552 42362 5580 44944
rect 6012 42362 6040 44944
rect 6472 42362 6500 44944
rect 6736 42560 6788 42566
rect 6736 42502 6788 42508
rect 1492 42356 1544 42362
rect 1492 42298 1544 42304
rect 1860 42356 1912 42362
rect 1860 42298 1912 42304
rect 2320 42356 2372 42362
rect 2320 42298 2372 42304
rect 2780 42356 2832 42362
rect 2780 42298 2832 42304
rect 3424 42356 3476 42362
rect 3424 42298 3476 42304
rect 3700 42356 3752 42362
rect 3700 42298 3752 42304
rect 4160 42356 4212 42362
rect 4160 42298 4212 42304
rect 4620 42356 4672 42362
rect 4620 42298 4672 42304
rect 5080 42356 5132 42362
rect 5080 42298 5132 42304
rect 5540 42356 5592 42362
rect 5540 42298 5592 42304
rect 6000 42356 6052 42362
rect 6000 42298 6052 42304
rect 6460 42356 6512 42362
rect 6460 42298 6512 42304
rect 3976 42288 4028 42294
rect 3976 42230 4028 42236
rect 2320 42220 2372 42226
rect 2320 42162 2372 42168
rect 1950 41916 2258 41925
rect 1950 41914 1956 41916
rect 2012 41914 2036 41916
rect 2092 41914 2116 41916
rect 2172 41914 2196 41916
rect 2252 41914 2258 41916
rect 2012 41862 2014 41914
rect 2194 41862 2196 41914
rect 1950 41860 1956 41862
rect 2012 41860 2036 41862
rect 2092 41860 2116 41862
rect 2172 41860 2196 41862
rect 2252 41860 2258 41862
rect 1950 41851 2258 41860
rect 1400 41812 1452 41818
rect 1400 41754 1452 41760
rect 1136 41386 1348 41414
rect 848 41064 900 41070
rect 848 41006 900 41012
rect 572 40112 624 40118
rect 572 40054 624 40060
rect 480 38004 532 38010
rect 480 37946 532 37952
rect 204 37460 256 37466
rect 204 37402 256 37408
rect 20 34196 72 34202
rect 20 34138 72 34144
rect 32 30138 60 34138
rect 216 31793 244 37402
rect 296 36032 348 36038
rect 296 35974 348 35980
rect 202 31784 258 31793
rect 202 31719 258 31728
rect 32 30110 244 30138
rect 112 30048 164 30054
rect 112 29990 164 29996
rect 18 28112 74 28121
rect 18 28047 74 28056
rect 32 23338 60 28047
rect 124 23458 152 29990
rect 216 26042 244 30110
rect 204 26036 256 26042
rect 204 25978 256 25984
rect 202 25800 258 25809
rect 202 25735 258 25744
rect 112 23452 164 23458
rect 112 23394 164 23400
rect 32 23310 152 23338
rect 18 23216 74 23225
rect 18 23151 74 23160
rect 32 7206 60 23151
rect 124 18170 152 23310
rect 216 22030 244 25735
rect 308 25498 336 35974
rect 388 34604 440 34610
rect 388 34546 440 34552
rect 400 33561 428 34546
rect 386 33552 442 33561
rect 386 33487 442 33496
rect 492 33436 520 37946
rect 400 33408 520 33436
rect 400 31754 428 33408
rect 400 31726 520 31754
rect 388 29164 440 29170
rect 388 29106 440 29112
rect 400 28665 428 29106
rect 386 28656 442 28665
rect 386 28591 442 28600
rect 388 28484 440 28490
rect 388 28426 440 28432
rect 296 25492 348 25498
rect 296 25434 348 25440
rect 400 25242 428 28426
rect 308 25214 428 25242
rect 204 22024 256 22030
rect 204 21966 256 21972
rect 308 18578 336 25214
rect 386 24984 442 24993
rect 386 24919 442 24928
rect 216 18550 336 18578
rect 216 18290 244 18550
rect 400 18442 428 24919
rect 492 23254 520 31726
rect 480 23248 532 23254
rect 480 23190 532 23196
rect 584 22094 612 40054
rect 756 38956 808 38962
rect 756 38898 808 38904
rect 768 38457 796 38898
rect 754 38448 810 38457
rect 754 38383 810 38392
rect 756 33516 808 33522
rect 756 33458 808 33464
rect 664 32768 716 32774
rect 768 32745 796 33458
rect 664 32710 716 32716
rect 754 32736 810 32745
rect 676 29306 704 32710
rect 754 32671 810 32680
rect 860 32586 888 41006
rect 1216 36236 1268 36242
rect 1216 36178 1268 36184
rect 1124 36168 1176 36174
rect 1124 36110 1176 36116
rect 1136 35154 1164 36110
rect 1124 35148 1176 35154
rect 1124 35090 1176 35096
rect 1122 35048 1178 35057
rect 1122 34983 1178 34992
rect 1032 34740 1084 34746
rect 1032 34682 1084 34688
rect 940 34672 992 34678
rect 940 34614 992 34620
rect 952 34377 980 34614
rect 938 34368 994 34377
rect 938 34303 994 34312
rect 768 32558 888 32586
rect 664 29300 716 29306
rect 664 29242 716 29248
rect 662 29064 718 29073
rect 662 28999 718 29008
rect 676 26489 704 28999
rect 662 26480 718 26489
rect 662 26415 718 26424
rect 664 26376 716 26382
rect 664 26318 716 26324
rect 676 26217 704 26318
rect 662 26208 718 26217
rect 662 26143 718 26152
rect 664 24744 716 24750
rect 664 24686 716 24692
rect 308 18414 428 18442
rect 492 22066 612 22094
rect 204 18284 256 18290
rect 204 18226 256 18232
rect 202 18184 258 18193
rect 124 18142 202 18170
rect 202 18119 258 18128
rect 204 18080 256 18086
rect 204 18022 256 18028
rect 216 13394 244 18022
rect 308 16590 336 18414
rect 388 18352 440 18358
rect 388 18294 440 18300
rect 296 16584 348 16590
rect 296 16526 348 16532
rect 296 16448 348 16454
rect 296 16390 348 16396
rect 204 13388 256 13394
rect 204 13330 256 13336
rect 308 8430 336 16390
rect 400 12442 428 18294
rect 388 12436 440 12442
rect 388 12378 440 12384
rect 492 9722 520 22066
rect 572 22024 624 22030
rect 572 21966 624 21972
rect 584 17082 612 21966
rect 676 18358 704 24686
rect 664 18352 716 18358
rect 664 18294 716 18300
rect 664 18216 716 18222
rect 664 18158 716 18164
rect 676 17241 704 18158
rect 662 17232 718 17241
rect 662 17167 718 17176
rect 584 17054 704 17082
rect 572 13252 624 13258
rect 572 13194 624 13200
rect 584 11626 612 13194
rect 572 11620 624 11626
rect 572 11562 624 11568
rect 480 9716 532 9722
rect 480 9658 532 9664
rect 296 8424 348 8430
rect 296 8366 348 8372
rect 20 7200 72 7206
rect 20 7142 72 7148
rect 676 2582 704 17054
rect 768 4282 796 32558
rect 940 31884 992 31890
rect 940 31826 992 31832
rect 848 31816 900 31822
rect 848 31758 900 31764
rect 860 31113 888 31758
rect 846 31104 902 31113
rect 846 31039 902 31048
rect 846 30016 902 30025
rect 846 29951 902 29960
rect 860 29073 888 29951
rect 846 29064 902 29073
rect 846 28999 902 29008
rect 848 27328 900 27334
rect 848 27270 900 27276
rect 860 21026 888 27270
rect 952 21162 980 31826
rect 1044 21350 1072 34682
rect 1136 34134 1164 34983
rect 1124 34128 1176 34134
rect 1124 34070 1176 34076
rect 1228 33590 1256 36178
rect 1320 34490 1348 41386
rect 1492 41132 1544 41138
rect 1492 41074 1544 41080
rect 1504 40905 1532 41074
rect 1860 40996 1912 41002
rect 1860 40938 1912 40944
rect 1490 40896 1546 40905
rect 1490 40831 1546 40840
rect 1492 40452 1544 40458
rect 1492 40394 1544 40400
rect 1768 40452 1820 40458
rect 1768 40394 1820 40400
rect 1504 40089 1532 40394
rect 1490 40080 1546 40089
rect 1490 40015 1546 40024
rect 1492 39364 1544 39370
rect 1492 39306 1544 39312
rect 1504 39273 1532 39306
rect 1490 39264 1546 39273
rect 1490 39199 1546 39208
rect 1584 38344 1636 38350
rect 1584 38286 1636 38292
rect 1492 38276 1544 38282
rect 1492 38218 1544 38224
rect 1504 37641 1532 38218
rect 1596 37874 1624 38286
rect 1780 37874 1808 40394
rect 1872 38282 1900 40938
rect 1950 40828 2258 40837
rect 1950 40826 1956 40828
rect 2012 40826 2036 40828
rect 2092 40826 2116 40828
rect 2172 40826 2196 40828
rect 2252 40826 2258 40828
rect 2012 40774 2014 40826
rect 2194 40774 2196 40826
rect 1950 40772 1956 40774
rect 2012 40772 2036 40774
rect 2092 40772 2116 40774
rect 2172 40772 2196 40774
rect 2252 40772 2258 40774
rect 1950 40763 2258 40772
rect 1950 39740 2258 39749
rect 1950 39738 1956 39740
rect 2012 39738 2036 39740
rect 2092 39738 2116 39740
rect 2172 39738 2196 39740
rect 2252 39738 2258 39740
rect 2012 39686 2014 39738
rect 2194 39686 2196 39738
rect 1950 39684 1956 39686
rect 2012 39684 2036 39686
rect 2092 39684 2116 39686
rect 2172 39684 2196 39686
rect 2252 39684 2258 39686
rect 1950 39675 2258 39684
rect 1950 38652 2258 38661
rect 1950 38650 1956 38652
rect 2012 38650 2036 38652
rect 2092 38650 2116 38652
rect 2172 38650 2196 38652
rect 2252 38650 2258 38652
rect 2012 38598 2014 38650
rect 2194 38598 2196 38650
rect 1950 38596 1956 38598
rect 2012 38596 2036 38598
rect 2092 38596 2116 38598
rect 2172 38596 2196 38598
rect 2252 38596 2258 38598
rect 1950 38587 2258 38596
rect 1860 38276 1912 38282
rect 1860 38218 1912 38224
rect 1584 37868 1636 37874
rect 1584 37810 1636 37816
rect 1768 37868 1820 37874
rect 1768 37810 1820 37816
rect 1490 37632 1546 37641
rect 1490 37567 1546 37576
rect 1596 37194 1624 37810
rect 1676 37256 1728 37262
rect 1780 37244 1808 37810
rect 1872 37346 1900 38218
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 1872 37318 2084 37346
rect 1860 37256 1912 37262
rect 1780 37216 1860 37244
rect 1676 37198 1728 37204
rect 1860 37198 1912 37204
rect 1492 37188 1544 37194
rect 1492 37130 1544 37136
rect 1584 37188 1636 37194
rect 1584 37130 1636 37136
rect 1504 36825 1532 37130
rect 1596 36922 1624 37130
rect 1584 36916 1636 36922
rect 1584 36858 1636 36864
rect 1490 36816 1546 36825
rect 1490 36751 1546 36760
rect 1596 36666 1624 36858
rect 1688 36825 1716 37198
rect 1768 36848 1820 36854
rect 1674 36816 1730 36825
rect 1768 36790 1820 36796
rect 1674 36751 1730 36760
rect 1504 36638 1624 36666
rect 1676 36712 1728 36718
rect 1676 36654 1728 36660
rect 1504 36242 1532 36638
rect 1584 36576 1636 36582
rect 1584 36518 1636 36524
rect 1492 36236 1544 36242
rect 1492 36178 1544 36184
rect 1492 36100 1544 36106
rect 1492 36042 1544 36048
rect 1504 36009 1532 36042
rect 1490 36000 1546 36009
rect 1490 35935 1546 35944
rect 1492 35692 1544 35698
rect 1492 35634 1544 35640
rect 1504 35193 1532 35634
rect 1490 35184 1546 35193
rect 1490 35119 1546 35128
rect 1320 34462 1440 34490
rect 1308 34400 1360 34406
rect 1308 34342 1360 34348
rect 1216 33584 1268 33590
rect 1216 33526 1268 33532
rect 1124 33380 1176 33386
rect 1124 33322 1176 33328
rect 1136 26897 1164 33322
rect 1228 32858 1256 33526
rect 1320 32978 1348 34342
rect 1308 32972 1360 32978
rect 1308 32914 1360 32920
rect 1228 32830 1348 32858
rect 1216 32224 1268 32230
rect 1216 32166 1268 32172
rect 1228 28694 1256 32166
rect 1320 31346 1348 32830
rect 1308 31340 1360 31346
rect 1308 31282 1360 31288
rect 1306 30288 1362 30297
rect 1306 30223 1362 30232
rect 1216 28688 1268 28694
rect 1216 28630 1268 28636
rect 1216 27668 1268 27674
rect 1216 27610 1268 27616
rect 1122 26888 1178 26897
rect 1122 26823 1178 26832
rect 1122 26344 1178 26353
rect 1122 26279 1178 26288
rect 1032 21344 1084 21350
rect 1032 21286 1084 21292
rect 952 21134 1072 21162
rect 860 20998 980 21026
rect 848 20868 900 20874
rect 848 20810 900 20816
rect 860 20505 888 20810
rect 846 20496 902 20505
rect 846 20431 902 20440
rect 952 17474 980 20998
rect 940 17468 992 17474
rect 940 17410 992 17416
rect 1044 17218 1072 21134
rect 860 17190 1072 17218
rect 860 11830 888 17190
rect 940 17128 992 17134
rect 1136 17082 1164 26279
rect 1228 17882 1256 27610
rect 1320 18426 1348 30223
rect 1412 29782 1440 34462
rect 1596 33454 1624 36518
rect 1688 36242 1716 36654
rect 1676 36236 1728 36242
rect 1676 36178 1728 36184
rect 1676 36100 1728 36106
rect 1676 36042 1728 36048
rect 1688 35601 1716 36042
rect 1780 35698 1808 36790
rect 1872 36009 1900 37198
rect 2056 37194 2084 37318
rect 2332 37210 2360 42162
rect 2412 42084 2464 42090
rect 2412 42026 2464 42032
rect 2044 37188 2096 37194
rect 2044 37130 2096 37136
rect 2240 37182 2360 37210
rect 2056 36582 2084 37130
rect 2240 37126 2268 37182
rect 2228 37120 2280 37126
rect 2228 37062 2280 37068
rect 2044 36576 2096 36582
rect 2044 36518 2096 36524
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 2320 36168 2372 36174
rect 2320 36110 2372 36116
rect 1858 36000 1914 36009
rect 1858 35935 1914 35944
rect 2332 35698 2360 36110
rect 1768 35692 1820 35698
rect 1768 35634 1820 35640
rect 2320 35692 2372 35698
rect 2320 35634 2372 35640
rect 1674 35592 1730 35601
rect 1674 35527 1730 35536
rect 1676 35148 1728 35154
rect 1676 35090 1728 35096
rect 1584 33448 1636 33454
rect 1584 33390 1636 33396
rect 1688 33386 1716 35090
rect 1780 34762 1808 35634
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 2332 35170 2360 35634
rect 2424 35290 2452 42026
rect 3792 41472 3844 41478
rect 3792 41414 3844 41420
rect 3010 41372 3318 41381
rect 3010 41370 3016 41372
rect 3072 41370 3096 41372
rect 3152 41370 3176 41372
rect 3232 41370 3256 41372
rect 3312 41370 3318 41372
rect 3072 41318 3074 41370
rect 3254 41318 3256 41370
rect 3010 41316 3016 41318
rect 3072 41316 3096 41318
rect 3152 41316 3176 41318
rect 3232 41316 3256 41318
rect 3312 41316 3318 41318
rect 3010 41307 3318 41316
rect 3010 40284 3318 40293
rect 3010 40282 3016 40284
rect 3072 40282 3096 40284
rect 3152 40282 3176 40284
rect 3232 40282 3256 40284
rect 3312 40282 3318 40284
rect 3072 40230 3074 40282
rect 3254 40230 3256 40282
rect 3010 40228 3016 40230
rect 3072 40228 3096 40230
rect 3152 40228 3176 40230
rect 3232 40228 3256 40230
rect 3312 40228 3318 40230
rect 3010 40219 3318 40228
rect 3700 39500 3752 39506
rect 3700 39442 3752 39448
rect 2780 39364 2832 39370
rect 2780 39306 2832 39312
rect 2596 38820 2648 38826
rect 2596 38762 2648 38768
rect 2504 38344 2556 38350
rect 2504 38286 2556 38292
rect 2516 37806 2544 38286
rect 2504 37800 2556 37806
rect 2504 37742 2556 37748
rect 2516 35698 2544 37742
rect 2504 35692 2556 35698
rect 2504 35634 2556 35640
rect 2412 35284 2464 35290
rect 2412 35226 2464 35232
rect 2332 35142 2544 35170
rect 1952 35012 2004 35018
rect 1952 34954 2004 34960
rect 1780 34734 1900 34762
rect 1768 34468 1820 34474
rect 1768 34410 1820 34416
rect 1780 33862 1808 34410
rect 1768 33856 1820 33862
rect 1768 33798 1820 33804
rect 1676 33380 1728 33386
rect 1676 33322 1728 33328
rect 1780 33266 1808 33798
rect 1688 33238 1808 33266
rect 1584 32972 1636 32978
rect 1584 32914 1636 32920
rect 1492 32428 1544 32434
rect 1492 32370 1544 32376
rect 1504 31929 1532 32370
rect 1490 31920 1546 31929
rect 1490 31855 1546 31864
rect 1492 31476 1544 31482
rect 1492 31418 1544 31424
rect 1504 30394 1532 31418
rect 1492 30388 1544 30394
rect 1492 30330 1544 30336
rect 1492 30252 1544 30258
rect 1492 30194 1544 30200
rect 1504 30161 1532 30194
rect 1490 30152 1546 30161
rect 1490 30087 1546 30096
rect 1400 29776 1452 29782
rect 1400 29718 1452 29724
rect 1400 29640 1452 29646
rect 1596 29594 1624 32914
rect 1688 32910 1716 33238
rect 1676 32904 1728 32910
rect 1674 32872 1676 32881
rect 1728 32872 1730 32881
rect 1674 32807 1730 32816
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1688 31686 1716 32506
rect 1768 32292 1820 32298
rect 1768 32234 1820 32240
rect 1780 32026 1808 32234
rect 1768 32020 1820 32026
rect 1768 31962 1820 31968
rect 1676 31680 1728 31686
rect 1676 31622 1728 31628
rect 1872 31464 1900 34734
rect 1964 34474 1992 34954
rect 1952 34468 2004 34474
rect 1952 34410 2004 34416
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 2320 33992 2372 33998
rect 2320 33934 2372 33940
rect 2412 33992 2464 33998
rect 2412 33934 2464 33940
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 1952 32904 2004 32910
rect 1952 32846 2004 32852
rect 1964 32570 1992 32846
rect 1952 32564 2004 32570
rect 1952 32506 2004 32512
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 2042 31920 2098 31929
rect 2042 31855 2098 31864
rect 2228 31884 2280 31890
rect 1952 31680 2004 31686
rect 1952 31622 2004 31628
rect 1780 31436 1900 31464
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 1688 30734 1716 31282
rect 1676 30728 1728 30734
rect 1676 30670 1728 30676
rect 1688 30054 1716 30670
rect 1780 30326 1808 31436
rect 1964 31362 1992 31622
rect 2056 31414 2084 31855
rect 2228 31826 2280 31832
rect 1872 31334 1992 31362
rect 2044 31408 2096 31414
rect 2044 31350 2096 31356
rect 1768 30320 1820 30326
rect 1768 30262 1820 30268
rect 1768 30184 1820 30190
rect 1768 30126 1820 30132
rect 1676 30048 1728 30054
rect 1676 29990 1728 29996
rect 1400 29582 1452 29588
rect 1412 29481 1440 29582
rect 1504 29566 1624 29594
rect 1398 29472 1454 29481
rect 1398 29407 1454 29416
rect 1398 29200 1454 29209
rect 1398 29135 1454 29144
rect 1412 28762 1440 29135
rect 1400 28756 1452 28762
rect 1400 28698 1452 28704
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27849 1440 28018
rect 1398 27840 1454 27849
rect 1398 27775 1454 27784
rect 1504 27441 1532 29566
rect 1584 29504 1636 29510
rect 1584 29446 1636 29452
rect 1490 27432 1546 27441
rect 1490 27367 1546 27376
rect 1492 27056 1544 27062
rect 1398 27024 1454 27033
rect 1492 26998 1544 27004
rect 1398 26959 1400 26968
rect 1452 26959 1454 26968
rect 1400 26930 1452 26936
rect 1398 25392 1454 25401
rect 1398 25327 1454 25336
rect 1412 25294 1440 25327
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 24585 1440 24754
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1504 24410 1532 26998
rect 1596 24682 1624 29446
rect 1780 29238 1808 30126
rect 1768 29232 1820 29238
rect 1688 29192 1768 29220
rect 1688 28937 1716 29192
rect 1768 29174 1820 29180
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 1674 28928 1730 28937
rect 1674 28863 1730 28872
rect 1780 28558 1808 29038
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1780 28150 1808 28494
rect 1768 28144 1820 28150
rect 1768 28086 1820 28092
rect 1676 27872 1728 27878
rect 1676 27814 1728 27820
rect 1688 26994 1716 27814
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 1688 26382 1716 26930
rect 1780 26926 1808 28086
rect 1872 27656 1900 31334
rect 2240 31249 2268 31826
rect 2226 31240 2282 31249
rect 2226 31175 2282 31184
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 2228 29776 2280 29782
rect 2228 29718 2280 29724
rect 2240 29322 2268 29718
rect 2332 29510 2360 33934
rect 2424 33590 2452 33934
rect 2412 33584 2464 33590
rect 2412 33526 2464 33532
rect 2412 33448 2464 33454
rect 2412 33390 2464 33396
rect 2424 31906 2452 33390
rect 2516 32026 2544 35142
rect 2504 32020 2556 32026
rect 2504 31962 2556 31968
rect 2424 31878 2544 31906
rect 2412 31816 2464 31822
rect 2412 31758 2464 31764
rect 2424 30938 2452 31758
rect 2412 30932 2464 30938
rect 2412 30874 2464 30880
rect 2412 30728 2464 30734
rect 2412 30670 2464 30676
rect 2424 29782 2452 30670
rect 2412 29776 2464 29782
rect 2412 29718 2464 29724
rect 2410 29608 2466 29617
rect 2410 29543 2466 29552
rect 2320 29504 2372 29510
rect 2320 29446 2372 29452
rect 2240 29306 2360 29322
rect 2240 29300 2372 29306
rect 2240 29294 2320 29300
rect 2320 29242 2372 29248
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 2332 28642 2360 29242
rect 2148 28614 2360 28642
rect 2148 28558 2176 28614
rect 2136 28552 2188 28558
rect 2424 28506 2452 29543
rect 2136 28494 2188 28500
rect 2148 27985 2176 28494
rect 2332 28478 2452 28506
rect 2134 27976 2190 27985
rect 2134 27911 2190 27920
rect 2332 27826 2360 28478
rect 2412 28416 2464 28422
rect 2412 28358 2464 28364
rect 2424 28218 2452 28358
rect 2412 28212 2464 28218
rect 2412 28154 2464 28160
rect 2332 27798 2452 27826
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 1872 27628 1992 27656
rect 1858 27568 1914 27577
rect 1858 27503 1914 27512
rect 1768 26920 1820 26926
rect 1768 26862 1820 26868
rect 1676 26376 1728 26382
rect 1780 26364 1808 26862
rect 1872 26466 1900 27503
rect 1964 27062 1992 27628
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2044 27328 2096 27334
rect 2044 27270 2096 27276
rect 2056 27130 2084 27270
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 1952 27056 2004 27062
rect 1952 26998 2004 27004
rect 2240 26994 2268 27406
rect 2320 27056 2372 27062
rect 2320 26998 2372 27004
rect 2228 26988 2280 26994
rect 2228 26930 2280 26936
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 1872 26438 1992 26466
rect 1860 26376 1912 26382
rect 1780 26336 1860 26364
rect 1676 26318 1728 26324
rect 1860 26318 1912 26324
rect 1584 24676 1636 24682
rect 1584 24618 1636 24624
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23769 1440 24142
rect 1398 23760 1454 23769
rect 1504 23730 1532 24346
rect 1398 23695 1454 23704
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22953 1440 23054
rect 1398 22944 1454 22953
rect 1504 22930 1532 23666
rect 1596 23050 1624 24618
rect 1584 23044 1636 23050
rect 1584 22986 1636 22992
rect 1504 22902 1624 22930
rect 1398 22879 1454 22888
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1492 22636 1544 22642
rect 1492 22578 1544 22584
rect 1412 22137 1440 22578
rect 1398 22128 1454 22137
rect 1504 22098 1532 22578
rect 1398 22063 1454 22072
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1490 21992 1546 22001
rect 1412 21554 1440 21966
rect 1596 21962 1624 22902
rect 1490 21927 1546 21936
rect 1584 21956 1636 21962
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 1412 20942 1440 21247
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1398 20632 1454 20641
rect 1398 20567 1454 20576
rect 1412 20058 1440 20567
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19689 1440 19790
rect 1398 19680 1454 19689
rect 1398 19615 1454 19624
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 18873 1440 19314
rect 1398 18864 1454 18873
rect 1398 18799 1454 18808
rect 1504 18698 1532 21927
rect 1584 21898 1636 21904
rect 1584 21616 1636 21622
rect 1584 21558 1636 21564
rect 1596 19258 1624 21558
rect 1688 21554 1716 26318
rect 1768 25968 1820 25974
rect 1768 25910 1820 25916
rect 1780 21622 1808 25910
rect 1872 24274 1900 26318
rect 1964 26246 1992 26438
rect 1952 26240 2004 26246
rect 1952 26182 2004 26188
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2148 24721 2176 24754
rect 2240 24750 2268 25094
rect 2228 24744 2280 24750
rect 2134 24712 2190 24721
rect 2228 24686 2280 24692
rect 2134 24647 2190 24656
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 2136 24268 2188 24274
rect 2136 24210 2188 24216
rect 2148 23798 2176 24210
rect 2332 24206 2360 26998
rect 2424 26738 2452 27798
rect 2516 27062 2544 31878
rect 2608 30870 2636 38762
rect 2688 38412 2740 38418
rect 2688 38354 2740 38360
rect 2700 37806 2728 38354
rect 2688 37800 2740 37806
rect 2688 37742 2740 37748
rect 2700 35630 2728 37742
rect 2792 35737 2820 39306
rect 3010 39196 3318 39205
rect 3010 39194 3016 39196
rect 3072 39194 3096 39196
rect 3152 39194 3176 39196
rect 3232 39194 3256 39196
rect 3312 39194 3318 39196
rect 3072 39142 3074 39194
rect 3254 39142 3256 39194
rect 3010 39140 3016 39142
rect 3072 39140 3096 39142
rect 3152 39140 3176 39142
rect 3232 39140 3256 39142
rect 3312 39140 3318 39142
rect 3010 39131 3318 39140
rect 3424 38548 3476 38554
rect 3424 38490 3476 38496
rect 3436 38282 3464 38490
rect 3424 38276 3476 38282
rect 3424 38218 3476 38224
rect 3516 38276 3568 38282
rect 3516 38218 3568 38224
rect 2872 38208 2924 38214
rect 2872 38150 2924 38156
rect 2884 37806 2912 38150
rect 3010 38108 3318 38117
rect 3010 38106 3016 38108
rect 3072 38106 3096 38108
rect 3152 38106 3176 38108
rect 3232 38106 3256 38108
rect 3312 38106 3318 38108
rect 3072 38054 3074 38106
rect 3254 38054 3256 38106
rect 3010 38052 3016 38054
rect 3072 38052 3096 38054
rect 3152 38052 3176 38054
rect 3232 38052 3256 38054
rect 3312 38052 3318 38054
rect 3010 38043 3318 38052
rect 3528 37806 3556 38218
rect 2872 37800 2924 37806
rect 2872 37742 2924 37748
rect 3424 37800 3476 37806
rect 3424 37742 3476 37748
rect 3516 37800 3568 37806
rect 3516 37742 3568 37748
rect 3010 37020 3318 37029
rect 3010 37018 3016 37020
rect 3072 37018 3096 37020
rect 3152 37018 3176 37020
rect 3232 37018 3256 37020
rect 3312 37018 3318 37020
rect 3072 36966 3074 37018
rect 3254 36966 3256 37018
rect 3010 36964 3016 36966
rect 3072 36964 3096 36966
rect 3152 36964 3176 36966
rect 3232 36964 3256 36966
rect 3312 36964 3318 36966
rect 3010 36955 3318 36964
rect 3436 36650 3464 37742
rect 3424 36644 3476 36650
rect 3424 36586 3476 36592
rect 2872 36032 2924 36038
rect 2872 35974 2924 35980
rect 2778 35728 2834 35737
rect 2778 35663 2834 35672
rect 2884 35630 2912 35974
rect 3010 35932 3318 35941
rect 3010 35930 3016 35932
rect 3072 35930 3096 35932
rect 3152 35930 3176 35932
rect 3232 35930 3256 35932
rect 3312 35930 3318 35932
rect 3072 35878 3074 35930
rect 3254 35878 3256 35930
rect 3010 35876 3016 35878
rect 3072 35876 3096 35878
rect 3152 35876 3176 35878
rect 3232 35876 3256 35878
rect 3312 35876 3318 35878
rect 3010 35867 3318 35876
rect 3436 35630 3464 36586
rect 3528 35630 3556 37742
rect 3608 36848 3660 36854
rect 3608 36790 3660 36796
rect 2688 35624 2740 35630
rect 2688 35566 2740 35572
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2872 35624 2924 35630
rect 2872 35566 2924 35572
rect 3424 35624 3476 35630
rect 3424 35566 3476 35572
rect 3516 35624 3568 35630
rect 3516 35566 3568 35572
rect 2596 30864 2648 30870
rect 2596 30806 2648 30812
rect 2596 30728 2648 30734
rect 2596 30670 2648 30676
rect 2608 30190 2636 30670
rect 2596 30184 2648 30190
rect 2700 30172 2728 35566
rect 2792 35476 2820 35566
rect 3240 35556 3292 35562
rect 3240 35498 3292 35504
rect 2792 35448 2912 35476
rect 2780 34604 2832 34610
rect 2780 34546 2832 34552
rect 2792 32774 2820 34546
rect 2780 32768 2832 32774
rect 2780 32710 2832 32716
rect 2884 32570 2912 35448
rect 3252 35193 3280 35498
rect 3238 35184 3294 35193
rect 3238 35119 3294 35128
rect 3010 34844 3318 34853
rect 3010 34842 3016 34844
rect 3072 34842 3096 34844
rect 3152 34842 3176 34844
rect 3232 34842 3256 34844
rect 3312 34842 3318 34844
rect 3072 34790 3074 34842
rect 3254 34790 3256 34842
rect 3010 34788 3016 34790
rect 3072 34788 3096 34790
rect 3152 34788 3176 34790
rect 3232 34788 3256 34790
rect 3312 34788 3318 34790
rect 3010 34779 3318 34788
rect 3436 34202 3464 35566
rect 3424 34196 3476 34202
rect 3424 34138 3476 34144
rect 3516 33992 3568 33998
rect 3436 33952 3516 33980
rect 3010 33756 3318 33765
rect 3010 33754 3016 33756
rect 3072 33754 3096 33756
rect 3152 33754 3176 33756
rect 3232 33754 3256 33756
rect 3312 33754 3318 33756
rect 3072 33702 3074 33754
rect 3254 33702 3256 33754
rect 3010 33700 3016 33702
rect 3072 33700 3096 33702
rect 3152 33700 3176 33702
rect 3232 33700 3256 33702
rect 3312 33700 3318 33702
rect 3010 33691 3318 33700
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 3240 33448 3292 33454
rect 3240 33390 3292 33396
rect 3332 33448 3384 33454
rect 3436 33436 3464 33952
rect 3516 33934 3568 33940
rect 3516 33856 3568 33862
rect 3516 33798 3568 33804
rect 3528 33454 3556 33798
rect 3384 33408 3464 33436
rect 3516 33448 3568 33454
rect 3332 33390 3384 33396
rect 3516 33390 3568 33396
rect 2964 33312 3016 33318
rect 2964 33254 3016 33260
rect 2976 32978 3004 33254
rect 3068 33114 3096 33390
rect 3252 33114 3280 33390
rect 3056 33108 3108 33114
rect 3056 33050 3108 33056
rect 3240 33108 3292 33114
rect 3240 33050 3292 33056
rect 2964 32972 3016 32978
rect 2964 32914 3016 32920
rect 3344 32722 3372 33390
rect 3620 33046 3648 36790
rect 3712 36718 3740 39442
rect 3700 36712 3752 36718
rect 3700 36654 3752 36660
rect 3700 36576 3752 36582
rect 3700 36518 3752 36524
rect 3712 35698 3740 36518
rect 3700 35692 3752 35698
rect 3700 35634 3752 35640
rect 3700 33856 3752 33862
rect 3700 33798 3752 33804
rect 3608 33040 3660 33046
rect 3608 32982 3660 32988
rect 3344 32694 3556 32722
rect 3010 32668 3318 32677
rect 3010 32666 3016 32668
rect 3072 32666 3096 32668
rect 3152 32666 3176 32668
rect 3232 32666 3256 32668
rect 3312 32666 3318 32668
rect 3072 32614 3074 32666
rect 3254 32614 3256 32666
rect 3010 32612 3016 32614
rect 3072 32612 3096 32614
rect 3152 32612 3176 32614
rect 3232 32612 3256 32614
rect 3312 32612 3318 32614
rect 3010 32603 3318 32612
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 3424 32564 3476 32570
rect 3424 32506 3476 32512
rect 3240 32360 3292 32366
rect 3240 32302 3292 32308
rect 2780 32224 2832 32230
rect 2780 32166 2832 32172
rect 2792 30297 2820 32166
rect 2884 32150 3096 32178
rect 2884 31482 2912 32150
rect 3068 31890 3096 32150
rect 3056 31884 3108 31890
rect 3056 31826 3108 31832
rect 3252 31686 3280 32302
rect 3240 31680 3292 31686
rect 3240 31622 3292 31628
rect 3010 31580 3318 31589
rect 3010 31578 3016 31580
rect 3072 31578 3096 31580
rect 3152 31578 3176 31580
rect 3232 31578 3256 31580
rect 3312 31578 3318 31580
rect 3072 31526 3074 31578
rect 3254 31526 3256 31578
rect 3010 31524 3016 31526
rect 3072 31524 3096 31526
rect 3152 31524 3176 31526
rect 3232 31524 3256 31526
rect 3312 31524 3318 31526
rect 3010 31515 3318 31524
rect 2872 31476 2924 31482
rect 2872 31418 2924 31424
rect 3332 31340 3384 31346
rect 3332 31282 3384 31288
rect 3344 30802 3372 31282
rect 3332 30796 3384 30802
rect 3332 30738 3384 30744
rect 2872 30592 2924 30598
rect 2872 30534 2924 30540
rect 2778 30288 2834 30297
rect 2778 30223 2834 30232
rect 2700 30144 2820 30172
rect 2596 30126 2648 30132
rect 2608 29646 2636 30126
rect 2688 29776 2740 29782
rect 2688 29718 2740 29724
rect 2596 29640 2648 29646
rect 2596 29582 2648 29588
rect 2608 27554 2636 29582
rect 2700 29073 2728 29718
rect 2686 29064 2742 29073
rect 2686 28999 2742 29008
rect 2688 28960 2740 28966
rect 2688 28902 2740 28908
rect 2700 28014 2728 28902
rect 2688 28008 2740 28014
rect 2688 27950 2740 27956
rect 2608 27526 2728 27554
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 2504 27056 2556 27062
rect 2504 26998 2556 27004
rect 2424 26710 2544 26738
rect 2412 26376 2464 26382
rect 2412 26318 2464 26324
rect 2424 25906 2452 26318
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2424 25378 2452 25842
rect 2516 25786 2544 26710
rect 2608 25906 2636 27406
rect 2700 26024 2728 27526
rect 2792 26976 2820 30144
rect 2884 28529 2912 30534
rect 3010 30492 3318 30501
rect 3010 30490 3016 30492
rect 3072 30490 3096 30492
rect 3152 30490 3176 30492
rect 3232 30490 3256 30492
rect 3312 30490 3318 30492
rect 3072 30438 3074 30490
rect 3254 30438 3256 30490
rect 3010 30436 3016 30438
rect 3072 30436 3096 30438
rect 3152 30436 3176 30438
rect 3232 30436 3256 30438
rect 3312 30436 3318 30438
rect 3010 30427 3318 30436
rect 3332 30320 3384 30326
rect 3332 30262 3384 30268
rect 3344 29458 3372 30262
rect 3436 29782 3464 32506
rect 3528 31822 3556 32694
rect 3608 32564 3660 32570
rect 3608 32506 3660 32512
rect 3516 31816 3568 31822
rect 3516 31758 3568 31764
rect 3516 31680 3568 31686
rect 3516 31622 3568 31628
rect 3528 30734 3556 31622
rect 3620 31482 3648 32506
rect 3608 31476 3660 31482
rect 3608 31418 3660 31424
rect 3608 31272 3660 31278
rect 3608 31214 3660 31220
rect 3620 30938 3648 31214
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3712 30818 3740 33798
rect 3804 33318 3832 41414
rect 3884 40996 3936 41002
rect 3884 40938 3936 40944
rect 3896 37126 3924 40938
rect 3988 39506 4016 42230
rect 4988 42220 5040 42226
rect 4988 42162 5040 42168
rect 5448 42220 5500 42226
rect 5448 42162 5500 42168
rect 6184 42220 6236 42226
rect 6184 42162 6236 42168
rect 6552 42220 6604 42226
rect 6552 42162 6604 42168
rect 5000 41546 5028 42162
rect 5460 41750 5488 42162
rect 5448 41744 5500 41750
rect 5448 41686 5500 41692
rect 6000 41676 6052 41682
rect 6000 41618 6052 41624
rect 5448 41608 5500 41614
rect 5448 41550 5500 41556
rect 4988 41540 5040 41546
rect 4988 41482 5040 41488
rect 4068 40180 4120 40186
rect 4068 40122 4120 40128
rect 3976 39500 4028 39506
rect 3976 39442 4028 39448
rect 3976 39364 4028 39370
rect 3976 39306 4028 39312
rect 3988 38010 4016 39306
rect 3976 38004 4028 38010
rect 3976 37946 4028 37952
rect 4080 37194 4108 40122
rect 5172 39432 5224 39438
rect 5172 39374 5224 39380
rect 4436 39296 4488 39302
rect 4436 39238 4488 39244
rect 4344 38956 4396 38962
rect 4344 38898 4396 38904
rect 4160 38208 4212 38214
rect 4160 38150 4212 38156
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3884 36712 3936 36718
rect 3884 36654 3936 36660
rect 3896 35873 3924 36654
rect 4068 36576 4120 36582
rect 4068 36518 4120 36524
rect 4080 36310 4108 36518
rect 4068 36304 4120 36310
rect 4068 36246 4120 36252
rect 3882 35864 3938 35873
rect 4172 35834 4200 38150
rect 4356 38010 4384 38898
rect 4448 38486 4476 39238
rect 4988 38956 5040 38962
rect 4988 38898 5040 38904
rect 4712 38548 4764 38554
rect 4712 38490 4764 38496
rect 4436 38480 4488 38486
rect 4436 38422 4488 38428
rect 4344 38004 4396 38010
rect 4344 37946 4396 37952
rect 4620 37868 4672 37874
rect 4620 37810 4672 37816
rect 4252 37800 4304 37806
rect 4252 37742 4304 37748
rect 4264 37262 4292 37742
rect 4252 37256 4304 37262
rect 4528 37256 4580 37262
rect 4252 37198 4304 37204
rect 4526 37224 4528 37233
rect 4580 37224 4582 37233
rect 4264 36922 4292 37198
rect 4526 37159 4582 37168
rect 4252 36916 4304 36922
rect 4252 36858 4304 36864
rect 4344 36780 4396 36786
rect 4344 36722 4396 36728
rect 4528 36780 4580 36786
rect 4528 36722 4580 36728
rect 4252 36712 4304 36718
rect 4252 36654 4304 36660
rect 4264 36378 4292 36654
rect 4252 36372 4304 36378
rect 4252 36314 4304 36320
rect 4356 35834 4384 36722
rect 4436 36236 4488 36242
rect 4436 36178 4488 36184
rect 3882 35799 3938 35808
rect 4160 35828 4212 35834
rect 4160 35770 4212 35776
rect 4344 35828 4396 35834
rect 4344 35770 4396 35776
rect 3884 35624 3936 35630
rect 3884 35566 3936 35572
rect 3792 33312 3844 33318
rect 3792 33254 3844 33260
rect 3792 33040 3844 33046
rect 3792 32982 3844 32988
rect 3896 32994 3924 35566
rect 4448 35034 4476 36178
rect 4540 35154 4568 36722
rect 4528 35148 4580 35154
rect 4528 35090 4580 35096
rect 4632 35034 4660 37810
rect 4356 35006 4476 35034
rect 4540 35006 4660 35034
rect 3976 34400 4028 34406
rect 3976 34342 4028 34348
rect 4068 34400 4120 34406
rect 4068 34342 4120 34348
rect 3988 34134 4016 34342
rect 3976 34128 4028 34134
rect 3976 34070 4028 34076
rect 3976 33992 4028 33998
rect 3976 33934 4028 33940
rect 3988 33114 4016 33934
rect 3976 33108 4028 33114
rect 3976 33050 4028 33056
rect 3620 30790 3740 30818
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3528 30190 3556 30670
rect 3516 30184 3568 30190
rect 3516 30126 3568 30132
rect 3424 29776 3476 29782
rect 3424 29718 3476 29724
rect 3344 29430 3464 29458
rect 3010 29404 3318 29413
rect 3010 29402 3016 29404
rect 3072 29402 3096 29404
rect 3152 29402 3176 29404
rect 3232 29402 3256 29404
rect 3312 29402 3318 29404
rect 3072 29350 3074 29402
rect 3254 29350 3256 29402
rect 3010 29348 3016 29350
rect 3072 29348 3096 29350
rect 3152 29348 3176 29350
rect 3232 29348 3256 29350
rect 3312 29348 3318 29350
rect 3010 29339 3318 29348
rect 3436 29322 3464 29430
rect 3344 29294 3464 29322
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 2870 28520 2926 28529
rect 2870 28455 2926 28464
rect 2976 28404 3004 29174
rect 3240 28756 3292 28762
rect 3240 28698 3292 28704
rect 3252 28490 3280 28698
rect 3344 28626 3372 29294
rect 3528 29238 3556 30126
rect 3620 29510 3648 30790
rect 3804 30682 3832 32982
rect 3896 32966 4016 32994
rect 3884 32224 3936 32230
rect 3884 32166 3936 32172
rect 3896 31958 3924 32166
rect 3884 31952 3936 31958
rect 3884 31894 3936 31900
rect 3884 31816 3936 31822
rect 3884 31758 3936 31764
rect 3712 30654 3832 30682
rect 3712 30297 3740 30654
rect 3790 30560 3846 30569
rect 3790 30495 3846 30504
rect 3698 30288 3754 30297
rect 3698 30223 3754 30232
rect 3700 30048 3752 30054
rect 3700 29990 3752 29996
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3516 29232 3568 29238
rect 3516 29174 3568 29180
rect 3608 29232 3660 29238
rect 3608 29174 3660 29180
rect 3422 29064 3478 29073
rect 3422 28999 3478 29008
rect 3332 28620 3384 28626
rect 3332 28562 3384 28568
rect 3240 28484 3292 28490
rect 3240 28426 3292 28432
rect 2884 28376 3004 28404
rect 2884 27674 2912 28376
rect 3010 28316 3318 28325
rect 3010 28314 3016 28316
rect 3072 28314 3096 28316
rect 3152 28314 3176 28316
rect 3232 28314 3256 28316
rect 3312 28314 3318 28316
rect 3072 28262 3074 28314
rect 3254 28262 3256 28314
rect 3010 28260 3016 28262
rect 3072 28260 3096 28262
rect 3152 28260 3176 28262
rect 3232 28260 3256 28262
rect 3312 28260 3318 28262
rect 3010 28251 3318 28260
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 3056 27872 3108 27878
rect 3054 27840 3056 27849
rect 3108 27840 3110 27849
rect 3054 27775 3110 27784
rect 3252 27674 3280 27950
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 3240 27668 3292 27674
rect 3240 27610 3292 27616
rect 3010 27228 3318 27237
rect 3010 27226 3016 27228
rect 3072 27226 3096 27228
rect 3152 27226 3176 27228
rect 3232 27226 3256 27228
rect 3312 27226 3318 27228
rect 3072 27174 3074 27226
rect 3254 27174 3256 27226
rect 3010 27172 3016 27174
rect 3072 27172 3096 27174
rect 3152 27172 3176 27174
rect 3232 27172 3256 27174
rect 3312 27172 3318 27174
rect 3010 27163 3318 27172
rect 2792 26948 3004 26976
rect 2870 26888 2926 26897
rect 2870 26823 2926 26832
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 2792 26382 2820 26726
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 2700 25996 2820 26024
rect 2686 25936 2742 25945
rect 2596 25900 2648 25906
rect 2686 25871 2742 25880
rect 2596 25842 2648 25848
rect 2516 25758 2636 25786
rect 2504 25696 2556 25702
rect 2504 25638 2556 25644
rect 2516 25537 2544 25638
rect 2502 25528 2558 25537
rect 2502 25463 2558 25472
rect 2424 25350 2544 25378
rect 2516 25294 2544 25350
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2424 24274 2452 24686
rect 2412 24268 2464 24274
rect 2412 24210 2464 24216
rect 2320 24200 2372 24206
rect 2372 24148 2452 24154
rect 2320 24142 2452 24148
rect 2228 24132 2280 24138
rect 2332 24126 2452 24142
rect 2228 24074 2280 24080
rect 2240 23866 2268 24074
rect 2320 24064 2372 24070
rect 2320 24006 2372 24012
rect 2228 23860 2280 23866
rect 2228 23802 2280 23808
rect 2136 23792 2188 23798
rect 2136 23734 2188 23740
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1872 23118 1900 23598
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 1952 23248 2004 23254
rect 1950 23216 1952 23225
rect 2004 23216 2006 23225
rect 1950 23151 2006 23160
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1768 21616 1820 21622
rect 1768 21558 1820 21564
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1688 19378 1716 21490
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 20602 1808 21286
rect 1872 21128 1900 23054
rect 2044 23044 2096 23050
rect 2044 22986 2096 22992
rect 2056 22642 2084 22986
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 2228 21956 2280 21962
rect 2228 21898 2280 21904
rect 2240 21457 2268 21898
rect 2226 21448 2282 21457
rect 2226 21383 2282 21392
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 1872 21100 1992 21128
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1768 20596 1820 20602
rect 1768 20538 1820 20544
rect 1872 20330 1900 20742
rect 1964 20466 1992 21100
rect 2042 21040 2098 21049
rect 2042 20975 2098 20984
rect 2228 21004 2280 21010
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 2056 20262 2084 20975
rect 2228 20946 2280 20952
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 2044 20256 2096 20262
rect 2240 20244 2268 20946
rect 2332 20369 2360 24006
rect 2318 20360 2374 20369
rect 2318 20295 2374 20304
rect 2240 20216 2360 20244
rect 2044 20198 2096 20204
rect 1780 19922 1808 20198
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 2332 20040 2360 20216
rect 2240 20012 2360 20040
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1596 19230 1716 19258
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1492 18692 1544 18698
rect 1492 18634 1544 18640
rect 1308 18420 1360 18426
rect 1308 18362 1360 18368
rect 1308 18284 1360 18290
rect 1308 18226 1360 18232
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1216 17876 1268 17882
rect 1216 17818 1268 17824
rect 1216 17672 1268 17678
rect 1216 17614 1268 17620
rect 940 17070 992 17076
rect 952 12220 980 17070
rect 1044 17054 1164 17082
rect 1044 15026 1072 17054
rect 1124 16584 1176 16590
rect 1124 16526 1176 16532
rect 1032 15020 1084 15026
rect 1032 14962 1084 14968
rect 1032 13456 1084 13462
rect 1032 13398 1084 13404
rect 1044 12345 1072 13398
rect 1030 12336 1086 12345
rect 1030 12271 1086 12280
rect 952 12192 1072 12220
rect 848 11824 900 11830
rect 848 11766 900 11772
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 848 11280 900 11286
rect 848 11222 900 11228
rect 860 10713 888 11222
rect 952 11218 980 11630
rect 940 11212 992 11218
rect 940 11154 992 11160
rect 940 11008 992 11014
rect 940 10950 992 10956
rect 846 10704 902 10713
rect 846 10639 902 10648
rect 848 8832 900 8838
rect 848 8774 900 8780
rect 860 8265 888 8774
rect 846 8256 902 8265
rect 846 8191 902 8200
rect 756 4276 808 4282
rect 756 4218 808 4224
rect 664 2576 716 2582
rect 664 2518 716 2524
rect 952 56 980 10950
rect 1044 10062 1072 12192
rect 1032 10056 1084 10062
rect 1032 9998 1084 10004
rect 1030 9752 1086 9761
rect 1030 9687 1086 9696
rect 1044 4690 1072 9687
rect 1032 4684 1084 4690
rect 1032 4626 1084 4632
rect 1136 4214 1164 16526
rect 1228 15609 1256 17614
rect 1214 15600 1270 15609
rect 1214 15535 1270 15544
rect 1320 15178 1348 18226
rect 1412 18057 1440 18226
rect 1492 18148 1544 18154
rect 1492 18090 1544 18096
rect 1398 18048 1454 18057
rect 1398 17983 1454 17992
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1412 17202 1440 17478
rect 1504 17270 1532 18090
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 16658 1440 17138
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1398 16416 1454 16425
rect 1398 16351 1454 16360
rect 1412 16114 1440 16351
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1320 15150 1440 15178
rect 1214 14920 1270 14929
rect 1214 14855 1270 14864
rect 1228 8634 1256 14855
rect 1308 12436 1360 12442
rect 1308 12378 1360 12384
rect 1320 11762 1348 12378
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1308 11620 1360 11626
rect 1308 11562 1360 11568
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 1320 6458 1348 11562
rect 1412 11014 1440 15150
rect 1504 15094 1532 17206
rect 1596 16590 1624 19110
rect 1688 18834 1716 19230
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1780 18578 1808 19654
rect 2240 19334 2268 20012
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 1688 18550 1808 18578
rect 1872 19306 2268 19334
rect 1688 18154 1716 18550
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1688 16114 1716 17818
rect 1780 17762 1808 18158
rect 1872 17864 1900 19306
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18290 1992 18770
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 1872 17836 1992 17864
rect 1780 17734 1900 17762
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1688 15570 1716 15914
rect 1676 15564 1728 15570
rect 1596 15524 1676 15552
rect 1492 15088 1544 15094
rect 1492 15030 1544 15036
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13977 1532 14214
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1596 13410 1624 15524
rect 1676 15506 1728 15512
rect 1780 14634 1808 17614
rect 1688 14606 1808 14634
rect 1688 14006 1716 14606
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 14000 1728 14006
rect 1676 13942 1728 13948
rect 1780 13938 1808 14418
rect 1872 14346 1900 17734
rect 1964 17678 1992 17836
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2240 16980 2268 17614
rect 2332 17105 2360 19751
rect 2424 18290 2452 24126
rect 2516 20942 2544 25230
rect 2608 24070 2636 25758
rect 2596 24064 2648 24070
rect 2596 24006 2648 24012
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2608 23186 2636 23734
rect 2700 23225 2728 25871
rect 2686 23216 2742 23225
rect 2596 23180 2648 23186
rect 2686 23151 2742 23160
rect 2596 23122 2648 23128
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2700 22556 2728 22918
rect 2792 22710 2820 25996
rect 2884 25498 2912 26823
rect 2976 26246 3004 26948
rect 3240 26920 3292 26926
rect 3240 26862 3292 26868
rect 3436 26874 3464 28999
rect 3620 28762 3648 29174
rect 3608 28756 3660 28762
rect 3608 28698 3660 28704
rect 3608 28620 3660 28626
rect 3608 28562 3660 28568
rect 3516 28416 3568 28422
rect 3516 28358 3568 28364
rect 3528 27946 3556 28358
rect 3516 27940 3568 27946
rect 3516 27882 3568 27888
rect 3516 27464 3568 27470
rect 3516 27406 3568 27412
rect 3528 27130 3556 27406
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3252 26586 3280 26862
rect 3436 26846 3556 26874
rect 3240 26580 3292 26586
rect 3240 26522 3292 26528
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 3010 26140 3318 26149
rect 3010 26138 3016 26140
rect 3072 26138 3096 26140
rect 3152 26138 3176 26140
rect 3232 26138 3256 26140
rect 3312 26138 3318 26140
rect 3072 26086 3074 26138
rect 3254 26086 3256 26138
rect 3010 26084 3016 26086
rect 3072 26084 3096 26086
rect 3152 26084 3176 26086
rect 3232 26084 3256 26086
rect 3312 26084 3318 26086
rect 3010 26075 3318 26084
rect 3424 26036 3476 26042
rect 3424 25978 3476 25984
rect 2964 25968 3016 25974
rect 2964 25910 3016 25916
rect 2872 25492 2924 25498
rect 2872 25434 2924 25440
rect 2976 25378 3004 25910
rect 3056 25492 3108 25498
rect 3056 25434 3108 25440
rect 2884 25350 3004 25378
rect 2884 23322 2912 25350
rect 3068 25226 3096 25434
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 3010 25052 3318 25061
rect 3010 25050 3016 25052
rect 3072 25050 3096 25052
rect 3152 25050 3176 25052
rect 3232 25050 3256 25052
rect 3312 25050 3318 25052
rect 3072 24998 3074 25050
rect 3254 24998 3256 25050
rect 3010 24996 3016 24998
rect 3072 24996 3096 24998
rect 3152 24996 3176 24998
rect 3232 24996 3256 24998
rect 3312 24996 3318 24998
rect 3010 24987 3318 24996
rect 2964 24948 3016 24954
rect 2964 24890 3016 24896
rect 2976 24177 3004 24890
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3160 24177 3188 24686
rect 2962 24168 3018 24177
rect 2962 24103 3018 24112
rect 3146 24168 3202 24177
rect 3146 24103 3202 24112
rect 3010 23964 3318 23973
rect 3010 23962 3016 23964
rect 3072 23962 3096 23964
rect 3152 23962 3176 23964
rect 3232 23962 3256 23964
rect 3312 23962 3318 23964
rect 3072 23910 3074 23962
rect 3254 23910 3256 23962
rect 3010 23908 3016 23910
rect 3072 23908 3096 23910
rect 3152 23908 3176 23910
rect 3232 23908 3256 23910
rect 3312 23908 3318 23910
rect 3010 23899 3318 23908
rect 3240 23792 3292 23798
rect 2962 23760 3018 23769
rect 2962 23695 3018 23704
rect 3238 23760 3240 23769
rect 3292 23760 3294 23769
rect 3238 23695 3294 23704
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2976 23202 3004 23695
rect 2884 23174 3004 23202
rect 2780 22704 2832 22710
rect 2780 22646 2832 22652
rect 2700 22528 2820 22556
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2608 21486 2636 22374
rect 2686 21992 2742 22001
rect 2686 21927 2742 21936
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2516 19854 2544 20878
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 2516 19446 2544 19654
rect 2504 19440 2556 19446
rect 2504 19382 2556 19388
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2424 17377 2452 18226
rect 2410 17368 2466 17377
rect 2410 17303 2466 17312
rect 2516 17218 2544 19382
rect 2608 18170 2636 19994
rect 2700 19334 2728 21927
rect 2792 19394 2820 22528
rect 2884 19961 2912 23174
rect 3010 22876 3318 22885
rect 3010 22874 3016 22876
rect 3072 22874 3096 22876
rect 3152 22874 3176 22876
rect 3232 22874 3256 22876
rect 3312 22874 3318 22876
rect 3072 22822 3074 22874
rect 3254 22822 3256 22874
rect 3010 22820 3016 22822
rect 3072 22820 3096 22822
rect 3152 22820 3176 22822
rect 3232 22820 3256 22822
rect 3312 22820 3318 22822
rect 3010 22811 3318 22820
rect 3238 22672 3294 22681
rect 3238 22607 3294 22616
rect 3252 22030 3280 22607
rect 3436 22438 3464 25978
rect 3424 22432 3476 22438
rect 3330 22400 3386 22409
rect 3424 22374 3476 22380
rect 3330 22335 3386 22344
rect 3344 22250 3372 22335
rect 3528 22273 3556 26846
rect 3620 26081 3648 28562
rect 3712 26586 3740 29990
rect 3804 28665 3832 30495
rect 3790 28656 3846 28665
rect 3790 28591 3846 28600
rect 3896 27962 3924 31758
rect 3804 27934 3924 27962
rect 3804 27674 3832 27934
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3792 27668 3844 27674
rect 3792 27610 3844 27616
rect 3804 27130 3832 27610
rect 3792 27124 3844 27130
rect 3792 27066 3844 27072
rect 3792 26920 3844 26926
rect 3792 26862 3844 26868
rect 3700 26580 3752 26586
rect 3700 26522 3752 26528
rect 3606 26072 3662 26081
rect 3606 26007 3662 26016
rect 3608 25900 3660 25906
rect 3608 25842 3660 25848
rect 3514 22264 3570 22273
rect 3344 22222 3464 22250
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3010 21788 3318 21797
rect 3010 21786 3016 21788
rect 3072 21786 3096 21788
rect 3152 21786 3176 21788
rect 3232 21786 3256 21788
rect 3312 21786 3318 21788
rect 3072 21734 3074 21786
rect 3254 21734 3256 21786
rect 3010 21732 3016 21734
rect 3072 21732 3096 21734
rect 3152 21732 3176 21734
rect 3232 21732 3256 21734
rect 3312 21732 3318 21734
rect 3010 21723 3318 21732
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3344 21078 3372 21422
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 3010 20700 3318 20709
rect 3010 20698 3016 20700
rect 3072 20698 3096 20700
rect 3152 20698 3176 20700
rect 3232 20698 3256 20700
rect 3312 20698 3318 20700
rect 3072 20646 3074 20698
rect 3254 20646 3256 20698
rect 3010 20644 3016 20646
rect 3072 20644 3096 20646
rect 3152 20644 3176 20646
rect 3232 20644 3256 20646
rect 3312 20644 3318 20646
rect 3010 20635 3318 20644
rect 2870 19952 2926 19961
rect 2870 19887 2926 19896
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2884 19514 2912 19790
rect 3010 19612 3318 19621
rect 3010 19610 3016 19612
rect 3072 19610 3096 19612
rect 3152 19610 3176 19612
rect 3232 19610 3256 19612
rect 3312 19610 3318 19612
rect 3072 19558 3074 19610
rect 3254 19558 3256 19610
rect 3010 19556 3016 19558
rect 3072 19556 3096 19558
rect 3152 19556 3176 19558
rect 3232 19556 3256 19558
rect 3312 19556 3318 19558
rect 3010 19547 3318 19556
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2962 19408 3018 19417
rect 2792 19366 2912 19394
rect 2700 19306 2820 19334
rect 2792 18358 2820 19306
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2608 18142 2820 18170
rect 2688 18080 2740 18086
rect 2424 17190 2544 17218
rect 2608 18040 2688 18068
rect 2318 17096 2374 17105
rect 2318 17031 2374 17040
rect 2240 16952 2360 16980
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 15910 2084 16526
rect 2148 15978 2176 16730
rect 2332 15994 2360 16952
rect 2424 16794 2452 17190
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2516 16250 2544 17070
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2516 16114 2544 16186
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2136 15972 2188 15978
rect 2332 15966 2544 15994
rect 2136 15914 2188 15920
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1964 15026 1992 15506
rect 2332 15502 2360 15846
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1596 13382 1716 13410
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1492 13184 1544 13190
rect 1490 13152 1492 13161
rect 1544 13152 1546 13161
rect 1490 13087 1546 13096
rect 1492 12912 1544 12918
rect 1492 12854 1544 12860
rect 1504 11694 1532 12854
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1492 11552 1544 11558
rect 1490 11520 1492 11529
rect 1544 11520 1546 11529
rect 1490 11455 1546 11464
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 6914 1440 10610
rect 1504 10266 1532 10911
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1492 9920 1544 9926
rect 1490 9888 1492 9897
rect 1544 9888 1546 9897
rect 1490 9823 1546 9832
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1504 9081 1532 9318
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1504 7449 1532 7482
rect 1490 7440 1546 7449
rect 1490 7375 1546 7384
rect 1412 6886 1532 6914
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1412 6322 1440 6559
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1504 5114 1532 6886
rect 1596 6474 1624 13262
rect 1688 12918 1716 13382
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 1676 12912 1728 12918
rect 1676 12854 1728 12860
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12306 1716 12718
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 8566 1716 12106
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1688 7886 1716 8502
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1780 6914 1808 13262
rect 1872 12850 1900 14282
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1860 12844 1912 12850
rect 1860 12786 1912 12792
rect 1872 8566 1900 12786
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2240 11558 2268 12106
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 2044 11144 2096 11150
rect 1950 11112 2006 11121
rect 2044 11086 2096 11092
rect 1950 11047 1952 11056
rect 2004 11047 2006 11056
rect 1952 11018 2004 11024
rect 1964 10810 1992 11018
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 2056 10577 2084 11086
rect 2042 10568 2098 10577
rect 2042 10503 2098 10512
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 1950 10160 2006 10169
rect 1950 10095 2006 10104
rect 1964 10062 1992 10095
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 1964 8378 1992 9114
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8430 2268 8774
rect 1688 6886 1808 6914
rect 1872 8350 1992 8378
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 1688 6662 1716 6886
rect 1872 6798 1900 8350
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2042 7984 2098 7993
rect 2042 7919 2098 7928
rect 2228 7948 2280 7954
rect 2056 7546 2084 7919
rect 2228 7890 2280 7896
rect 2240 7818 2268 7890
rect 2332 7818 2360 15438
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 12050 2452 14758
rect 2516 12918 2544 15966
rect 2608 14822 2636 18040
rect 2688 18022 2740 18028
rect 2686 17912 2742 17921
rect 2792 17882 2820 18142
rect 2686 17847 2742 17856
rect 2780 17876 2832 17882
rect 2700 15570 2728 17847
rect 2780 17818 2832 17824
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2792 16794 2820 17002
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2778 16688 2834 16697
rect 2778 16623 2834 16632
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2516 12374 2544 12854
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2608 12238 2636 13874
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2424 12022 2636 12050
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11150 2452 11494
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2424 10674 2452 11086
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2424 9178 2452 10610
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10130 2544 10406
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9586 2544 10066
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2410 8256 2466 8265
rect 2410 8191 2466 8200
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2240 7342 2268 7754
rect 2332 7478 2360 7754
rect 2424 7546 2452 8191
rect 2516 7954 2544 8774
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2608 6798 2636 12022
rect 2700 7478 2728 14962
rect 2792 10062 2820 16623
rect 2884 12306 2912 19366
rect 2962 19343 3018 19352
rect 2976 18630 3004 19343
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 3010 18524 3318 18533
rect 3010 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3176 18524
rect 3232 18522 3256 18524
rect 3312 18522 3318 18524
rect 3072 18470 3074 18522
rect 3254 18470 3256 18522
rect 3010 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3176 18470
rect 3232 18468 3256 18470
rect 3312 18468 3318 18470
rect 3010 18459 3318 18468
rect 3330 18048 3386 18057
rect 3330 17983 3386 17992
rect 3344 17610 3372 17983
rect 3436 17746 3464 22222
rect 3514 22199 3570 22208
rect 3516 22024 3568 22030
rect 3516 21966 3568 21972
rect 3528 17921 3556 21966
rect 3620 20534 3648 25842
rect 3712 25838 3740 26522
rect 3804 26382 3832 26862
rect 3792 26376 3844 26382
rect 3896 26353 3924 27814
rect 3792 26318 3844 26324
rect 3882 26344 3938 26353
rect 3882 26279 3938 26288
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3700 25832 3752 25838
rect 3700 25774 3752 25780
rect 3804 24834 3832 26182
rect 3896 26042 3924 26182
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3896 24954 3924 25978
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 3712 24806 3832 24834
rect 3712 22137 3740 24806
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3804 22982 3832 24686
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 23662 3924 24550
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3882 23488 3938 23497
rect 3882 23423 3938 23432
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3896 22234 3924 23423
rect 3884 22228 3936 22234
rect 3884 22170 3936 22176
rect 3698 22128 3754 22137
rect 3698 22063 3754 22072
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3712 21486 3740 21830
rect 3790 21720 3846 21729
rect 3790 21655 3846 21664
rect 3700 21480 3752 21486
rect 3700 21422 3752 21428
rect 3804 21298 3832 21655
rect 3712 21270 3832 21298
rect 3712 21078 3740 21270
rect 3790 21176 3846 21185
rect 3790 21111 3846 21120
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3608 20528 3660 20534
rect 3608 20470 3660 20476
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3620 18986 3648 19314
rect 3712 19174 3740 21014
rect 3804 20777 3832 21111
rect 3896 20806 3924 21966
rect 3988 21865 4016 32966
rect 4080 30433 4108 34342
rect 4160 33448 4212 33454
rect 4158 33416 4160 33425
rect 4252 33448 4304 33454
rect 4212 33416 4214 33425
rect 4252 33390 4304 33396
rect 4158 33351 4214 33360
rect 4160 33312 4212 33318
rect 4160 33254 4212 33260
rect 4066 30424 4122 30433
rect 4066 30359 4122 30368
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 4080 28098 4108 29446
rect 4172 29209 4200 33254
rect 4264 31249 4292 33390
rect 4356 33046 4384 35006
rect 4436 34944 4488 34950
rect 4436 34886 4488 34892
rect 4448 34134 4476 34886
rect 4436 34128 4488 34134
rect 4436 34070 4488 34076
rect 4436 33108 4488 33114
rect 4436 33050 4488 33056
rect 4344 33040 4396 33046
rect 4344 32982 4396 32988
rect 4344 32428 4396 32434
rect 4344 32370 4396 32376
rect 4356 32026 4384 32370
rect 4344 32020 4396 32026
rect 4344 31962 4396 31968
rect 4342 31920 4398 31929
rect 4448 31890 4476 33050
rect 4342 31855 4398 31864
rect 4436 31884 4488 31890
rect 4356 31754 4384 31855
rect 4436 31826 4488 31832
rect 4540 31793 4568 35006
rect 4724 34898 4752 38490
rect 4896 37664 4948 37670
rect 4896 37606 4948 37612
rect 4632 34870 4752 34898
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 4526 31784 4582 31793
rect 4356 31726 4476 31754
rect 4342 31648 4398 31657
rect 4342 31583 4398 31592
rect 4250 31240 4306 31249
rect 4250 31175 4306 31184
rect 4252 31136 4304 31142
rect 4252 31078 4304 31084
rect 4158 29200 4214 29209
rect 4158 29135 4214 29144
rect 4160 29096 4212 29102
rect 4264 29073 4292 31078
rect 4160 29038 4212 29044
rect 4250 29064 4306 29073
rect 4172 28558 4200 29038
rect 4250 28999 4306 29008
rect 4252 28960 4304 28966
rect 4252 28902 4304 28908
rect 4264 28558 4292 28902
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 4252 28552 4304 28558
rect 4252 28494 4304 28500
rect 4172 28218 4200 28494
rect 4160 28212 4212 28218
rect 4160 28154 4212 28160
rect 4080 28070 4200 28098
rect 4068 28008 4120 28014
rect 4068 27950 4120 27956
rect 4080 27713 4108 27950
rect 4066 27704 4122 27713
rect 4066 27639 4122 27648
rect 4172 27577 4200 28070
rect 4252 28008 4304 28014
rect 4252 27950 4304 27956
rect 4158 27568 4214 27577
rect 4158 27503 4214 27512
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4080 22273 4108 27066
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 4172 24138 4200 24618
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 4158 24032 4214 24041
rect 4264 24018 4292 27950
rect 4356 27334 4384 31583
rect 4448 28966 4476 31726
rect 4526 31719 4582 31728
rect 4528 31680 4580 31686
rect 4528 31622 4580 31628
rect 4540 31346 4568 31622
rect 4528 31340 4580 31346
rect 4528 31282 4580 31288
rect 4540 30870 4568 31282
rect 4528 30864 4580 30870
rect 4528 30806 4580 30812
rect 4528 30388 4580 30394
rect 4528 30330 4580 30336
rect 4436 28960 4488 28966
rect 4436 28902 4488 28908
rect 4436 28416 4488 28422
rect 4436 28358 4488 28364
rect 4448 27538 4476 28358
rect 4436 27532 4488 27538
rect 4436 27474 4488 27480
rect 4540 27418 4568 30330
rect 4448 27390 4568 27418
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4448 27146 4476 27390
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4356 27118 4476 27146
rect 4356 26081 4384 27118
rect 4436 26920 4488 26926
rect 4436 26862 4488 26868
rect 4448 26761 4476 26862
rect 4434 26752 4490 26761
rect 4434 26687 4490 26696
rect 4448 26353 4476 26687
rect 4434 26344 4490 26353
rect 4540 26314 4568 27270
rect 4632 27130 4660 34870
rect 4816 34610 4844 34886
rect 4804 34604 4856 34610
rect 4804 34546 4856 34552
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 4724 33998 4752 34342
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 4804 33992 4856 33998
rect 4804 33934 4856 33940
rect 4724 32230 4752 33934
rect 4816 33454 4844 33934
rect 4804 33448 4856 33454
rect 4804 33390 4856 33396
rect 4804 32972 4856 32978
rect 4804 32914 4856 32920
rect 4816 32298 4844 32914
rect 4804 32292 4856 32298
rect 4804 32234 4856 32240
rect 4712 32224 4764 32230
rect 4712 32166 4764 32172
rect 4724 31464 4752 32166
rect 4816 31929 4844 32234
rect 4802 31920 4858 31929
rect 4802 31855 4858 31864
rect 4908 31872 4936 37606
rect 5000 37262 5028 38898
rect 5080 38344 5132 38350
rect 5080 38286 5132 38292
rect 4988 37256 5040 37262
rect 4986 37224 4988 37233
rect 5040 37224 5042 37233
rect 4986 37159 5042 37168
rect 5092 35562 5120 38286
rect 5184 38010 5212 39374
rect 5264 38752 5316 38758
rect 5264 38694 5316 38700
rect 5356 38752 5408 38758
rect 5356 38694 5408 38700
rect 5460 38706 5488 41550
rect 5816 39432 5868 39438
rect 5816 39374 5868 39380
rect 5828 39030 5856 39374
rect 5816 39024 5868 39030
rect 5816 38966 5868 38972
rect 5724 38956 5776 38962
rect 5724 38898 5776 38904
rect 5172 38004 5224 38010
rect 5172 37946 5224 37952
rect 5276 37330 5304 38694
rect 5368 38418 5396 38694
rect 5460 38678 5580 38706
rect 5356 38412 5408 38418
rect 5356 38354 5408 38360
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 5552 36922 5580 38678
rect 5736 38554 5764 38898
rect 5724 38548 5776 38554
rect 5724 38490 5776 38496
rect 5632 37868 5684 37874
rect 5632 37810 5684 37816
rect 5644 37466 5672 37810
rect 5828 37738 5856 38966
rect 5908 37936 5960 37942
rect 5908 37878 5960 37884
rect 5816 37732 5868 37738
rect 5816 37674 5868 37680
rect 5632 37460 5684 37466
rect 5632 37402 5684 37408
rect 5632 37188 5684 37194
rect 5632 37130 5684 37136
rect 5724 37188 5776 37194
rect 5724 37130 5776 37136
rect 5540 36916 5592 36922
rect 5540 36858 5592 36864
rect 5644 36258 5672 37130
rect 5552 36230 5672 36258
rect 5080 35556 5132 35562
rect 5080 35498 5132 35504
rect 5356 35080 5408 35086
rect 5356 35022 5408 35028
rect 5172 34740 5224 34746
rect 5172 34682 5224 34688
rect 5184 34649 5212 34682
rect 5170 34640 5226 34649
rect 5368 34610 5396 35022
rect 5448 34672 5500 34678
rect 5448 34614 5500 34620
rect 5170 34575 5226 34584
rect 5356 34604 5408 34610
rect 5356 34546 5408 34552
rect 4988 31884 5040 31890
rect 4908 31844 4988 31872
rect 4988 31826 5040 31832
rect 5080 31816 5132 31822
rect 5080 31758 5132 31764
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5092 31668 5120 31758
rect 5276 31686 5304 31758
rect 5264 31680 5316 31686
rect 4986 31648 5042 31657
rect 5092 31640 5212 31668
rect 4986 31583 5042 31592
rect 4724 31436 4844 31464
rect 4816 31278 4844 31436
rect 4804 31272 4856 31278
rect 4804 31214 4856 31220
rect 4896 31204 4948 31210
rect 4896 31146 4948 31152
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4724 30258 4752 30670
rect 4802 30288 4858 30297
rect 4712 30252 4764 30258
rect 4802 30223 4858 30232
rect 4712 30194 4764 30200
rect 4712 29640 4764 29646
rect 4710 29608 4712 29617
rect 4764 29608 4766 29617
rect 4710 29543 4766 29552
rect 4710 29472 4766 29481
rect 4710 29407 4766 29416
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4632 26314 4660 26862
rect 4434 26279 4490 26288
rect 4528 26308 4580 26314
rect 4342 26072 4398 26081
rect 4342 26007 4398 26016
rect 4448 24177 4476 26279
rect 4528 26250 4580 26256
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 4434 24168 4490 24177
rect 4434 24103 4490 24112
rect 4436 24064 4488 24070
rect 4264 23990 4384 24018
rect 4436 24006 4488 24012
rect 4158 23967 4214 23976
rect 4172 23730 4200 23967
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4066 22264 4122 22273
rect 4066 22199 4122 22208
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 3974 21856 4030 21865
rect 3974 21791 4030 21800
rect 4080 21729 4108 22102
rect 4172 22098 4200 23666
rect 4356 23610 4384 23990
rect 4448 23730 4476 24006
rect 4436 23724 4488 23730
rect 4436 23666 4488 23672
rect 4540 23610 4568 26250
rect 4724 25378 4752 29407
rect 4816 28762 4844 30223
rect 4908 30122 4936 31146
rect 4896 30116 4948 30122
rect 4896 30058 4948 30064
rect 4894 30016 4950 30025
rect 4894 29951 4950 29960
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4804 28484 4856 28490
rect 4804 28426 4856 28432
rect 4816 28393 4844 28426
rect 4802 28384 4858 28393
rect 4802 28319 4858 28328
rect 4804 28144 4856 28150
rect 4804 28086 4856 28092
rect 4816 26246 4844 28086
rect 4908 27470 4936 29951
rect 5000 28994 5028 31583
rect 5184 31210 5212 31640
rect 5264 31622 5316 31628
rect 5262 31512 5318 31521
rect 5262 31447 5318 31456
rect 5172 31204 5224 31210
rect 5172 31146 5224 31152
rect 5080 31136 5132 31142
rect 5080 31078 5132 31084
rect 5092 30394 5120 31078
rect 5080 30388 5132 30394
rect 5080 30330 5132 30336
rect 5172 29708 5224 29714
rect 5172 29650 5224 29656
rect 5184 29306 5212 29650
rect 5172 29300 5224 29306
rect 5172 29242 5224 29248
rect 5000 28966 5120 28994
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 5000 27452 5028 28494
rect 5092 28422 5120 28966
rect 5172 28960 5224 28966
rect 5172 28902 5224 28908
rect 5080 28416 5132 28422
rect 5080 28358 5132 28364
rect 5080 27464 5132 27470
rect 5000 27424 5080 27452
rect 4908 27334 4936 27406
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 4908 26586 4936 26862
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 4894 26480 4950 26489
rect 4894 26415 4896 26424
rect 4948 26415 4950 26424
rect 4896 26386 4948 26392
rect 4804 26240 4856 26246
rect 4804 26182 4856 26188
rect 4908 26194 4936 26386
rect 5000 26382 5028 27424
rect 5080 27406 5132 27412
rect 5184 27316 5212 28902
rect 5092 27288 5212 27316
rect 5092 26586 5120 27288
rect 5276 27062 5304 31447
rect 5368 29850 5396 34546
rect 5460 34542 5488 34614
rect 5448 34536 5500 34542
rect 5448 34478 5500 34484
rect 5460 31793 5488 34478
rect 5552 31958 5580 36230
rect 5632 36100 5684 36106
rect 5632 36042 5684 36048
rect 5644 33289 5672 36042
rect 5630 33280 5686 33289
rect 5630 33215 5686 33224
rect 5632 32020 5684 32026
rect 5632 31962 5684 31968
rect 5540 31952 5592 31958
rect 5540 31894 5592 31900
rect 5446 31784 5502 31793
rect 5644 31754 5672 31962
rect 5446 31719 5502 31728
rect 5552 31726 5672 31754
rect 5448 31680 5500 31686
rect 5448 31622 5500 31628
rect 5460 31278 5488 31622
rect 5448 31272 5500 31278
rect 5448 31214 5500 31220
rect 5356 29844 5408 29850
rect 5356 29786 5408 29792
rect 5356 29708 5408 29714
rect 5356 29650 5408 29656
rect 5368 28762 5396 29650
rect 5460 29617 5488 31214
rect 5552 31142 5580 31726
rect 5632 31204 5684 31210
rect 5632 31146 5684 31152
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5540 30864 5592 30870
rect 5540 30806 5592 30812
rect 5552 29646 5580 30806
rect 5644 29646 5672 31146
rect 5540 29640 5592 29646
rect 5446 29608 5502 29617
rect 5540 29582 5592 29588
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5446 29543 5502 29552
rect 5552 29510 5580 29582
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5540 29504 5592 29510
rect 5540 29446 5592 29452
rect 5356 28756 5408 28762
rect 5356 28698 5408 28704
rect 5460 28626 5488 29446
rect 5538 29200 5594 29209
rect 5538 29135 5594 29144
rect 5448 28620 5500 28626
rect 5448 28562 5500 28568
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5460 28082 5488 28358
rect 5448 28076 5500 28082
rect 5448 28018 5500 28024
rect 5552 27985 5580 29135
rect 5538 27976 5594 27985
rect 5538 27911 5594 27920
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 5172 26988 5224 26994
rect 5172 26930 5224 26936
rect 5080 26580 5132 26586
rect 5080 26522 5132 26528
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 4816 25430 4844 26182
rect 4908 26166 5120 26194
rect 4632 25362 4752 25378
rect 4804 25424 4856 25430
rect 4804 25366 4856 25372
rect 4620 25356 4752 25362
rect 4672 25350 4752 25356
rect 4620 25298 4672 25304
rect 4988 25288 5040 25294
rect 4816 25248 4988 25276
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4632 24070 4660 24686
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4264 23582 4384 23610
rect 4448 23582 4568 23610
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4066 21720 4122 21729
rect 4066 21655 4122 21664
rect 4264 21570 4292 23582
rect 4342 22808 4398 22817
rect 4342 22743 4398 22752
rect 4356 22438 4384 22743
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 3988 21542 4292 21570
rect 3988 21010 4016 21542
rect 4160 21480 4212 21486
rect 4066 21448 4122 21457
rect 4122 21428 4160 21434
rect 4122 21422 4212 21428
rect 4250 21448 4306 21457
rect 4122 21406 4200 21422
rect 4066 21383 4122 21392
rect 4356 21418 4384 22374
rect 4250 21383 4306 21392
rect 4344 21412 4396 21418
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4080 20942 4108 21286
rect 4172 21146 4200 21286
rect 4264 21146 4292 21383
rect 4344 21354 4396 21360
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4252 21140 4304 21146
rect 4252 21082 4304 21088
rect 4356 21078 4384 21354
rect 4344 21072 4396 21078
rect 4344 21014 4396 21020
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3884 20800 3936 20806
rect 3790 20768 3846 20777
rect 4160 20800 4212 20806
rect 3884 20742 3936 20748
rect 3974 20768 4030 20777
rect 3790 20703 3846 20712
rect 4160 20742 4212 20748
rect 3974 20703 4030 20712
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 3620 18958 3740 18986
rect 3712 18834 3740 18958
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3608 18760 3660 18766
rect 3712 18737 3740 18770
rect 3608 18702 3660 18708
rect 3698 18728 3754 18737
rect 3514 17912 3570 17921
rect 3514 17847 3570 17856
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3620 17626 3648 18702
rect 3698 18663 3754 18672
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 3436 17598 3648 17626
rect 3010 17436 3318 17445
rect 3010 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3176 17436
rect 3232 17434 3256 17436
rect 3312 17434 3318 17436
rect 3072 17382 3074 17434
rect 3254 17382 3256 17434
rect 3010 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3176 17382
rect 3232 17380 3256 17382
rect 3312 17380 3318 17382
rect 3010 17371 3318 17380
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 2976 16969 3004 17274
rect 3238 17096 3294 17105
rect 3238 17031 3240 17040
rect 3292 17031 3294 17040
rect 3240 17002 3292 17008
rect 2962 16960 3018 16969
rect 2962 16895 3018 16904
rect 3010 16348 3318 16357
rect 3010 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3176 16348
rect 3232 16346 3256 16348
rect 3312 16346 3318 16348
rect 3072 16294 3074 16346
rect 3254 16294 3256 16346
rect 3010 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3176 16294
rect 3232 16292 3256 16294
rect 3312 16292 3318 16294
rect 3010 16283 3318 16292
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3056 15972 3108 15978
rect 3056 15914 3108 15920
rect 3068 15706 3096 15914
rect 3344 15881 3372 15982
rect 3330 15872 3386 15881
rect 3330 15807 3386 15816
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3010 15260 3318 15269
rect 3010 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3176 15260
rect 3232 15258 3256 15260
rect 3312 15258 3318 15260
rect 3072 15206 3074 15258
rect 3254 15206 3256 15258
rect 3010 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3176 15206
rect 3232 15204 3256 15206
rect 3312 15204 3318 15206
rect 3010 15195 3318 15204
rect 3010 14172 3318 14181
rect 3010 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3176 14172
rect 3232 14170 3256 14172
rect 3312 14170 3318 14172
rect 3072 14118 3074 14170
rect 3254 14118 3256 14170
rect 3010 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3176 14118
rect 3232 14116 3256 14118
rect 3312 14116 3318 14118
rect 3010 14107 3318 14116
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3068 13530 3096 13806
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3010 13084 3318 13093
rect 3010 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3176 13084
rect 3232 13082 3256 13084
rect 3312 13082 3318 13084
rect 3072 13030 3074 13082
rect 3254 13030 3256 13082
rect 3010 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3176 13030
rect 3232 13028 3256 13030
rect 3312 13028 3318 13030
rect 3010 13019 3318 13028
rect 2964 12776 3016 12782
rect 2962 12744 2964 12753
rect 3056 12776 3108 12782
rect 3016 12744 3018 12753
rect 3056 12718 3108 12724
rect 2962 12679 3018 12688
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 3068 12209 3096 12718
rect 3054 12200 3110 12209
rect 2872 12164 2924 12170
rect 3054 12135 3110 12144
rect 2872 12106 2924 12112
rect 2884 11778 2912 12106
rect 3010 11996 3318 12005
rect 3010 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3176 11996
rect 3232 11994 3256 11996
rect 3312 11994 3318 11996
rect 3072 11942 3074 11994
rect 3254 11942 3256 11994
rect 3010 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3176 11942
rect 3232 11940 3256 11942
rect 3312 11940 3318 11942
rect 3010 11931 3318 11940
rect 3054 11792 3110 11801
rect 2884 11750 3004 11778
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2884 11354 2912 11562
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2976 11098 3004 11750
rect 3054 11727 3110 11736
rect 3068 11694 3096 11727
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3068 11257 3096 11630
rect 3054 11248 3110 11257
rect 3252 11218 3280 11630
rect 3054 11183 3110 11192
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 2884 11070 3004 11098
rect 2884 10742 2912 11070
rect 3010 10908 3318 10917
rect 3010 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3176 10908
rect 3232 10906 3256 10908
rect 3312 10906 3318 10908
rect 3072 10854 3074 10906
rect 3254 10854 3256 10906
rect 3010 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3176 10854
rect 3232 10852 3256 10854
rect 3312 10852 3318 10854
rect 3010 10843 3318 10852
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2778 7848 2834 7857
rect 2778 7783 2834 7792
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1596 6458 1716 6474
rect 1596 6452 1728 6458
rect 1596 6446 1676 6452
rect 1676 6394 1728 6400
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5817 1900 6054
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2608 5914 2636 6734
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 1858 5808 1914 5817
rect 1858 5743 1914 5752
rect 1412 5086 1532 5114
rect 1124 4208 1176 4214
rect 1124 4150 1176 4156
rect 1412 56 1440 5086
rect 1492 5024 1544 5030
rect 1490 4992 1492 5001
rect 1544 4992 1546 5001
rect 1490 4927 1546 4936
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1504 4185 1532 4490
rect 1860 4208 1912 4214
rect 1490 4176 1546 4185
rect 1860 4150 1912 4156
rect 1490 4111 1546 4120
rect 1872 56 1900 4150
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2332 56 2360 2382
rect 2700 2106 2728 7142
rect 2792 5234 2820 7783
rect 2884 6458 2912 10406
rect 3010 9820 3318 9829
rect 3010 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3176 9820
rect 3232 9818 3256 9820
rect 3312 9818 3318 9820
rect 3072 9766 3074 9818
rect 3254 9766 3256 9818
rect 3010 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3176 9766
rect 3232 9764 3256 9766
rect 3312 9764 3318 9766
rect 3010 9755 3318 9764
rect 3436 9586 3464 17598
rect 3712 17524 3740 18566
rect 3620 17496 3740 17524
rect 3620 17134 3648 17496
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3608 17128 3660 17134
rect 3514 17096 3570 17105
rect 3608 17070 3660 17076
rect 3514 17031 3570 17040
rect 3528 14362 3556 17031
rect 3620 16289 3648 17070
rect 3606 16280 3662 16289
rect 3606 16215 3662 16224
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3620 15162 3648 16050
rect 3608 15156 3660 15162
rect 3608 15098 3660 15104
rect 3528 14334 3648 14362
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3528 13870 3556 14214
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3528 12986 3556 13670
rect 3620 13258 3648 14334
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3712 12434 3740 17274
rect 3804 15162 3832 20538
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 3896 19689 3924 20402
rect 3882 19680 3938 19689
rect 3882 19615 3938 19624
rect 3884 18896 3936 18902
rect 3882 18864 3884 18873
rect 3936 18864 3938 18873
rect 3882 18799 3938 18808
rect 3882 18592 3938 18601
rect 3882 18527 3938 18536
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3790 14784 3846 14793
rect 3896 14770 3924 18527
rect 3988 18057 4016 20703
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 19310 4108 19654
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3974 18048 4030 18057
rect 3974 17983 4030 17992
rect 4080 15706 4108 19110
rect 4172 16454 4200 20742
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4264 16046 4292 20946
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4356 18970 4384 19314
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4448 18850 4476 23582
rect 4632 23526 4660 24006
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4526 23352 4582 23361
rect 4724 23322 4752 24686
rect 4526 23287 4582 23296
rect 4712 23316 4764 23322
rect 4540 22166 4568 23287
rect 4712 23258 4764 23264
rect 4816 23202 4844 25248
rect 4988 25230 5040 25236
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4724 23174 4844 23202
rect 4632 22710 4660 23122
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4528 22160 4580 22166
rect 4528 22102 4580 22108
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4540 21026 4568 21966
rect 4632 21554 4660 22646
rect 4724 21570 4752 23174
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4816 22030 4844 22986
rect 4804 22024 4856 22030
rect 4908 22001 4936 24278
rect 5000 22642 5028 24890
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 4804 21966 4856 21972
rect 4894 21992 4950 22001
rect 4816 21865 4844 21966
rect 4894 21927 4950 21936
rect 5000 21876 5028 22442
rect 4802 21856 4858 21865
rect 4802 21791 4858 21800
rect 4908 21848 5028 21876
rect 4724 21554 4844 21570
rect 4620 21548 4672 21554
rect 4724 21548 4856 21554
rect 4724 21542 4804 21548
rect 4620 21490 4672 21496
rect 4804 21490 4856 21496
rect 4710 21312 4766 21321
rect 4710 21247 4766 21256
rect 4540 20998 4660 21026
rect 4528 20868 4580 20874
rect 4528 20810 4580 20816
rect 4540 20058 4568 20810
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4632 19394 4660 20998
rect 4356 18822 4476 18850
rect 4540 19366 4660 19394
rect 4356 17338 4384 18822
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4448 18154 4476 18702
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4172 15201 4200 15846
rect 4264 15745 4292 15982
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4250 15736 4306 15745
rect 4250 15671 4306 15680
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4158 15192 4214 15201
rect 4158 15127 4214 15136
rect 3846 14742 3924 14770
rect 3790 14719 3846 14728
rect 3804 13938 3832 14719
rect 4264 14618 4292 15506
rect 4356 15502 4384 15846
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4448 15366 4476 15982
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4158 14376 4214 14385
rect 3884 14340 3936 14346
rect 4158 14311 4214 14320
rect 3884 14282 3936 14288
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3804 13138 3832 13874
rect 3896 13258 3924 14282
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4080 13938 4108 14010
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3804 13110 4016 13138
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3620 12406 3740 12434
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5914 3096 6054
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5302 2912 5646
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 3436 5030 3464 8434
rect 3528 6322 3556 11834
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3620 2650 3648 12406
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3712 10742 3740 12174
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3698 9752 3754 9761
rect 3698 9687 3754 9696
rect 3712 9654 3740 9687
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3804 8786 3832 12922
rect 3884 12776 3936 12782
rect 3988 12764 4016 13110
rect 3936 12736 4016 12764
rect 3884 12718 3936 12724
rect 3988 11762 4016 12736
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4080 12050 4108 12679
rect 4172 12238 4200 14311
rect 4252 13864 4304 13870
rect 4356 13818 4384 14486
rect 4304 13812 4384 13818
rect 4252 13806 4384 13812
rect 4264 13790 4384 13806
rect 4264 13190 4292 13790
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 4080 12022 4200 12050
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4080 11762 4108 11834
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4172 11642 4200 12022
rect 4264 11898 4292 13126
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4080 11614 4200 11642
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3712 8758 3832 8786
rect 3712 5370 3740 8758
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3804 5234 3832 5510
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3896 2650 3924 9658
rect 3988 7274 4016 11290
rect 4080 10418 4108 11614
rect 4356 11506 4384 13194
rect 4448 12434 4476 15098
rect 4540 14550 4568 19366
rect 4724 19310 4752 21247
rect 4816 20942 4844 21490
rect 4804 20936 4856 20942
rect 4802 20904 4804 20913
rect 4856 20904 4858 20913
rect 4802 20839 4858 20848
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4632 18816 4660 19246
rect 4724 18970 4752 19246
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4607 18788 4660 18816
rect 4712 18828 4764 18834
rect 4607 18306 4635 18788
rect 4816 18816 4844 19178
rect 4764 18788 4844 18816
rect 4712 18770 4764 18776
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4607 18278 4660 18306
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 14074 4568 14350
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4448 12406 4568 12434
rect 4540 12050 4568 12406
rect 4632 12288 4660 18278
rect 4724 12986 4752 18566
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4816 12850 4844 18022
rect 4908 16697 4936 21848
rect 4986 21720 5042 21729
rect 4986 21655 5042 21664
rect 5000 21554 5028 21655
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 5092 21298 5120 26166
rect 5184 25294 5212 26930
rect 5276 26489 5304 26998
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5262 26480 5318 26489
rect 5262 26415 5318 26424
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5262 25120 5318 25129
rect 5262 25055 5318 25064
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5184 23730 5212 24550
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5000 21270 5120 21298
rect 5000 16810 5028 21270
rect 5078 21176 5134 21185
rect 5078 21111 5080 21120
rect 5132 21111 5134 21120
rect 5080 21082 5132 21088
rect 5184 20806 5212 22578
rect 5276 22574 5304 25055
rect 5368 24342 5396 26726
rect 5460 25294 5488 27270
rect 5552 25401 5580 27610
rect 5644 26625 5672 29582
rect 5736 26790 5764 37130
rect 5828 35018 5856 37674
rect 5920 35494 5948 37878
rect 6012 36242 6040 41618
rect 6196 41274 6224 42162
rect 6564 41818 6592 42162
rect 6748 41818 6776 42502
rect 6932 42362 6960 44944
rect 7392 42362 7420 44944
rect 7852 43518 7880 44944
rect 7840 43512 7892 43518
rect 7840 43454 7892 43460
rect 6920 42356 6972 42362
rect 6920 42298 6972 42304
rect 7380 42356 7432 42362
rect 7380 42298 7432 42304
rect 7196 42288 7248 42294
rect 7196 42230 7248 42236
rect 6920 42016 6972 42022
rect 6920 41958 6972 41964
rect 7012 42016 7064 42022
rect 7012 41958 7064 41964
rect 6552 41812 6604 41818
rect 6552 41754 6604 41760
rect 6736 41812 6788 41818
rect 6736 41754 6788 41760
rect 6932 41274 6960 41958
rect 7024 41614 7052 41958
rect 7012 41608 7064 41614
rect 7012 41550 7064 41556
rect 6184 41268 6236 41274
rect 6184 41210 6236 41216
rect 6920 41268 6972 41274
rect 6920 41210 6972 41216
rect 7024 41138 7052 41550
rect 6828 41132 6880 41138
rect 6828 41074 6880 41080
rect 7012 41132 7064 41138
rect 7012 41074 7064 41080
rect 6840 40390 6868 41074
rect 7024 41041 7052 41074
rect 7010 41032 7066 41041
rect 7010 40967 7066 40976
rect 7208 40730 7236 42230
rect 7472 42220 7524 42226
rect 7472 42162 7524 42168
rect 7840 42220 7892 42226
rect 7840 42162 7892 42168
rect 7380 42084 7432 42090
rect 7380 42026 7432 42032
rect 7288 42016 7340 42022
rect 7288 41958 7340 41964
rect 7196 40724 7248 40730
rect 7196 40666 7248 40672
rect 6828 40384 6880 40390
rect 6828 40326 6880 40332
rect 6276 38752 6328 38758
rect 6276 38694 6328 38700
rect 6184 38344 6236 38350
rect 6184 38286 6236 38292
rect 6196 38010 6224 38286
rect 6184 38004 6236 38010
rect 6184 37946 6236 37952
rect 6092 37392 6144 37398
rect 6092 37334 6144 37340
rect 6000 36236 6052 36242
rect 6000 36178 6052 36184
rect 6104 35850 6132 37334
rect 6184 36100 6236 36106
rect 6184 36042 6236 36048
rect 6012 35822 6132 35850
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 5816 35012 5868 35018
rect 5816 34954 5868 34960
rect 5828 34898 5856 34954
rect 5828 34870 5948 34898
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5828 30598 5856 31826
rect 5816 30592 5868 30598
rect 5816 30534 5868 30540
rect 5816 29504 5868 29510
rect 5816 29446 5868 29452
rect 5828 28370 5856 29446
rect 5920 28490 5948 34870
rect 6012 33017 6040 35822
rect 6092 35012 6144 35018
rect 6092 34954 6144 34960
rect 6104 34406 6132 34954
rect 6092 34400 6144 34406
rect 6092 34342 6144 34348
rect 5998 33008 6054 33017
rect 5998 32943 6054 32952
rect 6092 32224 6144 32230
rect 6092 32166 6144 32172
rect 6000 31816 6052 31822
rect 5998 31784 6000 31793
rect 6052 31784 6054 31793
rect 5998 31719 6054 31728
rect 6000 31476 6052 31482
rect 6000 31418 6052 31424
rect 6012 30938 6040 31418
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 6104 30546 6132 32166
rect 6196 30920 6224 36042
rect 6288 35193 6316 38694
rect 6460 38412 6512 38418
rect 6460 38354 6512 38360
rect 6368 37868 6420 37874
rect 6368 37810 6420 37816
rect 6380 37466 6408 37810
rect 6368 37460 6420 37466
rect 6368 37402 6420 37408
rect 6472 37233 6500 38354
rect 6644 38208 6696 38214
rect 6644 38150 6696 38156
rect 6458 37224 6514 37233
rect 6458 37159 6514 37168
rect 6552 37188 6604 37194
rect 6552 37130 6604 37136
rect 6366 35592 6422 35601
rect 6366 35527 6422 35536
rect 6274 35184 6330 35193
rect 6274 35119 6330 35128
rect 6276 34672 6328 34678
rect 6276 34614 6328 34620
rect 6288 34542 6316 34614
rect 6276 34536 6328 34542
rect 6276 34478 6328 34484
rect 6276 32836 6328 32842
rect 6276 32778 6328 32784
rect 6288 31090 6316 32778
rect 6380 32552 6408 35527
rect 6460 35284 6512 35290
rect 6460 35226 6512 35232
rect 6472 33674 6500 35226
rect 6564 34746 6592 37130
rect 6656 35018 6684 38150
rect 6736 36304 6788 36310
rect 6736 36246 6788 36252
rect 6748 35222 6776 36246
rect 6736 35216 6788 35222
rect 6736 35158 6788 35164
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 6644 35012 6696 35018
rect 6644 34954 6696 34960
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 6644 34604 6696 34610
rect 6644 34546 6696 34552
rect 6656 33998 6684 34546
rect 6748 34406 6776 35022
rect 6840 34513 6868 40326
rect 7012 37800 7064 37806
rect 7012 37742 7064 37748
rect 6920 37664 6972 37670
rect 6920 37606 6972 37612
rect 6932 36786 6960 37606
rect 6920 36780 6972 36786
rect 6920 36722 6972 36728
rect 7024 35834 7052 37742
rect 7104 36168 7156 36174
rect 7104 36110 7156 36116
rect 7012 35828 7064 35834
rect 7012 35770 7064 35776
rect 6920 35692 6972 35698
rect 6920 35634 6972 35640
rect 6932 34950 6960 35634
rect 7012 35556 7064 35562
rect 7012 35498 7064 35504
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 6932 34678 6960 34886
rect 6920 34672 6972 34678
rect 6920 34614 6972 34620
rect 6920 34536 6972 34542
rect 6826 34504 6882 34513
rect 6920 34478 6972 34484
rect 6826 34439 6882 34448
rect 6736 34400 6788 34406
rect 6932 34388 6960 34478
rect 6736 34342 6788 34348
rect 6840 34360 6960 34388
rect 6840 34241 6868 34360
rect 6826 34232 6882 34241
rect 6736 34196 6788 34202
rect 6826 34167 6882 34176
rect 6736 34138 6788 34144
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 6472 33646 6684 33674
rect 6552 33380 6604 33386
rect 6552 33322 6604 33328
rect 6564 32978 6592 33322
rect 6552 32972 6604 32978
rect 6552 32914 6604 32920
rect 6380 32524 6500 32552
rect 6472 31414 6500 32524
rect 6552 32428 6604 32434
rect 6552 32370 6604 32376
rect 6460 31408 6512 31414
rect 6460 31350 6512 31356
rect 6288 31062 6500 31090
rect 6196 30892 6408 30920
rect 6184 30796 6236 30802
rect 6184 30738 6236 30744
rect 6012 30518 6132 30546
rect 5908 28484 5960 28490
rect 5908 28426 5960 28432
rect 5828 28342 5948 28370
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5828 28082 5856 28154
rect 5816 28076 5868 28082
rect 5816 28018 5868 28024
rect 5828 27674 5856 28018
rect 5816 27668 5868 27674
rect 5816 27610 5868 27616
rect 5724 26784 5776 26790
rect 5724 26726 5776 26732
rect 5816 26784 5868 26790
rect 5816 26726 5868 26732
rect 5630 26616 5686 26625
rect 5828 26602 5856 26726
rect 5630 26551 5686 26560
rect 5736 26574 5856 26602
rect 5632 26512 5684 26518
rect 5736 26500 5764 26574
rect 5684 26472 5764 26500
rect 5632 26454 5684 26460
rect 5920 26432 5948 28342
rect 6012 27674 6040 30518
rect 6090 30424 6146 30433
rect 6090 30359 6146 30368
rect 6000 27668 6052 27674
rect 6000 27610 6052 27616
rect 6104 26625 6132 30359
rect 6196 29714 6224 30738
rect 6276 30660 6328 30666
rect 6276 30602 6328 30608
rect 6184 29708 6236 29714
rect 6184 29650 6236 29656
rect 6196 29345 6224 29650
rect 6182 29336 6238 29345
rect 6182 29271 6238 29280
rect 6196 28626 6224 29271
rect 6184 28620 6236 28626
rect 6184 28562 6236 28568
rect 6196 28082 6224 28562
rect 6184 28076 6236 28082
rect 6184 28018 6236 28024
rect 6288 27441 6316 30602
rect 6274 27432 6330 27441
rect 6274 27367 6330 27376
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6090 26616 6146 26625
rect 6090 26551 6146 26560
rect 6288 26450 6316 27270
rect 5736 26404 5948 26432
rect 6276 26444 6328 26450
rect 5630 26208 5686 26217
rect 5630 26143 5686 26152
rect 5538 25392 5594 25401
rect 5538 25327 5594 25336
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5460 24954 5488 25230
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5356 24336 5408 24342
rect 5356 24278 5408 24284
rect 5460 23866 5488 24754
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5448 23588 5500 23594
rect 5448 23530 5500 23536
rect 5356 22976 5408 22982
rect 5356 22918 5408 22924
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5276 22166 5304 22374
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5368 22012 5396 22918
rect 5276 21984 5396 22012
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5184 19854 5212 20266
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5080 18896 5132 18902
rect 5172 18896 5224 18902
rect 5080 18838 5132 18844
rect 5170 18864 5172 18873
rect 5224 18864 5226 18873
rect 5092 17338 5120 18838
rect 5170 18799 5226 18808
rect 5172 17604 5224 17610
rect 5172 17546 5224 17552
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5078 17096 5134 17105
rect 5078 17031 5080 17040
rect 5132 17031 5134 17040
rect 5080 17002 5132 17008
rect 5000 16794 5120 16810
rect 5000 16788 5132 16794
rect 5000 16782 5080 16788
rect 5080 16730 5132 16736
rect 4894 16688 4950 16697
rect 4894 16623 4950 16632
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 16046 5028 16390
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12442 4752 12650
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4712 12300 4764 12306
rect 4632 12260 4712 12288
rect 4764 12260 4844 12288
rect 4712 12242 4764 12248
rect 4540 12022 4660 12050
rect 4526 11928 4582 11937
rect 4526 11863 4582 11872
rect 4172 11478 4384 11506
rect 4172 11286 4200 11478
rect 4250 11384 4306 11393
rect 4250 11319 4306 11328
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4080 10390 4200 10418
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4080 10062 4108 10202
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4172 9874 4200 10390
rect 4080 9846 4200 9874
rect 4080 8498 4108 9846
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 4080 6662 4108 8298
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 7410 4200 8230
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4264 7290 4292 11319
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4172 7262 4292 7290
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4080 6254 4108 6394
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4172 5914 4200 7262
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4172 5710 4200 5850
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4264 4758 4292 5646
rect 4356 5098 4384 11222
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 6866 4476 11086
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4540 5370 4568 11863
rect 4632 11540 4660 12022
rect 4712 11552 4764 11558
rect 4632 11512 4712 11540
rect 4712 11494 4764 11500
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4724 9722 4752 9998
rect 4816 9897 4844 12260
rect 4908 11626 4936 15982
rect 4988 15904 5040 15910
rect 4986 15872 4988 15881
rect 5040 15872 5042 15881
rect 4986 15807 5042 15816
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5000 13705 5028 15438
rect 5184 15026 5212 17546
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5092 13938 5120 14282
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4986 13696 5042 13705
rect 4986 13631 5042 13640
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 4908 11150 4936 11562
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4908 9994 4936 10542
rect 5000 10266 5028 13330
rect 5092 12170 5120 13874
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 5092 10742 5120 11086
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4802 9888 4858 9897
rect 4802 9823 4858 9832
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4816 9654 4844 9823
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4618 9480 4674 9489
rect 4816 9466 4844 9590
rect 4908 9489 4936 9930
rect 5000 9586 5028 9930
rect 5092 9586 5120 10134
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4618 9415 4674 9424
rect 4724 9438 4844 9466
rect 4894 9480 4950 9489
rect 4632 9382 4660 9415
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4724 8820 4752 9438
rect 4894 9415 4950 9424
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4804 9376 4856 9382
rect 5092 9353 5120 9386
rect 4804 9318 4856 9324
rect 5078 9344 5134 9353
rect 4816 8974 4844 9318
rect 5078 9279 5134 9288
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4724 8792 4844 8820
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4618 7440 4674 7449
rect 4618 7375 4674 7384
rect 4632 7274 4660 7375
rect 4724 7342 4752 8366
rect 4816 8022 4844 8792
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 5184 7834 5212 12582
rect 5276 12374 5304 21984
rect 5460 21894 5488 23530
rect 5552 22216 5580 23802
rect 5644 22574 5672 26143
rect 5736 24052 5764 26404
rect 6000 26392 6052 26398
rect 5828 26353 6000 26364
rect 5814 26344 6000 26353
rect 5870 26340 6000 26344
rect 5870 26336 6052 26340
rect 6000 26334 6052 26336
rect 6092 26392 6144 26398
rect 6276 26386 6328 26392
rect 6092 26334 6144 26340
rect 5814 26279 5870 26288
rect 6104 26042 6132 26334
rect 6182 26208 6238 26217
rect 6182 26143 6238 26152
rect 6092 26036 6144 26042
rect 6092 25978 6144 25984
rect 5816 25152 5868 25158
rect 5816 25094 5868 25100
rect 5828 24206 5856 25094
rect 5906 24984 5962 24993
rect 5906 24919 5962 24928
rect 5816 24200 5868 24206
rect 5816 24142 5868 24148
rect 5736 24024 5856 24052
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 5552 22188 5672 22216
rect 5644 22098 5672 22188
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5632 22092 5684 22098
rect 5736 22094 5764 23054
rect 5828 22522 5856 24024
rect 5920 24018 5948 24919
rect 6196 24154 6224 26143
rect 6276 25968 6328 25974
rect 6276 25910 6328 25916
rect 6288 25401 6316 25910
rect 6274 25392 6330 25401
rect 6274 25327 6330 25336
rect 6276 24676 6328 24682
rect 6276 24618 6328 24624
rect 6288 24342 6316 24618
rect 6276 24336 6328 24342
rect 6276 24278 6328 24284
rect 6104 24126 6224 24154
rect 5920 23990 6040 24018
rect 5906 23896 5962 23905
rect 5906 23831 5962 23840
rect 5920 23730 5948 23831
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 6012 23089 6040 23990
rect 5998 23080 6054 23089
rect 5998 23015 6054 23024
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 6012 22642 6040 22918
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5828 22494 6040 22522
rect 5736 22066 5948 22094
rect 5632 22034 5684 22040
rect 5552 21978 5580 22034
rect 5816 22024 5868 22030
rect 5552 21950 5672 21978
rect 5816 21966 5868 21972
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5446 21720 5502 21729
rect 5446 21655 5448 21664
rect 5500 21655 5502 21664
rect 5448 21626 5500 21632
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5368 18737 5396 21422
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5552 19334 5580 21354
rect 5460 19306 5580 19334
rect 5354 18728 5410 18737
rect 5354 18663 5410 18672
rect 5368 18086 5396 18663
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5460 16969 5488 19306
rect 5538 17912 5594 17921
rect 5538 17847 5594 17856
rect 5446 16960 5502 16969
rect 5446 16895 5502 16904
rect 5552 16810 5580 17847
rect 5368 16782 5580 16810
rect 5368 15586 5396 16782
rect 5540 16652 5592 16658
rect 5460 16612 5540 16640
rect 5460 15706 5488 16612
rect 5540 16594 5592 16600
rect 5540 16108 5592 16114
rect 5540 16050 5592 16056
rect 5552 16017 5580 16050
rect 5538 16008 5594 16017
rect 5538 15943 5594 15952
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5368 15558 5488 15586
rect 5354 15056 5410 15065
rect 5354 14991 5410 15000
rect 5368 13938 5396 14991
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5460 12481 5488 15558
rect 5552 15434 5580 15846
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5446 12472 5502 12481
rect 5552 12442 5580 14214
rect 5644 12782 5672 21950
rect 5828 21865 5856 21966
rect 5814 21856 5870 21865
rect 5814 21791 5870 21800
rect 5920 21706 5948 22066
rect 5736 21678 5948 21706
rect 5736 16726 5764 21678
rect 6012 21604 6040 22494
rect 5920 21576 6040 21604
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 5828 21457 5856 21490
rect 5814 21448 5870 21457
rect 5814 21383 5870 21392
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5828 18766 5856 20742
rect 5920 19174 5948 21576
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5906 19000 5962 19009
rect 5906 18935 5908 18944
rect 5960 18935 5962 18944
rect 5908 18906 5960 18912
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5736 15745 5764 15982
rect 5722 15736 5778 15745
rect 5722 15671 5778 15680
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5736 12986 5764 15574
rect 5828 14414 5856 18702
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5632 12776 5684 12782
rect 5828 12753 5856 14214
rect 5920 13258 5948 18770
rect 6012 17678 6040 19790
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 16250 6040 17614
rect 6104 16561 6132 24126
rect 6288 23662 6316 24278
rect 6380 23798 6408 30892
rect 6472 30734 6500 31062
rect 6460 30728 6512 30734
rect 6460 30670 6512 30676
rect 6460 30252 6512 30258
rect 6460 30194 6512 30200
rect 6472 29850 6500 30194
rect 6460 29844 6512 29850
rect 6460 29786 6512 29792
rect 6458 28928 6514 28937
rect 6458 28863 6514 28872
rect 6472 27130 6500 28863
rect 6564 28665 6592 32370
rect 6550 28656 6606 28665
rect 6550 28591 6606 28600
rect 6552 28484 6604 28490
rect 6552 28426 6604 28432
rect 6460 27124 6512 27130
rect 6460 27066 6512 27072
rect 6460 26852 6512 26858
rect 6460 26794 6512 26800
rect 6472 24410 6500 26794
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6368 23792 6420 23798
rect 6368 23734 6420 23740
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6288 23089 6316 23598
rect 6368 23180 6420 23186
rect 6368 23122 6420 23128
rect 6274 23080 6330 23089
rect 6274 23015 6330 23024
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6288 22817 6316 22918
rect 6274 22808 6330 22817
rect 6380 22778 6408 23122
rect 6274 22743 6330 22752
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6196 18426 6224 22374
rect 6288 20874 6316 22646
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6276 20868 6328 20874
rect 6276 20810 6328 20816
rect 6380 20641 6408 22510
rect 6472 21146 6500 24006
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6366 20632 6422 20641
rect 6366 20567 6422 20576
rect 6276 20528 6328 20534
rect 6276 20470 6328 20476
rect 6288 19378 6316 20470
rect 6472 20466 6500 20946
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6380 19922 6408 20334
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6366 19816 6422 19825
rect 6366 19751 6422 19760
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6288 18034 6316 19314
rect 6380 18873 6408 19751
rect 6472 19718 6500 20402
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6366 18864 6422 18873
rect 6366 18799 6422 18808
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6380 18154 6408 18702
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6196 18006 6316 18034
rect 6196 16658 6224 18006
rect 6274 17912 6330 17921
rect 6274 17847 6276 17856
rect 6328 17847 6330 17856
rect 6276 17818 6328 17824
rect 6380 17746 6408 18090
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6380 16590 6408 17682
rect 6472 17678 6500 19654
rect 6564 18290 6592 28426
rect 6656 24614 6684 33646
rect 6748 32910 6776 34138
rect 6840 34134 6868 34167
rect 6828 34128 6880 34134
rect 6828 34070 6880 34076
rect 6736 32904 6788 32910
rect 6734 32872 6736 32881
rect 6788 32872 6790 32881
rect 6734 32807 6790 32816
rect 6840 32366 6868 34070
rect 6920 33652 6972 33658
rect 6920 33594 6972 33600
rect 6828 32360 6880 32366
rect 6828 32302 6880 32308
rect 6840 31890 6868 32302
rect 6828 31884 6880 31890
rect 6828 31826 6880 31832
rect 6932 31754 6960 33594
rect 7024 32178 7052 35498
rect 7116 35086 7144 36110
rect 7196 35216 7248 35222
rect 7196 35158 7248 35164
rect 7104 35080 7156 35086
rect 7104 35022 7156 35028
rect 7116 33114 7144 35022
rect 7104 33108 7156 33114
rect 7104 33050 7156 33056
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7116 32337 7144 32846
rect 7102 32328 7158 32337
rect 7102 32263 7158 32272
rect 7024 32150 7144 32178
rect 7010 32056 7066 32065
rect 7010 31991 7066 32000
rect 6748 31726 6960 31754
rect 6748 29492 6776 31726
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6840 29646 6868 30126
rect 6828 29640 6880 29646
rect 6828 29582 6880 29588
rect 6748 29464 6868 29492
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6748 25906 6776 28358
rect 6840 28218 6868 29464
rect 6828 28212 6880 28218
rect 6828 28154 6880 28160
rect 6932 28150 6960 31350
rect 7024 28234 7052 31991
rect 7116 30258 7144 32150
rect 7208 31793 7236 35158
rect 7300 34377 7328 41958
rect 7392 41274 7420 42026
rect 7484 41818 7512 42162
rect 7748 42016 7800 42022
rect 7748 41958 7800 41964
rect 7472 41812 7524 41818
rect 7472 41754 7524 41760
rect 7760 41698 7788 41958
rect 7852 41818 7880 42162
rect 8312 42090 8340 44944
rect 8392 43512 8444 43518
rect 8392 43454 8444 43460
rect 8404 42362 8432 43454
rect 8772 42362 8800 44944
rect 9232 42566 9260 44944
rect 9220 42560 9272 42566
rect 9220 42502 9272 42508
rect 9010 42460 9318 42469
rect 9010 42458 9016 42460
rect 9072 42458 9096 42460
rect 9152 42458 9176 42460
rect 9232 42458 9256 42460
rect 9312 42458 9318 42460
rect 9072 42406 9074 42458
rect 9254 42406 9256 42458
rect 9010 42404 9016 42406
rect 9072 42404 9096 42406
rect 9152 42404 9176 42406
rect 9232 42404 9256 42406
rect 9312 42404 9318 42406
rect 9010 42395 9318 42404
rect 8392 42356 8444 42362
rect 8392 42298 8444 42304
rect 8760 42356 8812 42362
rect 8760 42298 8812 42304
rect 8484 42288 8536 42294
rect 8484 42230 8536 42236
rect 8300 42084 8352 42090
rect 8300 42026 8352 42032
rect 7950 41916 8258 41925
rect 7950 41914 7956 41916
rect 8012 41914 8036 41916
rect 8092 41914 8116 41916
rect 8172 41914 8196 41916
rect 8252 41914 8258 41916
rect 8012 41862 8014 41914
rect 8194 41862 8196 41914
rect 7950 41860 7956 41862
rect 8012 41860 8036 41862
rect 8092 41860 8116 41862
rect 8172 41860 8196 41862
rect 8252 41860 8258 41862
rect 7950 41851 8258 41860
rect 7840 41812 7892 41818
rect 7840 41754 7892 41760
rect 7760 41670 8156 41698
rect 8128 41614 8156 41670
rect 8392 41676 8444 41682
rect 8392 41618 8444 41624
rect 8024 41608 8076 41614
rect 8024 41550 8076 41556
rect 8116 41608 8168 41614
rect 8116 41550 8168 41556
rect 8036 41274 8064 41550
rect 7380 41268 7432 41274
rect 7380 41210 7432 41216
rect 8024 41268 8076 41274
rect 8024 41210 8076 41216
rect 7748 41132 7800 41138
rect 7748 41074 7800 41080
rect 7840 41132 7892 41138
rect 7840 41074 7892 41080
rect 8300 41132 8352 41138
rect 8300 41074 8352 41080
rect 7380 40520 7432 40526
rect 7380 40462 7432 40468
rect 7392 39846 7420 40462
rect 7472 40452 7524 40458
rect 7472 40394 7524 40400
rect 7380 39840 7432 39846
rect 7380 39782 7432 39788
rect 7392 39545 7420 39782
rect 7378 39536 7434 39545
rect 7378 39471 7434 39480
rect 7484 37398 7512 40394
rect 7760 40390 7788 41074
rect 7852 40458 7880 41074
rect 7950 40828 8258 40837
rect 7950 40826 7956 40828
rect 8012 40826 8036 40828
rect 8092 40826 8116 40828
rect 8172 40826 8196 40828
rect 8252 40826 8258 40828
rect 8012 40774 8014 40826
rect 8194 40774 8196 40826
rect 7950 40772 7956 40774
rect 8012 40772 8036 40774
rect 8092 40772 8116 40774
rect 8172 40772 8196 40774
rect 8252 40772 8258 40774
rect 7950 40763 8258 40772
rect 7840 40452 7892 40458
rect 7840 40394 7892 40400
rect 8312 40390 8340 41074
rect 8404 40730 8432 41618
rect 8496 41002 8524 42230
rect 8576 42220 8628 42226
rect 8576 42162 8628 42168
rect 8588 41414 8616 42162
rect 8760 42152 8812 42158
rect 8760 42094 8812 42100
rect 9496 42152 9548 42158
rect 9496 42094 9548 42100
rect 8588 41386 8708 41414
rect 8484 40996 8536 41002
rect 8484 40938 8536 40944
rect 8576 40928 8628 40934
rect 8576 40870 8628 40876
rect 8392 40724 8444 40730
rect 8392 40666 8444 40672
rect 7748 40384 7800 40390
rect 7746 40352 7748 40361
rect 8300 40384 8352 40390
rect 7800 40352 7802 40361
rect 8300 40326 8352 40332
rect 7746 40287 7802 40296
rect 7950 39740 8258 39749
rect 7950 39738 7956 39740
rect 8012 39738 8036 39740
rect 8092 39738 8116 39740
rect 8172 39738 8196 39740
rect 8252 39738 8258 39740
rect 8012 39686 8014 39738
rect 8194 39686 8196 39738
rect 7950 39684 7956 39686
rect 8012 39684 8036 39686
rect 8092 39684 8116 39686
rect 8172 39684 8196 39686
rect 8252 39684 8258 39686
rect 7950 39675 8258 39684
rect 7950 38652 8258 38661
rect 7950 38650 7956 38652
rect 8012 38650 8036 38652
rect 8092 38650 8116 38652
rect 8172 38650 8196 38652
rect 8252 38650 8258 38652
rect 8012 38598 8014 38650
rect 8194 38598 8196 38650
rect 7950 38596 7956 38598
rect 8012 38596 8036 38598
rect 8092 38596 8116 38598
rect 8172 38596 8196 38598
rect 8252 38596 8258 38598
rect 7950 38587 8258 38596
rect 7840 38208 7892 38214
rect 7840 38150 7892 38156
rect 7472 37392 7524 37398
rect 7472 37334 7524 37340
rect 7380 37324 7432 37330
rect 7380 37266 7432 37272
rect 7564 37324 7616 37330
rect 7564 37266 7616 37272
rect 7286 34368 7342 34377
rect 7286 34303 7342 34312
rect 7288 33448 7340 33454
rect 7288 33390 7340 33396
rect 7194 31784 7250 31793
rect 7194 31719 7250 31728
rect 7196 31680 7248 31686
rect 7196 31622 7248 31628
rect 7208 30734 7236 31622
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7208 30297 7236 30670
rect 7194 30288 7250 30297
rect 7104 30252 7156 30258
rect 7194 30223 7250 30232
rect 7104 30194 7156 30200
rect 7116 29170 7144 30194
rect 7196 29844 7248 29850
rect 7196 29786 7248 29792
rect 7208 29238 7236 29786
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7104 29164 7156 29170
rect 7104 29106 7156 29112
rect 7104 29028 7156 29034
rect 7156 28976 7236 28994
rect 7104 28970 7236 28976
rect 7116 28966 7236 28970
rect 7208 28665 7236 28966
rect 7194 28656 7250 28665
rect 7194 28591 7250 28600
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 7116 28393 7144 28494
rect 7102 28384 7158 28393
rect 7102 28319 7158 28328
rect 7024 28206 7236 28234
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6840 25786 6868 27814
rect 6918 27568 6974 27577
rect 6918 27503 6974 27512
rect 6932 27334 6960 27503
rect 7012 27464 7064 27470
rect 7012 27406 7064 27412
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 6932 26586 6960 26930
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6748 25758 6868 25786
rect 6748 24954 6776 25758
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6736 24948 6788 24954
rect 6736 24890 6788 24896
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6656 21321 6684 24142
rect 6736 23792 6788 23798
rect 6736 23734 6788 23740
rect 6748 23202 6776 23734
rect 6840 23322 6868 25638
rect 6932 25294 6960 26318
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6932 24342 6960 25094
rect 6920 24336 6972 24342
rect 6920 24278 6972 24284
rect 6918 24168 6974 24177
rect 6918 24103 6974 24112
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6748 23174 6868 23202
rect 6734 22672 6790 22681
rect 6734 22607 6736 22616
rect 6788 22607 6790 22616
rect 6736 22578 6788 22584
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6748 22234 6776 22374
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 6840 22094 6868 23174
rect 6932 22420 6960 24103
rect 7024 23186 7052 27406
rect 7104 27396 7156 27402
rect 7104 27338 7156 27344
rect 7116 25945 7144 27338
rect 7102 25936 7158 25945
rect 7102 25871 7158 25880
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7116 24993 7144 25230
rect 7102 24984 7158 24993
rect 7208 24954 7236 28206
rect 7300 25906 7328 33390
rect 7392 32065 7420 37266
rect 7576 37233 7604 37266
rect 7562 37224 7618 37233
rect 7562 37159 7618 37168
rect 7852 36786 7880 38150
rect 7950 37564 8258 37573
rect 7950 37562 7956 37564
rect 8012 37562 8036 37564
rect 8092 37562 8116 37564
rect 8172 37562 8196 37564
rect 8252 37562 8258 37564
rect 8012 37510 8014 37562
rect 8194 37510 8196 37562
rect 7950 37508 7956 37510
rect 8012 37508 8036 37510
rect 8092 37508 8116 37510
rect 8172 37508 8196 37510
rect 8252 37508 8258 37510
rect 7950 37499 8258 37508
rect 7840 36780 7892 36786
rect 7840 36722 7892 36728
rect 7656 36712 7708 36718
rect 7562 36680 7618 36689
rect 8116 36712 8168 36718
rect 7656 36654 7708 36660
rect 8114 36680 8116 36689
rect 8168 36680 8170 36689
rect 7562 36615 7618 36624
rect 7472 36100 7524 36106
rect 7472 36042 7524 36048
rect 7484 35562 7512 36042
rect 7472 35556 7524 35562
rect 7472 35498 7524 35504
rect 7576 35442 7604 36615
rect 7668 35612 7696 36654
rect 8114 36615 8170 36624
rect 7950 36476 8258 36485
rect 7950 36474 7956 36476
rect 8012 36474 8036 36476
rect 8092 36474 8116 36476
rect 8172 36474 8196 36476
rect 8252 36474 8258 36476
rect 8012 36422 8014 36474
rect 8194 36422 8196 36474
rect 7950 36420 7956 36422
rect 8012 36420 8036 36422
rect 8092 36420 8116 36422
rect 8172 36420 8196 36422
rect 8252 36420 8258 36422
rect 7950 36411 8258 36420
rect 8312 36242 8340 40326
rect 8484 38344 8536 38350
rect 8484 38286 8536 38292
rect 8496 37777 8524 38286
rect 8482 37768 8538 37777
rect 8482 37703 8538 37712
rect 8484 37664 8536 37670
rect 8484 37606 8536 37612
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8404 36718 8432 37062
rect 8392 36712 8444 36718
rect 8392 36654 8444 36660
rect 8300 36236 8352 36242
rect 8300 36178 8352 36184
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 7760 35766 7788 36110
rect 8496 35986 8524 37606
rect 8220 35958 8524 35986
rect 7748 35760 7800 35766
rect 7748 35702 7800 35708
rect 7668 35584 7788 35612
rect 7484 35414 7604 35442
rect 7484 34950 7512 35414
rect 7564 35080 7616 35086
rect 7616 35040 7696 35068
rect 7564 35022 7616 35028
rect 7472 34944 7524 34950
rect 7472 34886 7524 34892
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 7484 33386 7512 34886
rect 7472 33380 7524 33386
rect 7472 33322 7524 33328
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7378 32056 7434 32065
rect 7378 31991 7434 32000
rect 7484 29850 7512 33050
rect 7576 30938 7604 34886
rect 7668 33998 7696 35040
rect 7760 34746 7788 35584
rect 7840 35556 7892 35562
rect 7840 35498 7892 35504
rect 7748 34740 7800 34746
rect 7748 34682 7800 34688
rect 7656 33992 7708 33998
rect 7656 33934 7708 33940
rect 7760 33844 7788 34682
rect 7852 34678 7880 35498
rect 8220 35494 8248 35958
rect 8588 35873 8616 40870
rect 8680 40730 8708 41386
rect 8668 40724 8720 40730
rect 8668 40666 8720 40672
rect 8668 40520 8720 40526
rect 8668 40462 8720 40468
rect 8680 39846 8708 40462
rect 8772 39914 8800 42094
rect 8852 41608 8904 41614
rect 8852 41550 8904 41556
rect 9404 41608 9456 41614
rect 9404 41550 9456 41556
rect 8864 41274 8892 41550
rect 9010 41372 9318 41381
rect 9010 41370 9016 41372
rect 9072 41370 9096 41372
rect 9152 41370 9176 41372
rect 9232 41370 9256 41372
rect 9312 41370 9318 41372
rect 9072 41318 9074 41370
rect 9254 41318 9256 41370
rect 9010 41316 9016 41318
rect 9072 41316 9096 41318
rect 9152 41316 9176 41318
rect 9232 41316 9256 41318
rect 9312 41316 9318 41318
rect 9010 41307 9318 41316
rect 9416 41274 9444 41550
rect 9508 41274 9536 42094
rect 9692 41614 9720 44944
rect 10152 41818 10180 44944
rect 10140 41812 10192 41818
rect 10140 41754 10192 41760
rect 9588 41608 9640 41614
rect 9586 41576 9588 41585
rect 9680 41608 9732 41614
rect 9640 41576 9642 41585
rect 9680 41550 9732 41556
rect 9586 41511 9642 41520
rect 9680 41472 9732 41478
rect 9680 41414 9732 41420
rect 8852 41268 8904 41274
rect 8852 41210 8904 41216
rect 9404 41268 9456 41274
rect 9404 41210 9456 41216
rect 9496 41268 9548 41274
rect 9496 41210 9548 41216
rect 9404 41132 9456 41138
rect 9404 41074 9456 41080
rect 9416 40390 9444 41074
rect 9588 40520 9640 40526
rect 9588 40462 9640 40468
rect 9404 40384 9456 40390
rect 9404 40326 9456 40332
rect 9010 40284 9318 40293
rect 9010 40282 9016 40284
rect 9072 40282 9096 40284
rect 9152 40282 9176 40284
rect 9232 40282 9256 40284
rect 9312 40282 9318 40284
rect 9072 40230 9074 40282
rect 9254 40230 9256 40282
rect 9010 40228 9016 40230
rect 9072 40228 9096 40230
rect 9152 40228 9176 40230
rect 9232 40228 9256 40230
rect 9312 40228 9318 40230
rect 9010 40219 9318 40228
rect 9416 40225 9444 40326
rect 9402 40216 9458 40225
rect 9402 40151 9458 40160
rect 9220 40112 9272 40118
rect 9218 40080 9220 40089
rect 9272 40080 9274 40089
rect 9218 40015 9274 40024
rect 8760 39908 8812 39914
rect 8760 39850 8812 39856
rect 8668 39840 8720 39846
rect 8668 39782 8720 39788
rect 8680 39681 8708 39782
rect 8666 39672 8722 39681
rect 8666 39607 8722 39616
rect 9496 39432 9548 39438
rect 9494 39400 9496 39409
rect 9548 39400 9550 39409
rect 9494 39335 9550 39344
rect 9010 39196 9318 39205
rect 9010 39194 9016 39196
rect 9072 39194 9096 39196
rect 9152 39194 9176 39196
rect 9232 39194 9256 39196
rect 9312 39194 9318 39196
rect 9072 39142 9074 39194
rect 9254 39142 9256 39194
rect 9010 39140 9016 39142
rect 9072 39140 9096 39142
rect 9152 39140 9176 39142
rect 9232 39140 9256 39142
rect 9312 39140 9318 39142
rect 9010 39131 9318 39140
rect 8760 38956 8812 38962
rect 8760 38898 8812 38904
rect 9128 38956 9180 38962
rect 9128 38898 9180 38904
rect 9496 38956 9548 38962
rect 9496 38898 9548 38904
rect 8772 38865 8800 38898
rect 8758 38856 8814 38865
rect 8758 38791 8814 38800
rect 8852 38752 8904 38758
rect 9140 38729 9168 38898
rect 8852 38694 8904 38700
rect 9126 38720 9182 38729
rect 8668 37868 8720 37874
rect 8668 37810 8720 37816
rect 8760 37868 8812 37874
rect 8760 37810 8812 37816
rect 8680 36922 8708 37810
rect 8772 37369 8800 37810
rect 8758 37360 8814 37369
rect 8758 37295 8814 37304
rect 8668 36916 8720 36922
rect 8668 36858 8720 36864
rect 8760 36712 8812 36718
rect 8760 36654 8812 36660
rect 8574 35864 8630 35873
rect 8392 35828 8444 35834
rect 8574 35799 8630 35808
rect 8392 35770 8444 35776
rect 8300 35692 8352 35698
rect 8300 35634 8352 35640
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 7950 35388 8258 35397
rect 7950 35386 7956 35388
rect 8012 35386 8036 35388
rect 8092 35386 8116 35388
rect 8172 35386 8196 35388
rect 8252 35386 8258 35388
rect 8012 35334 8014 35386
rect 8194 35334 8196 35386
rect 7950 35332 7956 35334
rect 8012 35332 8036 35334
rect 8092 35332 8116 35334
rect 8172 35332 8196 35334
rect 8252 35332 8258 35334
rect 7950 35323 8258 35332
rect 8312 35290 8340 35634
rect 8300 35284 8352 35290
rect 8300 35226 8352 35232
rect 7840 34672 7892 34678
rect 7840 34614 7892 34620
rect 7840 34400 7892 34406
rect 7840 34342 7892 34348
rect 7668 33816 7788 33844
rect 7668 32978 7696 33816
rect 7852 33454 7880 34342
rect 7950 34300 8258 34309
rect 7950 34298 7956 34300
rect 8012 34298 8036 34300
rect 8092 34298 8116 34300
rect 8172 34298 8196 34300
rect 8252 34298 8258 34300
rect 8012 34246 8014 34298
rect 8194 34246 8196 34298
rect 7950 34244 7956 34246
rect 8012 34244 8036 34246
rect 8092 34244 8116 34246
rect 8172 34244 8196 34246
rect 8252 34244 8258 34246
rect 7950 34235 8258 34244
rect 8208 33992 8260 33998
rect 8208 33934 8260 33940
rect 8300 33992 8352 33998
rect 8300 33934 8352 33940
rect 8220 33658 8248 33934
rect 8208 33652 8260 33658
rect 8208 33594 8260 33600
rect 7748 33448 7800 33454
rect 7748 33390 7800 33396
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7656 32972 7708 32978
rect 7656 32914 7708 32920
rect 7760 31346 7788 33390
rect 7950 33212 8258 33221
rect 7950 33210 7956 33212
rect 8012 33210 8036 33212
rect 8092 33210 8116 33212
rect 8172 33210 8196 33212
rect 8252 33210 8258 33212
rect 8012 33158 8014 33210
rect 8194 33158 8196 33210
rect 7950 33156 7956 33158
rect 8012 33156 8036 33158
rect 8092 33156 8116 33158
rect 8172 33156 8196 33158
rect 8252 33156 8258 33158
rect 7950 33147 8258 33156
rect 7838 33008 7894 33017
rect 7838 32943 7894 32952
rect 7748 31340 7800 31346
rect 7748 31282 7800 31288
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 7564 30932 7616 30938
rect 7564 30874 7616 30880
rect 7564 30116 7616 30122
rect 7564 30058 7616 30064
rect 7576 29850 7604 30058
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7564 29844 7616 29850
rect 7564 29786 7616 29792
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7102 24919 7158 24928
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 7104 24812 7156 24818
rect 7104 24754 7156 24760
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 7010 23080 7066 23089
rect 7010 23015 7066 23024
rect 7024 22817 7052 23015
rect 7010 22808 7066 22817
rect 7010 22743 7012 22752
rect 7064 22743 7066 22752
rect 7012 22714 7064 22720
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7024 22545 7052 22578
rect 7010 22536 7066 22545
rect 7010 22471 7066 22480
rect 6932 22392 7052 22420
rect 6918 22264 6974 22273
rect 7024 22234 7052 22392
rect 6918 22199 6974 22208
rect 7012 22228 7064 22234
rect 6748 22066 6868 22094
rect 6932 22080 6960 22199
rect 7012 22170 7064 22176
rect 6642 21312 6698 21321
rect 6642 21247 6698 21256
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6656 19961 6684 21082
rect 6642 19952 6698 19961
rect 6642 19887 6698 19896
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19378 6684 19790
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6656 17354 6684 18226
rect 6748 17882 6776 22066
rect 6932 22052 7052 22080
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6918 21992 6974 22001
rect 6840 18970 6868 21966
rect 6918 21927 6974 21936
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6932 18034 6960 21927
rect 7024 21894 7052 22052
rect 7116 22001 7144 24754
rect 7196 24744 7248 24750
rect 7194 24712 7196 24721
rect 7300 24732 7328 25842
rect 7248 24712 7328 24732
rect 7250 24704 7328 24712
rect 7194 24647 7250 24656
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7208 22273 7236 24550
rect 7300 24313 7328 24550
rect 7286 24304 7342 24313
rect 7286 24239 7342 24248
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7300 23662 7328 24142
rect 7392 23798 7420 28902
rect 7380 23792 7432 23798
rect 7380 23734 7432 23740
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7286 22944 7342 22953
rect 7286 22879 7342 22888
rect 7194 22264 7250 22273
rect 7194 22199 7250 22208
rect 7196 22160 7248 22166
rect 7196 22102 7248 22108
rect 7102 21992 7158 22001
rect 7102 21927 7158 21936
rect 7012 21888 7064 21894
rect 7012 21830 7064 21836
rect 7102 21856 7158 21865
rect 7102 21791 7158 21800
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 7024 18290 7052 21490
rect 7116 18766 7144 21791
rect 7208 21321 7236 22102
rect 7194 21312 7250 21321
rect 7194 21247 7250 21256
rect 7196 20952 7248 20958
rect 7196 20894 7248 20900
rect 7208 20466 7236 20894
rect 7300 20534 7328 22879
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7288 20392 7340 20398
rect 7194 20360 7250 20369
rect 7288 20334 7340 20340
rect 7194 20295 7250 20304
rect 7208 19334 7236 20295
rect 7300 19514 7328 20334
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7208 19306 7328 19334
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6840 18006 6960 18034
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6564 17326 6684 17354
rect 6368 16584 6420 16590
rect 6090 16552 6146 16561
rect 6368 16526 6420 16532
rect 6090 16487 6146 16496
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5998 15872 6054 15881
rect 5998 15807 6054 15816
rect 6012 15570 6040 15807
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5998 15464 6054 15473
rect 5998 15399 6054 15408
rect 6012 13394 6040 15399
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6104 13274 6132 16390
rect 6274 16144 6330 16153
rect 6274 16079 6330 16088
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15502 6224 15846
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6288 13297 6316 16079
rect 6380 16046 6408 16526
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6380 14958 6408 15982
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 6012 13246 6132 13274
rect 6274 13288 6330 13297
rect 5632 12718 5684 12724
rect 5814 12744 5870 12753
rect 5814 12679 5870 12688
rect 5828 12628 5856 12679
rect 5644 12600 5856 12628
rect 5446 12407 5502 12416
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5644 12306 5672 12600
rect 6012 12434 6040 13246
rect 6274 13223 6330 13232
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 5920 12406 6040 12434
rect 6184 12436 6236 12442
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5262 11928 5318 11937
rect 5262 11863 5264 11872
rect 5316 11863 5318 11872
rect 5264 11834 5316 11840
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 10198 5304 10406
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5276 9382 5304 10134
rect 5368 9625 5396 12174
rect 5644 11286 5672 12242
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 5460 9722 5488 10474
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5354 9616 5410 9625
rect 5354 9551 5410 9560
rect 5448 9580 5500 9586
rect 5368 9518 5396 9551
rect 5448 9522 5500 9528
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5000 7806 5212 7834
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7342 4844 7686
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 5000 5710 5028 7806
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 6118 5120 7686
rect 5276 7342 5304 7958
rect 5368 7954 5396 9454
rect 5460 9450 5488 9522
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5552 8294 5580 11154
rect 5736 10962 5764 12242
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 11150 5856 11562
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5644 10934 5764 10962
rect 5644 9722 5672 10934
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5644 7954 5672 9658
rect 5736 8362 5764 10746
rect 5828 10606 5856 11086
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5828 9654 5856 9998
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5828 9178 5856 9454
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5736 8022 5764 8298
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5356 7948 5408 7954
rect 5632 7948 5684 7954
rect 5408 7908 5488 7936
rect 5356 7890 5408 7896
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 7002 5396 7142
rect 5460 7002 5488 7908
rect 5632 7890 5684 7896
rect 5644 7449 5672 7890
rect 5630 7440 5686 7449
rect 5630 7375 5686 7384
rect 5828 7324 5856 8434
rect 5552 7296 5856 7324
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5552 6866 5580 7296
rect 5722 7168 5778 7177
rect 5722 7103 5778 7112
rect 5736 6866 5764 7103
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5644 6662 5672 6802
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6390 5764 6598
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5460 5914 5488 6054
rect 5722 5944 5778 5953
rect 5448 5908 5500 5914
rect 5722 5879 5778 5888
rect 5448 5850 5500 5856
rect 5736 5846 5764 5879
rect 5724 5840 5776 5846
rect 5538 5808 5594 5817
rect 5724 5782 5776 5788
rect 5538 5743 5594 5752
rect 5552 5710 5580 5743
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5920 5574 5948 12406
rect 6184 12378 6236 12384
rect 6196 12306 6224 12378
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6000 12232 6052 12238
rect 6288 12209 6316 12854
rect 6000 12174 6052 12180
rect 6274 12200 6330 12209
rect 6012 11665 6040 12174
rect 6274 12135 6330 12144
rect 6276 11688 6328 11694
rect 5998 11656 6054 11665
rect 6276 11630 6328 11636
rect 5998 11591 6054 11600
rect 6012 10674 6040 11591
rect 6288 11132 6316 11630
rect 6380 11234 6408 14894
rect 6472 14618 6500 15506
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6564 14414 6592 17326
rect 6840 17218 6868 18006
rect 7208 17542 7236 19110
rect 7300 18170 7328 19306
rect 7392 18290 7420 23258
rect 7484 22234 7512 29038
rect 7576 26042 7604 29106
rect 7564 26036 7616 26042
rect 7564 25978 7616 25984
rect 7668 25922 7696 31214
rect 7760 30394 7788 31282
rect 7748 30388 7800 30394
rect 7748 30330 7800 30336
rect 7748 30184 7800 30190
rect 7748 30126 7800 30132
rect 7760 29034 7788 30126
rect 7852 29832 7880 32943
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8128 32570 8156 32846
rect 8208 32768 8260 32774
rect 8208 32710 8260 32716
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 8220 32434 8248 32710
rect 8208 32428 8260 32434
rect 8208 32370 8260 32376
rect 8312 32230 8340 33934
rect 8404 32502 8432 35770
rect 8588 35698 8708 35714
rect 8576 35692 8708 35698
rect 8628 35686 8708 35692
rect 8576 35634 8628 35640
rect 8484 35624 8536 35630
rect 8574 35592 8630 35601
rect 8536 35572 8574 35578
rect 8484 35566 8574 35572
rect 8496 35550 8574 35566
rect 8574 35527 8630 35536
rect 8484 35488 8536 35494
rect 8484 35430 8536 35436
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8300 32224 8352 32230
rect 8300 32166 8352 32172
rect 7950 32124 8258 32133
rect 7950 32122 7956 32124
rect 8012 32122 8036 32124
rect 8092 32122 8116 32124
rect 8172 32122 8196 32124
rect 8252 32122 8258 32124
rect 8012 32070 8014 32122
rect 8194 32070 8196 32122
rect 7950 32068 7956 32070
rect 8012 32068 8036 32070
rect 8092 32068 8116 32070
rect 8172 32068 8196 32070
rect 8252 32068 8258 32070
rect 7950 32059 8258 32068
rect 8116 31748 8168 31754
rect 8116 31690 8168 31696
rect 8128 31482 8156 31690
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8116 31476 8168 31482
rect 8116 31418 8168 31424
rect 8312 31278 8340 31622
rect 8404 31385 8432 32302
rect 8390 31376 8446 31385
rect 8390 31311 8446 31320
rect 8300 31272 8352 31278
rect 8300 31214 8352 31220
rect 8392 31272 8444 31278
rect 8392 31214 8444 31220
rect 7950 31036 8258 31045
rect 7950 31034 7956 31036
rect 8012 31034 8036 31036
rect 8092 31034 8116 31036
rect 8172 31034 8196 31036
rect 8252 31034 8258 31036
rect 8012 30982 8014 31034
rect 8194 30982 8196 31034
rect 7950 30980 7956 30982
rect 8012 30980 8036 30982
rect 8092 30980 8116 30982
rect 8172 30980 8196 30982
rect 8252 30980 8258 30982
rect 7950 30971 8258 30980
rect 8404 30818 8432 31214
rect 8128 30790 8432 30818
rect 8128 30258 8156 30790
rect 8392 30728 8444 30734
rect 8496 30716 8524 35430
rect 8680 34746 8708 35686
rect 8772 35601 8800 36654
rect 8864 36174 8892 38694
rect 9126 38655 9182 38664
rect 9128 38344 9180 38350
rect 9126 38312 9128 38321
rect 9180 38312 9182 38321
rect 9126 38247 9182 38256
rect 9010 38108 9318 38117
rect 9010 38106 9016 38108
rect 9072 38106 9096 38108
rect 9152 38106 9176 38108
rect 9232 38106 9256 38108
rect 9312 38106 9318 38108
rect 9072 38054 9074 38106
rect 9254 38054 9256 38106
rect 9010 38052 9016 38054
rect 9072 38052 9096 38054
rect 9152 38052 9176 38054
rect 9232 38052 9256 38054
rect 9312 38052 9318 38054
rect 9010 38043 9318 38052
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 9010 37020 9318 37029
rect 9010 37018 9016 37020
rect 9072 37018 9096 37020
rect 9152 37018 9176 37020
rect 9232 37018 9256 37020
rect 9312 37018 9318 37020
rect 9072 36966 9074 37018
rect 9254 36966 9256 37018
rect 9010 36964 9016 36966
rect 9072 36964 9096 36966
rect 9152 36964 9176 36966
rect 9232 36964 9256 36966
rect 9312 36964 9318 36966
rect 9010 36955 9318 36964
rect 9312 36848 9364 36854
rect 9312 36790 9364 36796
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 8852 36168 8904 36174
rect 9140 36145 9168 36722
rect 9324 36258 9352 36790
rect 9416 36378 9444 37198
rect 9404 36372 9456 36378
rect 9404 36314 9456 36320
rect 9508 36310 9536 38898
rect 9496 36304 9548 36310
rect 9324 36230 9444 36258
rect 9496 36246 9548 36252
rect 8852 36110 8904 36116
rect 9126 36136 9182 36145
rect 9126 36071 9182 36080
rect 8852 36032 8904 36038
rect 8852 35974 8904 35980
rect 8864 35630 8892 35974
rect 9010 35932 9318 35941
rect 9010 35930 9016 35932
rect 9072 35930 9096 35932
rect 9152 35930 9176 35932
rect 9232 35930 9256 35932
rect 9312 35930 9318 35932
rect 9072 35878 9074 35930
rect 9254 35878 9256 35930
rect 9010 35876 9016 35878
rect 9072 35876 9096 35878
rect 9152 35876 9176 35878
rect 9232 35876 9256 35878
rect 9312 35876 9318 35878
rect 9010 35867 9318 35876
rect 9416 35630 9444 36230
rect 9600 36122 9628 40462
rect 9692 39273 9720 41414
rect 9772 41132 9824 41138
rect 9772 41074 9824 41080
rect 9784 40390 9812 41074
rect 10416 40928 10468 40934
rect 10416 40870 10468 40876
rect 9772 40384 9824 40390
rect 9770 40352 9772 40361
rect 9824 40352 9826 40361
rect 9770 40287 9826 40296
rect 10428 39817 10456 40870
rect 10600 39908 10652 39914
rect 10600 39850 10652 39856
rect 10414 39808 10470 39817
rect 10414 39743 10470 39752
rect 10232 39568 10284 39574
rect 10612 39545 10640 39850
rect 10784 39840 10836 39846
rect 10784 39782 10836 39788
rect 10232 39510 10284 39516
rect 10598 39536 10654 39545
rect 9678 39264 9734 39273
rect 9678 39199 9734 39208
rect 10244 39001 10272 39510
rect 10598 39471 10654 39480
rect 10416 39296 10468 39302
rect 10416 39238 10468 39244
rect 10324 39092 10376 39098
rect 10324 39034 10376 39040
rect 10230 38992 10286 39001
rect 10230 38927 10286 38936
rect 10140 38820 10192 38826
rect 10140 38762 10192 38768
rect 10048 38480 10100 38486
rect 10152 38457 10180 38762
rect 10048 38422 10100 38428
rect 10138 38448 10194 38457
rect 9956 38276 10008 38282
rect 9956 38218 10008 38224
rect 9968 37369 9996 38218
rect 9954 37360 10010 37369
rect 9954 37295 10010 37304
rect 9680 37120 9732 37126
rect 10060 37097 10088 38422
rect 10138 38383 10194 38392
rect 10140 38004 10192 38010
rect 10140 37946 10192 37952
rect 9680 37062 9732 37068
rect 10046 37088 10102 37097
rect 9508 36094 9628 36122
rect 8852 35624 8904 35630
rect 8758 35592 8814 35601
rect 8852 35566 8904 35572
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 8758 35527 8814 35536
rect 8772 35476 8800 35527
rect 8772 35448 8892 35476
rect 8668 34740 8720 34746
rect 8668 34682 8720 34688
rect 8760 33924 8812 33930
rect 8760 33866 8812 33872
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8680 31822 8708 33798
rect 8772 33522 8800 33866
rect 8760 33516 8812 33522
rect 8760 33458 8812 33464
rect 8864 32910 8892 35448
rect 9324 35290 9352 35566
rect 9312 35284 9364 35290
rect 9312 35226 9364 35232
rect 8944 35080 8996 35086
rect 8942 35048 8944 35057
rect 8996 35048 8998 35057
rect 8942 34983 8998 34992
rect 9010 34844 9318 34853
rect 9010 34842 9016 34844
rect 9072 34842 9096 34844
rect 9152 34842 9176 34844
rect 9232 34842 9256 34844
rect 9312 34842 9318 34844
rect 9072 34790 9074 34842
rect 9254 34790 9256 34842
rect 9010 34788 9016 34790
rect 9072 34788 9096 34790
rect 9152 34788 9176 34790
rect 9232 34788 9256 34790
rect 9312 34788 9318 34790
rect 9010 34779 9318 34788
rect 9416 34202 9444 35566
rect 9404 34196 9456 34202
rect 9404 34138 9456 34144
rect 9508 34082 9536 36094
rect 9588 36032 9640 36038
rect 9588 35974 9640 35980
rect 9600 34649 9628 35974
rect 9692 35193 9720 37062
rect 10046 37023 10102 37032
rect 10152 36553 10180 37946
rect 10336 37913 10364 39034
rect 10428 38185 10456 39238
rect 10508 38752 10560 38758
rect 10796 38729 10824 39782
rect 10508 38694 10560 38700
rect 10782 38720 10838 38729
rect 10414 38176 10470 38185
rect 10414 38111 10470 38120
rect 10322 37904 10378 37913
rect 10322 37839 10378 37848
rect 10232 37732 10284 37738
rect 10232 37674 10284 37680
rect 10244 37641 10272 37674
rect 10230 37632 10286 37641
rect 10230 37567 10286 37576
rect 10324 37188 10376 37194
rect 10324 37130 10376 37136
rect 10138 36544 10194 36553
rect 10138 36479 10194 36488
rect 10232 36304 10284 36310
rect 10232 36246 10284 36252
rect 10140 36032 10192 36038
rect 10140 35974 10192 35980
rect 9956 35216 10008 35222
rect 9678 35184 9734 35193
rect 9956 35158 10008 35164
rect 9678 35119 9734 35128
rect 9968 34921 9996 35158
rect 9954 34912 10010 34921
rect 9954 34847 10010 34856
rect 9586 34640 9642 34649
rect 9586 34575 9642 34584
rect 9416 34054 9536 34082
rect 9956 34128 10008 34134
rect 9956 34070 10008 34076
rect 9128 33992 9180 33998
rect 9126 33960 9128 33969
rect 9180 33960 9182 33969
rect 9126 33895 9182 33904
rect 9010 33756 9318 33765
rect 9010 33754 9016 33756
rect 9072 33754 9096 33756
rect 9152 33754 9176 33756
rect 9232 33754 9256 33756
rect 9312 33754 9318 33756
rect 9072 33702 9074 33754
rect 9254 33702 9256 33754
rect 9010 33700 9016 33702
rect 9072 33700 9096 33702
rect 9152 33700 9176 33702
rect 9232 33700 9256 33702
rect 9312 33700 9318 33702
rect 9010 33691 9318 33700
rect 8852 32904 8904 32910
rect 8852 32846 8904 32852
rect 8852 32768 8904 32774
rect 8850 32736 8852 32745
rect 8904 32736 8906 32745
rect 8850 32671 8906 32680
rect 9010 32668 9318 32677
rect 9010 32666 9016 32668
rect 9072 32666 9096 32668
rect 9152 32666 9176 32668
rect 9232 32666 9256 32668
rect 9312 32666 9318 32668
rect 9072 32614 9074 32666
rect 9254 32614 9256 32666
rect 9010 32612 9016 32614
rect 9072 32612 9096 32614
rect 9152 32612 9176 32614
rect 9232 32612 9256 32614
rect 9312 32612 9318 32614
rect 9010 32603 9318 32612
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8852 32292 8904 32298
rect 8852 32234 8904 32240
rect 8576 31816 8628 31822
rect 8576 31758 8628 31764
rect 8668 31816 8720 31822
rect 8668 31758 8720 31764
rect 8588 31482 8616 31758
rect 8760 31680 8812 31686
rect 8760 31622 8812 31628
rect 8576 31476 8628 31482
rect 8576 31418 8628 31424
rect 8574 31376 8630 31385
rect 8574 31311 8576 31320
rect 8628 31311 8630 31320
rect 8576 31282 8628 31288
rect 8668 31272 8720 31278
rect 8666 31240 8668 31249
rect 8720 31240 8722 31249
rect 8666 31175 8722 31184
rect 8576 31136 8628 31142
rect 8576 31078 8628 31084
rect 8444 30688 8524 30716
rect 8392 30670 8444 30676
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8404 30258 8432 30534
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 8392 30252 8444 30258
rect 8392 30194 8444 30200
rect 8588 30190 8616 31078
rect 8680 30977 8708 31175
rect 8666 30968 8722 30977
rect 8666 30903 8722 30912
rect 8668 30796 8720 30802
rect 8668 30738 8720 30744
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 7950 29948 8258 29957
rect 7950 29946 7956 29948
rect 8012 29946 8036 29948
rect 8092 29946 8116 29948
rect 8172 29946 8196 29948
rect 8252 29946 8258 29948
rect 8012 29894 8014 29946
rect 8194 29894 8196 29946
rect 7950 29892 7956 29894
rect 8012 29892 8036 29894
rect 8092 29892 8116 29894
rect 8172 29892 8196 29894
rect 8252 29892 8258 29894
rect 7950 29883 8258 29892
rect 8312 29832 8340 30126
rect 8680 29866 8708 30738
rect 8772 30734 8800 31622
rect 8864 31346 8892 32234
rect 8956 31754 8984 32370
rect 9416 32314 9444 34054
rect 9496 33992 9548 33998
rect 9496 33934 9548 33940
rect 9508 33425 9536 33934
rect 9680 33856 9732 33862
rect 9968 33833 9996 34070
rect 9680 33798 9732 33804
rect 9954 33824 10010 33833
rect 9494 33416 9550 33425
rect 9494 33351 9496 33360
rect 9548 33351 9550 33360
rect 9496 33322 9548 33328
rect 9692 32745 9720 33798
rect 9954 33759 10010 33768
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9678 32736 9734 32745
rect 9678 32671 9734 32680
rect 9864 32564 9916 32570
rect 9864 32506 9916 32512
rect 9140 32286 9444 32314
rect 9140 31958 9168 32286
rect 9220 32224 9272 32230
rect 9220 32166 9272 32172
rect 9404 32224 9456 32230
rect 9404 32166 9456 32172
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9232 32026 9260 32166
rect 9220 32020 9272 32026
rect 9220 31962 9272 31968
rect 9128 31952 9180 31958
rect 9128 31894 9180 31900
rect 9312 31816 9364 31822
rect 9416 31793 9444 32166
rect 9496 31952 9548 31958
rect 9496 31894 9548 31900
rect 9588 31952 9640 31958
rect 9588 31894 9640 31900
rect 9312 31758 9364 31764
rect 9402 31784 9458 31793
rect 8944 31748 8996 31754
rect 8944 31690 8996 31696
rect 9324 31668 9352 31758
rect 9402 31719 9458 31728
rect 9324 31640 9444 31668
rect 9010 31580 9318 31589
rect 9010 31578 9016 31580
rect 9072 31578 9096 31580
rect 9152 31578 9176 31580
rect 9232 31578 9256 31580
rect 9312 31578 9318 31580
rect 9072 31526 9074 31578
rect 9254 31526 9256 31578
rect 9010 31524 9016 31526
rect 9072 31524 9096 31526
rect 9152 31524 9176 31526
rect 9232 31524 9256 31526
rect 9312 31524 9318 31526
rect 9010 31515 9318 31524
rect 9034 31376 9090 31385
rect 8852 31340 8904 31346
rect 9416 31362 9444 31640
rect 9034 31311 9090 31320
rect 9324 31334 9444 31362
rect 8852 31282 8904 31288
rect 9048 31278 9076 31311
rect 9036 31272 9088 31278
rect 9036 31214 9088 31220
rect 8852 31136 8904 31142
rect 8852 31078 8904 31084
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 8758 30424 8814 30433
rect 8758 30359 8814 30368
rect 7852 29804 7972 29832
rect 7748 29028 7800 29034
rect 7748 28970 7800 28976
rect 7840 29028 7892 29034
rect 7840 28970 7892 28976
rect 7576 25894 7696 25922
rect 7576 25498 7604 25894
rect 7656 25832 7708 25838
rect 7656 25774 7708 25780
rect 7564 25492 7616 25498
rect 7564 25434 7616 25440
rect 7564 25220 7616 25226
rect 7564 25162 7616 25168
rect 7576 23322 7604 25162
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7564 22704 7616 22710
rect 7564 22646 7616 22652
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7470 22128 7526 22137
rect 7470 22063 7526 22072
rect 7484 21622 7512 22063
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7576 21486 7604 22646
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7484 19378 7512 21422
rect 7668 21185 7696 25774
rect 7760 23866 7788 28970
rect 7852 28218 7880 28970
rect 7944 28966 7972 29804
rect 8220 29804 8340 29832
rect 8404 29838 8708 29866
rect 8024 29776 8076 29782
rect 8022 29744 8024 29753
rect 8076 29744 8078 29753
rect 8022 29679 8078 29688
rect 8024 29640 8076 29646
rect 8024 29582 8076 29588
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8036 29152 8064 29582
rect 8128 29345 8156 29582
rect 8114 29336 8170 29345
rect 8114 29271 8170 29280
rect 8116 29164 8168 29170
rect 8036 29124 8116 29152
rect 8116 29106 8168 29112
rect 8220 29102 8248 29804
rect 8404 29288 8432 29838
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8666 29608 8722 29617
rect 8312 29260 8432 29288
rect 8208 29096 8260 29102
rect 8208 29038 8260 29044
rect 7932 28960 7984 28966
rect 7932 28902 7984 28908
rect 7950 28860 8258 28869
rect 7950 28858 7956 28860
rect 8012 28858 8036 28860
rect 8092 28858 8116 28860
rect 8172 28858 8196 28860
rect 8252 28858 8258 28860
rect 8012 28806 8014 28858
rect 8194 28806 8196 28858
rect 7950 28804 7956 28806
rect 8012 28804 8036 28806
rect 8092 28804 8116 28806
rect 8172 28804 8196 28806
rect 8252 28804 8258 28806
rect 7950 28795 8258 28804
rect 7932 28688 7984 28694
rect 7932 28630 7984 28636
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7852 27470 7880 28018
rect 7944 27878 7972 28630
rect 8114 28248 8170 28257
rect 8114 28183 8116 28192
rect 8168 28183 8170 28192
rect 8116 28154 8168 28160
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7950 27772 8258 27781
rect 7950 27770 7956 27772
rect 8012 27770 8036 27772
rect 8092 27770 8116 27772
rect 8172 27770 8196 27772
rect 8252 27770 8258 27772
rect 8012 27718 8014 27770
rect 8194 27718 8196 27770
rect 7950 27716 7956 27718
rect 8012 27716 8036 27718
rect 8092 27716 8116 27718
rect 8172 27716 8196 27718
rect 8252 27716 8258 27718
rect 7950 27707 8258 27716
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7852 26246 7880 27066
rect 7950 26684 8258 26693
rect 7950 26682 7956 26684
rect 8012 26682 8036 26684
rect 8092 26682 8116 26684
rect 8172 26682 8196 26684
rect 8252 26682 8258 26684
rect 8012 26630 8014 26682
rect 8194 26630 8196 26682
rect 7950 26628 7956 26630
rect 8012 26628 8036 26630
rect 8092 26628 8116 26630
rect 8172 26628 8196 26630
rect 8252 26628 8258 26630
rect 7950 26619 8258 26628
rect 8312 26466 8340 29260
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8404 28762 8432 29038
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8404 26897 8432 27610
rect 8390 26888 8446 26897
rect 8390 26823 8446 26832
rect 8496 26625 8524 29582
rect 8666 29543 8722 29552
rect 8680 29073 8708 29543
rect 8772 29102 8800 30359
rect 8760 29096 8812 29102
rect 8666 29064 8722 29073
rect 8760 29038 8812 29044
rect 8666 28999 8722 29008
rect 8576 28960 8628 28966
rect 8576 28902 8628 28908
rect 8588 28558 8616 28902
rect 8576 28552 8628 28558
rect 8576 28494 8628 28500
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 8588 27470 8616 28018
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8482 26616 8538 26625
rect 8482 26551 8538 26560
rect 8484 26512 8536 26518
rect 8312 26438 8432 26466
rect 8484 26454 8536 26460
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7852 24970 7880 25978
rect 7944 25809 7972 26318
rect 8220 26217 8248 26318
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 8206 26208 8262 26217
rect 8206 26143 8262 26152
rect 7930 25800 7986 25809
rect 8312 25770 8340 26250
rect 7930 25735 7986 25744
rect 8300 25764 8352 25770
rect 8300 25706 8352 25712
rect 7950 25596 8258 25605
rect 7950 25594 7956 25596
rect 8012 25594 8036 25596
rect 8092 25594 8116 25596
rect 8172 25594 8196 25596
rect 8252 25594 8258 25596
rect 8012 25542 8014 25594
rect 8194 25542 8196 25594
rect 7950 25540 7956 25542
rect 8012 25540 8036 25542
rect 8092 25540 8116 25542
rect 8172 25540 8196 25542
rect 8252 25540 8258 25542
rect 7950 25531 8258 25540
rect 7932 25492 7984 25498
rect 8312 25480 8340 25706
rect 7932 25434 7984 25440
rect 8128 25452 8340 25480
rect 7944 25158 7972 25434
rect 8022 25392 8078 25401
rect 8022 25327 8078 25336
rect 8036 25294 8064 25327
rect 8024 25288 8076 25294
rect 8024 25230 8076 25236
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7852 24942 7972 24970
rect 7944 24750 7972 24942
rect 8128 24818 8156 25452
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8220 25158 8248 25230
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8220 24857 8248 25094
rect 8206 24848 8262 24857
rect 8116 24812 8168 24818
rect 8206 24783 8208 24792
rect 8116 24754 8168 24760
rect 8260 24783 8262 24792
rect 8208 24754 8260 24760
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7840 24676 7892 24682
rect 7840 24618 7892 24624
rect 7852 23866 7880 24618
rect 8128 24614 8156 24754
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 7950 24508 8258 24517
rect 7950 24506 7956 24508
rect 8012 24506 8036 24508
rect 8092 24506 8116 24508
rect 8172 24506 8196 24508
rect 8252 24506 8258 24508
rect 8012 24454 8014 24506
rect 8194 24454 8196 24506
rect 7950 24452 7956 24454
rect 8012 24452 8036 24454
rect 8092 24452 8116 24454
rect 8172 24452 8196 24454
rect 8252 24452 8258 24454
rect 7950 24443 8258 24452
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7760 23474 7788 23802
rect 7944 23769 7972 24074
rect 7930 23760 7986 23769
rect 7930 23695 7986 23704
rect 8036 23633 8064 24142
rect 8312 24018 8340 25094
rect 8404 24834 8432 26438
rect 8496 26042 8524 26454
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 8588 25786 8616 27406
rect 8680 27402 8708 28494
rect 8760 28416 8812 28422
rect 8760 28358 8812 28364
rect 8772 28082 8800 28358
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 8760 27600 8812 27606
rect 8758 27568 8760 27577
rect 8812 27568 8814 27577
rect 8758 27503 8814 27512
rect 8668 27396 8720 27402
rect 8668 27338 8720 27344
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8666 26616 8722 26625
rect 8666 26551 8722 26560
rect 8496 25758 8616 25786
rect 8496 25140 8524 25758
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8588 25294 8616 25638
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8496 25112 8616 25140
rect 8404 24806 8524 24834
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8404 24410 8432 24686
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8312 23990 8432 24018
rect 8298 23896 8354 23905
rect 8298 23831 8354 23840
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8220 23633 8248 23666
rect 8022 23624 8078 23633
rect 8022 23559 8078 23568
rect 8206 23624 8262 23633
rect 8206 23559 8262 23568
rect 7760 23446 7880 23474
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7760 21729 7788 23258
rect 7746 21720 7802 21729
rect 7746 21655 7802 21664
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7654 21176 7710 21185
rect 7654 21111 7710 21120
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 7576 20058 7604 20946
rect 7760 20466 7788 21354
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7576 19689 7604 19722
rect 7562 19680 7618 19689
rect 7562 19615 7618 19624
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7300 18142 7420 18170
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 6656 17190 6868 17218
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6472 12102 6500 12786
rect 6656 12434 6684 17190
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6748 15706 6776 16662
rect 7024 16590 7052 17478
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 14521 6776 14962
rect 6920 14544 6972 14550
rect 6734 14512 6790 14521
rect 6920 14486 6972 14492
rect 6734 14447 6790 14456
rect 6828 14408 6880 14414
rect 6748 14356 6828 14362
rect 6748 14350 6880 14356
rect 6748 14334 6868 14350
rect 6748 13870 6776 14334
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6748 13326 6776 13670
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12986 6776 13262
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6840 12850 6868 13398
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6748 12442 6776 12582
rect 6564 12406 6684 12434
rect 6736 12436 6788 12442
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6472 11762 6500 12038
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6564 11626 6592 12406
rect 6736 12378 6788 12384
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6380 11206 6592 11234
rect 6656 11218 6684 12310
rect 6840 12238 6868 12650
rect 6828 12232 6880 12238
rect 6734 12200 6790 12209
rect 6828 12174 6880 12180
rect 6734 12135 6736 12144
rect 6788 12135 6790 12144
rect 6736 12106 6788 12112
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6460 11144 6512 11150
rect 6288 11104 6460 11132
rect 6460 11086 6512 11092
rect 6472 11014 6500 11086
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6012 7936 6040 10610
rect 6564 10606 6592 11206
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6748 10674 6776 11494
rect 6840 11354 6868 12038
rect 6932 11558 6960 14486
rect 7024 12782 7052 15030
rect 7116 13870 7144 17138
rect 7300 17134 7328 18022
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 14482 7236 15982
rect 7300 15586 7328 17070
rect 7392 16046 7420 18142
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7378 15736 7434 15745
rect 7378 15671 7380 15680
rect 7432 15671 7434 15680
rect 7380 15642 7432 15648
rect 7300 15558 7420 15586
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 11762 7052 12718
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6932 11098 6960 11494
rect 6840 11070 6960 11098
rect 6840 10810 6868 11070
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6090 9480 6146 9489
rect 6090 9415 6092 9424
rect 6144 9415 6146 9424
rect 6092 9386 6144 9392
rect 6092 7948 6144 7954
rect 6012 7908 6092 7936
rect 6012 7177 6040 7908
rect 6092 7890 6144 7896
rect 5998 7168 6054 7177
rect 5998 7103 6054 7112
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6012 6866 6040 6938
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6092 6180 6144 6186
rect 6092 6122 6144 6128
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 5920 5234 5948 5510
rect 6104 5234 6132 6122
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 5920 4622 5948 5170
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 2792 56 2820 2518
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3252 56 3280 2042
rect 3698 1320 3754 1329
rect 3698 1255 3754 1264
rect 3712 56 3740 1255
rect 4172 56 4200 4218
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5078 1320 5134 1329
rect 5078 1255 5134 1264
rect 4618 1184 4674 1193
rect 4618 1119 4674 1128
rect 4632 56 4660 1119
rect 5092 56 5120 1255
rect 5552 56 5580 2586
rect 6012 56 6132 82
rect 938 0 994 56
rect 1398 0 1454 56
rect 1858 0 1914 56
rect 2318 0 2374 56
rect 2778 0 2834 56
rect 3238 0 3294 56
rect 3698 0 3754 56
rect 4158 0 4214 56
rect 4618 0 4674 56
rect 5078 0 5134 56
rect 5538 0 5594 56
rect 5998 54 6132 56
rect 5998 0 6054 54
rect 6104 42 6132 54
rect 6196 42 6224 10202
rect 6380 9926 6408 10542
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6276 9376 6328 9382
rect 6274 9344 6276 9353
rect 6328 9344 6330 9353
rect 6274 9279 6330 9288
rect 6274 8664 6330 8673
rect 6274 8599 6330 8608
rect 6288 7886 6316 8599
rect 6380 8498 6408 9862
rect 6472 9586 6500 10066
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6472 9178 6500 9522
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6564 8838 6592 10542
rect 6748 9489 6776 10610
rect 6826 10568 6882 10577
rect 6826 10503 6882 10512
rect 6840 10130 6868 10503
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9518 6868 10066
rect 6828 9512 6880 9518
rect 6734 9480 6790 9489
rect 6828 9454 6880 9460
rect 6734 9415 6790 9424
rect 6932 9382 6960 10950
rect 7010 10160 7066 10169
rect 7010 10095 7066 10104
rect 7024 10062 7052 10095
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7024 9194 7052 9998
rect 6748 9166 7052 9194
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7750 6316 7822
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6380 6866 6408 8026
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6656 7002 6684 7346
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6748 6322 6776 9166
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6826 8392 6882 8401
rect 6826 8327 6882 8336
rect 6840 7274 6868 8327
rect 6932 8090 6960 9046
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8430 7052 8774
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6918 7576 6974 7585
rect 6918 7511 6920 7520
rect 6972 7511 6974 7520
rect 6920 7482 6972 7488
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 7116 6662 7144 13806
rect 7208 7546 7236 14010
rect 7300 13462 7328 15302
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7392 12850 7420 15558
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7300 11354 7328 12786
rect 7378 12744 7434 12753
rect 7378 12679 7380 12688
rect 7432 12679 7434 12688
rect 7380 12650 7432 12656
rect 7484 12434 7512 19314
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7576 18222 7604 18634
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7564 17876 7616 17882
rect 7668 17864 7696 20266
rect 7760 19446 7788 20402
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7760 18222 7788 19246
rect 7852 18970 7880 23446
rect 7950 23420 8258 23429
rect 7950 23418 7956 23420
rect 8012 23418 8036 23420
rect 8092 23418 8116 23420
rect 8172 23418 8196 23420
rect 8252 23418 8258 23420
rect 8012 23366 8014 23418
rect 8194 23366 8196 23418
rect 7950 23364 7956 23366
rect 8012 23364 8036 23366
rect 8092 23364 8116 23366
rect 8172 23364 8196 23366
rect 8252 23364 8258 23366
rect 7950 23355 8258 23364
rect 8022 23216 8078 23225
rect 8022 23151 8078 23160
rect 8036 23118 8064 23151
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7944 22574 7972 23054
rect 7932 22568 7984 22574
rect 8036 22545 8064 23054
rect 7932 22510 7984 22516
rect 8022 22536 8078 22545
rect 8022 22471 8078 22480
rect 7950 22332 8258 22341
rect 7950 22330 7956 22332
rect 8012 22330 8036 22332
rect 8092 22330 8116 22332
rect 8172 22330 8196 22332
rect 8252 22330 8258 22332
rect 8012 22278 8014 22330
rect 8194 22278 8196 22330
rect 7950 22276 7956 22278
rect 8012 22276 8036 22278
rect 8092 22276 8116 22278
rect 8172 22276 8196 22278
rect 8252 22276 8258 22278
rect 7950 22267 8258 22276
rect 8312 22234 8340 23831
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 7944 21729 7972 22034
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 7930 21720 7986 21729
rect 8220 21690 8248 21966
rect 7930 21655 7986 21664
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8208 21412 8260 21418
rect 8260 21372 8340 21400
rect 8208 21354 8260 21360
rect 7950 21244 8258 21253
rect 7950 21242 7956 21244
rect 8012 21242 8036 21244
rect 8092 21242 8116 21244
rect 8172 21242 8196 21244
rect 8252 21242 8258 21244
rect 8012 21190 8014 21242
rect 8194 21190 8196 21242
rect 7950 21188 7956 21190
rect 8012 21188 8036 21190
rect 8092 21188 8116 21190
rect 8172 21188 8196 21190
rect 8252 21188 8258 21190
rect 7950 21179 8258 21188
rect 8312 21146 8340 21372
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 7930 21040 7986 21049
rect 7930 20975 7932 20984
rect 7984 20975 7986 20984
rect 7932 20946 7984 20952
rect 7944 20330 7972 20946
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8128 20602 8156 20878
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8220 20346 8248 20742
rect 7932 20324 7984 20330
rect 8220 20318 8340 20346
rect 7932 20266 7984 20272
rect 7950 20156 8258 20165
rect 7950 20154 7956 20156
rect 8012 20154 8036 20156
rect 8092 20154 8116 20156
rect 8172 20154 8196 20156
rect 8252 20154 8258 20156
rect 8012 20102 8014 20154
rect 8194 20102 8196 20154
rect 7950 20100 7956 20102
rect 8012 20100 8036 20102
rect 8092 20100 8116 20102
rect 8172 20100 8196 20102
rect 8252 20100 8258 20102
rect 7950 20091 8258 20100
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7944 19514 7972 19722
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7932 19304 7984 19310
rect 7930 19272 7932 19281
rect 7984 19272 7986 19281
rect 7930 19207 7986 19216
rect 7950 19068 8258 19077
rect 7950 19066 7956 19068
rect 8012 19066 8036 19068
rect 8092 19066 8116 19068
rect 8172 19066 8196 19068
rect 8252 19066 8258 19068
rect 8012 19014 8014 19066
rect 8194 19014 8196 19066
rect 7950 19012 7956 19014
rect 8012 19012 8036 19014
rect 8092 19012 8116 19014
rect 8172 19012 8196 19014
rect 8252 19012 8258 19014
rect 7950 19003 8258 19012
rect 8312 18970 8340 20318
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 8114 18184 8170 18193
rect 7616 17836 7696 17864
rect 7564 17818 7616 17824
rect 7654 17776 7710 17785
rect 7654 17711 7710 17720
rect 7668 17678 7696 17711
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7576 16726 7604 17274
rect 7760 17202 7788 18158
rect 8114 18119 8116 18128
rect 8168 18119 8170 18128
rect 8116 18090 8168 18096
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7852 17134 7880 18022
rect 7950 17980 8258 17989
rect 7950 17978 7956 17980
rect 8012 17978 8036 17980
rect 8092 17978 8116 17980
rect 8172 17978 8196 17980
rect 8252 17978 8258 17980
rect 8012 17926 8014 17978
rect 8194 17926 8196 17978
rect 7950 17924 7956 17926
rect 8012 17924 8036 17926
rect 8092 17924 8116 17926
rect 8172 17924 8196 17926
rect 8252 17924 8258 17926
rect 7950 17915 8258 17924
rect 8312 17864 8340 18906
rect 8220 17836 8340 17864
rect 8220 17218 8248 17836
rect 8404 17678 8432 23990
rect 8496 23746 8524 24806
rect 8588 24750 8616 25112
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8588 24206 8616 24550
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8680 23866 8708 26551
rect 8772 24154 8800 26726
rect 8864 26382 8892 31078
rect 9324 30598 9352 31334
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9010 30492 9318 30501
rect 9010 30490 9016 30492
rect 9072 30490 9096 30492
rect 9152 30490 9176 30492
rect 9232 30490 9256 30492
rect 9312 30490 9318 30492
rect 9072 30438 9074 30490
rect 9254 30438 9256 30490
rect 9010 30436 9016 30438
rect 9072 30436 9096 30438
rect 9152 30436 9176 30438
rect 9232 30436 9256 30438
rect 9312 30436 9318 30438
rect 9010 30427 9318 30436
rect 9220 30388 9272 30394
rect 9220 30330 9272 30336
rect 9034 29744 9090 29753
rect 9034 29679 9090 29688
rect 9048 29646 9076 29679
rect 9036 29640 9088 29646
rect 9036 29582 9088 29588
rect 9232 29510 9260 30330
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 9220 29504 9272 29510
rect 9324 29492 9352 30194
rect 9416 29714 9444 31214
rect 9508 31113 9536 31894
rect 9494 31104 9550 31113
rect 9494 31039 9550 31048
rect 9600 30841 9628 31894
rect 9692 31385 9720 32166
rect 9678 31376 9734 31385
rect 9678 31311 9734 31320
rect 9772 31340 9824 31346
rect 9772 31282 9824 31288
rect 9680 30864 9732 30870
rect 9586 30832 9642 30841
rect 9680 30806 9732 30812
rect 9586 30767 9642 30776
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 9588 30592 9640 30598
rect 9692 30569 9720 30806
rect 9588 30534 9640 30540
rect 9678 30560 9734 30569
rect 9508 29889 9536 30534
rect 9494 29880 9550 29889
rect 9494 29815 9550 29824
rect 9600 29753 9628 30534
rect 9678 30495 9734 30504
rect 9784 30326 9812 31282
rect 9772 30320 9824 30326
rect 9772 30262 9824 30268
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9586 29744 9642 29753
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 9496 29708 9548 29714
rect 9586 29679 9642 29688
rect 9496 29650 9548 29656
rect 9324 29464 9444 29492
rect 9220 29446 9272 29452
rect 9010 29404 9318 29413
rect 9010 29402 9016 29404
rect 9072 29402 9096 29404
rect 9152 29402 9176 29404
rect 9232 29402 9256 29404
rect 9312 29402 9318 29404
rect 9072 29350 9074 29402
rect 9254 29350 9256 29402
rect 9010 29348 9016 29350
rect 9072 29348 9096 29350
rect 9152 29348 9176 29350
rect 9232 29348 9256 29350
rect 9312 29348 9318 29350
rect 9010 29339 9318 29348
rect 9220 29164 9272 29170
rect 9220 29106 9272 29112
rect 8942 29064 8998 29073
rect 8942 28999 8998 29008
rect 8956 28665 8984 28999
rect 8942 28656 8998 28665
rect 8942 28591 8998 28600
rect 9232 28529 9260 29106
rect 9416 28762 9444 29464
rect 9404 28756 9456 28762
rect 9404 28698 9456 28704
rect 9404 28552 9456 28558
rect 9218 28520 9274 28529
rect 9404 28494 9456 28500
rect 9218 28455 9274 28464
rect 9010 28316 9318 28325
rect 9010 28314 9016 28316
rect 9072 28314 9096 28316
rect 9152 28314 9176 28316
rect 9232 28314 9256 28316
rect 9312 28314 9318 28316
rect 9072 28262 9074 28314
rect 9254 28262 9256 28314
rect 9010 28260 9016 28262
rect 9072 28260 9096 28262
rect 9152 28260 9176 28262
rect 9232 28260 9256 28262
rect 9312 28260 9318 28262
rect 9010 28251 9318 28260
rect 9416 27713 9444 28494
rect 9508 28218 9536 29650
rect 9588 29504 9640 29510
rect 9588 29446 9640 29452
rect 9600 29209 9628 29446
rect 9586 29200 9642 29209
rect 9692 29170 9720 30126
rect 9772 29776 9824 29782
rect 9772 29718 9824 29724
rect 9784 29481 9812 29718
rect 9770 29472 9826 29481
rect 9770 29407 9826 29416
rect 9876 29186 9904 32506
rect 9968 30802 9996 33390
rect 10048 33312 10100 33318
rect 10152 33289 10180 35974
rect 10244 35306 10272 36246
rect 10336 36009 10364 37130
rect 10520 36825 10548 38694
rect 10782 38655 10838 38664
rect 10968 38208 11020 38214
rect 10968 38150 11020 38156
rect 10600 37664 10652 37670
rect 10600 37606 10652 37612
rect 10506 36816 10562 36825
rect 10506 36751 10562 36760
rect 10508 36644 10560 36650
rect 10508 36586 10560 36592
rect 10416 36576 10468 36582
rect 10416 36518 10468 36524
rect 10322 36000 10378 36009
rect 10322 35935 10378 35944
rect 10244 35278 10364 35306
rect 10232 35012 10284 35018
rect 10232 34954 10284 34960
rect 10244 34377 10272 34954
rect 10230 34368 10286 34377
rect 10230 34303 10286 34312
rect 10048 33254 10100 33260
rect 10138 33280 10194 33289
rect 10060 33130 10088 33254
rect 10138 33215 10194 33224
rect 10060 33102 10180 33130
rect 10152 31278 10180 33102
rect 10232 33040 10284 33046
rect 10232 32982 10284 32988
rect 10244 32473 10272 32982
rect 10230 32464 10286 32473
rect 10230 32399 10286 32408
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 10244 32201 10272 32234
rect 10230 32192 10286 32201
rect 10230 32127 10286 32136
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10244 31668 10272 31962
rect 10336 31754 10364 35278
rect 10428 34105 10456 36518
rect 10520 35465 10548 36586
rect 10612 35737 10640 37606
rect 10980 36281 11008 38150
rect 10966 36272 11022 36281
rect 10876 36236 10928 36242
rect 10966 36207 11022 36216
rect 10876 36178 10928 36184
rect 10598 35728 10654 35737
rect 10598 35663 10654 35672
rect 10506 35456 10562 35465
rect 10506 35391 10562 35400
rect 10600 34944 10652 34950
rect 10600 34886 10652 34892
rect 10414 34096 10470 34105
rect 10414 34031 10470 34040
rect 10612 33561 10640 34886
rect 10784 34060 10836 34066
rect 10784 34002 10836 34008
rect 10692 33924 10744 33930
rect 10692 33866 10744 33872
rect 10598 33552 10654 33561
rect 10598 33487 10654 33496
rect 10704 33017 10732 33866
rect 10690 33008 10746 33017
rect 10690 32943 10746 32952
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 10428 31929 10456 32710
rect 10414 31920 10470 31929
rect 10414 31855 10470 31864
rect 10796 31754 10824 34002
rect 10336 31726 10456 31754
rect 10244 31640 10364 31668
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 9956 30796 10008 30802
rect 9956 30738 10008 30744
rect 9956 30660 10008 30666
rect 9956 30602 10008 30608
rect 10048 30660 10100 30666
rect 10048 30602 10100 30608
rect 9968 30297 9996 30602
rect 9954 30288 10010 30297
rect 9954 30223 10010 30232
rect 9956 29572 10008 29578
rect 9956 29514 10008 29520
rect 9968 29209 9996 29514
rect 9586 29135 9642 29144
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 9784 29158 9904 29186
rect 9954 29200 10010 29209
rect 9588 29028 9640 29034
rect 9588 28970 9640 28976
rect 9680 29028 9732 29034
rect 9680 28970 9732 28976
rect 9600 28393 9628 28970
rect 9586 28384 9642 28393
rect 9586 28319 9642 28328
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 9692 28121 9720 28970
rect 9494 28112 9550 28121
rect 9494 28047 9550 28056
rect 9678 28112 9734 28121
rect 9678 28047 9734 28056
rect 9402 27704 9458 27713
rect 9402 27639 9458 27648
rect 9508 27588 9536 28047
rect 9784 27962 9812 29158
rect 9954 29135 10010 29144
rect 9864 29096 9916 29102
rect 9864 29038 9916 29044
rect 9956 29096 10008 29102
rect 9956 29038 10008 29044
rect 9416 27560 9536 27588
rect 9600 27934 9812 27962
rect 9128 27464 9180 27470
rect 9126 27432 9128 27441
rect 9180 27432 9182 27441
rect 9126 27367 9182 27376
rect 9010 27228 9318 27237
rect 9010 27226 9016 27228
rect 9072 27226 9096 27228
rect 9152 27226 9176 27228
rect 9232 27226 9256 27228
rect 9312 27226 9318 27228
rect 9072 27174 9074 27226
rect 9254 27174 9256 27226
rect 9010 27172 9016 27174
rect 9072 27172 9096 27174
rect 9152 27172 9176 27174
rect 9232 27172 9256 27174
rect 9312 27172 9318 27174
rect 9010 27163 9318 27172
rect 9416 26994 9444 27560
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9508 26994 9536 27270
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9324 26761 9352 26794
rect 9310 26752 9366 26761
rect 9600 26738 9628 27934
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9692 27305 9720 27814
rect 9678 27296 9734 27305
rect 9678 27231 9734 27240
rect 9772 26920 9824 26926
rect 9772 26862 9824 26868
rect 9310 26687 9366 26696
rect 9416 26710 9628 26738
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8956 26194 8984 26318
rect 8910 26166 8984 26194
rect 8910 26058 8938 26166
rect 9010 26140 9318 26149
rect 9010 26138 9016 26140
rect 9072 26138 9096 26140
rect 9152 26138 9176 26140
rect 9232 26138 9256 26140
rect 9312 26138 9318 26140
rect 9072 26086 9074 26138
rect 9254 26086 9256 26138
rect 9010 26084 9016 26086
rect 9072 26084 9096 26086
rect 9152 26084 9176 26086
rect 9232 26084 9256 26086
rect 9312 26084 9318 26086
rect 9010 26075 9318 26084
rect 8910 26030 8984 26058
rect 8850 25936 8906 25945
rect 8956 25922 8984 26030
rect 8956 25894 9076 25922
rect 8850 25871 8906 25880
rect 8864 24274 8892 25871
rect 8944 25832 8996 25838
rect 8944 25774 8996 25780
rect 8956 25430 8984 25774
rect 8944 25424 8996 25430
rect 8944 25366 8996 25372
rect 9048 25294 9076 25894
rect 9416 25378 9444 26710
rect 9588 26580 9640 26586
rect 9588 26522 9640 26528
rect 9496 26376 9548 26382
rect 9494 26344 9496 26353
rect 9548 26344 9550 26353
rect 9494 26279 9550 26288
rect 9496 25764 9548 25770
rect 9496 25706 9548 25712
rect 9508 25498 9536 25706
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9600 25401 9628 26522
rect 9692 25945 9720 26726
rect 9678 25936 9734 25945
rect 9678 25871 9734 25880
rect 9586 25392 9642 25401
rect 9416 25350 9536 25378
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9010 25052 9318 25061
rect 9010 25050 9016 25052
rect 9072 25050 9096 25052
rect 9152 25050 9176 25052
rect 9232 25050 9256 25052
rect 9312 25050 9318 25052
rect 9072 24998 9074 25050
rect 9254 24998 9256 25050
rect 9010 24996 9016 24998
rect 9072 24996 9096 24998
rect 9152 24996 9176 24998
rect 9232 24996 9256 24998
rect 9312 24996 9318 24998
rect 9010 24987 9318 24996
rect 9416 24886 9444 25230
rect 9404 24880 9456 24886
rect 9310 24848 9366 24857
rect 9404 24822 9456 24828
rect 9508 24834 9536 25350
rect 9586 25327 9642 25336
rect 9680 25152 9732 25158
rect 9678 25120 9680 25129
rect 9732 25120 9734 25129
rect 9678 25055 9734 25064
rect 9508 24806 9628 24834
rect 9310 24783 9366 24792
rect 8944 24744 8996 24750
rect 8944 24686 8996 24692
rect 8956 24342 8984 24686
rect 8944 24336 8996 24342
rect 8944 24278 8996 24284
rect 9126 24304 9182 24313
rect 8852 24268 8904 24274
rect 9126 24239 9182 24248
rect 8852 24210 8904 24216
rect 9140 24206 9168 24239
rect 9128 24200 9180 24206
rect 8772 24126 8892 24154
rect 9128 24142 9180 24148
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8496 23718 8708 23746
rect 8772 23730 8800 24006
rect 8864 23798 8892 24126
rect 9324 24052 9352 24783
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9324 24024 9444 24052
rect 9010 23964 9318 23973
rect 9010 23962 9016 23964
rect 9072 23962 9096 23964
rect 9152 23962 9176 23964
rect 9232 23962 9256 23964
rect 9312 23962 9318 23964
rect 9072 23910 9074 23962
rect 9254 23910 9256 23962
rect 9010 23908 9016 23910
rect 9072 23908 9096 23910
rect 9152 23908 9176 23910
rect 9232 23908 9256 23910
rect 9312 23908 9318 23910
rect 9010 23899 9318 23908
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8496 22030 8524 23462
rect 8576 23044 8628 23050
rect 8576 22986 8628 22992
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8482 21856 8538 21865
rect 8482 21791 8538 21800
rect 8496 21486 8524 21791
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8496 21049 8524 21422
rect 8482 21040 8538 21049
rect 8482 20975 8538 20984
rect 8588 20890 8616 22986
rect 8496 20862 8616 20890
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8312 17338 8340 17614
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8220 17190 8340 17218
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 8114 17096 8170 17105
rect 8114 17031 8116 17040
rect 8168 17031 8170 17040
rect 8116 17002 8168 17008
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 7562 16144 7618 16153
rect 7618 16088 7788 16096
rect 7562 16079 7564 16088
rect 7616 16068 7788 16088
rect 7564 16050 7616 16056
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7668 15609 7696 15642
rect 7654 15600 7710 15609
rect 7654 15535 7710 15544
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 15162 7696 15438
rect 7760 15162 7788 16068
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7392 12406 7512 12434
rect 7392 11354 7420 12406
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11898 7512 12174
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 9994 7328 10950
rect 7392 10674 7420 11290
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7484 10130 7512 11630
rect 7576 10810 7604 14894
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 13938 7696 14418
rect 7852 14414 7880 16934
rect 7950 16892 8258 16901
rect 7950 16890 7956 16892
rect 8012 16890 8036 16892
rect 8092 16890 8116 16892
rect 8172 16890 8196 16892
rect 8252 16890 8258 16892
rect 8012 16838 8014 16890
rect 8194 16838 8196 16890
rect 7950 16836 7956 16838
rect 8012 16836 8036 16838
rect 8092 16836 8116 16838
rect 8172 16836 8196 16838
rect 8252 16836 8258 16838
rect 7950 16827 8258 16836
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8022 16144 8078 16153
rect 8022 16079 8078 16088
rect 8036 15978 8064 16079
rect 8128 16046 8156 16390
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 7950 15804 8258 15813
rect 7950 15802 7956 15804
rect 8012 15802 8036 15804
rect 8092 15802 8116 15804
rect 8172 15802 8196 15804
rect 8252 15802 8258 15804
rect 8012 15750 8014 15802
rect 8194 15750 8196 15802
rect 7950 15748 7956 15750
rect 8012 15748 8036 15750
rect 8092 15748 8116 15750
rect 8172 15748 8196 15750
rect 8252 15748 8258 15750
rect 7950 15739 8258 15748
rect 7950 14716 8258 14725
rect 7950 14714 7956 14716
rect 8012 14714 8036 14716
rect 8092 14714 8116 14716
rect 8172 14714 8196 14716
rect 8252 14714 8258 14716
rect 8012 14662 8014 14714
rect 8194 14662 8196 14714
rect 7950 14660 7956 14662
rect 8012 14660 8036 14662
rect 8092 14660 8116 14662
rect 8172 14660 8196 14662
rect 8252 14660 8258 14662
rect 7950 14651 8258 14660
rect 7840 14408 7892 14414
rect 7760 14368 7840 14396
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7760 13818 7788 14368
rect 7840 14350 7892 14356
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8036 14074 8064 14350
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8128 13841 8156 14350
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8220 13870 8248 14010
rect 8208 13864 8260 13870
rect 7668 13790 7788 13818
rect 8114 13832 8170 13841
rect 7840 13796 7892 13802
rect 7668 13734 7696 13790
rect 8208 13806 8260 13812
rect 8114 13767 8170 13776
rect 7840 13738 7892 13744
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13530 7696 13670
rect 7746 13560 7802 13569
rect 7656 13524 7708 13530
rect 7746 13495 7748 13504
rect 7656 13466 7708 13472
rect 7800 13495 7802 13504
rect 7748 13466 7800 13472
rect 7668 13410 7696 13466
rect 7668 13382 7788 13410
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7668 12442 7696 13194
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7760 12322 7788 13382
rect 7852 12753 7880 13738
rect 7950 13628 8258 13637
rect 7950 13626 7956 13628
rect 8012 13626 8036 13628
rect 8092 13626 8116 13628
rect 8172 13626 8196 13628
rect 8252 13626 8258 13628
rect 8012 13574 8014 13626
rect 8194 13574 8196 13626
rect 7950 13572 7956 13574
rect 8012 13572 8036 13574
rect 8092 13572 8116 13574
rect 8172 13572 8196 13574
rect 8252 13572 8258 13574
rect 7950 13563 8258 13572
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 8208 13456 8260 13462
rect 8312 13444 8340 17190
rect 8404 16250 8432 17478
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8390 15192 8446 15201
rect 8390 15127 8446 15136
rect 8404 15026 8432 15127
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8404 14074 8432 14962
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8404 13734 8432 13874
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8390 13560 8446 13569
rect 8390 13495 8446 13504
rect 8260 13416 8340 13444
rect 8208 13398 8260 13404
rect 7944 12889 7972 13398
rect 8312 13138 8340 13416
rect 8404 13258 8432 13495
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8312 13110 8432 13138
rect 8298 13016 8354 13025
rect 8298 12951 8354 12960
rect 7930 12880 7986 12889
rect 8312 12850 8340 12951
rect 7930 12815 7986 12824
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7932 12776 7984 12782
rect 7838 12744 7894 12753
rect 8116 12776 8168 12782
rect 7932 12718 7984 12724
rect 8114 12744 8116 12753
rect 8168 12744 8170 12753
rect 7838 12679 7894 12688
rect 7944 12628 7972 12718
rect 8114 12679 8170 12688
rect 7852 12600 7972 12628
rect 7852 12434 7880 12600
rect 7950 12540 8258 12549
rect 7950 12538 7956 12540
rect 8012 12538 8036 12540
rect 8092 12538 8116 12540
rect 8172 12538 8196 12540
rect 8252 12538 8258 12540
rect 8012 12486 8014 12538
rect 8194 12486 8196 12538
rect 7950 12484 7956 12486
rect 8012 12484 8036 12486
rect 8092 12484 8116 12486
rect 8172 12484 8196 12486
rect 8252 12484 8258 12486
rect 7950 12475 8258 12484
rect 7852 12406 7972 12434
rect 7668 12294 7788 12322
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7300 7818 7328 9930
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7484 9489 7512 9522
rect 7470 9480 7526 9489
rect 7470 9415 7526 9424
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8537 7420 9318
rect 7378 8528 7434 8537
rect 7378 8463 7434 8472
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7993 7420 8366
rect 7378 7984 7434 7993
rect 7378 7919 7434 7928
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7286 7576 7342 7585
rect 7196 7540 7248 7546
rect 7286 7511 7342 7520
rect 7196 7482 7248 7488
rect 7300 7410 7328 7511
rect 7378 7440 7434 7449
rect 7288 7404 7340 7410
rect 7378 7375 7380 7384
rect 7288 7346 7340 7352
rect 7432 7375 7434 7384
rect 7380 7346 7432 7352
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6458 5944 6514 5953
rect 6564 5914 6592 6258
rect 6458 5879 6514 5888
rect 6552 5908 6604 5914
rect 6472 5846 6500 5879
rect 6552 5850 6604 5856
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6564 5778 6592 5850
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6748 5642 6776 6258
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 7300 5302 7328 7210
rect 7392 6934 7420 7346
rect 7484 7274 7512 9415
rect 7576 8838 7604 10542
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 7750 7604 8230
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7392 6458 7420 6870
rect 7576 6662 7604 7686
rect 7668 7546 7696 12294
rect 7838 11792 7894 11801
rect 7748 11756 7800 11762
rect 7838 11727 7894 11736
rect 7748 11698 7800 11704
rect 7760 8022 7788 11698
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7852 7834 7880 11727
rect 7944 11626 7972 12406
rect 8208 12368 8260 12374
rect 8206 12336 8208 12345
rect 8260 12336 8262 12345
rect 8206 12271 8262 12280
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11898 8248 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8312 11694 8340 12786
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7950 11452 8258 11461
rect 7950 11450 7956 11452
rect 8012 11450 8036 11452
rect 8092 11450 8116 11452
rect 8172 11450 8196 11452
rect 8252 11450 8258 11452
rect 8012 11398 8014 11450
rect 8194 11398 8196 11450
rect 7950 11396 7956 11398
rect 8012 11396 8036 11398
rect 8092 11396 8116 11398
rect 8172 11396 8196 11398
rect 8252 11396 8258 11398
rect 7950 11387 8258 11396
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10810 8340 11086
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8404 10656 8432 13110
rect 8496 11354 8524 20862
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8588 20466 8616 20742
rect 8680 20602 8708 23718
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8760 23316 8812 23322
rect 8760 23258 8812 23264
rect 8772 22030 8800 23258
rect 9324 23066 9352 23802
rect 9416 23186 9444 24024
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9324 23038 9444 23066
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 8864 22574 8892 22918
rect 9010 22876 9318 22885
rect 9010 22874 9016 22876
rect 9072 22874 9096 22876
rect 9152 22874 9176 22876
rect 9232 22874 9256 22876
rect 9312 22874 9318 22876
rect 9072 22822 9074 22874
rect 9254 22822 9256 22874
rect 9010 22820 9016 22822
rect 9072 22820 9096 22822
rect 9152 22820 9176 22822
rect 9232 22820 9256 22822
rect 9312 22820 9318 22822
rect 9010 22811 9318 22820
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 9416 22098 9444 23038
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9402 21992 9458 22001
rect 9232 21894 9260 21966
rect 9402 21927 9458 21936
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 8772 21146 8800 21830
rect 9010 21788 9318 21797
rect 9010 21786 9016 21788
rect 9072 21786 9096 21788
rect 9152 21786 9176 21788
rect 9232 21786 9256 21788
rect 9312 21786 9318 21788
rect 9072 21734 9074 21786
rect 9254 21734 9256 21786
rect 9010 21732 9016 21734
rect 9072 21732 9096 21734
rect 9152 21732 9176 21734
rect 9232 21732 9256 21734
rect 9312 21732 9318 21734
rect 9010 21723 9318 21732
rect 9416 21554 9444 21927
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9036 21480 9088 21486
rect 9034 21448 9036 21457
rect 9088 21448 9090 21457
rect 9034 21383 9090 21392
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8666 20496 8722 20505
rect 8576 20460 8628 20466
rect 8666 20431 8722 20440
rect 8576 20402 8628 20408
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8588 19514 8616 19790
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8588 18970 8616 19246
rect 8680 19174 8708 20431
rect 8772 20058 8800 20878
rect 9010 20700 9318 20709
rect 9010 20698 9016 20700
rect 9072 20698 9096 20700
rect 9152 20698 9176 20700
rect 9232 20698 9256 20700
rect 9312 20698 9318 20700
rect 9072 20646 9074 20698
rect 9254 20646 9256 20698
rect 9010 20644 9016 20646
rect 9072 20644 9096 20646
rect 9152 20644 9176 20646
rect 9232 20644 9256 20646
rect 9312 20644 9318 20646
rect 9010 20635 9318 20644
rect 9126 20496 9182 20505
rect 9036 20460 9088 20466
rect 9126 20431 9182 20440
rect 9220 20460 9272 20466
rect 9036 20402 9088 20408
rect 8944 20392 8996 20398
rect 8942 20360 8944 20369
rect 8996 20360 8998 20369
rect 8942 20295 8998 20304
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 9048 19825 9076 20402
rect 9140 19854 9168 20431
rect 9220 20402 9272 20408
rect 9128 19848 9180 19854
rect 9034 19816 9090 19825
rect 9128 19790 9180 19796
rect 9232 19786 9260 20402
rect 9034 19751 9090 19760
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8772 19496 8800 19654
rect 9010 19612 9318 19621
rect 9010 19610 9016 19612
rect 9072 19610 9096 19612
rect 9152 19610 9176 19612
rect 9232 19610 9256 19612
rect 9312 19610 9318 19612
rect 9072 19558 9074 19610
rect 9254 19558 9256 19610
rect 9010 19556 9016 19558
rect 9072 19556 9096 19558
rect 9152 19556 9176 19558
rect 9232 19556 9256 19558
rect 9312 19556 9318 19558
rect 9010 19547 9318 19556
rect 9416 19496 9444 21082
rect 8772 19468 9076 19496
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8772 18290 8800 18634
rect 8956 18578 8984 19343
rect 9048 19292 9076 19468
rect 9324 19468 9444 19496
rect 9128 19304 9180 19310
rect 9048 19264 9128 19292
rect 9128 19246 9180 19252
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 9048 18766 9076 18838
rect 9036 18760 9088 18766
rect 9324 18737 9352 19468
rect 9508 19378 9536 24618
rect 9600 23322 9628 24806
rect 9784 24682 9812 26862
rect 9772 24676 9824 24682
rect 9772 24618 9824 24624
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9770 24576 9826 24585
rect 9692 24313 9720 24550
rect 9770 24511 9826 24520
rect 9784 24410 9812 24511
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9678 24304 9734 24313
rect 9678 24239 9734 24248
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9692 23769 9720 23802
rect 9678 23760 9734 23769
rect 9678 23695 9734 23704
rect 9876 23594 9904 29038
rect 9968 26330 9996 29038
rect 10060 26926 10088 30602
rect 10140 30592 10192 30598
rect 10140 30534 10192 30540
rect 10152 27470 10180 30534
rect 10244 30025 10272 30874
rect 10336 30666 10364 31640
rect 10324 30660 10376 30666
rect 10324 30602 10376 30608
rect 10324 30116 10376 30122
rect 10324 30058 10376 30064
rect 10230 30016 10286 30025
rect 10230 29951 10286 29960
rect 10336 28937 10364 30058
rect 10428 29345 10456 31726
rect 10520 31726 10824 31754
rect 10414 29336 10470 29345
rect 10414 29271 10470 29280
rect 10322 28928 10378 28937
rect 10322 28863 10378 28872
rect 10232 28688 10284 28694
rect 10232 28630 10284 28636
rect 10244 27849 10272 28630
rect 10324 28620 10376 28626
rect 10324 28562 10376 28568
rect 10230 27840 10286 27849
rect 10230 27775 10286 27784
rect 10232 27600 10284 27606
rect 10232 27542 10284 27548
rect 10140 27464 10192 27470
rect 10140 27406 10192 27412
rect 10244 27033 10272 27542
rect 10336 27418 10364 28562
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10428 27577 10456 28358
rect 10414 27568 10470 27577
rect 10414 27503 10470 27512
rect 10336 27390 10456 27418
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10230 27024 10286 27033
rect 10230 26959 10286 26968
rect 10048 26920 10100 26926
rect 10048 26862 10100 26868
rect 10232 26512 10284 26518
rect 10232 26454 10284 26460
rect 9968 26302 10088 26330
rect 9954 26208 10010 26217
rect 9954 26143 10010 26152
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9680 23248 9732 23254
rect 9678 23216 9680 23225
rect 9732 23216 9734 23225
rect 9588 23180 9640 23186
rect 9678 23151 9734 23160
rect 9588 23122 9640 23128
rect 9600 22166 9628 23122
rect 9770 22672 9826 22681
rect 9770 22607 9826 22616
rect 9678 22400 9734 22409
rect 9678 22335 9734 22344
rect 9588 22160 9640 22166
rect 9588 22102 9640 22108
rect 9692 21978 9720 22335
rect 9600 21950 9720 21978
rect 9600 21894 9628 21950
rect 9784 21894 9812 22607
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9876 22137 9904 22442
rect 9862 22128 9918 22137
rect 9862 22063 9918 22072
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9588 21888 9640 21894
rect 9772 21888 9824 21894
rect 9588 21830 9640 21836
rect 9678 21856 9734 21865
rect 9772 21830 9824 21836
rect 9678 21791 9734 21800
rect 9692 21690 9720 21791
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9876 21593 9904 21898
rect 9862 21584 9918 21593
rect 9862 21519 9918 21528
rect 9678 21312 9734 21321
rect 9678 21247 9734 21256
rect 9692 21146 9720 21247
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9678 20768 9734 20777
rect 9678 20703 9734 20712
rect 9692 20602 9720 20703
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9404 19304 9456 19310
rect 9600 19258 9628 20470
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9678 20224 9734 20233
rect 9678 20159 9734 20168
rect 9692 20058 9720 20159
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9692 19417 9720 19450
rect 9678 19408 9734 19417
rect 9678 19343 9734 19352
rect 9404 19246 9456 19252
rect 9036 18702 9088 18708
rect 9310 18728 9366 18737
rect 9310 18663 9366 18672
rect 8864 18550 8984 18578
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8576 18216 8628 18222
rect 8864 18170 8892 18550
rect 9010 18524 9318 18533
rect 9010 18522 9016 18524
rect 9072 18522 9096 18524
rect 9152 18522 9176 18524
rect 9232 18522 9256 18524
rect 9312 18522 9318 18524
rect 9072 18470 9074 18522
rect 9254 18470 9256 18522
rect 9010 18468 9016 18470
rect 9072 18468 9096 18470
rect 9152 18468 9176 18470
rect 9232 18468 9256 18470
rect 9312 18468 9318 18470
rect 9010 18459 9318 18468
rect 9034 18320 9090 18329
rect 9034 18255 9090 18264
rect 8628 18164 8641 18170
rect 8576 18158 8641 18164
rect 8588 18142 8641 18158
rect 8864 18142 8984 18170
rect 8613 18136 8641 18142
rect 8613 18108 8708 18136
rect 8680 17524 8708 18108
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8588 17496 8708 17524
rect 8588 17134 8616 17496
rect 8772 17202 8800 17750
rect 8864 17678 8892 18022
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8956 17490 8984 18142
rect 9048 17746 9076 18255
rect 9416 17882 9444 19246
rect 9508 19230 9628 19258
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8864 17462 8984 17490
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16998 8616 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8588 16153 8616 16662
rect 8574 16144 8630 16153
rect 8574 16079 8630 16088
rect 8668 16108 8720 16114
rect 8588 14940 8616 16079
rect 8668 16050 8720 16056
rect 8680 15201 8708 16050
rect 8864 15638 8892 17462
rect 9010 17436 9318 17445
rect 9010 17434 9016 17436
rect 9072 17434 9096 17436
rect 9152 17434 9176 17436
rect 9232 17434 9256 17436
rect 9312 17434 9318 17436
rect 9072 17382 9074 17434
rect 9254 17382 9256 17434
rect 9010 17380 9016 17382
rect 9072 17380 9096 17382
rect 9152 17380 9176 17382
rect 9232 17380 9256 17382
rect 9312 17380 9318 17382
rect 9010 17371 9318 17380
rect 9508 17270 9536 19230
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9678 19136 9734 19145
rect 9600 17377 9628 19110
rect 9678 19071 9734 19080
rect 9692 18970 9720 19071
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9680 18760 9732 18766
rect 9678 18728 9680 18737
rect 9732 18728 9734 18737
rect 9678 18663 9734 18672
rect 9678 18592 9734 18601
rect 9678 18527 9734 18536
rect 9692 18426 9720 18527
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 17898 9812 20334
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9876 19174 9904 19722
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9876 18057 9904 18770
rect 9968 18766 9996 26143
rect 10060 26081 10088 26302
rect 10046 26072 10102 26081
rect 10046 26007 10102 26016
rect 10244 25673 10272 26454
rect 10336 26217 10364 27066
rect 10322 26208 10378 26217
rect 10322 26143 10378 26152
rect 10230 25664 10286 25673
rect 10230 25599 10286 25608
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10324 25424 10376 25430
rect 10324 25366 10376 25372
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 10060 20942 10088 25162
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10060 19961 10088 20198
rect 10046 19952 10102 19961
rect 10046 19887 10102 19896
rect 10048 19236 10100 19242
rect 10048 19178 10100 19184
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18329 9996 18566
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 9862 18048 9918 18057
rect 9862 17983 9918 17992
rect 9784 17870 9996 17898
rect 9770 17776 9826 17785
rect 9770 17711 9772 17720
rect 9824 17711 9826 17720
rect 9772 17682 9824 17688
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9692 17513 9720 17614
rect 9678 17504 9734 17513
rect 9678 17439 9734 17448
rect 9586 17368 9642 17377
rect 9586 17303 9642 17312
rect 9496 17264 9548 17270
rect 9310 17232 9366 17241
rect 9496 17206 9548 17212
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9770 17232 9826 17241
rect 9310 17167 9366 17176
rect 9324 16454 9352 17167
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9010 16348 9318 16357
rect 9010 16346 9016 16348
rect 9072 16346 9096 16348
rect 9152 16346 9176 16348
rect 9232 16346 9256 16348
rect 9312 16346 9318 16348
rect 9072 16294 9074 16346
rect 9254 16294 9256 16346
rect 9010 16292 9016 16294
rect 9072 16292 9096 16294
rect 9152 16292 9176 16294
rect 9232 16292 9256 16294
rect 9312 16292 9318 16294
rect 9010 16283 9318 16292
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8666 15192 8722 15201
rect 8666 15127 8722 15136
rect 8772 15065 8800 15438
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8758 15056 8814 15065
rect 8758 14991 8814 15000
rect 8668 14952 8720 14958
rect 8588 14912 8668 14940
rect 8588 12753 8616 14912
rect 8668 14894 8720 14900
rect 8864 14521 8892 15370
rect 9010 15260 9318 15269
rect 9010 15258 9016 15260
rect 9072 15258 9096 15260
rect 9152 15258 9176 15260
rect 9232 15258 9256 15260
rect 9312 15258 9318 15260
rect 9072 15206 9074 15258
rect 9254 15206 9256 15258
rect 9010 15204 9016 15206
rect 9072 15204 9096 15206
rect 9152 15204 9176 15206
rect 9232 15204 9256 15206
rect 9312 15204 9318 15206
rect 9010 15195 9318 15204
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 8666 14512 8722 14521
rect 8666 14447 8722 14456
rect 8850 14512 8906 14521
rect 9232 14482 9260 14894
rect 9310 14648 9366 14657
rect 9310 14583 9312 14592
rect 9364 14583 9366 14592
rect 9312 14554 9364 14560
rect 8850 14447 8906 14456
rect 9220 14476 9272 14482
rect 8680 14074 8708 14447
rect 9220 14418 9272 14424
rect 9416 14414 9444 15846
rect 9494 14920 9550 14929
rect 9494 14855 9496 14864
rect 9548 14855 9550 14864
rect 9496 14826 9548 14832
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8574 12744 8630 12753
rect 8574 12679 8630 12688
rect 8588 11694 8616 12679
rect 8680 12102 8708 13126
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8588 11014 8616 11630
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8680 10826 8708 11494
rect 8772 11014 8800 14214
rect 9010 14172 9318 14181
rect 9010 14170 9016 14172
rect 9072 14170 9096 14172
rect 9152 14170 9176 14172
rect 9232 14170 9256 14172
rect 9312 14170 9318 14172
rect 9072 14118 9074 14170
rect 9254 14118 9256 14170
rect 9010 14116 9016 14118
rect 9072 14116 9096 14118
rect 9152 14116 9176 14118
rect 9232 14116 9256 14118
rect 9312 14116 9318 14118
rect 9010 14107 9318 14116
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 13002 8892 13806
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9232 13326 9260 13398
rect 9324 13326 9352 13670
rect 9402 13560 9458 13569
rect 9402 13495 9458 13504
rect 9416 13326 9444 13495
rect 9600 13394 9628 17206
rect 9680 17196 9732 17202
rect 9770 17167 9826 17176
rect 9680 17138 9732 17144
rect 9692 16969 9720 17138
rect 9678 16960 9734 16969
rect 9678 16895 9734 16904
rect 9678 16688 9734 16697
rect 9784 16658 9812 17167
rect 9678 16623 9734 16632
rect 9772 16652 9824 16658
rect 9692 16182 9720 16623
rect 9772 16594 9824 16600
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9784 16425 9812 16458
rect 9770 16416 9826 16425
rect 9770 16351 9826 16360
rect 9680 16176 9732 16182
rect 9876 16153 9904 16526
rect 9680 16118 9732 16124
rect 9862 16144 9918 16153
rect 9862 16079 9918 16088
rect 9678 15872 9734 15881
rect 9678 15807 9734 15816
rect 9692 15094 9720 15807
rect 9968 15638 9996 17870
rect 9956 15632 10008 15638
rect 9770 15600 9826 15609
rect 9956 15574 10008 15580
rect 9770 15535 9772 15544
rect 9824 15535 9826 15544
rect 9772 15506 9824 15512
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9770 14784 9826 14793
rect 9770 14719 9826 14728
rect 9784 13938 9812 14719
rect 10060 14634 10088 19178
rect 9968 14618 10088 14634
rect 9956 14612 10088 14618
rect 10008 14606 10088 14612
rect 9956 14554 10008 14560
rect 9772 13932 9824 13938
rect 9968 13920 9996 14554
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 9772 13874 9824 13880
rect 9876 13892 9996 13920
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9010 13084 9318 13093
rect 9010 13082 9016 13084
rect 9072 13082 9096 13084
rect 9152 13082 9176 13084
rect 9232 13082 9256 13084
rect 9312 13082 9318 13084
rect 9072 13030 9074 13082
rect 9254 13030 9256 13082
rect 9010 13028 9016 13030
rect 9072 13028 9096 13030
rect 9152 13028 9176 13030
rect 9232 13028 9256 13030
rect 9312 13028 9318 13030
rect 9010 13019 9318 13028
rect 8864 12974 8984 13002
rect 9416 12986 9444 13126
rect 8850 12880 8906 12889
rect 8850 12815 8906 12824
rect 8864 11354 8892 12815
rect 8956 12782 8984 12974
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9508 12866 9536 13330
rect 9586 13288 9642 13297
rect 9586 13223 9642 13232
rect 9416 12850 9536 12866
rect 9404 12844 9536 12850
rect 9456 12838 9536 12844
rect 9404 12786 9456 12792
rect 8944 12776 8996 12782
rect 9600 12764 9628 13223
rect 9692 13161 9720 13466
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9678 13152 9734 13161
rect 9678 13087 9734 13096
rect 9784 12889 9812 13262
rect 9770 12880 9826 12889
rect 9770 12815 9826 12824
rect 8944 12718 8996 12724
rect 9508 12736 9628 12764
rect 8956 12442 8984 12718
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 9128 12368 9180 12374
rect 9126 12336 9128 12345
rect 9180 12336 9182 12345
rect 9126 12271 9182 12280
rect 9508 12238 9536 12736
rect 9876 12628 9904 13892
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9968 13462 9996 13631
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9954 13288 10010 13297
rect 9954 13223 10010 13232
rect 9600 12600 9904 12628
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 8944 12164 8996 12170
rect 9128 12164 9180 12170
rect 8996 12124 9128 12152
rect 8944 12106 8996 12112
rect 9128 12106 9180 12112
rect 9404 12164 9456 12170
rect 9404 12106 9456 12112
rect 9010 11996 9318 12005
rect 9010 11994 9016 11996
rect 9072 11994 9096 11996
rect 9152 11994 9176 11996
rect 9232 11994 9256 11996
rect 9312 11994 9318 11996
rect 9072 11942 9074 11994
rect 9254 11942 9256 11994
rect 9010 11940 9016 11942
rect 9072 11940 9096 11942
rect 9152 11940 9176 11942
rect 9232 11940 9256 11942
rect 9312 11940 9318 11942
rect 9010 11931 9318 11940
rect 9416 11898 9444 12106
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 8944 11688 8996 11694
rect 9128 11688 9180 11694
rect 8944 11630 8996 11636
rect 9126 11656 9128 11665
rect 9180 11656 9182 11665
rect 8956 11529 8984 11630
rect 9126 11591 9182 11600
rect 9220 11552 9272 11558
rect 8942 11520 8998 11529
rect 9220 11494 9272 11500
rect 8942 11455 8998 11464
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 9232 11218 9260 11494
rect 9494 11248 9550 11257
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9220 11212 9272 11218
rect 9494 11183 9550 11192
rect 9220 11154 9272 11160
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8680 10798 8800 10826
rect 8668 10668 8720 10674
rect 8404 10628 8668 10656
rect 8668 10610 8720 10616
rect 8482 10568 8538 10577
rect 8300 10532 8352 10538
rect 8482 10503 8538 10512
rect 8300 10474 8352 10480
rect 7950 10364 8258 10373
rect 7950 10362 7956 10364
rect 8012 10362 8036 10364
rect 8092 10362 8116 10364
rect 8172 10362 8196 10364
rect 8252 10362 8258 10364
rect 8012 10310 8014 10362
rect 8194 10310 8196 10362
rect 7950 10308 7956 10310
rect 8012 10308 8036 10310
rect 8092 10308 8116 10310
rect 8172 10308 8196 10310
rect 8252 10308 8258 10310
rect 7950 10299 8258 10308
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8024 9920 8076 9926
rect 8022 9888 8024 9897
rect 8076 9888 8078 9897
rect 8022 9823 8078 9832
rect 8128 9722 8156 9930
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9602 8248 10066
rect 8312 9722 8340 10474
rect 8496 10198 8524 10503
rect 8484 10192 8536 10198
rect 8536 10152 8708 10180
rect 8484 10134 8536 10140
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8220 9574 8340 9602
rect 7950 9276 8258 9285
rect 7950 9274 7956 9276
rect 8012 9274 8036 9276
rect 8092 9274 8116 9276
rect 8172 9274 8196 9276
rect 8252 9274 8258 9276
rect 8012 9222 8014 9274
rect 8194 9222 8196 9274
rect 7950 9220 7956 9222
rect 8012 9220 8036 9222
rect 8092 9220 8116 9222
rect 8172 9220 8196 9222
rect 8252 9220 8258 9222
rect 7950 9211 8258 9220
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8634 8248 8774
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8206 8528 8262 8537
rect 8206 8463 8262 8472
rect 8220 8430 8248 8463
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7760 7806 7880 7834
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 6934 7696 7210
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7392 5778 7420 6122
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7392 5234 7420 5714
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7484 2774 7512 6394
rect 7760 6322 7788 7806
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7840 7200 7892 7206
rect 8220 7188 8248 7346
rect 8312 7313 8340 9574
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8404 8974 8432 9522
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8298 7304 8354 7313
rect 8298 7239 8354 7248
rect 8220 7160 8340 7188
rect 7840 7142 7892 7148
rect 7852 6866 7880 7142
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8312 6882 8340 7160
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 8220 6854 8340 6882
rect 8220 6798 8248 6854
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7392 2746 7512 2774
rect 6918 2680 6974 2689
rect 6918 2615 6974 2624
rect 6458 1184 6514 1193
rect 6458 1119 6514 1128
rect 6472 56 6500 1119
rect 6932 56 6960 2615
rect 7392 56 7420 2746
rect 7852 56 7880 6054
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8404 5914 8432 8910
rect 8496 8673 8524 9046
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8496 8430 8524 8599
rect 8484 8424 8536 8430
rect 8588 8401 8616 9658
rect 8680 9625 8708 10152
rect 8772 9654 8800 10798
rect 8864 10713 8892 11154
rect 9140 11098 9168 11154
rect 9140 11070 9444 11098
rect 9010 10908 9318 10917
rect 9010 10906 9016 10908
rect 9072 10906 9096 10908
rect 9152 10906 9176 10908
rect 9232 10906 9256 10908
rect 9312 10906 9318 10908
rect 9072 10854 9074 10906
rect 9254 10854 9256 10906
rect 9010 10852 9016 10854
rect 9072 10852 9096 10854
rect 9152 10852 9176 10854
rect 9232 10852 9256 10854
rect 9312 10852 9318 10854
rect 9010 10843 9318 10852
rect 8850 10704 8906 10713
rect 8850 10639 8906 10648
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8864 10266 8892 10542
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8850 10160 8906 10169
rect 8850 10095 8906 10104
rect 8760 9648 8812 9654
rect 8666 9616 8722 9625
rect 8760 9590 8812 9596
rect 8666 9551 8722 9560
rect 8772 8922 8800 9590
rect 8864 9110 8892 10095
rect 9010 9820 9318 9829
rect 9010 9818 9016 9820
rect 9072 9818 9096 9820
rect 9152 9818 9176 9820
rect 9232 9818 9256 9820
rect 9312 9818 9318 9820
rect 9072 9766 9074 9818
rect 9254 9766 9256 9818
rect 9010 9764 9016 9766
rect 9072 9764 9096 9766
rect 9152 9764 9176 9766
rect 9232 9764 9256 9766
rect 9312 9764 9318 9766
rect 9010 9755 9318 9764
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9324 8945 9352 9046
rect 9416 8974 9444 11070
rect 9508 10606 9536 11183
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9496 10464 9548 10470
rect 9600 10452 9628 12600
rect 9968 12434 9996 13223
rect 10060 12646 10088 14486
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9968 12406 10088 12434
rect 9862 12336 9918 12345
rect 9862 12271 9864 12280
rect 9916 12271 9918 12280
rect 9864 12242 9916 12248
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 12073 9720 12106
rect 9678 12064 9734 12073
rect 9678 11999 9734 12008
rect 9784 11801 9812 12174
rect 9770 11792 9826 11801
rect 9770 11727 9826 11736
rect 9770 11520 9826 11529
rect 9770 11455 9826 11464
rect 9784 10674 9812 11455
rect 9954 11248 10010 11257
rect 9954 11183 10010 11192
rect 9968 11150 9996 11183
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10985 9904 11018
rect 9862 10976 9918 10985
rect 9862 10911 9918 10920
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9548 10424 9628 10452
rect 9770 10432 9826 10441
rect 9496 10406 9548 10412
rect 9770 10367 9826 10376
rect 9784 10130 9812 10367
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9772 10124 9824 10130
rect 10060 10112 10088 12406
rect 9772 10066 9824 10072
rect 9968 10084 10088 10112
rect 9496 9920 9548 9926
rect 9692 9897 9720 10066
rect 9496 9862 9548 9868
rect 9678 9888 9734 9897
rect 9508 9489 9536 9862
rect 9678 9823 9734 9832
rect 9772 9512 9824 9518
rect 9494 9480 9550 9489
rect 9772 9454 9824 9460
rect 9494 9415 9550 9424
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 8968 9456 8974
rect 8680 8894 8800 8922
rect 9310 8936 9366 8945
rect 8852 8900 8904 8906
rect 8680 8430 8708 8894
rect 9404 8910 9456 8916
rect 9310 8871 9366 8880
rect 8852 8842 8904 8848
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8668 8424 8720 8430
rect 8484 8366 8536 8372
rect 8574 8392 8630 8401
rect 8668 8366 8720 8372
rect 8574 8327 8630 8336
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 7478 8524 8230
rect 8680 8090 8708 8366
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8772 7886 8800 8774
rect 8864 8634 8892 8842
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9310 8528 9366 8537
rect 9310 8463 9366 8472
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8574 7576 8630 7585
rect 8574 7511 8630 7520
rect 8588 7478 8616 7511
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8576 7472 8628 7478
rect 8864 7449 8892 8298
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7857 8984 8026
rect 9232 7886 9260 8230
rect 9324 7993 9352 8463
rect 9416 8294 9444 8774
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9220 7880 9272 7886
rect 8942 7848 8998 7857
rect 9220 7822 9272 7828
rect 8942 7783 8998 7792
rect 9324 7732 9352 7919
rect 9416 7886 9444 8026
rect 9508 7886 9536 9318
rect 9784 9081 9812 9454
rect 9770 9072 9826 9081
rect 9770 9007 9826 9016
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9324 7704 9444 7732
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 8576 7414 8628 7420
rect 8850 7440 8906 7449
rect 8668 7404 8720 7410
rect 9416 7410 9444 7704
rect 9494 7712 9550 7721
rect 9494 7647 9550 7656
rect 9508 7410 9536 7647
rect 8850 7375 8852 7384
rect 8668 7346 8720 7352
rect 8904 7375 8906 7384
rect 9404 7404 9456 7410
rect 8852 7346 8904 7352
rect 9404 7346 9456 7352
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8496 5370 8524 6734
rect 8588 6662 8616 7142
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8680 6186 8708 7346
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9494 7304 9550 7313
rect 8772 6798 8800 7278
rect 9232 7206 9260 7278
rect 9494 7239 9496 7248
rect 9548 7239 9550 7248
rect 9496 7210 9548 7216
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8864 7002 8892 7142
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8298 5128 8354 5137
rect 8298 5063 8354 5072
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8312 56 8340 5063
rect 8772 56 8800 6598
rect 8864 6458 8892 6938
rect 9324 6866 9352 7142
rect 9402 6896 9458 6905
rect 9312 6860 9364 6866
rect 9402 6831 9458 6840
rect 9312 6802 9364 6808
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8864 6322 8892 6394
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9416 5370 9444 6831
rect 9494 6760 9550 6769
rect 9494 6695 9550 6704
rect 9508 5778 9536 6695
rect 9600 5914 9628 8910
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8537 9720 8842
rect 9876 8809 9904 8978
rect 9862 8800 9918 8809
rect 9862 8735 9918 8744
rect 9678 8528 9734 8537
rect 9678 8463 9734 8472
rect 9968 8378 9996 10084
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 9625 10088 9930
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 9968 8350 10088 8378
rect 9954 8256 10010 8265
rect 9954 8191 10010 8200
rect 9864 8016 9916 8022
rect 9678 7984 9734 7993
rect 9864 7958 9916 7964
rect 9678 7919 9680 7928
rect 9732 7919 9734 7928
rect 9680 7890 9732 7896
rect 9770 7712 9826 7721
rect 9770 7647 9826 7656
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9692 7177 9720 7482
rect 9784 7410 9812 7647
rect 9876 7449 9904 7958
rect 9968 7818 9996 8191
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 9956 7472 10008 7478
rect 9862 7440 9918 7449
rect 9772 7404 9824 7410
rect 9956 7414 10008 7420
rect 9862 7375 9918 7384
rect 9772 7346 9824 7352
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9968 6905 9996 7414
rect 9954 6896 10010 6905
rect 9954 6831 10010 6840
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6633 9720 6666
rect 9678 6624 9734 6633
rect 9678 6559 9734 6568
rect 9784 6361 9812 6734
rect 9770 6352 9826 6361
rect 9770 6287 9826 6296
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 6089 9812 6190
rect 10060 6118 10088 8350
rect 10048 6112 10100 6118
rect 9770 6080 9826 6089
rect 10048 6054 10100 6060
rect 9770 6015 9826 6024
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9678 5536 9734 5545
rect 9678 5471 9734 5480
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9692 5234 9720 5471
rect 9784 5273 9812 5646
rect 9770 5264 9826 5273
rect 9680 5228 9732 5234
rect 9770 5199 9826 5208
rect 9680 5170 9732 5176
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 10152 2774 10180 25298
rect 10244 24857 10272 25366
rect 10230 24848 10286 24857
rect 10230 24783 10286 24792
rect 10232 24336 10284 24342
rect 10232 24278 10284 24284
rect 10244 24041 10272 24278
rect 10230 24032 10286 24041
rect 10230 23967 10286 23976
rect 10232 23520 10284 23526
rect 10230 23488 10232 23497
rect 10284 23488 10286 23497
rect 10230 23423 10286 23432
rect 10232 22976 10284 22982
rect 10230 22944 10232 22953
rect 10284 22944 10286 22953
rect 10230 22879 10286 22888
rect 10232 22840 10284 22846
rect 10232 22782 10284 22788
rect 10244 21214 10272 22782
rect 10232 21208 10284 21214
rect 10232 21150 10284 21156
rect 10232 21072 10284 21078
rect 10230 21040 10232 21049
rect 10284 21040 10286 21049
rect 10230 20975 10286 20984
rect 10230 20496 10286 20505
rect 10230 20431 10286 20440
rect 10244 20330 10272 20431
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 10244 19689 10272 19926
rect 10230 19680 10286 19689
rect 10336 19666 10364 25366
rect 10428 19786 10456 27390
rect 10520 27062 10548 31726
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10612 28665 10640 29990
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10598 28656 10654 28665
rect 10598 28591 10654 28600
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10508 27056 10560 27062
rect 10508 26998 10560 27004
rect 10508 26920 10560 26926
rect 10508 26862 10560 26868
rect 10520 19854 10548 26862
rect 10612 26314 10640 27406
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10600 26172 10652 26178
rect 10600 26114 10652 26120
rect 10612 22846 10640 26114
rect 10600 22840 10652 22846
rect 10600 22782 10652 22788
rect 10600 22160 10652 22166
rect 10600 22102 10652 22108
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10336 19638 10548 19666
rect 10230 19615 10286 19624
rect 10414 19544 10470 19553
rect 10414 19479 10470 19488
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10232 18896 10284 18902
rect 10230 18864 10232 18873
rect 10284 18864 10286 18873
rect 10230 18799 10286 18808
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10244 12730 10272 18702
rect 10336 15473 10364 19314
rect 10322 15464 10378 15473
rect 10322 15399 10378 15408
rect 10322 13968 10378 13977
rect 10322 13903 10378 13912
rect 10336 12918 10364 13903
rect 10428 13297 10456 19479
rect 10520 15450 10548 19638
rect 10612 16794 10640 22102
rect 10704 21729 10732 29582
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10796 26489 10824 27270
rect 10782 26480 10838 26489
rect 10782 26415 10838 26424
rect 10888 25362 10916 36178
rect 11152 32836 11204 32842
rect 11152 32778 11204 32784
rect 11060 28484 11112 28490
rect 11060 28426 11112 28432
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10980 25242 11008 27338
rect 10888 25214 11008 25242
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10690 21720 10746 21729
rect 10690 21655 10746 21664
rect 10692 21208 10744 21214
rect 10692 21150 10744 21156
rect 10704 19378 10732 21150
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10690 19272 10746 19281
rect 10690 19207 10746 19216
rect 10704 17116 10732 19207
rect 10796 17218 10824 24754
rect 10888 19310 10916 25214
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10980 17270 11008 23598
rect 10968 17264 11020 17270
rect 10796 17190 10916 17218
rect 10968 17206 11020 17212
rect 10704 17088 10824 17116
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10520 15422 10640 15450
rect 10506 15328 10562 15337
rect 10506 15263 10562 15272
rect 10520 14414 10548 15263
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10414 13288 10470 13297
rect 10414 13223 10470 13232
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10244 12702 10364 12730
rect 10230 12608 10286 12617
rect 10230 12543 10286 12552
rect 10244 12102 10272 12543
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10244 8090 10272 11222
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10336 6662 10364 12702
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10520 6390 10548 13330
rect 10612 12714 10640 15422
rect 10690 14240 10746 14249
rect 10690 14175 10746 14184
rect 10704 12850 10732 14175
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10796 12730 10824 17088
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10704 12702 10824 12730
rect 10704 12434 10732 12702
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10612 12406 10732 12434
rect 10612 11354 10640 12406
rect 10796 11914 10824 12582
rect 10704 11886 10824 11914
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10704 6934 10732 11886
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 10169 10824 11698
rect 10782 10160 10838 10169
rect 10782 10095 10838 10104
rect 10888 9722 10916 17190
rect 11072 16726 11100 28426
rect 11164 25430 11192 32778
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11164 15706 11192 22034
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10966 13424 11022 13433
rect 10966 13359 11022 13368
rect 10980 13258 11008 13359
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10966 9344 11022 9353
rect 10966 9279 11022 9288
rect 10980 7886 11008 9279
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10690 5808 10746 5817
rect 10690 5743 10746 5752
rect 10704 5234 10732 5743
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10060 2746 10180 2774
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9218 1184 9274 1193
rect 9218 1119 9274 1128
rect 9232 56 9260 1119
rect 9692 56 9812 82
rect 6104 14 6224 42
rect 6458 0 6514 56
rect 6918 0 6974 56
rect 7378 0 7434 56
rect 7838 0 7894 56
rect 8298 0 8354 56
rect 8758 0 8814 56
rect 9218 0 9274 56
rect 9678 54 9812 56
rect 9678 0 9734 54
rect 9784 42 9812 54
rect 10060 42 10088 2746
rect 10138 1320 10194 1329
rect 10138 1255 10194 1264
rect 10152 56 10180 1255
rect 9784 14 10088 42
rect 10138 0 10194 56
<< via2 >>
rect 3016 42458 3072 42460
rect 3096 42458 3152 42460
rect 3176 42458 3232 42460
rect 3256 42458 3312 42460
rect 3016 42406 3062 42458
rect 3062 42406 3072 42458
rect 3096 42406 3126 42458
rect 3126 42406 3138 42458
rect 3138 42406 3152 42458
rect 3176 42406 3190 42458
rect 3190 42406 3202 42458
rect 3202 42406 3232 42458
rect 3256 42406 3266 42458
rect 3266 42406 3312 42458
rect 3016 42404 3072 42406
rect 3096 42404 3152 42406
rect 3176 42404 3232 42406
rect 3256 42404 3312 42406
rect 1956 41914 2012 41916
rect 2036 41914 2092 41916
rect 2116 41914 2172 41916
rect 2196 41914 2252 41916
rect 1956 41862 2002 41914
rect 2002 41862 2012 41914
rect 2036 41862 2066 41914
rect 2066 41862 2078 41914
rect 2078 41862 2092 41914
rect 2116 41862 2130 41914
rect 2130 41862 2142 41914
rect 2142 41862 2172 41914
rect 2196 41862 2206 41914
rect 2206 41862 2252 41914
rect 1956 41860 2012 41862
rect 2036 41860 2092 41862
rect 2116 41860 2172 41862
rect 2196 41860 2252 41862
rect 202 31728 258 31784
rect 18 28056 74 28112
rect 202 25744 258 25800
rect 18 23160 74 23216
rect 386 33496 442 33552
rect 386 28600 442 28656
rect 386 24928 442 24984
rect 754 38392 810 38448
rect 754 32680 810 32736
rect 1122 34992 1178 35048
rect 938 34312 994 34368
rect 662 29008 718 29064
rect 662 26424 718 26480
rect 662 26152 718 26208
rect 202 18128 258 18184
rect 662 17176 718 17232
rect 846 31048 902 31104
rect 846 29960 902 30016
rect 846 29008 902 29064
rect 1490 40840 1546 40896
rect 1490 40024 1546 40080
rect 1490 39208 1546 39264
rect 1956 40826 2012 40828
rect 2036 40826 2092 40828
rect 2116 40826 2172 40828
rect 2196 40826 2252 40828
rect 1956 40774 2002 40826
rect 2002 40774 2012 40826
rect 2036 40774 2066 40826
rect 2066 40774 2078 40826
rect 2078 40774 2092 40826
rect 2116 40774 2130 40826
rect 2130 40774 2142 40826
rect 2142 40774 2172 40826
rect 2196 40774 2206 40826
rect 2206 40774 2252 40826
rect 1956 40772 2012 40774
rect 2036 40772 2092 40774
rect 2116 40772 2172 40774
rect 2196 40772 2252 40774
rect 1956 39738 2012 39740
rect 2036 39738 2092 39740
rect 2116 39738 2172 39740
rect 2196 39738 2252 39740
rect 1956 39686 2002 39738
rect 2002 39686 2012 39738
rect 2036 39686 2066 39738
rect 2066 39686 2078 39738
rect 2078 39686 2092 39738
rect 2116 39686 2130 39738
rect 2130 39686 2142 39738
rect 2142 39686 2172 39738
rect 2196 39686 2206 39738
rect 2206 39686 2252 39738
rect 1956 39684 2012 39686
rect 2036 39684 2092 39686
rect 2116 39684 2172 39686
rect 2196 39684 2252 39686
rect 1956 38650 2012 38652
rect 2036 38650 2092 38652
rect 2116 38650 2172 38652
rect 2196 38650 2252 38652
rect 1956 38598 2002 38650
rect 2002 38598 2012 38650
rect 2036 38598 2066 38650
rect 2066 38598 2078 38650
rect 2078 38598 2092 38650
rect 2116 38598 2130 38650
rect 2130 38598 2142 38650
rect 2142 38598 2172 38650
rect 2196 38598 2206 38650
rect 2206 38598 2252 38650
rect 1956 38596 2012 38598
rect 2036 38596 2092 38598
rect 2116 38596 2172 38598
rect 2196 38596 2252 38598
rect 1490 37576 1546 37632
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 1490 36760 1546 36816
rect 1674 36760 1730 36816
rect 1490 35944 1546 36000
rect 1490 35128 1546 35184
rect 1306 30232 1362 30288
rect 1122 26832 1178 26888
rect 1122 26288 1178 26344
rect 846 20440 902 20496
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 1858 35944 1914 36000
rect 1674 35536 1730 35592
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 3016 41370 3072 41372
rect 3096 41370 3152 41372
rect 3176 41370 3232 41372
rect 3256 41370 3312 41372
rect 3016 41318 3062 41370
rect 3062 41318 3072 41370
rect 3096 41318 3126 41370
rect 3126 41318 3138 41370
rect 3138 41318 3152 41370
rect 3176 41318 3190 41370
rect 3190 41318 3202 41370
rect 3202 41318 3232 41370
rect 3256 41318 3266 41370
rect 3266 41318 3312 41370
rect 3016 41316 3072 41318
rect 3096 41316 3152 41318
rect 3176 41316 3232 41318
rect 3256 41316 3312 41318
rect 3016 40282 3072 40284
rect 3096 40282 3152 40284
rect 3176 40282 3232 40284
rect 3256 40282 3312 40284
rect 3016 40230 3062 40282
rect 3062 40230 3072 40282
rect 3096 40230 3126 40282
rect 3126 40230 3138 40282
rect 3138 40230 3152 40282
rect 3176 40230 3190 40282
rect 3190 40230 3202 40282
rect 3202 40230 3232 40282
rect 3256 40230 3266 40282
rect 3266 40230 3312 40282
rect 3016 40228 3072 40230
rect 3096 40228 3152 40230
rect 3176 40228 3232 40230
rect 3256 40228 3312 40230
rect 1490 31864 1546 31920
rect 1490 30096 1546 30152
rect 1674 32852 1676 32872
rect 1676 32852 1728 32872
rect 1728 32852 1730 32872
rect 1674 32816 1730 32852
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 2042 31864 2098 31920
rect 1398 29416 1454 29472
rect 1398 29144 1454 29200
rect 1398 27784 1454 27840
rect 1490 27376 1546 27432
rect 1398 26988 1454 27024
rect 1398 26968 1400 26988
rect 1400 26968 1452 26988
rect 1452 26968 1454 26988
rect 1398 25336 1454 25392
rect 1398 24520 1454 24576
rect 1674 28872 1730 28928
rect 2226 31184 2282 31240
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 2410 29552 2466 29608
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 2134 27920 2190 27976
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 1858 27512 1914 27568
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 1398 23704 1454 23760
rect 1398 22888 1454 22944
rect 1398 22072 1454 22128
rect 1490 21936 1546 21992
rect 1398 21256 1454 21312
rect 1398 20576 1454 20632
rect 1398 19624 1454 19680
rect 1398 18808 1454 18864
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 2134 24656 2190 24712
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 3016 39194 3072 39196
rect 3096 39194 3152 39196
rect 3176 39194 3232 39196
rect 3256 39194 3312 39196
rect 3016 39142 3062 39194
rect 3062 39142 3072 39194
rect 3096 39142 3126 39194
rect 3126 39142 3138 39194
rect 3138 39142 3152 39194
rect 3176 39142 3190 39194
rect 3190 39142 3202 39194
rect 3202 39142 3232 39194
rect 3256 39142 3266 39194
rect 3266 39142 3312 39194
rect 3016 39140 3072 39142
rect 3096 39140 3152 39142
rect 3176 39140 3232 39142
rect 3256 39140 3312 39142
rect 3016 38106 3072 38108
rect 3096 38106 3152 38108
rect 3176 38106 3232 38108
rect 3256 38106 3312 38108
rect 3016 38054 3062 38106
rect 3062 38054 3072 38106
rect 3096 38054 3126 38106
rect 3126 38054 3138 38106
rect 3138 38054 3152 38106
rect 3176 38054 3190 38106
rect 3190 38054 3202 38106
rect 3202 38054 3232 38106
rect 3256 38054 3266 38106
rect 3266 38054 3312 38106
rect 3016 38052 3072 38054
rect 3096 38052 3152 38054
rect 3176 38052 3232 38054
rect 3256 38052 3312 38054
rect 3016 37018 3072 37020
rect 3096 37018 3152 37020
rect 3176 37018 3232 37020
rect 3256 37018 3312 37020
rect 3016 36966 3062 37018
rect 3062 36966 3072 37018
rect 3096 36966 3126 37018
rect 3126 36966 3138 37018
rect 3138 36966 3152 37018
rect 3176 36966 3190 37018
rect 3190 36966 3202 37018
rect 3202 36966 3232 37018
rect 3256 36966 3266 37018
rect 3266 36966 3312 37018
rect 3016 36964 3072 36966
rect 3096 36964 3152 36966
rect 3176 36964 3232 36966
rect 3256 36964 3312 36966
rect 2778 35672 2834 35728
rect 3016 35930 3072 35932
rect 3096 35930 3152 35932
rect 3176 35930 3232 35932
rect 3256 35930 3312 35932
rect 3016 35878 3062 35930
rect 3062 35878 3072 35930
rect 3096 35878 3126 35930
rect 3126 35878 3138 35930
rect 3138 35878 3152 35930
rect 3176 35878 3190 35930
rect 3190 35878 3202 35930
rect 3202 35878 3232 35930
rect 3256 35878 3266 35930
rect 3266 35878 3312 35930
rect 3016 35876 3072 35878
rect 3096 35876 3152 35878
rect 3176 35876 3232 35878
rect 3256 35876 3312 35878
rect 3238 35128 3294 35184
rect 3016 34842 3072 34844
rect 3096 34842 3152 34844
rect 3176 34842 3232 34844
rect 3256 34842 3312 34844
rect 3016 34790 3062 34842
rect 3062 34790 3072 34842
rect 3096 34790 3126 34842
rect 3126 34790 3138 34842
rect 3138 34790 3152 34842
rect 3176 34790 3190 34842
rect 3190 34790 3202 34842
rect 3202 34790 3232 34842
rect 3256 34790 3266 34842
rect 3266 34790 3312 34842
rect 3016 34788 3072 34790
rect 3096 34788 3152 34790
rect 3176 34788 3232 34790
rect 3256 34788 3312 34790
rect 3016 33754 3072 33756
rect 3096 33754 3152 33756
rect 3176 33754 3232 33756
rect 3256 33754 3312 33756
rect 3016 33702 3062 33754
rect 3062 33702 3072 33754
rect 3096 33702 3126 33754
rect 3126 33702 3138 33754
rect 3138 33702 3152 33754
rect 3176 33702 3190 33754
rect 3190 33702 3202 33754
rect 3202 33702 3232 33754
rect 3256 33702 3266 33754
rect 3266 33702 3312 33754
rect 3016 33700 3072 33702
rect 3096 33700 3152 33702
rect 3176 33700 3232 33702
rect 3256 33700 3312 33702
rect 3016 32666 3072 32668
rect 3096 32666 3152 32668
rect 3176 32666 3232 32668
rect 3256 32666 3312 32668
rect 3016 32614 3062 32666
rect 3062 32614 3072 32666
rect 3096 32614 3126 32666
rect 3126 32614 3138 32666
rect 3138 32614 3152 32666
rect 3176 32614 3190 32666
rect 3190 32614 3202 32666
rect 3202 32614 3232 32666
rect 3256 32614 3266 32666
rect 3266 32614 3312 32666
rect 3016 32612 3072 32614
rect 3096 32612 3152 32614
rect 3176 32612 3232 32614
rect 3256 32612 3312 32614
rect 3016 31578 3072 31580
rect 3096 31578 3152 31580
rect 3176 31578 3232 31580
rect 3256 31578 3312 31580
rect 3016 31526 3062 31578
rect 3062 31526 3072 31578
rect 3096 31526 3126 31578
rect 3126 31526 3138 31578
rect 3138 31526 3152 31578
rect 3176 31526 3190 31578
rect 3190 31526 3202 31578
rect 3202 31526 3232 31578
rect 3256 31526 3266 31578
rect 3266 31526 3312 31578
rect 3016 31524 3072 31526
rect 3096 31524 3152 31526
rect 3176 31524 3232 31526
rect 3256 31524 3312 31526
rect 2778 30232 2834 30288
rect 2686 29008 2742 29064
rect 3016 30490 3072 30492
rect 3096 30490 3152 30492
rect 3176 30490 3232 30492
rect 3256 30490 3312 30492
rect 3016 30438 3062 30490
rect 3062 30438 3072 30490
rect 3096 30438 3126 30490
rect 3126 30438 3138 30490
rect 3138 30438 3152 30490
rect 3176 30438 3190 30490
rect 3190 30438 3202 30490
rect 3202 30438 3232 30490
rect 3256 30438 3266 30490
rect 3266 30438 3312 30490
rect 3016 30436 3072 30438
rect 3096 30436 3152 30438
rect 3176 30436 3232 30438
rect 3256 30436 3312 30438
rect 3882 35808 3938 35864
rect 4526 37204 4528 37224
rect 4528 37204 4580 37224
rect 4580 37204 4582 37224
rect 4526 37168 4582 37204
rect 3016 29402 3072 29404
rect 3096 29402 3152 29404
rect 3176 29402 3232 29404
rect 3256 29402 3312 29404
rect 3016 29350 3062 29402
rect 3062 29350 3072 29402
rect 3096 29350 3126 29402
rect 3126 29350 3138 29402
rect 3138 29350 3152 29402
rect 3176 29350 3190 29402
rect 3190 29350 3202 29402
rect 3202 29350 3232 29402
rect 3256 29350 3266 29402
rect 3266 29350 3312 29402
rect 3016 29348 3072 29350
rect 3096 29348 3152 29350
rect 3176 29348 3232 29350
rect 3256 29348 3312 29350
rect 2870 28464 2926 28520
rect 3790 30504 3846 30560
rect 3698 30232 3754 30288
rect 3422 29008 3478 29064
rect 3016 28314 3072 28316
rect 3096 28314 3152 28316
rect 3176 28314 3232 28316
rect 3256 28314 3312 28316
rect 3016 28262 3062 28314
rect 3062 28262 3072 28314
rect 3096 28262 3126 28314
rect 3126 28262 3138 28314
rect 3138 28262 3152 28314
rect 3176 28262 3190 28314
rect 3190 28262 3202 28314
rect 3202 28262 3232 28314
rect 3256 28262 3266 28314
rect 3266 28262 3312 28314
rect 3016 28260 3072 28262
rect 3096 28260 3152 28262
rect 3176 28260 3232 28262
rect 3256 28260 3312 28262
rect 3054 27820 3056 27840
rect 3056 27820 3108 27840
rect 3108 27820 3110 27840
rect 3054 27784 3110 27820
rect 3016 27226 3072 27228
rect 3096 27226 3152 27228
rect 3176 27226 3232 27228
rect 3256 27226 3312 27228
rect 3016 27174 3062 27226
rect 3062 27174 3072 27226
rect 3096 27174 3126 27226
rect 3126 27174 3138 27226
rect 3138 27174 3152 27226
rect 3176 27174 3190 27226
rect 3190 27174 3202 27226
rect 3202 27174 3232 27226
rect 3256 27174 3266 27226
rect 3266 27174 3312 27226
rect 3016 27172 3072 27174
rect 3096 27172 3152 27174
rect 3176 27172 3232 27174
rect 3256 27172 3312 27174
rect 2870 26832 2926 26888
rect 2686 25880 2742 25936
rect 2502 25472 2558 25528
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 1950 23196 1952 23216
rect 1952 23196 2004 23216
rect 2004 23196 2006 23216
rect 1950 23160 2006 23196
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 2226 21392 2282 21448
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 2042 20984 2098 21040
rect 2318 20304 2374 20360
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 1030 12280 1086 12336
rect 846 10648 902 10704
rect 846 8200 902 8256
rect 1030 9696 1086 9752
rect 1214 15544 1270 15600
rect 1398 17992 1454 18048
rect 1398 16360 1454 16416
rect 1214 14864 1270 14920
rect 2318 19760 2374 19816
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1490 13912 1546 13968
rect 2686 23160 2742 23216
rect 3016 26138 3072 26140
rect 3096 26138 3152 26140
rect 3176 26138 3232 26140
rect 3256 26138 3312 26140
rect 3016 26086 3062 26138
rect 3062 26086 3072 26138
rect 3096 26086 3126 26138
rect 3126 26086 3138 26138
rect 3138 26086 3152 26138
rect 3176 26086 3190 26138
rect 3190 26086 3202 26138
rect 3202 26086 3232 26138
rect 3256 26086 3266 26138
rect 3266 26086 3312 26138
rect 3016 26084 3072 26086
rect 3096 26084 3152 26086
rect 3176 26084 3232 26086
rect 3256 26084 3312 26086
rect 3016 25050 3072 25052
rect 3096 25050 3152 25052
rect 3176 25050 3232 25052
rect 3256 25050 3312 25052
rect 3016 24998 3062 25050
rect 3062 24998 3072 25050
rect 3096 24998 3126 25050
rect 3126 24998 3138 25050
rect 3138 24998 3152 25050
rect 3176 24998 3190 25050
rect 3190 24998 3202 25050
rect 3202 24998 3232 25050
rect 3256 24998 3266 25050
rect 3266 24998 3312 25050
rect 3016 24996 3072 24998
rect 3096 24996 3152 24998
rect 3176 24996 3232 24998
rect 3256 24996 3312 24998
rect 2962 24112 3018 24168
rect 3146 24112 3202 24168
rect 3016 23962 3072 23964
rect 3096 23962 3152 23964
rect 3176 23962 3232 23964
rect 3256 23962 3312 23964
rect 3016 23910 3062 23962
rect 3062 23910 3072 23962
rect 3096 23910 3126 23962
rect 3126 23910 3138 23962
rect 3138 23910 3152 23962
rect 3176 23910 3190 23962
rect 3190 23910 3202 23962
rect 3202 23910 3232 23962
rect 3256 23910 3266 23962
rect 3266 23910 3312 23962
rect 3016 23908 3072 23910
rect 3096 23908 3152 23910
rect 3176 23908 3232 23910
rect 3256 23908 3312 23910
rect 2962 23704 3018 23760
rect 3238 23740 3240 23760
rect 3240 23740 3292 23760
rect 3292 23740 3294 23760
rect 3238 23704 3294 23740
rect 2686 21936 2742 21992
rect 2410 17312 2466 17368
rect 3016 22874 3072 22876
rect 3096 22874 3152 22876
rect 3176 22874 3232 22876
rect 3256 22874 3312 22876
rect 3016 22822 3062 22874
rect 3062 22822 3072 22874
rect 3096 22822 3126 22874
rect 3126 22822 3138 22874
rect 3138 22822 3152 22874
rect 3176 22822 3190 22874
rect 3190 22822 3202 22874
rect 3202 22822 3232 22874
rect 3256 22822 3266 22874
rect 3266 22822 3312 22874
rect 3016 22820 3072 22822
rect 3096 22820 3152 22822
rect 3176 22820 3232 22822
rect 3256 22820 3312 22822
rect 3238 22616 3294 22672
rect 3330 22344 3386 22400
rect 3790 28600 3846 28656
rect 3606 26016 3662 26072
rect 3016 21786 3072 21788
rect 3096 21786 3152 21788
rect 3176 21786 3232 21788
rect 3256 21786 3312 21788
rect 3016 21734 3062 21786
rect 3062 21734 3072 21786
rect 3096 21734 3126 21786
rect 3126 21734 3138 21786
rect 3138 21734 3152 21786
rect 3176 21734 3190 21786
rect 3190 21734 3202 21786
rect 3202 21734 3232 21786
rect 3256 21734 3266 21786
rect 3266 21734 3312 21786
rect 3016 21732 3072 21734
rect 3096 21732 3152 21734
rect 3176 21732 3232 21734
rect 3256 21732 3312 21734
rect 3016 20698 3072 20700
rect 3096 20698 3152 20700
rect 3176 20698 3232 20700
rect 3256 20698 3312 20700
rect 3016 20646 3062 20698
rect 3062 20646 3072 20698
rect 3096 20646 3126 20698
rect 3126 20646 3138 20698
rect 3138 20646 3152 20698
rect 3176 20646 3190 20698
rect 3190 20646 3202 20698
rect 3202 20646 3232 20698
rect 3256 20646 3266 20698
rect 3266 20646 3312 20698
rect 3016 20644 3072 20646
rect 3096 20644 3152 20646
rect 3176 20644 3232 20646
rect 3256 20644 3312 20646
rect 2870 19896 2926 19952
rect 3016 19610 3072 19612
rect 3096 19610 3152 19612
rect 3176 19610 3232 19612
rect 3256 19610 3312 19612
rect 3016 19558 3062 19610
rect 3062 19558 3072 19610
rect 3096 19558 3126 19610
rect 3126 19558 3138 19610
rect 3138 19558 3152 19610
rect 3176 19558 3190 19610
rect 3190 19558 3202 19610
rect 3202 19558 3232 19610
rect 3256 19558 3266 19610
rect 3266 19558 3312 19610
rect 3016 19556 3072 19558
rect 3096 19556 3152 19558
rect 3176 19556 3232 19558
rect 3256 19556 3312 19558
rect 2318 17040 2374 17096
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1490 13132 1492 13152
rect 1492 13132 1544 13152
rect 1544 13132 1546 13152
rect 1490 13096 1546 13132
rect 1490 11500 1492 11520
rect 1492 11500 1544 11520
rect 1544 11500 1546 11520
rect 1490 11464 1546 11500
rect 1490 10920 1546 10976
rect 1490 9868 1492 9888
rect 1492 9868 1544 9888
rect 1544 9868 1546 9888
rect 1490 9832 1546 9868
rect 1490 9016 1546 9072
rect 1490 7384 1546 7440
rect 1398 6568 1454 6624
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1950 11076 2006 11112
rect 1950 11056 1952 11076
rect 1952 11056 2004 11076
rect 2004 11056 2006 11076
rect 2042 10512 2098 10568
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1950 10104 2006 10160
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2042 7928 2098 7984
rect 2686 17856 2742 17912
rect 2778 16632 2834 16688
rect 2410 8200 2466 8256
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2962 19352 3018 19408
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 3176 18522 3232 18524
rect 3256 18522 3312 18524
rect 3016 18470 3062 18522
rect 3062 18470 3072 18522
rect 3096 18470 3126 18522
rect 3126 18470 3138 18522
rect 3138 18470 3152 18522
rect 3176 18470 3190 18522
rect 3190 18470 3202 18522
rect 3202 18470 3232 18522
rect 3256 18470 3266 18522
rect 3266 18470 3312 18522
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 3176 18468 3232 18470
rect 3256 18468 3312 18470
rect 3330 17992 3386 18048
rect 3514 22208 3570 22264
rect 3882 26288 3938 26344
rect 3882 23432 3938 23488
rect 3698 22072 3754 22128
rect 3790 21664 3846 21720
rect 3790 21120 3846 21176
rect 4158 33396 4160 33416
rect 4160 33396 4212 33416
rect 4212 33396 4214 33416
rect 4158 33360 4214 33396
rect 4066 30368 4122 30424
rect 4342 31864 4398 31920
rect 4342 31592 4398 31648
rect 4250 31184 4306 31240
rect 4158 29144 4214 29200
rect 4250 29008 4306 29064
rect 4066 27648 4122 27704
rect 4158 27512 4214 27568
rect 4158 23976 4214 24032
rect 4526 31728 4582 31784
rect 4434 26696 4490 26752
rect 4434 26288 4490 26344
rect 4802 31864 4858 31920
rect 4986 37204 4988 37224
rect 4988 37204 5040 37224
rect 5040 37204 5042 37224
rect 4986 37168 5042 37204
rect 5170 34584 5226 34640
rect 4986 31592 5042 31648
rect 4802 30232 4858 30288
rect 4710 29588 4712 29608
rect 4712 29588 4764 29608
rect 4764 29588 4766 29608
rect 4710 29552 4766 29588
rect 4710 29416 4766 29472
rect 4342 26016 4398 26072
rect 4434 24112 4490 24168
rect 4066 22208 4122 22264
rect 3974 21800 4030 21856
rect 4894 29960 4950 30016
rect 4802 28328 4858 28384
rect 5262 31456 5318 31512
rect 4894 26444 4950 26480
rect 4894 26424 4896 26444
rect 4896 26424 4948 26444
rect 4948 26424 4950 26444
rect 5630 33224 5686 33280
rect 5446 31728 5502 31784
rect 5446 29552 5502 29608
rect 5538 29144 5594 29200
rect 5538 27920 5594 27976
rect 4066 21664 4122 21720
rect 4342 22752 4398 22808
rect 4066 21392 4122 21448
rect 4250 21392 4306 21448
rect 3790 20712 3846 20768
rect 3974 20712 4030 20768
rect 3514 17856 3570 17912
rect 3698 18672 3754 18728
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 3176 17434 3232 17436
rect 3256 17434 3312 17436
rect 3016 17382 3062 17434
rect 3062 17382 3072 17434
rect 3096 17382 3126 17434
rect 3126 17382 3138 17434
rect 3138 17382 3152 17434
rect 3176 17382 3190 17434
rect 3190 17382 3202 17434
rect 3202 17382 3232 17434
rect 3256 17382 3266 17434
rect 3266 17382 3312 17434
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 3176 17380 3232 17382
rect 3256 17380 3312 17382
rect 3238 17060 3294 17096
rect 3238 17040 3240 17060
rect 3240 17040 3292 17060
rect 3292 17040 3294 17060
rect 2962 16904 3018 16960
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 3176 16346 3232 16348
rect 3256 16346 3312 16348
rect 3016 16294 3062 16346
rect 3062 16294 3072 16346
rect 3096 16294 3126 16346
rect 3126 16294 3138 16346
rect 3138 16294 3152 16346
rect 3176 16294 3190 16346
rect 3190 16294 3202 16346
rect 3202 16294 3232 16346
rect 3256 16294 3266 16346
rect 3266 16294 3312 16346
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 3176 16292 3232 16294
rect 3256 16292 3312 16294
rect 3330 15816 3386 15872
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 3176 15258 3232 15260
rect 3256 15258 3312 15260
rect 3016 15206 3062 15258
rect 3062 15206 3072 15258
rect 3096 15206 3126 15258
rect 3126 15206 3138 15258
rect 3138 15206 3152 15258
rect 3176 15206 3190 15258
rect 3190 15206 3202 15258
rect 3202 15206 3232 15258
rect 3256 15206 3266 15258
rect 3266 15206 3312 15258
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 3176 15204 3232 15206
rect 3256 15204 3312 15206
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 3176 14170 3232 14172
rect 3256 14170 3312 14172
rect 3016 14118 3062 14170
rect 3062 14118 3072 14170
rect 3096 14118 3126 14170
rect 3126 14118 3138 14170
rect 3138 14118 3152 14170
rect 3176 14118 3190 14170
rect 3190 14118 3202 14170
rect 3202 14118 3232 14170
rect 3256 14118 3266 14170
rect 3266 14118 3312 14170
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 3176 14116 3232 14118
rect 3256 14116 3312 14118
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 3176 13082 3232 13084
rect 3256 13082 3312 13084
rect 3016 13030 3062 13082
rect 3062 13030 3072 13082
rect 3096 13030 3126 13082
rect 3126 13030 3138 13082
rect 3138 13030 3152 13082
rect 3176 13030 3190 13082
rect 3190 13030 3202 13082
rect 3202 13030 3232 13082
rect 3256 13030 3266 13082
rect 3266 13030 3312 13082
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 3176 13028 3232 13030
rect 3256 13028 3312 13030
rect 2962 12724 2964 12744
rect 2964 12724 3016 12744
rect 3016 12724 3018 12744
rect 2962 12688 3018 12724
rect 3054 12144 3110 12200
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 3176 11994 3232 11996
rect 3256 11994 3312 11996
rect 3016 11942 3062 11994
rect 3062 11942 3072 11994
rect 3096 11942 3126 11994
rect 3126 11942 3138 11994
rect 3138 11942 3152 11994
rect 3176 11942 3190 11994
rect 3190 11942 3202 11994
rect 3202 11942 3232 11994
rect 3256 11942 3266 11994
rect 3266 11942 3312 11994
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 3176 11940 3232 11942
rect 3256 11940 3312 11942
rect 3054 11736 3110 11792
rect 3054 11192 3110 11248
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 3176 10906 3232 10908
rect 3256 10906 3312 10908
rect 3016 10854 3062 10906
rect 3062 10854 3072 10906
rect 3096 10854 3126 10906
rect 3126 10854 3138 10906
rect 3138 10854 3152 10906
rect 3176 10854 3190 10906
rect 3190 10854 3202 10906
rect 3202 10854 3232 10906
rect 3256 10854 3266 10906
rect 3266 10854 3312 10906
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 3176 10852 3232 10854
rect 3256 10852 3312 10854
rect 2778 7792 2834 7848
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1858 5752 1914 5808
rect 1490 4972 1492 4992
rect 1492 4972 1544 4992
rect 1544 4972 1546 4992
rect 1490 4936 1546 4972
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1490 4120 1546 4176
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 3176 9818 3232 9820
rect 3256 9818 3312 9820
rect 3016 9766 3062 9818
rect 3062 9766 3072 9818
rect 3096 9766 3126 9818
rect 3126 9766 3138 9818
rect 3138 9766 3152 9818
rect 3176 9766 3190 9818
rect 3190 9766 3202 9818
rect 3202 9766 3232 9818
rect 3256 9766 3266 9818
rect 3266 9766 3312 9818
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 3176 9764 3232 9766
rect 3256 9764 3312 9766
rect 3514 17040 3570 17096
rect 3606 16224 3662 16280
rect 3882 19624 3938 19680
rect 3882 18844 3884 18864
rect 3884 18844 3936 18864
rect 3936 18844 3938 18864
rect 3882 18808 3938 18844
rect 3882 18536 3938 18592
rect 3790 14728 3846 14784
rect 3974 17992 4030 18048
rect 4526 23296 4582 23352
rect 4894 21936 4950 21992
rect 4802 21800 4858 21856
rect 4710 21256 4766 21312
rect 4250 15680 4306 15736
rect 4158 15136 4214 15192
rect 4158 14320 4214 14376
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3698 9696 3754 9752
rect 4066 12688 4122 12744
rect 4802 20884 4804 20904
rect 4804 20884 4856 20904
rect 4856 20884 4858 20904
rect 4802 20848 4858 20884
rect 4986 21664 5042 21720
rect 5262 26424 5318 26480
rect 5262 25064 5318 25120
rect 5078 21140 5134 21176
rect 5078 21120 5080 21140
rect 5080 21120 5132 21140
rect 5132 21120 5134 21140
rect 7010 40976 7066 41032
rect 5998 32952 6054 33008
rect 5998 31764 6000 31784
rect 6000 31764 6052 31784
rect 6052 31764 6054 31784
rect 5998 31728 6054 31764
rect 6458 37168 6514 37224
rect 6366 35536 6422 35592
rect 6274 35128 6330 35184
rect 6826 34448 6882 34504
rect 6826 34176 6882 34232
rect 5630 26560 5686 26616
rect 6090 30368 6146 30424
rect 6182 29280 6238 29336
rect 6274 27376 6330 27432
rect 6090 26560 6146 26616
rect 5630 26152 5686 26208
rect 5538 25336 5594 25392
rect 5170 18844 5172 18864
rect 5172 18844 5224 18864
rect 5224 18844 5226 18864
rect 5170 18808 5226 18844
rect 5078 17060 5134 17096
rect 5078 17040 5080 17060
rect 5080 17040 5132 17060
rect 5132 17040 5134 17060
rect 4894 16632 4950 16688
rect 4526 11872 4582 11928
rect 4250 11328 4306 11384
rect 4986 15852 4988 15872
rect 4988 15852 5040 15872
rect 5040 15852 5042 15872
rect 4986 15816 5042 15852
rect 4986 13640 5042 13696
rect 4802 9832 4858 9888
rect 4618 9424 4674 9480
rect 4894 9424 4950 9480
rect 5078 9288 5134 9344
rect 4618 7384 4674 7440
rect 5814 26288 5870 26344
rect 6182 26152 6238 26208
rect 5906 24928 5962 24984
rect 6274 25336 6330 25392
rect 5906 23840 5962 23896
rect 5998 23024 6054 23080
rect 5446 21684 5502 21720
rect 5446 21664 5448 21684
rect 5448 21664 5500 21684
rect 5500 21664 5502 21684
rect 5354 18672 5410 18728
rect 5538 17856 5594 17912
rect 5446 16904 5502 16960
rect 5538 15952 5594 16008
rect 5354 15000 5410 15056
rect 5446 12416 5502 12472
rect 5814 21800 5870 21856
rect 5814 21392 5870 21448
rect 5906 18964 5962 19000
rect 5906 18944 5908 18964
rect 5908 18944 5960 18964
rect 5960 18944 5962 18964
rect 5722 15680 5778 15736
rect 6458 28872 6514 28928
rect 6550 28600 6606 28656
rect 6274 23024 6330 23080
rect 6274 22752 6330 22808
rect 6366 20576 6422 20632
rect 6366 19760 6422 19816
rect 6366 18808 6422 18864
rect 6274 17876 6330 17912
rect 6274 17856 6276 17876
rect 6276 17856 6328 17876
rect 6328 17856 6330 17876
rect 6734 32852 6736 32872
rect 6736 32852 6788 32872
rect 6788 32852 6790 32872
rect 6734 32816 6790 32852
rect 7102 32272 7158 32328
rect 7010 32000 7066 32056
rect 9016 42458 9072 42460
rect 9096 42458 9152 42460
rect 9176 42458 9232 42460
rect 9256 42458 9312 42460
rect 9016 42406 9062 42458
rect 9062 42406 9072 42458
rect 9096 42406 9126 42458
rect 9126 42406 9138 42458
rect 9138 42406 9152 42458
rect 9176 42406 9190 42458
rect 9190 42406 9202 42458
rect 9202 42406 9232 42458
rect 9256 42406 9266 42458
rect 9266 42406 9312 42458
rect 9016 42404 9072 42406
rect 9096 42404 9152 42406
rect 9176 42404 9232 42406
rect 9256 42404 9312 42406
rect 7956 41914 8012 41916
rect 8036 41914 8092 41916
rect 8116 41914 8172 41916
rect 8196 41914 8252 41916
rect 7956 41862 8002 41914
rect 8002 41862 8012 41914
rect 8036 41862 8066 41914
rect 8066 41862 8078 41914
rect 8078 41862 8092 41914
rect 8116 41862 8130 41914
rect 8130 41862 8142 41914
rect 8142 41862 8172 41914
rect 8196 41862 8206 41914
rect 8206 41862 8252 41914
rect 7956 41860 8012 41862
rect 8036 41860 8092 41862
rect 8116 41860 8172 41862
rect 8196 41860 8252 41862
rect 7378 39480 7434 39536
rect 7956 40826 8012 40828
rect 8036 40826 8092 40828
rect 8116 40826 8172 40828
rect 8196 40826 8252 40828
rect 7956 40774 8002 40826
rect 8002 40774 8012 40826
rect 8036 40774 8066 40826
rect 8066 40774 8078 40826
rect 8078 40774 8092 40826
rect 8116 40774 8130 40826
rect 8130 40774 8142 40826
rect 8142 40774 8172 40826
rect 8196 40774 8206 40826
rect 8206 40774 8252 40826
rect 7956 40772 8012 40774
rect 8036 40772 8092 40774
rect 8116 40772 8172 40774
rect 8196 40772 8252 40774
rect 7746 40332 7748 40352
rect 7748 40332 7800 40352
rect 7800 40332 7802 40352
rect 7746 40296 7802 40332
rect 7956 39738 8012 39740
rect 8036 39738 8092 39740
rect 8116 39738 8172 39740
rect 8196 39738 8252 39740
rect 7956 39686 8002 39738
rect 8002 39686 8012 39738
rect 8036 39686 8066 39738
rect 8066 39686 8078 39738
rect 8078 39686 8092 39738
rect 8116 39686 8130 39738
rect 8130 39686 8142 39738
rect 8142 39686 8172 39738
rect 8196 39686 8206 39738
rect 8206 39686 8252 39738
rect 7956 39684 8012 39686
rect 8036 39684 8092 39686
rect 8116 39684 8172 39686
rect 8196 39684 8252 39686
rect 7956 38650 8012 38652
rect 8036 38650 8092 38652
rect 8116 38650 8172 38652
rect 8196 38650 8252 38652
rect 7956 38598 8002 38650
rect 8002 38598 8012 38650
rect 8036 38598 8066 38650
rect 8066 38598 8078 38650
rect 8078 38598 8092 38650
rect 8116 38598 8130 38650
rect 8130 38598 8142 38650
rect 8142 38598 8172 38650
rect 8196 38598 8206 38650
rect 8206 38598 8252 38650
rect 7956 38596 8012 38598
rect 8036 38596 8092 38598
rect 8116 38596 8172 38598
rect 8196 38596 8252 38598
rect 7286 34312 7342 34368
rect 7194 31728 7250 31784
rect 7194 30232 7250 30288
rect 7194 28600 7250 28656
rect 7102 28328 7158 28384
rect 6918 27512 6974 27568
rect 6918 24112 6974 24168
rect 6734 22636 6790 22672
rect 6734 22616 6736 22636
rect 6736 22616 6788 22636
rect 6788 22616 6790 22636
rect 7102 25880 7158 25936
rect 7102 24928 7158 24984
rect 7562 37168 7618 37224
rect 7956 37562 8012 37564
rect 8036 37562 8092 37564
rect 8116 37562 8172 37564
rect 8196 37562 8252 37564
rect 7956 37510 8002 37562
rect 8002 37510 8012 37562
rect 8036 37510 8066 37562
rect 8066 37510 8078 37562
rect 8078 37510 8092 37562
rect 8116 37510 8130 37562
rect 8130 37510 8142 37562
rect 8142 37510 8172 37562
rect 8196 37510 8206 37562
rect 8206 37510 8252 37562
rect 7956 37508 8012 37510
rect 8036 37508 8092 37510
rect 8116 37508 8172 37510
rect 8196 37508 8252 37510
rect 7562 36624 7618 36680
rect 8114 36660 8116 36680
rect 8116 36660 8168 36680
rect 8168 36660 8170 36680
rect 8114 36624 8170 36660
rect 7956 36474 8012 36476
rect 8036 36474 8092 36476
rect 8116 36474 8172 36476
rect 8196 36474 8252 36476
rect 7956 36422 8002 36474
rect 8002 36422 8012 36474
rect 8036 36422 8066 36474
rect 8066 36422 8078 36474
rect 8078 36422 8092 36474
rect 8116 36422 8130 36474
rect 8130 36422 8142 36474
rect 8142 36422 8172 36474
rect 8196 36422 8206 36474
rect 8206 36422 8252 36474
rect 7956 36420 8012 36422
rect 8036 36420 8092 36422
rect 8116 36420 8172 36422
rect 8196 36420 8252 36422
rect 8482 37712 8538 37768
rect 7378 32000 7434 32056
rect 9016 41370 9072 41372
rect 9096 41370 9152 41372
rect 9176 41370 9232 41372
rect 9256 41370 9312 41372
rect 9016 41318 9062 41370
rect 9062 41318 9072 41370
rect 9096 41318 9126 41370
rect 9126 41318 9138 41370
rect 9138 41318 9152 41370
rect 9176 41318 9190 41370
rect 9190 41318 9202 41370
rect 9202 41318 9232 41370
rect 9256 41318 9266 41370
rect 9266 41318 9312 41370
rect 9016 41316 9072 41318
rect 9096 41316 9152 41318
rect 9176 41316 9232 41318
rect 9256 41316 9312 41318
rect 9586 41556 9588 41576
rect 9588 41556 9640 41576
rect 9640 41556 9642 41576
rect 9586 41520 9642 41556
rect 9016 40282 9072 40284
rect 9096 40282 9152 40284
rect 9176 40282 9232 40284
rect 9256 40282 9312 40284
rect 9016 40230 9062 40282
rect 9062 40230 9072 40282
rect 9096 40230 9126 40282
rect 9126 40230 9138 40282
rect 9138 40230 9152 40282
rect 9176 40230 9190 40282
rect 9190 40230 9202 40282
rect 9202 40230 9232 40282
rect 9256 40230 9266 40282
rect 9266 40230 9312 40282
rect 9016 40228 9072 40230
rect 9096 40228 9152 40230
rect 9176 40228 9232 40230
rect 9256 40228 9312 40230
rect 9402 40160 9458 40216
rect 9218 40060 9220 40080
rect 9220 40060 9272 40080
rect 9272 40060 9274 40080
rect 9218 40024 9274 40060
rect 8666 39616 8722 39672
rect 9494 39380 9496 39400
rect 9496 39380 9548 39400
rect 9548 39380 9550 39400
rect 9494 39344 9550 39380
rect 9016 39194 9072 39196
rect 9096 39194 9152 39196
rect 9176 39194 9232 39196
rect 9256 39194 9312 39196
rect 9016 39142 9062 39194
rect 9062 39142 9072 39194
rect 9096 39142 9126 39194
rect 9126 39142 9138 39194
rect 9138 39142 9152 39194
rect 9176 39142 9190 39194
rect 9190 39142 9202 39194
rect 9202 39142 9232 39194
rect 9256 39142 9266 39194
rect 9266 39142 9312 39194
rect 9016 39140 9072 39142
rect 9096 39140 9152 39142
rect 9176 39140 9232 39142
rect 9256 39140 9312 39142
rect 8758 38800 8814 38856
rect 8758 37304 8814 37360
rect 8574 35808 8630 35864
rect 7956 35386 8012 35388
rect 8036 35386 8092 35388
rect 8116 35386 8172 35388
rect 8196 35386 8252 35388
rect 7956 35334 8002 35386
rect 8002 35334 8012 35386
rect 8036 35334 8066 35386
rect 8066 35334 8078 35386
rect 8078 35334 8092 35386
rect 8116 35334 8130 35386
rect 8130 35334 8142 35386
rect 8142 35334 8172 35386
rect 8196 35334 8206 35386
rect 8206 35334 8252 35386
rect 7956 35332 8012 35334
rect 8036 35332 8092 35334
rect 8116 35332 8172 35334
rect 8196 35332 8252 35334
rect 7956 34298 8012 34300
rect 8036 34298 8092 34300
rect 8116 34298 8172 34300
rect 8196 34298 8252 34300
rect 7956 34246 8002 34298
rect 8002 34246 8012 34298
rect 8036 34246 8066 34298
rect 8066 34246 8078 34298
rect 8078 34246 8092 34298
rect 8116 34246 8130 34298
rect 8130 34246 8142 34298
rect 8142 34246 8172 34298
rect 8196 34246 8206 34298
rect 8206 34246 8252 34298
rect 7956 34244 8012 34246
rect 8036 34244 8092 34246
rect 8116 34244 8172 34246
rect 8196 34244 8252 34246
rect 7956 33210 8012 33212
rect 8036 33210 8092 33212
rect 8116 33210 8172 33212
rect 8196 33210 8252 33212
rect 7956 33158 8002 33210
rect 8002 33158 8012 33210
rect 8036 33158 8066 33210
rect 8066 33158 8078 33210
rect 8078 33158 8092 33210
rect 8116 33158 8130 33210
rect 8130 33158 8142 33210
rect 8142 33158 8172 33210
rect 8196 33158 8206 33210
rect 8206 33158 8252 33210
rect 7956 33156 8012 33158
rect 8036 33156 8092 33158
rect 8116 33156 8172 33158
rect 8196 33156 8252 33158
rect 7838 32952 7894 33008
rect 7010 23024 7066 23080
rect 7010 22772 7066 22808
rect 7010 22752 7012 22772
rect 7012 22752 7064 22772
rect 7064 22752 7066 22772
rect 7010 22480 7066 22536
rect 6918 22208 6974 22264
rect 6642 21256 6698 21312
rect 6642 19896 6698 19952
rect 6918 21936 6974 21992
rect 7194 24692 7196 24712
rect 7196 24692 7248 24712
rect 7248 24692 7250 24712
rect 7194 24656 7250 24692
rect 7286 24248 7342 24304
rect 7286 22888 7342 22944
rect 7194 22208 7250 22264
rect 7102 21936 7158 21992
rect 7102 21800 7158 21856
rect 7194 21256 7250 21312
rect 7194 20304 7250 20360
rect 6090 16496 6146 16552
rect 5998 15816 6054 15872
rect 5998 15408 6054 15464
rect 6274 16088 6330 16144
rect 5814 12688 5870 12744
rect 6274 13232 6330 13288
rect 5262 11892 5318 11928
rect 5262 11872 5264 11892
rect 5264 11872 5316 11892
rect 5316 11872 5318 11892
rect 5354 9560 5410 9616
rect 5630 7384 5686 7440
rect 5722 7112 5778 7168
rect 5722 5888 5778 5944
rect 5538 5752 5594 5808
rect 6274 12144 6330 12200
rect 5998 11600 6054 11656
rect 8574 35536 8630 35592
rect 7956 32122 8012 32124
rect 8036 32122 8092 32124
rect 8116 32122 8172 32124
rect 8196 32122 8252 32124
rect 7956 32070 8002 32122
rect 8002 32070 8012 32122
rect 8036 32070 8066 32122
rect 8066 32070 8078 32122
rect 8078 32070 8092 32122
rect 8116 32070 8130 32122
rect 8130 32070 8142 32122
rect 8142 32070 8172 32122
rect 8196 32070 8206 32122
rect 8206 32070 8252 32122
rect 7956 32068 8012 32070
rect 8036 32068 8092 32070
rect 8116 32068 8172 32070
rect 8196 32068 8252 32070
rect 8390 31320 8446 31376
rect 7956 31034 8012 31036
rect 8036 31034 8092 31036
rect 8116 31034 8172 31036
rect 8196 31034 8252 31036
rect 7956 30982 8002 31034
rect 8002 30982 8012 31034
rect 8036 30982 8066 31034
rect 8066 30982 8078 31034
rect 8078 30982 8092 31034
rect 8116 30982 8130 31034
rect 8130 30982 8142 31034
rect 8142 30982 8172 31034
rect 8196 30982 8206 31034
rect 8206 30982 8252 31034
rect 7956 30980 8012 30982
rect 8036 30980 8092 30982
rect 8116 30980 8172 30982
rect 8196 30980 8252 30982
rect 9126 38664 9182 38720
rect 9126 38292 9128 38312
rect 9128 38292 9180 38312
rect 9180 38292 9182 38312
rect 9126 38256 9182 38292
rect 9016 38106 9072 38108
rect 9096 38106 9152 38108
rect 9176 38106 9232 38108
rect 9256 38106 9312 38108
rect 9016 38054 9062 38106
rect 9062 38054 9072 38106
rect 9096 38054 9126 38106
rect 9126 38054 9138 38106
rect 9138 38054 9152 38106
rect 9176 38054 9190 38106
rect 9190 38054 9202 38106
rect 9202 38054 9232 38106
rect 9256 38054 9266 38106
rect 9266 38054 9312 38106
rect 9016 38052 9072 38054
rect 9096 38052 9152 38054
rect 9176 38052 9232 38054
rect 9256 38052 9312 38054
rect 9016 37018 9072 37020
rect 9096 37018 9152 37020
rect 9176 37018 9232 37020
rect 9256 37018 9312 37020
rect 9016 36966 9062 37018
rect 9062 36966 9072 37018
rect 9096 36966 9126 37018
rect 9126 36966 9138 37018
rect 9138 36966 9152 37018
rect 9176 36966 9190 37018
rect 9190 36966 9202 37018
rect 9202 36966 9232 37018
rect 9256 36966 9266 37018
rect 9266 36966 9312 37018
rect 9016 36964 9072 36966
rect 9096 36964 9152 36966
rect 9176 36964 9232 36966
rect 9256 36964 9312 36966
rect 9126 36080 9182 36136
rect 9016 35930 9072 35932
rect 9096 35930 9152 35932
rect 9176 35930 9232 35932
rect 9256 35930 9312 35932
rect 9016 35878 9062 35930
rect 9062 35878 9072 35930
rect 9096 35878 9126 35930
rect 9126 35878 9138 35930
rect 9138 35878 9152 35930
rect 9176 35878 9190 35930
rect 9190 35878 9202 35930
rect 9202 35878 9232 35930
rect 9256 35878 9266 35930
rect 9266 35878 9312 35930
rect 9016 35876 9072 35878
rect 9096 35876 9152 35878
rect 9176 35876 9232 35878
rect 9256 35876 9312 35878
rect 9770 40332 9772 40352
rect 9772 40332 9824 40352
rect 9824 40332 9826 40352
rect 9770 40296 9826 40332
rect 10414 39752 10470 39808
rect 9678 39208 9734 39264
rect 10598 39480 10654 39536
rect 10230 38936 10286 38992
rect 9954 37304 10010 37360
rect 10138 38392 10194 38448
rect 8758 35536 8814 35592
rect 8942 35028 8944 35048
rect 8944 35028 8996 35048
rect 8996 35028 8998 35048
rect 8942 34992 8998 35028
rect 9016 34842 9072 34844
rect 9096 34842 9152 34844
rect 9176 34842 9232 34844
rect 9256 34842 9312 34844
rect 9016 34790 9062 34842
rect 9062 34790 9072 34842
rect 9096 34790 9126 34842
rect 9126 34790 9138 34842
rect 9138 34790 9152 34842
rect 9176 34790 9190 34842
rect 9190 34790 9202 34842
rect 9202 34790 9232 34842
rect 9256 34790 9266 34842
rect 9266 34790 9312 34842
rect 9016 34788 9072 34790
rect 9096 34788 9152 34790
rect 9176 34788 9232 34790
rect 9256 34788 9312 34790
rect 10046 37032 10102 37088
rect 10414 38120 10470 38176
rect 10322 37848 10378 37904
rect 10230 37576 10286 37632
rect 10138 36488 10194 36544
rect 9678 35128 9734 35184
rect 9954 34856 10010 34912
rect 9586 34584 9642 34640
rect 9126 33940 9128 33960
rect 9128 33940 9180 33960
rect 9180 33940 9182 33960
rect 9126 33904 9182 33940
rect 9016 33754 9072 33756
rect 9096 33754 9152 33756
rect 9176 33754 9232 33756
rect 9256 33754 9312 33756
rect 9016 33702 9062 33754
rect 9062 33702 9072 33754
rect 9096 33702 9126 33754
rect 9126 33702 9138 33754
rect 9138 33702 9152 33754
rect 9176 33702 9190 33754
rect 9190 33702 9202 33754
rect 9202 33702 9232 33754
rect 9256 33702 9266 33754
rect 9266 33702 9312 33754
rect 9016 33700 9072 33702
rect 9096 33700 9152 33702
rect 9176 33700 9232 33702
rect 9256 33700 9312 33702
rect 8850 32716 8852 32736
rect 8852 32716 8904 32736
rect 8904 32716 8906 32736
rect 8850 32680 8906 32716
rect 9016 32666 9072 32668
rect 9096 32666 9152 32668
rect 9176 32666 9232 32668
rect 9256 32666 9312 32668
rect 9016 32614 9062 32666
rect 9062 32614 9072 32666
rect 9096 32614 9126 32666
rect 9126 32614 9138 32666
rect 9138 32614 9152 32666
rect 9176 32614 9190 32666
rect 9190 32614 9202 32666
rect 9202 32614 9232 32666
rect 9256 32614 9266 32666
rect 9266 32614 9312 32666
rect 9016 32612 9072 32614
rect 9096 32612 9152 32614
rect 9176 32612 9232 32614
rect 9256 32612 9312 32614
rect 8574 31340 8630 31376
rect 8574 31320 8576 31340
rect 8576 31320 8628 31340
rect 8628 31320 8630 31340
rect 8666 31220 8668 31240
rect 8668 31220 8720 31240
rect 8720 31220 8722 31240
rect 8666 31184 8722 31220
rect 8666 30912 8722 30968
rect 7956 29946 8012 29948
rect 8036 29946 8092 29948
rect 8116 29946 8172 29948
rect 8196 29946 8252 29948
rect 7956 29894 8002 29946
rect 8002 29894 8012 29946
rect 8036 29894 8066 29946
rect 8066 29894 8078 29946
rect 8078 29894 8092 29946
rect 8116 29894 8130 29946
rect 8130 29894 8142 29946
rect 8142 29894 8172 29946
rect 8196 29894 8206 29946
rect 8206 29894 8252 29946
rect 7956 29892 8012 29894
rect 8036 29892 8092 29894
rect 8116 29892 8172 29894
rect 8196 29892 8252 29894
rect 9494 33380 9550 33416
rect 9494 33360 9496 33380
rect 9496 33360 9548 33380
rect 9548 33360 9550 33380
rect 9954 33768 10010 33824
rect 9678 32680 9734 32736
rect 9402 31728 9458 31784
rect 9016 31578 9072 31580
rect 9096 31578 9152 31580
rect 9176 31578 9232 31580
rect 9256 31578 9312 31580
rect 9016 31526 9062 31578
rect 9062 31526 9072 31578
rect 9096 31526 9126 31578
rect 9126 31526 9138 31578
rect 9138 31526 9152 31578
rect 9176 31526 9190 31578
rect 9190 31526 9202 31578
rect 9202 31526 9232 31578
rect 9256 31526 9266 31578
rect 9266 31526 9312 31578
rect 9016 31524 9072 31526
rect 9096 31524 9152 31526
rect 9176 31524 9232 31526
rect 9256 31524 9312 31526
rect 9034 31320 9090 31376
rect 8758 30368 8814 30424
rect 7470 22072 7526 22128
rect 8022 29724 8024 29744
rect 8024 29724 8076 29744
rect 8076 29724 8078 29744
rect 8022 29688 8078 29724
rect 8114 29280 8170 29336
rect 7956 28858 8012 28860
rect 8036 28858 8092 28860
rect 8116 28858 8172 28860
rect 8196 28858 8252 28860
rect 7956 28806 8002 28858
rect 8002 28806 8012 28858
rect 8036 28806 8066 28858
rect 8066 28806 8078 28858
rect 8078 28806 8092 28858
rect 8116 28806 8130 28858
rect 8130 28806 8142 28858
rect 8142 28806 8172 28858
rect 8196 28806 8206 28858
rect 8206 28806 8252 28858
rect 7956 28804 8012 28806
rect 8036 28804 8092 28806
rect 8116 28804 8172 28806
rect 8196 28804 8252 28806
rect 8114 28212 8170 28248
rect 8114 28192 8116 28212
rect 8116 28192 8168 28212
rect 8168 28192 8170 28212
rect 7956 27770 8012 27772
rect 8036 27770 8092 27772
rect 8116 27770 8172 27772
rect 8196 27770 8252 27772
rect 7956 27718 8002 27770
rect 8002 27718 8012 27770
rect 8036 27718 8066 27770
rect 8066 27718 8078 27770
rect 8078 27718 8092 27770
rect 8116 27718 8130 27770
rect 8130 27718 8142 27770
rect 8142 27718 8172 27770
rect 8196 27718 8206 27770
rect 8206 27718 8252 27770
rect 7956 27716 8012 27718
rect 8036 27716 8092 27718
rect 8116 27716 8172 27718
rect 8196 27716 8252 27718
rect 7956 26682 8012 26684
rect 8036 26682 8092 26684
rect 8116 26682 8172 26684
rect 8196 26682 8252 26684
rect 7956 26630 8002 26682
rect 8002 26630 8012 26682
rect 8036 26630 8066 26682
rect 8066 26630 8078 26682
rect 8078 26630 8092 26682
rect 8116 26630 8130 26682
rect 8130 26630 8142 26682
rect 8142 26630 8172 26682
rect 8196 26630 8206 26682
rect 8206 26630 8252 26682
rect 7956 26628 8012 26630
rect 8036 26628 8092 26630
rect 8116 26628 8172 26630
rect 8196 26628 8252 26630
rect 8390 26832 8446 26888
rect 8666 29552 8722 29608
rect 8666 29008 8722 29064
rect 8482 26560 8538 26616
rect 8206 26152 8262 26208
rect 7930 25744 7986 25800
rect 7956 25594 8012 25596
rect 8036 25594 8092 25596
rect 8116 25594 8172 25596
rect 8196 25594 8252 25596
rect 7956 25542 8002 25594
rect 8002 25542 8012 25594
rect 8036 25542 8066 25594
rect 8066 25542 8078 25594
rect 8078 25542 8092 25594
rect 8116 25542 8130 25594
rect 8130 25542 8142 25594
rect 8142 25542 8172 25594
rect 8196 25542 8206 25594
rect 8206 25542 8252 25594
rect 7956 25540 8012 25542
rect 8036 25540 8092 25542
rect 8116 25540 8172 25542
rect 8196 25540 8252 25542
rect 8022 25336 8078 25392
rect 8206 24812 8262 24848
rect 8206 24792 8208 24812
rect 8208 24792 8260 24812
rect 8260 24792 8262 24812
rect 7956 24506 8012 24508
rect 8036 24506 8092 24508
rect 8116 24506 8172 24508
rect 8196 24506 8252 24508
rect 7956 24454 8002 24506
rect 8002 24454 8012 24506
rect 8036 24454 8066 24506
rect 8066 24454 8078 24506
rect 8078 24454 8092 24506
rect 8116 24454 8130 24506
rect 8130 24454 8142 24506
rect 8142 24454 8172 24506
rect 8196 24454 8206 24506
rect 8206 24454 8252 24506
rect 7956 24452 8012 24454
rect 8036 24452 8092 24454
rect 8116 24452 8172 24454
rect 8196 24452 8252 24454
rect 7930 23704 7986 23760
rect 8758 27548 8760 27568
rect 8760 27548 8812 27568
rect 8812 27548 8814 27568
rect 8758 27512 8814 27548
rect 8666 26560 8722 26616
rect 8298 23840 8354 23896
rect 8022 23568 8078 23624
rect 8206 23568 8262 23624
rect 7746 21664 7802 21720
rect 7654 21120 7710 21176
rect 7562 19624 7618 19680
rect 6734 14456 6790 14512
rect 6734 12164 6790 12200
rect 6734 12144 6736 12164
rect 6736 12144 6788 12164
rect 6788 12144 6790 12164
rect 7378 15700 7434 15736
rect 7378 15680 7380 15700
rect 7380 15680 7432 15700
rect 7432 15680 7434 15700
rect 6090 9444 6146 9480
rect 6090 9424 6092 9444
rect 6092 9424 6144 9444
rect 6144 9424 6146 9444
rect 5998 7112 6054 7168
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 3698 1264 3754 1320
rect 5078 1264 5134 1320
rect 4618 1128 4674 1184
rect 6274 9324 6276 9344
rect 6276 9324 6328 9344
rect 6328 9324 6330 9344
rect 6274 9288 6330 9324
rect 6274 8608 6330 8664
rect 6826 10512 6882 10568
rect 6734 9424 6790 9480
rect 7010 10104 7066 10160
rect 6826 8336 6882 8392
rect 6918 7540 6974 7576
rect 6918 7520 6920 7540
rect 6920 7520 6972 7540
rect 6972 7520 6974 7540
rect 7378 12708 7434 12744
rect 7378 12688 7380 12708
rect 7380 12688 7432 12708
rect 7432 12688 7434 12708
rect 7956 23418 8012 23420
rect 8036 23418 8092 23420
rect 8116 23418 8172 23420
rect 8196 23418 8252 23420
rect 7956 23366 8002 23418
rect 8002 23366 8012 23418
rect 8036 23366 8066 23418
rect 8066 23366 8078 23418
rect 8078 23366 8092 23418
rect 8116 23366 8130 23418
rect 8130 23366 8142 23418
rect 8142 23366 8172 23418
rect 8196 23366 8206 23418
rect 8206 23366 8252 23418
rect 7956 23364 8012 23366
rect 8036 23364 8092 23366
rect 8116 23364 8172 23366
rect 8196 23364 8252 23366
rect 8022 23160 8078 23216
rect 8022 22480 8078 22536
rect 7956 22330 8012 22332
rect 8036 22330 8092 22332
rect 8116 22330 8172 22332
rect 8196 22330 8252 22332
rect 7956 22278 8002 22330
rect 8002 22278 8012 22330
rect 8036 22278 8066 22330
rect 8066 22278 8078 22330
rect 8078 22278 8092 22330
rect 8116 22278 8130 22330
rect 8130 22278 8142 22330
rect 8142 22278 8172 22330
rect 8196 22278 8206 22330
rect 8206 22278 8252 22330
rect 7956 22276 8012 22278
rect 8036 22276 8092 22278
rect 8116 22276 8172 22278
rect 8196 22276 8252 22278
rect 7930 21664 7986 21720
rect 7956 21242 8012 21244
rect 8036 21242 8092 21244
rect 8116 21242 8172 21244
rect 8196 21242 8252 21244
rect 7956 21190 8002 21242
rect 8002 21190 8012 21242
rect 8036 21190 8066 21242
rect 8066 21190 8078 21242
rect 8078 21190 8092 21242
rect 8116 21190 8130 21242
rect 8130 21190 8142 21242
rect 8142 21190 8172 21242
rect 8196 21190 8206 21242
rect 8206 21190 8252 21242
rect 7956 21188 8012 21190
rect 8036 21188 8092 21190
rect 8116 21188 8172 21190
rect 8196 21188 8252 21190
rect 7930 21004 7986 21040
rect 7930 20984 7932 21004
rect 7932 20984 7984 21004
rect 7984 20984 7986 21004
rect 7956 20154 8012 20156
rect 8036 20154 8092 20156
rect 8116 20154 8172 20156
rect 8196 20154 8252 20156
rect 7956 20102 8002 20154
rect 8002 20102 8012 20154
rect 8036 20102 8066 20154
rect 8066 20102 8078 20154
rect 8078 20102 8092 20154
rect 8116 20102 8130 20154
rect 8130 20102 8142 20154
rect 8142 20102 8172 20154
rect 8196 20102 8206 20154
rect 8206 20102 8252 20154
rect 7956 20100 8012 20102
rect 8036 20100 8092 20102
rect 8116 20100 8172 20102
rect 8196 20100 8252 20102
rect 7930 19252 7932 19272
rect 7932 19252 7984 19272
rect 7984 19252 7986 19272
rect 7930 19216 7986 19252
rect 7956 19066 8012 19068
rect 8036 19066 8092 19068
rect 8116 19066 8172 19068
rect 8196 19066 8252 19068
rect 7956 19014 8002 19066
rect 8002 19014 8012 19066
rect 8036 19014 8066 19066
rect 8066 19014 8078 19066
rect 8078 19014 8092 19066
rect 8116 19014 8130 19066
rect 8130 19014 8142 19066
rect 8142 19014 8172 19066
rect 8196 19014 8206 19066
rect 8206 19014 8252 19066
rect 7956 19012 8012 19014
rect 8036 19012 8092 19014
rect 8116 19012 8172 19014
rect 8196 19012 8252 19014
rect 7654 17720 7710 17776
rect 8114 18148 8170 18184
rect 8114 18128 8116 18148
rect 8116 18128 8168 18148
rect 8168 18128 8170 18148
rect 7956 17978 8012 17980
rect 8036 17978 8092 17980
rect 8116 17978 8172 17980
rect 8196 17978 8252 17980
rect 7956 17926 8002 17978
rect 8002 17926 8012 17978
rect 8036 17926 8066 17978
rect 8066 17926 8078 17978
rect 8078 17926 8092 17978
rect 8116 17926 8130 17978
rect 8130 17926 8142 17978
rect 8142 17926 8172 17978
rect 8196 17926 8206 17978
rect 8206 17926 8252 17978
rect 7956 17924 8012 17926
rect 8036 17924 8092 17926
rect 8116 17924 8172 17926
rect 8196 17924 8252 17926
rect 9016 30490 9072 30492
rect 9096 30490 9152 30492
rect 9176 30490 9232 30492
rect 9256 30490 9312 30492
rect 9016 30438 9062 30490
rect 9062 30438 9072 30490
rect 9096 30438 9126 30490
rect 9126 30438 9138 30490
rect 9138 30438 9152 30490
rect 9176 30438 9190 30490
rect 9190 30438 9202 30490
rect 9202 30438 9232 30490
rect 9256 30438 9266 30490
rect 9266 30438 9312 30490
rect 9016 30436 9072 30438
rect 9096 30436 9152 30438
rect 9176 30436 9232 30438
rect 9256 30436 9312 30438
rect 9034 29688 9090 29744
rect 9494 31048 9550 31104
rect 9678 31320 9734 31376
rect 9586 30776 9642 30832
rect 9494 29824 9550 29880
rect 9678 30504 9734 30560
rect 9586 29688 9642 29744
rect 9016 29402 9072 29404
rect 9096 29402 9152 29404
rect 9176 29402 9232 29404
rect 9256 29402 9312 29404
rect 9016 29350 9062 29402
rect 9062 29350 9072 29402
rect 9096 29350 9126 29402
rect 9126 29350 9138 29402
rect 9138 29350 9152 29402
rect 9176 29350 9190 29402
rect 9190 29350 9202 29402
rect 9202 29350 9232 29402
rect 9256 29350 9266 29402
rect 9266 29350 9312 29402
rect 9016 29348 9072 29350
rect 9096 29348 9152 29350
rect 9176 29348 9232 29350
rect 9256 29348 9312 29350
rect 8942 29008 8998 29064
rect 8942 28600 8998 28656
rect 9218 28464 9274 28520
rect 9016 28314 9072 28316
rect 9096 28314 9152 28316
rect 9176 28314 9232 28316
rect 9256 28314 9312 28316
rect 9016 28262 9062 28314
rect 9062 28262 9072 28314
rect 9096 28262 9126 28314
rect 9126 28262 9138 28314
rect 9138 28262 9152 28314
rect 9176 28262 9190 28314
rect 9190 28262 9202 28314
rect 9202 28262 9232 28314
rect 9256 28262 9266 28314
rect 9266 28262 9312 28314
rect 9016 28260 9072 28262
rect 9096 28260 9152 28262
rect 9176 28260 9232 28262
rect 9256 28260 9312 28262
rect 9586 29144 9642 29200
rect 9770 29416 9826 29472
rect 10782 38664 10838 38720
rect 10506 36760 10562 36816
rect 10322 35944 10378 36000
rect 10230 34312 10286 34368
rect 10138 33224 10194 33280
rect 10230 32408 10286 32464
rect 10230 32136 10286 32192
rect 10966 36216 11022 36272
rect 10598 35672 10654 35728
rect 10506 35400 10562 35456
rect 10414 34040 10470 34096
rect 10598 33496 10654 33552
rect 10690 32952 10746 33008
rect 10414 31864 10470 31920
rect 9954 30232 10010 30288
rect 9586 28328 9642 28384
rect 9494 28056 9550 28112
rect 9678 28056 9734 28112
rect 9402 27648 9458 27704
rect 9954 29144 10010 29200
rect 9126 27412 9128 27432
rect 9128 27412 9180 27432
rect 9180 27412 9182 27432
rect 9126 27376 9182 27412
rect 9016 27226 9072 27228
rect 9096 27226 9152 27228
rect 9176 27226 9232 27228
rect 9256 27226 9312 27228
rect 9016 27174 9062 27226
rect 9062 27174 9072 27226
rect 9096 27174 9126 27226
rect 9126 27174 9138 27226
rect 9138 27174 9152 27226
rect 9176 27174 9190 27226
rect 9190 27174 9202 27226
rect 9202 27174 9232 27226
rect 9256 27174 9266 27226
rect 9266 27174 9312 27226
rect 9016 27172 9072 27174
rect 9096 27172 9152 27174
rect 9176 27172 9232 27174
rect 9256 27172 9312 27174
rect 9310 26696 9366 26752
rect 9678 27240 9734 27296
rect 9016 26138 9072 26140
rect 9096 26138 9152 26140
rect 9176 26138 9232 26140
rect 9256 26138 9312 26140
rect 9016 26086 9062 26138
rect 9062 26086 9072 26138
rect 9096 26086 9126 26138
rect 9126 26086 9138 26138
rect 9138 26086 9152 26138
rect 9176 26086 9190 26138
rect 9190 26086 9202 26138
rect 9202 26086 9232 26138
rect 9256 26086 9266 26138
rect 9266 26086 9312 26138
rect 9016 26084 9072 26086
rect 9096 26084 9152 26086
rect 9176 26084 9232 26086
rect 9256 26084 9312 26086
rect 8850 25880 8906 25936
rect 9494 26324 9496 26344
rect 9496 26324 9548 26344
rect 9548 26324 9550 26344
rect 9494 26288 9550 26324
rect 9678 25880 9734 25936
rect 9016 25050 9072 25052
rect 9096 25050 9152 25052
rect 9176 25050 9232 25052
rect 9256 25050 9312 25052
rect 9016 24998 9062 25050
rect 9062 24998 9072 25050
rect 9096 24998 9126 25050
rect 9126 24998 9138 25050
rect 9138 24998 9152 25050
rect 9176 24998 9190 25050
rect 9190 24998 9202 25050
rect 9202 24998 9232 25050
rect 9256 24998 9266 25050
rect 9266 24998 9312 25050
rect 9016 24996 9072 24998
rect 9096 24996 9152 24998
rect 9176 24996 9232 24998
rect 9256 24996 9312 24998
rect 9310 24792 9366 24848
rect 9586 25336 9642 25392
rect 9678 25100 9680 25120
rect 9680 25100 9732 25120
rect 9732 25100 9734 25120
rect 9678 25064 9734 25100
rect 9126 24248 9182 24304
rect 9016 23962 9072 23964
rect 9096 23962 9152 23964
rect 9176 23962 9232 23964
rect 9256 23962 9312 23964
rect 9016 23910 9062 23962
rect 9062 23910 9072 23962
rect 9096 23910 9126 23962
rect 9126 23910 9138 23962
rect 9138 23910 9152 23962
rect 9176 23910 9190 23962
rect 9190 23910 9202 23962
rect 9202 23910 9232 23962
rect 9256 23910 9266 23962
rect 9266 23910 9312 23962
rect 9016 23908 9072 23910
rect 9096 23908 9152 23910
rect 9176 23908 9232 23910
rect 9256 23908 9312 23910
rect 8482 21800 8538 21856
rect 8482 20984 8538 21040
rect 8114 17060 8170 17096
rect 8114 17040 8116 17060
rect 8116 17040 8168 17060
rect 8168 17040 8170 17060
rect 7562 16108 7618 16144
rect 7562 16088 7564 16108
rect 7564 16088 7616 16108
rect 7616 16088 7618 16108
rect 7654 15544 7710 15600
rect 7956 16890 8012 16892
rect 8036 16890 8092 16892
rect 8116 16890 8172 16892
rect 8196 16890 8252 16892
rect 7956 16838 8002 16890
rect 8002 16838 8012 16890
rect 8036 16838 8066 16890
rect 8066 16838 8078 16890
rect 8078 16838 8092 16890
rect 8116 16838 8130 16890
rect 8130 16838 8142 16890
rect 8142 16838 8172 16890
rect 8196 16838 8206 16890
rect 8206 16838 8252 16890
rect 7956 16836 8012 16838
rect 8036 16836 8092 16838
rect 8116 16836 8172 16838
rect 8196 16836 8252 16838
rect 8022 16088 8078 16144
rect 7956 15802 8012 15804
rect 8036 15802 8092 15804
rect 8116 15802 8172 15804
rect 8196 15802 8252 15804
rect 7956 15750 8002 15802
rect 8002 15750 8012 15802
rect 8036 15750 8066 15802
rect 8066 15750 8078 15802
rect 8078 15750 8092 15802
rect 8116 15750 8130 15802
rect 8130 15750 8142 15802
rect 8142 15750 8172 15802
rect 8196 15750 8206 15802
rect 8206 15750 8252 15802
rect 7956 15748 8012 15750
rect 8036 15748 8092 15750
rect 8116 15748 8172 15750
rect 8196 15748 8252 15750
rect 7956 14714 8012 14716
rect 8036 14714 8092 14716
rect 8116 14714 8172 14716
rect 8196 14714 8252 14716
rect 7956 14662 8002 14714
rect 8002 14662 8012 14714
rect 8036 14662 8066 14714
rect 8066 14662 8078 14714
rect 8078 14662 8092 14714
rect 8116 14662 8130 14714
rect 8130 14662 8142 14714
rect 8142 14662 8172 14714
rect 8196 14662 8206 14714
rect 8206 14662 8252 14714
rect 7956 14660 8012 14662
rect 8036 14660 8092 14662
rect 8116 14660 8172 14662
rect 8196 14660 8252 14662
rect 8114 13776 8170 13832
rect 7746 13524 7802 13560
rect 7746 13504 7748 13524
rect 7748 13504 7800 13524
rect 7800 13504 7802 13524
rect 7956 13626 8012 13628
rect 8036 13626 8092 13628
rect 8116 13626 8172 13628
rect 8196 13626 8252 13628
rect 7956 13574 8002 13626
rect 8002 13574 8012 13626
rect 8036 13574 8066 13626
rect 8066 13574 8078 13626
rect 8078 13574 8092 13626
rect 8116 13574 8130 13626
rect 8130 13574 8142 13626
rect 8142 13574 8172 13626
rect 8196 13574 8206 13626
rect 8206 13574 8252 13626
rect 7956 13572 8012 13574
rect 8036 13572 8092 13574
rect 8116 13572 8172 13574
rect 8196 13572 8252 13574
rect 8390 15136 8446 15192
rect 8390 13504 8446 13560
rect 8298 12960 8354 13016
rect 7930 12824 7986 12880
rect 7838 12688 7894 12744
rect 8114 12724 8116 12744
rect 8116 12724 8168 12744
rect 8168 12724 8170 12744
rect 8114 12688 8170 12724
rect 7956 12538 8012 12540
rect 8036 12538 8092 12540
rect 8116 12538 8172 12540
rect 8196 12538 8252 12540
rect 7956 12486 8002 12538
rect 8002 12486 8012 12538
rect 8036 12486 8066 12538
rect 8066 12486 8078 12538
rect 8078 12486 8092 12538
rect 8116 12486 8130 12538
rect 8130 12486 8142 12538
rect 8142 12486 8172 12538
rect 8196 12486 8206 12538
rect 8206 12486 8252 12538
rect 7956 12484 8012 12486
rect 8036 12484 8092 12486
rect 8116 12484 8172 12486
rect 8196 12484 8252 12486
rect 7470 9424 7526 9480
rect 7378 8472 7434 8528
rect 7378 7928 7434 7984
rect 7286 7520 7342 7576
rect 7378 7404 7434 7440
rect 7378 7384 7380 7404
rect 7380 7384 7432 7404
rect 7432 7384 7434 7404
rect 6458 5888 6514 5944
rect 7838 11736 7894 11792
rect 8206 12316 8208 12336
rect 8208 12316 8260 12336
rect 8260 12316 8262 12336
rect 8206 12280 8262 12316
rect 7956 11450 8012 11452
rect 8036 11450 8092 11452
rect 8116 11450 8172 11452
rect 8196 11450 8252 11452
rect 7956 11398 8002 11450
rect 8002 11398 8012 11450
rect 8036 11398 8066 11450
rect 8066 11398 8078 11450
rect 8078 11398 8092 11450
rect 8116 11398 8130 11450
rect 8130 11398 8142 11450
rect 8142 11398 8172 11450
rect 8196 11398 8206 11450
rect 8206 11398 8252 11450
rect 7956 11396 8012 11398
rect 8036 11396 8092 11398
rect 8116 11396 8172 11398
rect 8196 11396 8252 11398
rect 9016 22874 9072 22876
rect 9096 22874 9152 22876
rect 9176 22874 9232 22876
rect 9256 22874 9312 22876
rect 9016 22822 9062 22874
rect 9062 22822 9072 22874
rect 9096 22822 9126 22874
rect 9126 22822 9138 22874
rect 9138 22822 9152 22874
rect 9176 22822 9190 22874
rect 9190 22822 9202 22874
rect 9202 22822 9232 22874
rect 9256 22822 9266 22874
rect 9266 22822 9312 22874
rect 9016 22820 9072 22822
rect 9096 22820 9152 22822
rect 9176 22820 9232 22822
rect 9256 22820 9312 22822
rect 9402 21936 9458 21992
rect 9016 21786 9072 21788
rect 9096 21786 9152 21788
rect 9176 21786 9232 21788
rect 9256 21786 9312 21788
rect 9016 21734 9062 21786
rect 9062 21734 9072 21786
rect 9096 21734 9126 21786
rect 9126 21734 9138 21786
rect 9138 21734 9152 21786
rect 9176 21734 9190 21786
rect 9190 21734 9202 21786
rect 9202 21734 9232 21786
rect 9256 21734 9266 21786
rect 9266 21734 9312 21786
rect 9016 21732 9072 21734
rect 9096 21732 9152 21734
rect 9176 21732 9232 21734
rect 9256 21732 9312 21734
rect 9034 21428 9036 21448
rect 9036 21428 9088 21448
rect 9088 21428 9090 21448
rect 9034 21392 9090 21428
rect 8666 20440 8722 20496
rect 9016 20698 9072 20700
rect 9096 20698 9152 20700
rect 9176 20698 9232 20700
rect 9256 20698 9312 20700
rect 9016 20646 9062 20698
rect 9062 20646 9072 20698
rect 9096 20646 9126 20698
rect 9126 20646 9138 20698
rect 9138 20646 9152 20698
rect 9176 20646 9190 20698
rect 9190 20646 9202 20698
rect 9202 20646 9232 20698
rect 9256 20646 9266 20698
rect 9266 20646 9312 20698
rect 9016 20644 9072 20646
rect 9096 20644 9152 20646
rect 9176 20644 9232 20646
rect 9256 20644 9312 20646
rect 9126 20440 9182 20496
rect 8942 20340 8944 20360
rect 8944 20340 8996 20360
rect 8996 20340 8998 20360
rect 8942 20304 8998 20340
rect 9034 19760 9090 19816
rect 9016 19610 9072 19612
rect 9096 19610 9152 19612
rect 9176 19610 9232 19612
rect 9256 19610 9312 19612
rect 9016 19558 9062 19610
rect 9062 19558 9072 19610
rect 9096 19558 9126 19610
rect 9126 19558 9138 19610
rect 9138 19558 9152 19610
rect 9176 19558 9190 19610
rect 9190 19558 9202 19610
rect 9202 19558 9232 19610
rect 9256 19558 9266 19610
rect 9266 19558 9312 19610
rect 9016 19556 9072 19558
rect 9096 19556 9152 19558
rect 9176 19556 9232 19558
rect 9256 19556 9312 19558
rect 8942 19352 8998 19408
rect 9770 24520 9826 24576
rect 9678 24248 9734 24304
rect 9678 23704 9734 23760
rect 10230 29960 10286 30016
rect 10414 29280 10470 29336
rect 10322 28872 10378 28928
rect 10230 27784 10286 27840
rect 10414 27512 10470 27568
rect 10230 26968 10286 27024
rect 9954 26152 10010 26208
rect 9678 23196 9680 23216
rect 9680 23196 9732 23216
rect 9732 23196 9734 23216
rect 9678 23160 9734 23196
rect 9770 22616 9826 22672
rect 9678 22344 9734 22400
rect 9862 22072 9918 22128
rect 9678 21800 9734 21856
rect 9862 21528 9918 21584
rect 9678 21256 9734 21312
rect 9678 20712 9734 20768
rect 9678 20168 9734 20224
rect 9678 19352 9734 19408
rect 9310 18672 9366 18728
rect 9016 18522 9072 18524
rect 9096 18522 9152 18524
rect 9176 18522 9232 18524
rect 9256 18522 9312 18524
rect 9016 18470 9062 18522
rect 9062 18470 9072 18522
rect 9096 18470 9126 18522
rect 9126 18470 9138 18522
rect 9138 18470 9152 18522
rect 9176 18470 9190 18522
rect 9190 18470 9202 18522
rect 9202 18470 9232 18522
rect 9256 18470 9266 18522
rect 9266 18470 9312 18522
rect 9016 18468 9072 18470
rect 9096 18468 9152 18470
rect 9176 18468 9232 18470
rect 9256 18468 9312 18470
rect 9034 18264 9090 18320
rect 8574 16088 8630 16144
rect 9016 17434 9072 17436
rect 9096 17434 9152 17436
rect 9176 17434 9232 17436
rect 9256 17434 9312 17436
rect 9016 17382 9062 17434
rect 9062 17382 9072 17434
rect 9096 17382 9126 17434
rect 9126 17382 9138 17434
rect 9138 17382 9152 17434
rect 9176 17382 9190 17434
rect 9190 17382 9202 17434
rect 9202 17382 9232 17434
rect 9256 17382 9266 17434
rect 9266 17382 9312 17434
rect 9016 17380 9072 17382
rect 9096 17380 9152 17382
rect 9176 17380 9232 17382
rect 9256 17380 9312 17382
rect 9678 19080 9734 19136
rect 9678 18708 9680 18728
rect 9680 18708 9732 18728
rect 9732 18708 9734 18728
rect 9678 18672 9734 18708
rect 9678 18536 9734 18592
rect 10046 26016 10102 26072
rect 10322 26152 10378 26208
rect 10230 25608 10286 25664
rect 10046 19896 10102 19952
rect 9954 18264 10010 18320
rect 9862 17992 9918 18048
rect 9770 17740 9826 17776
rect 9770 17720 9772 17740
rect 9772 17720 9824 17740
rect 9824 17720 9826 17740
rect 9678 17448 9734 17504
rect 9586 17312 9642 17368
rect 9310 17176 9366 17232
rect 9016 16346 9072 16348
rect 9096 16346 9152 16348
rect 9176 16346 9232 16348
rect 9256 16346 9312 16348
rect 9016 16294 9062 16346
rect 9062 16294 9072 16346
rect 9096 16294 9126 16346
rect 9126 16294 9138 16346
rect 9138 16294 9152 16346
rect 9176 16294 9190 16346
rect 9190 16294 9202 16346
rect 9202 16294 9232 16346
rect 9256 16294 9266 16346
rect 9266 16294 9312 16346
rect 9016 16292 9072 16294
rect 9096 16292 9152 16294
rect 9176 16292 9232 16294
rect 9256 16292 9312 16294
rect 8666 15136 8722 15192
rect 8758 15000 8814 15056
rect 9016 15258 9072 15260
rect 9096 15258 9152 15260
rect 9176 15258 9232 15260
rect 9256 15258 9312 15260
rect 9016 15206 9062 15258
rect 9062 15206 9072 15258
rect 9096 15206 9126 15258
rect 9126 15206 9138 15258
rect 9138 15206 9152 15258
rect 9176 15206 9190 15258
rect 9190 15206 9202 15258
rect 9202 15206 9232 15258
rect 9256 15206 9266 15258
rect 9266 15206 9312 15258
rect 9016 15204 9072 15206
rect 9096 15204 9152 15206
rect 9176 15204 9232 15206
rect 9256 15204 9312 15206
rect 8666 14456 8722 14512
rect 8850 14456 8906 14512
rect 9310 14612 9366 14648
rect 9310 14592 9312 14612
rect 9312 14592 9364 14612
rect 9364 14592 9366 14612
rect 9494 14884 9550 14920
rect 9494 14864 9496 14884
rect 9496 14864 9548 14884
rect 9548 14864 9550 14884
rect 8574 12688 8630 12744
rect 9016 14170 9072 14172
rect 9096 14170 9152 14172
rect 9176 14170 9232 14172
rect 9256 14170 9312 14172
rect 9016 14118 9062 14170
rect 9062 14118 9072 14170
rect 9096 14118 9126 14170
rect 9126 14118 9138 14170
rect 9138 14118 9152 14170
rect 9176 14118 9190 14170
rect 9190 14118 9202 14170
rect 9202 14118 9232 14170
rect 9256 14118 9266 14170
rect 9266 14118 9312 14170
rect 9016 14116 9072 14118
rect 9096 14116 9152 14118
rect 9176 14116 9232 14118
rect 9256 14116 9312 14118
rect 9402 13504 9458 13560
rect 9770 17176 9826 17232
rect 9678 16904 9734 16960
rect 9678 16632 9734 16688
rect 9770 16360 9826 16416
rect 9862 16088 9918 16144
rect 9678 15816 9734 15872
rect 9770 15564 9826 15600
rect 9770 15544 9772 15564
rect 9772 15544 9824 15564
rect 9824 15544 9826 15564
rect 9770 14728 9826 14784
rect 9016 13082 9072 13084
rect 9096 13082 9152 13084
rect 9176 13082 9232 13084
rect 9256 13082 9312 13084
rect 9016 13030 9062 13082
rect 9062 13030 9072 13082
rect 9096 13030 9126 13082
rect 9126 13030 9138 13082
rect 9138 13030 9152 13082
rect 9176 13030 9190 13082
rect 9190 13030 9202 13082
rect 9202 13030 9232 13082
rect 9256 13030 9266 13082
rect 9266 13030 9312 13082
rect 9016 13028 9072 13030
rect 9096 13028 9152 13030
rect 9176 13028 9232 13030
rect 9256 13028 9312 13030
rect 8850 12824 8906 12880
rect 9586 13232 9642 13288
rect 9678 13096 9734 13152
rect 9770 12824 9826 12880
rect 9126 12316 9128 12336
rect 9128 12316 9180 12336
rect 9180 12316 9182 12336
rect 9126 12280 9182 12316
rect 9954 13640 10010 13696
rect 9954 13232 10010 13288
rect 9016 11994 9072 11996
rect 9096 11994 9152 11996
rect 9176 11994 9232 11996
rect 9256 11994 9312 11996
rect 9016 11942 9062 11994
rect 9062 11942 9072 11994
rect 9096 11942 9126 11994
rect 9126 11942 9138 11994
rect 9138 11942 9152 11994
rect 9176 11942 9190 11994
rect 9190 11942 9202 11994
rect 9202 11942 9232 11994
rect 9256 11942 9266 11994
rect 9266 11942 9312 11994
rect 9016 11940 9072 11942
rect 9096 11940 9152 11942
rect 9176 11940 9232 11942
rect 9256 11940 9312 11942
rect 9126 11636 9128 11656
rect 9128 11636 9180 11656
rect 9180 11636 9182 11656
rect 9126 11600 9182 11636
rect 8942 11464 8998 11520
rect 9494 11192 9550 11248
rect 8482 10512 8538 10568
rect 7956 10362 8012 10364
rect 8036 10362 8092 10364
rect 8116 10362 8172 10364
rect 8196 10362 8252 10364
rect 7956 10310 8002 10362
rect 8002 10310 8012 10362
rect 8036 10310 8066 10362
rect 8066 10310 8078 10362
rect 8078 10310 8092 10362
rect 8116 10310 8130 10362
rect 8130 10310 8142 10362
rect 8142 10310 8172 10362
rect 8196 10310 8206 10362
rect 8206 10310 8252 10362
rect 7956 10308 8012 10310
rect 8036 10308 8092 10310
rect 8116 10308 8172 10310
rect 8196 10308 8252 10310
rect 8022 9868 8024 9888
rect 8024 9868 8076 9888
rect 8076 9868 8078 9888
rect 8022 9832 8078 9868
rect 7956 9274 8012 9276
rect 8036 9274 8092 9276
rect 8116 9274 8172 9276
rect 8196 9274 8252 9276
rect 7956 9222 8002 9274
rect 8002 9222 8012 9274
rect 8036 9222 8066 9274
rect 8066 9222 8078 9274
rect 8078 9222 8092 9274
rect 8116 9222 8130 9274
rect 8130 9222 8142 9274
rect 8142 9222 8172 9274
rect 8196 9222 8206 9274
rect 8206 9222 8252 9274
rect 7956 9220 8012 9222
rect 8036 9220 8092 9222
rect 8116 9220 8172 9222
rect 8196 9220 8252 9222
rect 8206 8472 8262 8528
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 8298 7248 8354 7304
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 6918 2624 6974 2680
rect 6458 1128 6514 1184
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8482 8608 8538 8664
rect 9016 10906 9072 10908
rect 9096 10906 9152 10908
rect 9176 10906 9232 10908
rect 9256 10906 9312 10908
rect 9016 10854 9062 10906
rect 9062 10854 9072 10906
rect 9096 10854 9126 10906
rect 9126 10854 9138 10906
rect 9138 10854 9152 10906
rect 9176 10854 9190 10906
rect 9190 10854 9202 10906
rect 9202 10854 9232 10906
rect 9256 10854 9266 10906
rect 9266 10854 9312 10906
rect 9016 10852 9072 10854
rect 9096 10852 9152 10854
rect 9176 10852 9232 10854
rect 9256 10852 9312 10854
rect 8850 10648 8906 10704
rect 8850 10104 8906 10160
rect 8666 9560 8722 9616
rect 9016 9818 9072 9820
rect 9096 9818 9152 9820
rect 9176 9818 9232 9820
rect 9256 9818 9312 9820
rect 9016 9766 9062 9818
rect 9062 9766 9072 9818
rect 9096 9766 9126 9818
rect 9126 9766 9138 9818
rect 9138 9766 9152 9818
rect 9176 9766 9190 9818
rect 9190 9766 9202 9818
rect 9202 9766 9232 9818
rect 9256 9766 9266 9818
rect 9266 9766 9312 9818
rect 9016 9764 9072 9766
rect 9096 9764 9152 9766
rect 9176 9764 9232 9766
rect 9256 9764 9312 9766
rect 9862 12300 9918 12336
rect 9862 12280 9864 12300
rect 9864 12280 9916 12300
rect 9916 12280 9918 12300
rect 9678 12008 9734 12064
rect 9770 11736 9826 11792
rect 9770 11464 9826 11520
rect 9954 11192 10010 11248
rect 9862 10920 9918 10976
rect 9770 10376 9826 10432
rect 9678 9832 9734 9888
rect 9494 9424 9550 9480
rect 9310 8880 9366 8936
rect 8574 8336 8630 8392
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 9310 8472 9366 8528
rect 8574 7520 8630 7576
rect 9310 7928 9366 7984
rect 8942 7792 8998 7848
rect 9770 9016 9826 9072
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 8850 7404 8906 7440
rect 9494 7656 9550 7712
rect 8850 7384 8852 7404
rect 8852 7384 8904 7404
rect 8904 7384 8906 7404
rect 9494 7268 9550 7304
rect 9494 7248 9496 7268
rect 9496 7248 9548 7268
rect 9548 7248 9550 7268
rect 8298 5072 8354 5128
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9402 6840 9458 6896
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9494 6704 9550 6760
rect 9862 8744 9918 8800
rect 9678 8472 9734 8528
rect 10046 9560 10102 9616
rect 9954 8200 10010 8256
rect 9678 7948 9734 7984
rect 9678 7928 9680 7948
rect 9680 7928 9732 7948
rect 9732 7928 9734 7948
rect 9770 7656 9826 7712
rect 9862 7384 9918 7440
rect 9678 7112 9734 7168
rect 9954 6840 10010 6896
rect 9678 6568 9734 6624
rect 9770 6296 9826 6352
rect 9770 6024 9826 6080
rect 9678 5480 9734 5536
rect 9770 5208 9826 5264
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 10230 24792 10286 24848
rect 10230 23976 10286 24032
rect 10230 23468 10232 23488
rect 10232 23468 10284 23488
rect 10284 23468 10286 23488
rect 10230 23432 10286 23468
rect 10230 22924 10232 22944
rect 10232 22924 10284 22944
rect 10284 22924 10286 22944
rect 10230 22888 10286 22924
rect 10230 21020 10232 21040
rect 10232 21020 10284 21040
rect 10284 21020 10286 21040
rect 10230 20984 10286 21020
rect 10230 20440 10286 20496
rect 10230 19624 10286 19680
rect 10598 28600 10654 28656
rect 10414 19488 10470 19544
rect 10230 18844 10232 18864
rect 10232 18844 10284 18864
rect 10284 18844 10286 18864
rect 10230 18808 10286 18844
rect 10322 15408 10378 15464
rect 10322 13912 10378 13968
rect 10782 26424 10838 26480
rect 10690 21664 10746 21720
rect 10690 19216 10746 19272
rect 10506 15272 10562 15328
rect 10414 13232 10470 13288
rect 10230 12552 10286 12608
rect 10690 14184 10746 14240
rect 10782 10104 10838 10160
rect 10966 13368 11022 13424
rect 10966 9288 11022 9344
rect 10690 5752 10746 5808
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9218 1128 9274 1184
rect 10138 1264 10194 1320
<< metal3 >>
rect 3006 42464 3322 42465
rect 3006 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3322 42464
rect 3006 42399 3322 42400
rect 9006 42464 9322 42465
rect 9006 42400 9012 42464
rect 9076 42400 9092 42464
rect 9156 42400 9172 42464
rect 9236 42400 9252 42464
rect 9316 42400 9322 42464
rect 9006 42399 9322 42400
rect 1946 41920 2262 41921
rect 1946 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2262 41920
rect 1946 41855 2262 41856
rect 7946 41920 8262 41921
rect 7946 41856 7952 41920
rect 8016 41856 8032 41920
rect 8096 41856 8112 41920
rect 8176 41856 8192 41920
rect 8256 41856 8262 41920
rect 7946 41855 8262 41856
rect 790 41516 796 41580
rect 860 41578 866 41580
rect 9581 41578 9647 41581
rect 860 41576 9647 41578
rect 860 41520 9586 41576
rect 9642 41520 9647 41576
rect 860 41518 9647 41520
rect 860 41516 866 41518
rect 9581 41515 9647 41518
rect 3006 41376 3322 41377
rect 3006 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3322 41376
rect 3006 41311 3322 41312
rect 9006 41376 9322 41377
rect 9006 41312 9012 41376
rect 9076 41312 9092 41376
rect 9156 41312 9172 41376
rect 9236 41312 9252 41376
rect 9316 41312 9322 41376
rect 9006 41311 9322 41312
rect 606 40972 612 41036
rect 676 41034 682 41036
rect 7005 41034 7071 41037
rect 676 41032 7071 41034
rect 676 40976 7010 41032
rect 7066 40976 7071 41032
rect 676 40974 7071 40976
rect 676 40972 682 40974
rect 7005 40971 7071 40974
rect 0 40898 120 40928
rect 1485 40898 1551 40901
rect 0 40896 1551 40898
rect 0 40840 1490 40896
rect 1546 40840 1551 40896
rect 0 40838 1551 40840
rect 0 40808 120 40838
rect 1485 40835 1551 40838
rect 1946 40832 2262 40833
rect 1946 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2262 40832
rect 1946 40767 2262 40768
rect 7946 40832 8262 40833
rect 7946 40768 7952 40832
rect 8016 40768 8032 40832
rect 8096 40768 8112 40832
rect 8176 40768 8192 40832
rect 8256 40768 8262 40832
rect 7946 40767 8262 40768
rect 7741 40356 7807 40357
rect 9765 40356 9831 40357
rect 7741 40354 7788 40356
rect 7696 40352 7788 40354
rect 7696 40296 7746 40352
rect 7696 40294 7788 40296
rect 7741 40292 7788 40294
rect 7852 40292 7858 40356
rect 9765 40354 9812 40356
rect 9720 40352 9812 40354
rect 9720 40296 9770 40352
rect 9720 40294 9812 40296
rect 9765 40292 9812 40294
rect 9876 40292 9882 40356
rect 7741 40291 7807 40292
rect 9765 40291 9831 40292
rect 3006 40288 3322 40289
rect 3006 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3322 40288
rect 3006 40223 3322 40224
rect 9006 40288 9322 40289
rect 9006 40224 9012 40288
rect 9076 40224 9092 40288
rect 9156 40224 9172 40288
rect 9236 40224 9252 40288
rect 9316 40224 9322 40288
rect 9006 40223 9322 40224
rect 9397 40218 9463 40221
rect 10174 40218 10180 40220
rect 9397 40216 10180 40218
rect 9397 40160 9402 40216
rect 9458 40160 10180 40216
rect 9397 40158 10180 40160
rect 9397 40155 9463 40158
rect 10174 40156 10180 40158
rect 10244 40156 10250 40220
rect 0 40082 120 40112
rect 1485 40082 1551 40085
rect 0 40080 1551 40082
rect 0 40024 1490 40080
rect 1546 40024 1551 40080
rect 0 40022 1551 40024
rect 0 39992 120 40022
rect 1485 40019 1551 40022
rect 5206 40020 5212 40084
rect 5276 40082 5282 40084
rect 9213 40082 9279 40085
rect 5276 40080 9279 40082
rect 5276 40024 9218 40080
rect 9274 40024 9279 40080
rect 5276 40022 9279 40024
rect 5276 40020 5282 40022
rect 9213 40019 9279 40022
rect 10409 39810 10475 39813
rect 11130 39810 11250 39840
rect 10409 39808 11250 39810
rect 10409 39752 10414 39808
rect 10470 39752 11250 39808
rect 10409 39750 11250 39752
rect 10409 39747 10475 39750
rect 1946 39744 2262 39745
rect 1946 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2262 39744
rect 1946 39679 2262 39680
rect 7946 39744 8262 39745
rect 7946 39680 7952 39744
rect 8016 39680 8032 39744
rect 8096 39680 8112 39744
rect 8176 39680 8192 39744
rect 8256 39680 8262 39744
rect 11130 39720 11250 39750
rect 7946 39679 8262 39680
rect 8661 39674 8727 39677
rect 10542 39674 10548 39676
rect 8661 39672 10548 39674
rect 8661 39616 8666 39672
rect 8722 39616 10548 39672
rect 8661 39614 10548 39616
rect 8661 39611 8727 39614
rect 10542 39612 10548 39614
rect 10612 39612 10618 39676
rect 974 39476 980 39540
rect 1044 39538 1050 39540
rect 7373 39538 7439 39541
rect 1044 39536 7439 39538
rect 1044 39480 7378 39536
rect 7434 39480 7439 39536
rect 1044 39478 7439 39480
rect 1044 39476 1050 39478
rect 7373 39475 7439 39478
rect 10593 39538 10659 39541
rect 11130 39538 11250 39568
rect 10593 39536 11250 39538
rect 10593 39480 10598 39536
rect 10654 39480 11250 39536
rect 10593 39478 11250 39480
rect 10593 39475 10659 39478
rect 11130 39448 11250 39478
rect 8702 39340 8708 39404
rect 8772 39402 8778 39404
rect 9489 39402 9555 39405
rect 8772 39400 9555 39402
rect 8772 39344 9494 39400
rect 9550 39344 9555 39400
rect 8772 39342 9555 39344
rect 8772 39340 8778 39342
rect 9489 39339 9555 39342
rect 0 39266 120 39296
rect 1485 39266 1551 39269
rect 0 39264 1551 39266
rect 0 39208 1490 39264
rect 1546 39208 1551 39264
rect 0 39206 1551 39208
rect 0 39176 120 39206
rect 1485 39203 1551 39206
rect 9673 39266 9739 39269
rect 11130 39266 11250 39296
rect 9673 39264 11250 39266
rect 9673 39208 9678 39264
rect 9734 39208 11250 39264
rect 9673 39206 11250 39208
rect 9673 39203 9739 39206
rect 3006 39200 3322 39201
rect 3006 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3322 39200
rect 3006 39135 3322 39136
rect 9006 39200 9322 39201
rect 9006 39136 9012 39200
rect 9076 39136 9092 39200
rect 9156 39136 9172 39200
rect 9236 39136 9252 39200
rect 9316 39136 9322 39200
rect 11130 39176 11250 39206
rect 9006 39135 9322 39136
rect 10225 38994 10291 38997
rect 11130 38994 11250 39024
rect 10225 38992 11250 38994
rect 10225 38936 10230 38992
rect 10286 38936 11250 38992
rect 10225 38934 11250 38936
rect 10225 38931 10291 38934
rect 11130 38904 11250 38934
rect 5942 38796 5948 38860
rect 6012 38858 6018 38860
rect 8753 38858 8819 38861
rect 6012 38856 8819 38858
rect 6012 38800 8758 38856
rect 8814 38800 8819 38856
rect 6012 38798 8819 38800
rect 6012 38796 6018 38798
rect 8753 38795 8819 38798
rect 8334 38660 8340 38724
rect 8404 38722 8410 38724
rect 9121 38722 9187 38725
rect 8404 38720 9187 38722
rect 8404 38664 9126 38720
rect 9182 38664 9187 38720
rect 8404 38662 9187 38664
rect 8404 38660 8410 38662
rect 9121 38659 9187 38662
rect 10777 38722 10843 38725
rect 11130 38722 11250 38752
rect 10777 38720 11250 38722
rect 10777 38664 10782 38720
rect 10838 38664 11250 38720
rect 10777 38662 11250 38664
rect 10777 38659 10843 38662
rect 1946 38656 2262 38657
rect 1946 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2262 38656
rect 1946 38591 2262 38592
rect 7946 38656 8262 38657
rect 7946 38592 7952 38656
rect 8016 38592 8032 38656
rect 8096 38592 8112 38656
rect 8176 38592 8192 38656
rect 8256 38592 8262 38656
rect 11130 38632 11250 38662
rect 7946 38591 8262 38592
rect 0 38450 120 38480
rect 749 38450 815 38453
rect 0 38448 815 38450
rect 0 38392 754 38448
rect 810 38392 815 38448
rect 0 38390 815 38392
rect 0 38360 120 38390
rect 749 38387 815 38390
rect 10133 38450 10199 38453
rect 11130 38450 11250 38480
rect 10133 38448 11250 38450
rect 10133 38392 10138 38448
rect 10194 38392 11250 38448
rect 10133 38390 11250 38392
rect 10133 38387 10199 38390
rect 11130 38360 11250 38390
rect 9121 38314 9187 38317
rect 10358 38314 10364 38316
rect 9121 38312 10364 38314
rect 9121 38256 9126 38312
rect 9182 38256 10364 38312
rect 9121 38254 10364 38256
rect 9121 38251 9187 38254
rect 10358 38252 10364 38254
rect 10428 38252 10434 38316
rect 10409 38178 10475 38181
rect 11130 38178 11250 38208
rect 10409 38176 11250 38178
rect 10409 38120 10414 38176
rect 10470 38120 11250 38176
rect 10409 38118 11250 38120
rect 10409 38115 10475 38118
rect 3006 38112 3322 38113
rect 3006 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3322 38112
rect 3006 38047 3322 38048
rect 9006 38112 9322 38113
rect 9006 38048 9012 38112
rect 9076 38048 9092 38112
rect 9156 38048 9172 38112
rect 9236 38048 9252 38112
rect 9316 38048 9322 38112
rect 11130 38088 11250 38118
rect 9006 38047 9322 38048
rect 10317 37906 10383 37909
rect 11130 37906 11250 37936
rect 10317 37904 11250 37906
rect 10317 37848 10322 37904
rect 10378 37848 11250 37904
rect 10317 37846 11250 37848
rect 10317 37843 10383 37846
rect 11130 37816 11250 37846
rect 4470 37708 4476 37772
rect 4540 37770 4546 37772
rect 8477 37770 8543 37773
rect 4540 37768 8543 37770
rect 4540 37712 8482 37768
rect 8538 37712 8543 37768
rect 4540 37710 8543 37712
rect 4540 37708 4546 37710
rect 8477 37707 8543 37710
rect 0 37634 120 37664
rect 1485 37634 1551 37637
rect 0 37632 1551 37634
rect 0 37576 1490 37632
rect 1546 37576 1551 37632
rect 0 37574 1551 37576
rect 0 37544 120 37574
rect 1485 37571 1551 37574
rect 10225 37634 10291 37637
rect 11130 37634 11250 37664
rect 10225 37632 11250 37634
rect 10225 37576 10230 37632
rect 10286 37576 11250 37632
rect 10225 37574 11250 37576
rect 10225 37571 10291 37574
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 7946 37568 8262 37569
rect 7946 37504 7952 37568
rect 8016 37504 8032 37568
rect 8096 37504 8112 37568
rect 8176 37504 8192 37568
rect 8256 37504 8262 37568
rect 11130 37544 11250 37574
rect 7946 37503 8262 37504
rect 6494 37300 6500 37364
rect 6564 37362 6570 37364
rect 8753 37362 8819 37365
rect 6564 37360 8819 37362
rect 6564 37304 8758 37360
rect 8814 37304 8819 37360
rect 6564 37302 8819 37304
rect 6564 37300 6570 37302
rect 8753 37299 8819 37302
rect 9949 37362 10015 37365
rect 11130 37362 11250 37392
rect 9949 37360 11250 37362
rect 9949 37304 9954 37360
rect 10010 37304 11250 37360
rect 9949 37302 11250 37304
rect 9949 37299 10015 37302
rect 11130 37272 11250 37302
rect 4521 37226 4587 37229
rect 4981 37228 5047 37229
rect 4981 37226 5028 37228
rect 4521 37224 5028 37226
rect 4521 37168 4526 37224
rect 4582 37168 4986 37224
rect 4521 37166 5028 37168
rect 4521 37163 4587 37166
rect 4981 37164 5028 37166
rect 5092 37164 5098 37228
rect 6453 37226 6519 37229
rect 6862 37226 6868 37228
rect 6453 37224 6868 37226
rect 6453 37168 6458 37224
rect 6514 37168 6868 37224
rect 6453 37166 6868 37168
rect 4981 37163 5047 37164
rect 6453 37163 6519 37166
rect 6862 37164 6868 37166
rect 6932 37226 6938 37228
rect 7557 37226 7623 37229
rect 6932 37224 7623 37226
rect 6932 37168 7562 37224
rect 7618 37168 7623 37224
rect 6932 37166 7623 37168
rect 6932 37164 6938 37166
rect 7557 37163 7623 37166
rect 10041 37090 10107 37093
rect 11130 37090 11250 37120
rect 10041 37088 11250 37090
rect 10041 37032 10046 37088
rect 10102 37032 11250 37088
rect 10041 37030 11250 37032
rect 10041 37027 10107 37030
rect 3006 37024 3322 37025
rect 3006 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3322 37024
rect 3006 36959 3322 36960
rect 9006 37024 9322 37025
rect 9006 36960 9012 37024
rect 9076 36960 9092 37024
rect 9156 36960 9172 37024
rect 9236 36960 9252 37024
rect 9316 36960 9322 37024
rect 11130 37000 11250 37030
rect 9006 36959 9322 36960
rect 0 36818 120 36848
rect 1485 36818 1551 36821
rect 0 36816 1551 36818
rect 0 36760 1490 36816
rect 1546 36760 1551 36816
rect 0 36758 1551 36760
rect 0 36728 120 36758
rect 1485 36755 1551 36758
rect 1669 36818 1735 36821
rect 4654 36818 4660 36820
rect 1669 36816 4660 36818
rect 1669 36760 1674 36816
rect 1730 36760 4660 36816
rect 1669 36758 4660 36760
rect 1669 36755 1735 36758
rect 4654 36756 4660 36758
rect 4724 36756 4730 36820
rect 10501 36818 10567 36821
rect 11130 36818 11250 36848
rect 10501 36816 11250 36818
rect 10501 36760 10506 36816
rect 10562 36760 11250 36816
rect 10501 36758 11250 36760
rect 10501 36755 10567 36758
rect 11130 36728 11250 36758
rect 7557 36682 7623 36685
rect 8109 36682 8175 36685
rect 7557 36680 8175 36682
rect 7557 36624 7562 36680
rect 7618 36624 8114 36680
rect 8170 36624 8175 36680
rect 7557 36622 8175 36624
rect 7557 36619 7623 36622
rect 8109 36619 8175 36622
rect 10133 36546 10199 36549
rect 11130 36546 11250 36576
rect 10133 36544 11250 36546
rect 10133 36488 10138 36544
rect 10194 36488 11250 36544
rect 10133 36486 11250 36488
rect 10133 36483 10199 36486
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 7946 36480 8262 36481
rect 7946 36416 7952 36480
rect 8016 36416 8032 36480
rect 8096 36416 8112 36480
rect 8176 36416 8192 36480
rect 8256 36416 8262 36480
rect 11130 36456 11250 36486
rect 7946 36415 8262 36416
rect 10961 36274 11027 36277
rect 11130 36274 11250 36304
rect 10961 36272 11250 36274
rect 10961 36216 10966 36272
rect 11022 36216 11250 36272
rect 10961 36214 11250 36216
rect 10961 36211 11027 36214
rect 11130 36184 11250 36214
rect 3734 36076 3740 36140
rect 3804 36138 3810 36140
rect 9121 36138 9187 36141
rect 3804 36136 9187 36138
rect 3804 36080 9126 36136
rect 9182 36080 9187 36136
rect 3804 36078 9187 36080
rect 3804 36076 3810 36078
rect 9121 36075 9187 36078
rect 0 36002 120 36032
rect 1485 36002 1551 36005
rect 0 36000 1551 36002
rect 0 35944 1490 36000
rect 1546 35944 1551 36000
rect 0 35942 1551 35944
rect 0 35912 120 35942
rect 1485 35939 1551 35942
rect 1853 36002 1919 36005
rect 10317 36002 10383 36005
rect 11130 36002 11250 36032
rect 1853 36000 1962 36002
rect 1853 35944 1858 36000
rect 1914 35944 1962 36000
rect 1853 35939 1962 35944
rect 10317 36000 11250 36002
rect 10317 35944 10322 36000
rect 10378 35944 11250 36000
rect 10317 35942 11250 35944
rect 10317 35939 10383 35942
rect 1526 35804 1532 35868
rect 1596 35866 1602 35868
rect 1902 35866 1962 35939
rect 3006 35936 3322 35937
rect 3006 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3322 35936
rect 3006 35871 3322 35872
rect 9006 35936 9322 35937
rect 9006 35872 9012 35936
rect 9076 35872 9092 35936
rect 9156 35872 9172 35936
rect 9236 35872 9252 35936
rect 9316 35872 9322 35936
rect 11130 35912 11250 35942
rect 9006 35871 9322 35872
rect 1596 35806 1962 35866
rect 3877 35866 3943 35869
rect 8569 35868 8635 35869
rect 7414 35866 7420 35868
rect 3877 35864 7420 35866
rect 3877 35808 3882 35864
rect 3938 35808 7420 35864
rect 3877 35806 7420 35808
rect 1596 35804 1602 35806
rect 3877 35803 3943 35806
rect 7414 35804 7420 35806
rect 7484 35804 7490 35868
rect 8518 35866 8524 35868
rect 8478 35806 8524 35866
rect 8588 35864 8635 35868
rect 8630 35808 8635 35864
rect 8518 35804 8524 35806
rect 8588 35804 8635 35808
rect 8569 35803 8635 35804
rect 2630 35668 2636 35732
rect 2700 35730 2706 35732
rect 2773 35730 2839 35733
rect 2700 35728 2839 35730
rect 2700 35672 2778 35728
rect 2834 35672 2839 35728
rect 2700 35670 2839 35672
rect 2700 35668 2706 35670
rect 2773 35667 2839 35670
rect 7782 35668 7788 35732
rect 7852 35730 7858 35732
rect 9990 35730 9996 35732
rect 7852 35670 9996 35730
rect 7852 35668 7858 35670
rect 9990 35668 9996 35670
rect 10060 35668 10066 35732
rect 10593 35730 10659 35733
rect 11130 35730 11250 35760
rect 10593 35728 11250 35730
rect 10593 35672 10598 35728
rect 10654 35672 11250 35728
rect 10593 35670 11250 35672
rect 10593 35667 10659 35670
rect 11130 35640 11250 35670
rect 1669 35594 1735 35597
rect 6361 35594 6427 35597
rect 1669 35592 6427 35594
rect 1669 35536 1674 35592
rect 1730 35536 6366 35592
rect 6422 35536 6427 35592
rect 1669 35534 6427 35536
rect 1669 35531 1735 35534
rect 6361 35531 6427 35534
rect 8569 35594 8635 35597
rect 8753 35594 8819 35597
rect 8569 35592 8819 35594
rect 8569 35536 8574 35592
rect 8630 35536 8758 35592
rect 8814 35536 8819 35592
rect 8569 35534 8819 35536
rect 8569 35531 8635 35534
rect 8753 35531 8819 35534
rect 10501 35458 10567 35461
rect 11130 35458 11250 35488
rect 10501 35456 11250 35458
rect 10501 35400 10506 35456
rect 10562 35400 11250 35456
rect 10501 35398 11250 35400
rect 10501 35395 10567 35398
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 7946 35392 8262 35393
rect 7946 35328 7952 35392
rect 8016 35328 8032 35392
rect 8096 35328 8112 35392
rect 8176 35328 8192 35392
rect 8256 35328 8262 35392
rect 11130 35368 11250 35398
rect 7946 35327 8262 35328
rect 0 35186 120 35216
rect 1485 35186 1551 35189
rect 0 35184 1551 35186
rect 0 35128 1490 35184
rect 1546 35128 1551 35184
rect 0 35126 1551 35128
rect 0 35096 120 35126
rect 1485 35123 1551 35126
rect 3233 35186 3299 35189
rect 5390 35186 5396 35188
rect 3233 35184 5396 35186
rect 3233 35128 3238 35184
rect 3294 35128 5396 35184
rect 3233 35126 5396 35128
rect 3233 35123 3299 35126
rect 5390 35124 5396 35126
rect 5460 35124 5466 35188
rect 6269 35186 6335 35189
rect 9438 35186 9444 35188
rect 6269 35184 9444 35186
rect 6269 35128 6274 35184
rect 6330 35128 9444 35184
rect 6269 35126 9444 35128
rect 6269 35123 6335 35126
rect 9438 35124 9444 35126
rect 9508 35124 9514 35188
rect 9673 35186 9739 35189
rect 11130 35186 11250 35216
rect 9673 35184 11250 35186
rect 9673 35128 9678 35184
rect 9734 35128 11250 35184
rect 9673 35126 11250 35128
rect 9673 35123 9739 35126
rect 11130 35096 11250 35126
rect 1117 35050 1183 35053
rect 8937 35050 9003 35053
rect 1117 35048 9003 35050
rect 1117 34992 1122 35048
rect 1178 34992 8942 35048
rect 8998 34992 9003 35048
rect 1117 34990 9003 34992
rect 1117 34987 1183 34990
rect 8937 34987 9003 34990
rect 9949 34914 10015 34917
rect 11130 34914 11250 34944
rect 9949 34912 11250 34914
rect 9949 34856 9954 34912
rect 10010 34856 11250 34912
rect 9949 34854 11250 34856
rect 9949 34851 10015 34854
rect 3006 34848 3322 34849
rect 3006 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3322 34848
rect 3006 34783 3322 34784
rect 9006 34848 9322 34849
rect 9006 34784 9012 34848
rect 9076 34784 9092 34848
rect 9156 34784 9172 34848
rect 9236 34784 9252 34848
rect 9316 34784 9322 34848
rect 11130 34824 11250 34854
rect 9006 34783 9322 34784
rect 3550 34580 3556 34644
rect 3620 34642 3626 34644
rect 5165 34642 5231 34645
rect 3620 34640 5231 34642
rect 3620 34584 5170 34640
rect 5226 34584 5231 34640
rect 3620 34582 5231 34584
rect 3620 34580 3626 34582
rect 5165 34579 5231 34582
rect 9581 34642 9647 34645
rect 11130 34642 11250 34672
rect 9581 34640 11250 34642
rect 9581 34584 9586 34640
rect 9642 34584 11250 34640
rect 9581 34582 11250 34584
rect 9581 34579 9647 34582
rect 11130 34552 11250 34582
rect 2446 34444 2452 34508
rect 2516 34506 2522 34508
rect 6821 34506 6887 34509
rect 7046 34506 7052 34508
rect 2516 34446 2790 34506
rect 2516 34444 2522 34446
rect 0 34370 120 34400
rect 933 34370 999 34373
rect 0 34368 999 34370
rect 0 34312 938 34368
rect 994 34312 999 34368
rect 0 34310 999 34312
rect 2730 34370 2790 34446
rect 6821 34504 7052 34506
rect 6821 34448 6826 34504
rect 6882 34448 7052 34504
rect 6821 34446 7052 34448
rect 6821 34443 6887 34446
rect 7046 34444 7052 34446
rect 7116 34444 7122 34508
rect 7281 34370 7347 34373
rect 2730 34368 7347 34370
rect 2730 34312 7286 34368
rect 7342 34312 7347 34368
rect 2730 34310 7347 34312
rect 0 34280 120 34310
rect 933 34307 999 34310
rect 7281 34307 7347 34310
rect 10225 34370 10291 34373
rect 11130 34370 11250 34400
rect 10225 34368 11250 34370
rect 10225 34312 10230 34368
rect 10286 34312 11250 34368
rect 10225 34310 11250 34312
rect 10225 34307 10291 34310
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 7946 34304 8262 34305
rect 7946 34240 7952 34304
rect 8016 34240 8032 34304
rect 8096 34240 8112 34304
rect 8176 34240 8192 34304
rect 8256 34240 8262 34304
rect 11130 34280 11250 34310
rect 7946 34239 8262 34240
rect 6821 34236 6887 34237
rect 6821 34232 6868 34236
rect 6932 34234 6938 34236
rect 6821 34176 6826 34232
rect 6821 34172 6868 34176
rect 6932 34174 6978 34234
rect 6932 34172 6938 34174
rect 6821 34171 6887 34172
rect 10409 34098 10475 34101
rect 11130 34098 11250 34128
rect 10409 34096 11250 34098
rect 10409 34040 10414 34096
rect 10470 34040 11250 34096
rect 10409 34038 11250 34040
rect 10409 34035 10475 34038
rect 11130 34008 11250 34038
rect 6310 33900 6316 33964
rect 6380 33962 6386 33964
rect 9121 33962 9187 33965
rect 6380 33960 9187 33962
rect 6380 33904 9126 33960
rect 9182 33904 9187 33960
rect 6380 33902 9187 33904
rect 6380 33900 6386 33902
rect 9121 33899 9187 33902
rect 9949 33826 10015 33829
rect 11130 33826 11250 33856
rect 9949 33824 11250 33826
rect 9949 33768 9954 33824
rect 10010 33768 11250 33824
rect 9949 33766 11250 33768
rect 9949 33763 10015 33766
rect 3006 33760 3322 33761
rect 3006 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3322 33760
rect 3006 33695 3322 33696
rect 9006 33760 9322 33761
rect 9006 33696 9012 33760
rect 9076 33696 9092 33760
rect 9156 33696 9172 33760
rect 9236 33696 9252 33760
rect 9316 33696 9322 33760
rect 11130 33736 11250 33766
rect 9006 33695 9322 33696
rect 0 33554 120 33584
rect 381 33554 447 33557
rect 0 33552 447 33554
rect 0 33496 386 33552
rect 442 33496 447 33552
rect 0 33494 447 33496
rect 0 33464 120 33494
rect 381 33491 447 33494
rect 10593 33554 10659 33557
rect 11130 33554 11250 33584
rect 10593 33552 11250 33554
rect 10593 33496 10598 33552
rect 10654 33496 11250 33552
rect 10593 33494 11250 33496
rect 10593 33491 10659 33494
rect 11130 33464 11250 33494
rect 4153 33418 4219 33421
rect 4286 33418 4292 33420
rect 4153 33416 4292 33418
rect 4153 33360 4158 33416
rect 4214 33360 4292 33416
rect 4153 33358 4292 33360
rect 4153 33355 4219 33358
rect 4286 33356 4292 33358
rect 4356 33356 4362 33420
rect 5574 33356 5580 33420
rect 5644 33418 5650 33420
rect 9489 33418 9555 33421
rect 5644 33416 9555 33418
rect 5644 33360 9494 33416
rect 9550 33360 9555 33416
rect 5644 33358 9555 33360
rect 5644 33356 5650 33358
rect 9489 33355 9555 33358
rect 5625 33282 5691 33285
rect 4110 33280 5691 33282
rect 4110 33224 5630 33280
rect 5686 33224 5691 33280
rect 4110 33222 5691 33224
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 2814 33084 2820 33148
rect 2884 33146 2890 33148
rect 4110 33146 4170 33222
rect 5625 33219 5691 33222
rect 10133 33282 10199 33285
rect 11130 33282 11250 33312
rect 10133 33280 11250 33282
rect 10133 33224 10138 33280
rect 10194 33224 11250 33280
rect 10133 33222 11250 33224
rect 10133 33219 10199 33222
rect 7946 33216 8262 33217
rect 7946 33152 7952 33216
rect 8016 33152 8032 33216
rect 8096 33152 8112 33216
rect 8176 33152 8192 33216
rect 8256 33152 8262 33216
rect 11130 33192 11250 33222
rect 7946 33151 8262 33152
rect 2884 33086 4170 33146
rect 2884 33084 2890 33086
rect 3918 32948 3924 33012
rect 3988 33010 3994 33012
rect 5993 33010 6059 33013
rect 3988 33008 6059 33010
rect 3988 32952 5998 33008
rect 6054 32952 6059 33008
rect 3988 32950 6059 32952
rect 3988 32948 3994 32950
rect 5993 32947 6059 32950
rect 7833 33010 7899 33013
rect 8518 33010 8524 33012
rect 7833 33008 8524 33010
rect 7833 32952 7838 33008
rect 7894 32952 8524 33008
rect 7833 32950 8524 32952
rect 7833 32947 7899 32950
rect 8518 32948 8524 32950
rect 8588 32948 8594 33012
rect 10685 33010 10751 33013
rect 11130 33010 11250 33040
rect 10685 33008 11250 33010
rect 10685 32952 10690 33008
rect 10746 32952 11250 33008
rect 10685 32950 11250 32952
rect 10685 32947 10751 32950
rect 11130 32920 11250 32950
rect 1669 32876 1735 32877
rect 1669 32874 1716 32876
rect 1624 32872 1716 32874
rect 1624 32816 1674 32872
rect 1624 32814 1716 32816
rect 1669 32812 1716 32814
rect 1780 32812 1786 32876
rect 5758 32812 5764 32876
rect 5828 32874 5834 32876
rect 6729 32874 6795 32877
rect 5828 32872 6795 32874
rect 5828 32816 6734 32872
rect 6790 32816 6795 32872
rect 5828 32814 6795 32816
rect 5828 32812 5834 32814
rect 1669 32811 1735 32812
rect 6729 32811 6795 32814
rect 0 32738 120 32768
rect 749 32738 815 32741
rect 0 32736 815 32738
rect 0 32680 754 32736
rect 810 32680 815 32736
rect 0 32678 815 32680
rect 0 32648 120 32678
rect 749 32675 815 32678
rect 7782 32676 7788 32740
rect 7852 32738 7858 32740
rect 8845 32738 8911 32741
rect 7852 32736 8911 32738
rect 7852 32680 8850 32736
rect 8906 32680 8911 32736
rect 7852 32678 8911 32680
rect 7852 32676 7858 32678
rect 8845 32675 8911 32678
rect 9673 32738 9739 32741
rect 11130 32738 11250 32768
rect 9673 32736 11250 32738
rect 9673 32680 9678 32736
rect 9734 32680 11250 32736
rect 9673 32678 11250 32680
rect 9673 32675 9739 32678
rect 3006 32672 3322 32673
rect 3006 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3322 32672
rect 3006 32607 3322 32608
rect 9006 32672 9322 32673
rect 9006 32608 9012 32672
rect 9076 32608 9092 32672
rect 9156 32608 9172 32672
rect 9236 32608 9252 32672
rect 9316 32608 9322 32672
rect 11130 32648 11250 32678
rect 9006 32607 9322 32608
rect 10225 32466 10291 32469
rect 11130 32466 11250 32496
rect 10225 32464 11250 32466
rect 10225 32408 10230 32464
rect 10286 32408 11250 32464
rect 10225 32406 11250 32408
rect 10225 32403 10291 32406
rect 11130 32376 11250 32406
rect 7097 32330 7163 32333
rect 7598 32330 7604 32332
rect 7097 32328 7604 32330
rect 7097 32272 7102 32328
rect 7158 32272 7604 32328
rect 7097 32270 7604 32272
rect 7097 32267 7163 32270
rect 7598 32268 7604 32270
rect 7668 32268 7674 32332
rect 10225 32194 10291 32197
rect 11130 32194 11250 32224
rect 10225 32192 11250 32194
rect 10225 32136 10230 32192
rect 10286 32136 11250 32192
rect 10225 32134 11250 32136
rect 10225 32131 10291 32134
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 7946 32128 8262 32129
rect 7946 32064 7952 32128
rect 8016 32064 8032 32128
rect 8096 32064 8112 32128
rect 8176 32064 8192 32128
rect 8256 32064 8262 32128
rect 11130 32104 11250 32134
rect 7946 32063 8262 32064
rect 7005 32058 7071 32061
rect 7373 32058 7439 32061
rect 7005 32056 7439 32058
rect 7005 32000 7010 32056
rect 7066 32000 7378 32056
rect 7434 32000 7439 32056
rect 7005 31998 7439 32000
rect 7005 31995 7071 31998
rect 7373 31995 7439 31998
rect 0 31922 120 31952
rect 1485 31922 1551 31925
rect 0 31920 1551 31922
rect 0 31864 1490 31920
rect 1546 31864 1551 31920
rect 0 31862 1551 31864
rect 0 31832 120 31862
rect 1485 31859 1551 31862
rect 2037 31922 2103 31925
rect 2630 31922 2636 31924
rect 2037 31920 2636 31922
rect 2037 31864 2042 31920
rect 2098 31864 2636 31920
rect 2037 31862 2636 31864
rect 2037 31859 2103 31862
rect 2630 31860 2636 31862
rect 2700 31860 2706 31924
rect 4337 31922 4403 31925
rect 4797 31922 4863 31925
rect 4337 31920 4863 31922
rect 4337 31864 4342 31920
rect 4398 31864 4802 31920
rect 4858 31864 4863 31920
rect 4337 31862 4863 31864
rect 4337 31859 4403 31862
rect 4797 31859 4863 31862
rect 10409 31922 10475 31925
rect 11130 31922 11250 31952
rect 10409 31920 11250 31922
rect 10409 31864 10414 31920
rect 10470 31864 11250 31920
rect 10409 31862 11250 31864
rect 10409 31859 10475 31862
rect 11130 31832 11250 31862
rect 197 31786 263 31789
rect 4521 31786 4587 31789
rect 197 31784 306 31786
rect 197 31728 202 31784
rect 258 31728 306 31784
rect 197 31723 306 31728
rect 246 31652 306 31723
rect 4478 31784 4587 31786
rect 4478 31728 4526 31784
rect 4582 31728 4587 31784
rect 4478 31723 4587 31728
rect 5441 31784 5507 31789
rect 5441 31728 5446 31784
rect 5502 31728 5507 31784
rect 5441 31723 5507 31728
rect 5993 31786 6059 31789
rect 7189 31788 7255 31789
rect 6126 31786 6132 31788
rect 5993 31784 6132 31786
rect 5993 31728 5998 31784
rect 6054 31728 6132 31784
rect 5993 31726 6132 31728
rect 5993 31723 6059 31726
rect 6126 31724 6132 31726
rect 6196 31724 6202 31788
rect 7189 31784 7236 31788
rect 7300 31786 7306 31788
rect 9397 31786 9463 31789
rect 7189 31728 7194 31784
rect 7189 31724 7236 31728
rect 7300 31726 7346 31786
rect 9397 31784 9690 31786
rect 9397 31728 9402 31784
rect 9458 31728 9690 31784
rect 9397 31726 9690 31728
rect 7300 31724 7306 31726
rect 7189 31723 7255 31724
rect 9397 31723 9463 31726
rect 238 31588 244 31652
rect 308 31588 314 31652
rect 4337 31650 4403 31653
rect 4478 31650 4538 31723
rect 4337 31648 4538 31650
rect 4337 31592 4342 31648
rect 4398 31592 4538 31648
rect 4337 31590 4538 31592
rect 4981 31650 5047 31653
rect 5444 31650 5504 31723
rect 4981 31648 5504 31650
rect 4981 31592 4986 31648
rect 5042 31592 5504 31648
rect 4981 31590 5504 31592
rect 9630 31650 9690 31726
rect 11130 31650 11250 31680
rect 9630 31590 11250 31650
rect 4337 31587 4403 31590
rect 4981 31587 5047 31590
rect 3006 31584 3322 31585
rect 3006 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3322 31584
rect 3006 31519 3322 31520
rect 9006 31584 9322 31585
rect 9006 31520 9012 31584
rect 9076 31520 9092 31584
rect 9156 31520 9172 31584
rect 9236 31520 9252 31584
rect 9316 31520 9322 31584
rect 11130 31560 11250 31590
rect 9006 31519 9322 31520
rect 4286 31452 4292 31516
rect 4356 31514 4362 31516
rect 5257 31514 5323 31517
rect 4356 31512 5323 31514
rect 4356 31456 5262 31512
rect 5318 31456 5323 31512
rect 4356 31454 5323 31456
rect 4356 31452 4362 31454
rect 5257 31451 5323 31454
rect 7230 31452 7236 31516
rect 7300 31514 7306 31516
rect 8518 31514 8524 31516
rect 7300 31454 8524 31514
rect 7300 31452 7306 31454
rect 8518 31452 8524 31454
rect 8588 31452 8594 31516
rect 4838 31316 4844 31380
rect 4908 31378 4914 31380
rect 8385 31378 8451 31381
rect 4908 31376 8451 31378
rect 4908 31320 8390 31376
rect 8446 31320 8451 31376
rect 4908 31318 8451 31320
rect 4908 31316 4914 31318
rect 8385 31315 8451 31318
rect 8569 31378 8635 31381
rect 9029 31378 9095 31381
rect 8569 31376 9095 31378
rect 8569 31320 8574 31376
rect 8630 31320 9034 31376
rect 9090 31320 9095 31376
rect 8569 31318 9095 31320
rect 8569 31315 8635 31318
rect 9029 31315 9095 31318
rect 9673 31378 9739 31381
rect 11130 31378 11250 31408
rect 9673 31376 11250 31378
rect 9673 31320 9678 31376
rect 9734 31320 11250 31376
rect 9673 31318 11250 31320
rect 9673 31315 9739 31318
rect 11130 31288 11250 31318
rect 2221 31242 2287 31245
rect 4245 31242 4311 31245
rect 8661 31242 8727 31245
rect 2221 31240 8727 31242
rect 2221 31184 2226 31240
rect 2282 31184 4250 31240
rect 4306 31184 8666 31240
rect 8722 31184 8727 31240
rect 2221 31182 8727 31184
rect 2221 31179 2287 31182
rect 4245 31179 4311 31182
rect 8661 31179 8727 31182
rect 0 31106 120 31136
rect 841 31106 907 31109
rect 0 31104 907 31106
rect 0 31048 846 31104
rect 902 31048 907 31104
rect 0 31046 907 31048
rect 0 31016 120 31046
rect 841 31043 907 31046
rect 9489 31106 9555 31109
rect 11130 31106 11250 31136
rect 9489 31104 11250 31106
rect 9489 31048 9494 31104
rect 9550 31048 11250 31104
rect 9489 31046 11250 31048
rect 9489 31043 9555 31046
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 7946 31040 8262 31041
rect 7946 30976 7952 31040
rect 8016 30976 8032 31040
rect 8096 30976 8112 31040
rect 8176 30976 8192 31040
rect 8256 30976 8262 31040
rect 11130 31016 11250 31046
rect 7946 30975 8262 30976
rect 8661 30970 8727 30973
rect 9622 30970 9628 30972
rect 8661 30968 9628 30970
rect 8661 30912 8666 30968
rect 8722 30912 9628 30968
rect 8661 30910 9628 30912
rect 8661 30907 8727 30910
rect 9622 30908 9628 30910
rect 9692 30908 9698 30972
rect 9581 30834 9647 30837
rect 11130 30834 11250 30864
rect 9581 30832 11250 30834
rect 9581 30776 9586 30832
rect 9642 30776 11250 30832
rect 9581 30774 11250 30776
rect 9581 30771 9647 30774
rect 11130 30744 11250 30774
rect 3785 30562 3851 30565
rect 5574 30562 5580 30564
rect 3785 30560 5580 30562
rect 3785 30504 3790 30560
rect 3846 30504 5580 30560
rect 3785 30502 5580 30504
rect 3785 30499 3851 30502
rect 5574 30500 5580 30502
rect 5644 30500 5650 30564
rect 9673 30562 9739 30565
rect 11130 30562 11250 30592
rect 9673 30560 11250 30562
rect 9673 30504 9678 30560
rect 9734 30504 11250 30560
rect 9673 30502 11250 30504
rect 9673 30499 9739 30502
rect 3006 30496 3322 30497
rect 3006 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3322 30496
rect 3006 30431 3322 30432
rect 9006 30496 9322 30497
rect 9006 30432 9012 30496
rect 9076 30432 9092 30496
rect 9156 30432 9172 30496
rect 9236 30432 9252 30496
rect 9316 30432 9322 30496
rect 11130 30472 11250 30502
rect 9006 30431 9322 30432
rect 4061 30428 4127 30429
rect 2814 30426 2820 30428
rect 1350 30366 2820 30426
rect 0 30290 120 30320
rect 1350 30293 1410 30366
rect 2814 30364 2820 30366
rect 2884 30364 2890 30428
rect 4061 30424 4108 30428
rect 4172 30426 4178 30428
rect 6085 30426 6151 30429
rect 6494 30426 6500 30428
rect 4061 30368 4066 30424
rect 4061 30364 4108 30368
rect 4172 30366 4218 30426
rect 6085 30424 6500 30426
rect 6085 30368 6090 30424
rect 6146 30368 6500 30424
rect 6085 30366 6500 30368
rect 4172 30364 4178 30366
rect 4061 30363 4127 30364
rect 6085 30363 6151 30366
rect 6494 30364 6500 30366
rect 6564 30364 6570 30428
rect 8334 30364 8340 30428
rect 8404 30426 8410 30428
rect 8753 30426 8819 30429
rect 8404 30424 8819 30426
rect 8404 30368 8758 30424
rect 8814 30368 8819 30424
rect 8404 30366 8819 30368
rect 8404 30364 8410 30366
rect 8753 30363 8819 30366
rect 0 30230 858 30290
rect 0 30200 120 30230
rect 798 30154 858 30230
rect 1301 30288 1410 30293
rect 1301 30232 1306 30288
rect 1362 30232 1410 30288
rect 1301 30230 1410 30232
rect 1301 30227 1367 30230
rect 2446 30228 2452 30292
rect 2516 30290 2522 30292
rect 2773 30290 2839 30293
rect 2516 30288 2839 30290
rect 2516 30232 2778 30288
rect 2834 30232 2839 30288
rect 2516 30230 2839 30232
rect 2516 30228 2522 30230
rect 2773 30227 2839 30230
rect 3693 30290 3759 30293
rect 4286 30290 4292 30292
rect 3693 30288 4292 30290
rect 3693 30232 3698 30288
rect 3754 30232 4292 30288
rect 3693 30230 4292 30232
rect 3693 30227 3759 30230
rect 4286 30228 4292 30230
rect 4356 30228 4362 30292
rect 4797 30290 4863 30293
rect 7046 30290 7052 30292
rect 4797 30288 7052 30290
rect 4797 30232 4802 30288
rect 4858 30232 7052 30288
rect 4797 30230 7052 30232
rect 4797 30227 4863 30230
rect 7046 30228 7052 30230
rect 7116 30228 7122 30292
rect 7189 30288 7255 30293
rect 7189 30232 7194 30288
rect 7250 30232 7255 30288
rect 7189 30227 7255 30232
rect 9949 30290 10015 30293
rect 11130 30290 11250 30320
rect 9949 30288 11250 30290
rect 9949 30232 9954 30288
rect 10010 30232 11250 30288
rect 9949 30230 11250 30232
rect 9949 30227 10015 30230
rect 1485 30154 1551 30157
rect 3918 30154 3924 30156
rect 798 30152 1551 30154
rect 798 30096 1490 30152
rect 1546 30096 1551 30152
rect 798 30094 1551 30096
rect 1485 30091 1551 30094
rect 1718 30094 3924 30154
rect 841 30018 907 30021
rect 1718 30018 1778 30094
rect 3918 30092 3924 30094
rect 3988 30092 3994 30156
rect 7046 30092 7052 30156
rect 7116 30154 7122 30156
rect 7192 30154 7252 30227
rect 11130 30200 11250 30230
rect 7116 30094 7252 30154
rect 7116 30092 7122 30094
rect 841 30016 1778 30018
rect 841 29960 846 30016
rect 902 29960 1778 30016
rect 841 29958 1778 29960
rect 841 29955 907 29958
rect 4654 29956 4660 30020
rect 4724 30018 4730 30020
rect 4889 30018 4955 30021
rect 4724 30016 4955 30018
rect 4724 29960 4894 30016
rect 4950 29960 4955 30016
rect 4724 29958 4955 29960
rect 4724 29956 4730 29958
rect 4889 29955 4955 29958
rect 10225 30018 10291 30021
rect 11130 30018 11250 30048
rect 10225 30016 11250 30018
rect 10225 29960 10230 30016
rect 10286 29960 11250 30016
rect 10225 29958 11250 29960
rect 10225 29955 10291 29958
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 7946 29952 8262 29953
rect 7946 29888 7952 29952
rect 8016 29888 8032 29952
rect 8096 29888 8112 29952
rect 8176 29888 8192 29952
rect 8256 29888 8262 29952
rect 11130 29928 11250 29958
rect 7946 29887 8262 29888
rect 9489 29882 9555 29885
rect 9262 29880 9555 29882
rect 9262 29824 9494 29880
rect 9550 29824 9555 29880
rect 9262 29822 9555 29824
rect 7782 29746 7788 29748
rect 2730 29686 7788 29746
rect 2405 29610 2471 29613
rect 2730 29610 2790 29686
rect 7782 29684 7788 29686
rect 7852 29684 7858 29748
rect 8017 29746 8083 29749
rect 9029 29746 9095 29749
rect 8017 29744 9095 29746
rect 8017 29688 8022 29744
rect 8078 29688 9034 29744
rect 9090 29688 9095 29744
rect 8017 29686 9095 29688
rect 8017 29683 8083 29686
rect 9029 29683 9095 29686
rect 4705 29612 4771 29613
rect 2405 29608 2790 29610
rect 2405 29552 2410 29608
rect 2466 29552 2790 29608
rect 2405 29550 2790 29552
rect 2405 29547 2471 29550
rect 4654 29548 4660 29612
rect 4724 29610 4771 29612
rect 5441 29610 5507 29613
rect 4724 29608 5507 29610
rect 4766 29552 5446 29608
rect 5502 29552 5507 29608
rect 4724 29550 5507 29552
rect 4724 29548 4771 29550
rect 4705 29547 4771 29548
rect 5441 29547 5507 29550
rect 8661 29610 8727 29613
rect 9262 29610 9322 29822
rect 9489 29819 9555 29822
rect 9581 29746 9647 29749
rect 11130 29746 11250 29776
rect 9581 29744 11250 29746
rect 9581 29688 9586 29744
rect 9642 29688 11250 29744
rect 9581 29686 11250 29688
rect 9581 29683 9647 29686
rect 11130 29656 11250 29686
rect 8661 29608 9322 29610
rect 8661 29552 8666 29608
rect 8722 29552 9322 29608
rect 8661 29550 9322 29552
rect 8661 29547 8727 29550
rect 0 29474 120 29504
rect 1393 29474 1459 29477
rect 0 29472 1459 29474
rect 0 29416 1398 29472
rect 1454 29416 1459 29472
rect 0 29414 1459 29416
rect 0 29384 120 29414
rect 1393 29411 1459 29414
rect 4705 29474 4771 29477
rect 5022 29474 5028 29476
rect 4705 29472 5028 29474
rect 4705 29416 4710 29472
rect 4766 29416 5028 29472
rect 4705 29414 5028 29416
rect 4705 29411 4771 29414
rect 5022 29412 5028 29414
rect 5092 29412 5098 29476
rect 9765 29474 9831 29477
rect 11130 29474 11250 29504
rect 9765 29472 11250 29474
rect 9765 29416 9770 29472
rect 9826 29416 11250 29472
rect 9765 29414 11250 29416
rect 9765 29411 9831 29414
rect 3006 29408 3322 29409
rect 3006 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3322 29408
rect 3006 29343 3322 29344
rect 9006 29408 9322 29409
rect 9006 29344 9012 29408
rect 9076 29344 9092 29408
rect 9156 29344 9172 29408
rect 9236 29344 9252 29408
rect 9316 29344 9322 29408
rect 11130 29384 11250 29414
rect 9006 29343 9322 29344
rect 6177 29338 6243 29341
rect 3558 29336 6243 29338
rect 3558 29280 6182 29336
rect 6238 29280 6243 29336
rect 3558 29278 6243 29280
rect 1393 29202 1459 29205
rect 1710 29202 1716 29204
rect 1393 29200 1716 29202
rect 1393 29144 1398 29200
rect 1454 29144 1716 29200
rect 1393 29142 1716 29144
rect 1393 29139 1459 29142
rect 1710 29140 1716 29142
rect 1780 29202 1786 29204
rect 3558 29202 3618 29278
rect 6177 29275 6243 29278
rect 6862 29276 6868 29340
rect 6932 29338 6938 29340
rect 8109 29338 8175 29341
rect 10409 29338 10475 29341
rect 6932 29336 8175 29338
rect 6932 29280 8114 29336
rect 8170 29280 8175 29336
rect 6932 29278 8175 29280
rect 6932 29276 6938 29278
rect 8109 29275 8175 29278
rect 9400 29336 10475 29338
rect 9400 29280 10414 29336
rect 10470 29280 10475 29336
rect 9400 29278 10475 29280
rect 1780 29142 3618 29202
rect 4153 29202 4219 29205
rect 5533 29202 5599 29205
rect 9400 29202 9460 29278
rect 10409 29275 10475 29278
rect 4153 29200 5274 29202
rect 4153 29144 4158 29200
rect 4214 29144 5274 29200
rect 4153 29142 5274 29144
rect 1780 29140 1786 29142
rect 4153 29139 4219 29142
rect 657 29066 723 29069
rect 841 29066 907 29069
rect 657 29064 907 29066
rect 657 29008 662 29064
rect 718 29008 846 29064
rect 902 29008 907 29064
rect 657 29006 907 29008
rect 657 29003 723 29006
rect 841 29003 907 29006
rect 2681 29066 2747 29069
rect 3417 29066 3483 29069
rect 2681 29064 3483 29066
rect 2681 29008 2686 29064
rect 2742 29008 3422 29064
rect 3478 29008 3483 29064
rect 2681 29006 3483 29008
rect 2681 29003 2747 29006
rect 3417 29003 3483 29006
rect 4245 29064 4311 29069
rect 4245 29008 4250 29064
rect 4306 29008 4311 29064
rect 4245 29003 4311 29008
rect 1669 28932 1735 28933
rect 1669 28930 1716 28932
rect 1624 28928 1716 28930
rect 1624 28872 1674 28928
rect 1624 28870 1716 28872
rect 1669 28868 1716 28870
rect 1780 28868 1786 28932
rect 1669 28867 1735 28868
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 0 28658 120 28688
rect 381 28658 447 28661
rect 0 28656 447 28658
rect 0 28600 386 28656
rect 442 28600 447 28656
rect 0 28598 447 28600
rect 0 28568 120 28598
rect 381 28595 447 28598
rect 1158 28596 1164 28660
rect 1228 28658 1234 28660
rect 3785 28658 3851 28661
rect 1228 28656 3851 28658
rect 1228 28600 3790 28656
rect 3846 28600 3851 28656
rect 1228 28598 3851 28600
rect 1228 28596 1234 28598
rect 3785 28595 3851 28598
rect 1342 28460 1348 28524
rect 1412 28522 1418 28524
rect 2865 28522 2931 28525
rect 1412 28520 2931 28522
rect 1412 28464 2870 28520
rect 2926 28464 2931 28520
rect 1412 28462 2931 28464
rect 1412 28460 1418 28462
rect 2865 28459 2931 28462
rect 3006 28320 3322 28321
rect 3006 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3322 28320
rect 3006 28255 3322 28256
rect 13 28114 79 28117
rect 2630 28114 2636 28116
rect 13 28112 2636 28114
rect 13 28056 18 28112
rect 74 28056 2636 28112
rect 13 28054 2636 28056
rect 13 28051 79 28054
rect 2630 28052 2636 28054
rect 2700 28052 2706 28116
rect 2129 27978 2195 27981
rect 2630 27978 2636 27980
rect 2129 27976 2636 27978
rect 2129 27920 2134 27976
rect 2190 27920 2636 27976
rect 2129 27918 2636 27920
rect 2129 27915 2195 27918
rect 2630 27916 2636 27918
rect 2700 27916 2706 27980
rect 0 27842 120 27872
rect 1393 27842 1459 27845
rect 0 27840 1459 27842
rect 0 27784 1398 27840
rect 1454 27784 1459 27840
rect 0 27782 1459 27784
rect 0 27752 120 27782
rect 1393 27779 1459 27782
rect 3049 27842 3115 27845
rect 4248 27842 4308 29003
rect 5214 28930 5274 29142
rect 5533 29200 9460 29202
rect 5533 29144 5538 29200
rect 5594 29144 9460 29200
rect 5533 29142 9460 29144
rect 9581 29202 9647 29205
rect 9949 29202 10015 29205
rect 11130 29202 11250 29232
rect 9581 29200 9690 29202
rect 9581 29144 9586 29200
rect 9642 29144 9690 29200
rect 5533 29139 5599 29142
rect 9581 29139 9690 29144
rect 9949 29200 11250 29202
rect 9949 29144 9954 29200
rect 10010 29144 11250 29200
rect 9949 29142 11250 29144
rect 9949 29139 10015 29142
rect 8661 29066 8727 29069
rect 8937 29066 9003 29069
rect 8661 29064 9003 29066
rect 8661 29008 8666 29064
rect 8722 29008 8942 29064
rect 8998 29008 9003 29064
rect 8661 29006 9003 29008
rect 8661 29003 8727 29006
rect 8937 29003 9003 29006
rect 6453 28930 6519 28933
rect 5214 28928 6519 28930
rect 5214 28872 6458 28928
rect 6514 28872 6519 28928
rect 5214 28870 6519 28872
rect 6453 28867 6519 28870
rect 7946 28864 8262 28865
rect 7946 28800 7952 28864
rect 8016 28800 8032 28864
rect 8096 28800 8112 28864
rect 8176 28800 8192 28864
rect 8256 28800 8262 28864
rect 7946 28799 8262 28800
rect 9630 28794 9690 29139
rect 11130 29112 11250 29142
rect 10317 28930 10383 28933
rect 11130 28930 11250 28960
rect 10317 28928 11250 28930
rect 10317 28872 10322 28928
rect 10378 28872 11250 28928
rect 10317 28870 11250 28872
rect 10317 28867 10383 28870
rect 11130 28840 11250 28870
rect 10910 28794 10916 28796
rect 9630 28734 10916 28794
rect 10910 28732 10916 28734
rect 10980 28732 10986 28796
rect 6545 28660 6611 28661
rect 6494 28596 6500 28660
rect 6564 28658 6611 28660
rect 7189 28660 7255 28661
rect 6564 28656 6656 28658
rect 6606 28600 6656 28656
rect 6564 28598 6656 28600
rect 7189 28656 7236 28660
rect 7300 28658 7306 28660
rect 7189 28600 7194 28656
rect 6564 28596 6611 28598
rect 6545 28595 6611 28596
rect 7189 28596 7236 28600
rect 7300 28598 7346 28658
rect 7300 28596 7306 28598
rect 8334 28596 8340 28660
rect 8404 28658 8410 28660
rect 8937 28658 9003 28661
rect 8404 28656 9003 28658
rect 8404 28600 8942 28656
rect 8998 28600 9003 28656
rect 8404 28598 9003 28600
rect 8404 28596 8410 28598
rect 7189 28595 7255 28596
rect 8937 28595 9003 28598
rect 10593 28658 10659 28661
rect 11130 28658 11250 28688
rect 10593 28656 11250 28658
rect 10593 28600 10598 28656
rect 10654 28600 11250 28656
rect 10593 28598 11250 28600
rect 10593 28595 10659 28598
rect 11130 28568 11250 28598
rect 6678 28460 6684 28524
rect 6748 28522 6754 28524
rect 9213 28522 9279 28525
rect 6748 28520 9279 28522
rect 6748 28464 9218 28520
rect 9274 28464 9279 28520
rect 6748 28462 9279 28464
rect 6748 28460 6754 28462
rect 9213 28459 9279 28462
rect 4797 28386 4863 28389
rect 7097 28386 7163 28389
rect 4797 28384 7163 28386
rect 4797 28328 4802 28384
rect 4858 28328 7102 28384
rect 7158 28328 7163 28384
rect 4797 28326 7163 28328
rect 4797 28323 4863 28326
rect 7097 28323 7163 28326
rect 9581 28386 9647 28389
rect 11130 28386 11250 28416
rect 9581 28384 11250 28386
rect 9581 28328 9586 28384
rect 9642 28328 11250 28384
rect 9581 28326 11250 28328
rect 9581 28323 9647 28326
rect 9006 28320 9322 28321
rect 9006 28256 9012 28320
rect 9076 28256 9092 28320
rect 9156 28256 9172 28320
rect 9236 28256 9252 28320
rect 9316 28256 9322 28320
rect 11130 28296 11250 28326
rect 9006 28255 9322 28256
rect 7414 28188 7420 28252
rect 7484 28250 7490 28252
rect 8109 28250 8175 28253
rect 7484 28248 8175 28250
rect 7484 28192 8114 28248
rect 8170 28192 8175 28248
rect 7484 28190 8175 28192
rect 7484 28188 7490 28190
rect 8109 28187 8175 28190
rect 9489 28116 9555 28117
rect 9438 28114 9444 28116
rect 9398 28054 9444 28114
rect 9508 28112 9555 28116
rect 9550 28056 9555 28112
rect 9438 28052 9444 28054
rect 9508 28052 9555 28056
rect 9489 28051 9555 28052
rect 9673 28114 9739 28117
rect 11130 28114 11250 28144
rect 9673 28112 11250 28114
rect 9673 28056 9678 28112
rect 9734 28056 11250 28112
rect 9673 28054 11250 28056
rect 9673 28051 9739 28054
rect 11130 28024 11250 28054
rect 5533 27980 5599 27981
rect 5533 27976 5580 27980
rect 5644 27978 5650 27980
rect 5533 27920 5538 27976
rect 5533 27916 5580 27920
rect 5644 27918 5690 27978
rect 5644 27916 5650 27918
rect 7782 27916 7788 27980
rect 7852 27978 7858 27980
rect 9622 27978 9628 27980
rect 7852 27918 9628 27978
rect 7852 27916 7858 27918
rect 9622 27916 9628 27918
rect 9692 27916 9698 27980
rect 5533 27915 5599 27916
rect 7230 27842 7236 27844
rect 3049 27840 7236 27842
rect 3049 27784 3054 27840
rect 3110 27784 7236 27840
rect 3049 27782 7236 27784
rect 3049 27779 3115 27782
rect 7230 27780 7236 27782
rect 7300 27780 7306 27844
rect 10225 27842 10291 27845
rect 11130 27842 11250 27872
rect 10225 27840 11250 27842
rect 10225 27784 10230 27840
rect 10286 27784 11250 27840
rect 10225 27782 11250 27784
rect 10225 27779 10291 27782
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 7946 27776 8262 27777
rect 7946 27712 7952 27776
rect 8016 27712 8032 27776
rect 8096 27712 8112 27776
rect 8176 27712 8192 27776
rect 8256 27712 8262 27776
rect 11130 27752 11250 27782
rect 7946 27711 8262 27712
rect 3918 27644 3924 27708
rect 3988 27706 3994 27708
rect 4061 27706 4127 27709
rect 3988 27704 4127 27706
rect 3988 27648 4066 27704
rect 4122 27648 4127 27704
rect 3988 27646 4127 27648
rect 3988 27644 3994 27646
rect 4061 27643 4127 27646
rect 9397 27708 9463 27709
rect 9397 27704 9444 27708
rect 9508 27706 9514 27708
rect 9397 27648 9402 27704
rect 9397 27644 9444 27648
rect 9508 27646 9554 27706
rect 9508 27644 9514 27646
rect 9397 27643 9463 27644
rect 1853 27570 1919 27573
rect 3734 27570 3740 27572
rect 1853 27568 3740 27570
rect 1853 27512 1858 27568
rect 1914 27512 3740 27568
rect 1853 27510 3740 27512
rect 1853 27507 1919 27510
rect 3734 27508 3740 27510
rect 3804 27508 3810 27572
rect 4153 27570 4219 27573
rect 6913 27570 6979 27573
rect 8753 27572 8819 27573
rect 4153 27568 6979 27570
rect 4153 27512 4158 27568
rect 4214 27512 6918 27568
rect 6974 27512 6979 27568
rect 4153 27510 6979 27512
rect 4153 27507 4219 27510
rect 6913 27507 6979 27510
rect 8702 27508 8708 27572
rect 8772 27570 8819 27572
rect 10409 27570 10475 27573
rect 11130 27570 11250 27600
rect 8772 27568 8864 27570
rect 8814 27512 8864 27568
rect 8772 27510 8864 27512
rect 10409 27568 11250 27570
rect 10409 27512 10414 27568
rect 10470 27512 11250 27568
rect 10409 27510 11250 27512
rect 8772 27508 8819 27510
rect 8753 27507 8819 27508
rect 10409 27507 10475 27510
rect 11130 27480 11250 27510
rect 1485 27434 1551 27437
rect 2814 27434 2820 27436
rect 1485 27432 2820 27434
rect 1485 27376 1490 27432
rect 1546 27376 2820 27432
rect 1485 27374 2820 27376
rect 1485 27371 1551 27374
rect 2814 27372 2820 27374
rect 2884 27372 2890 27436
rect 5022 27372 5028 27436
rect 5092 27434 5098 27436
rect 6269 27434 6335 27437
rect 5092 27432 6335 27434
rect 5092 27376 6274 27432
rect 6330 27376 6335 27432
rect 5092 27374 6335 27376
rect 5092 27372 5098 27374
rect 6269 27371 6335 27374
rect 8518 27372 8524 27436
rect 8588 27434 8594 27436
rect 9121 27434 9187 27437
rect 8588 27432 9187 27434
rect 8588 27376 9126 27432
rect 9182 27376 9187 27432
rect 8588 27374 9187 27376
rect 8588 27372 8594 27374
rect 9121 27371 9187 27374
rect 9673 27298 9739 27301
rect 11130 27298 11250 27328
rect 9673 27296 11250 27298
rect 9673 27240 9678 27296
rect 9734 27240 11250 27296
rect 9673 27238 11250 27240
rect 9673 27235 9739 27238
rect 3006 27232 3322 27233
rect 3006 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3322 27232
rect 3006 27167 3322 27168
rect 9006 27232 9322 27233
rect 9006 27168 9012 27232
rect 9076 27168 9092 27232
rect 9156 27168 9172 27232
rect 9236 27168 9252 27232
rect 9316 27168 9322 27232
rect 11130 27208 11250 27238
rect 9006 27167 9322 27168
rect 0 27026 120 27056
rect 1393 27026 1459 27029
rect 3550 27026 3556 27028
rect 0 27024 1459 27026
rect 0 26968 1398 27024
rect 1454 26968 1459 27024
rect 0 26966 1459 26968
rect 0 26936 120 26966
rect 1393 26963 1459 26966
rect 2868 26966 3556 27026
rect 2868 26893 2928 26966
rect 3550 26964 3556 26966
rect 3620 26964 3626 27028
rect 10225 27026 10291 27029
rect 11130 27026 11250 27056
rect 10225 27024 11250 27026
rect 10225 26968 10230 27024
rect 10286 26968 11250 27024
rect 10225 26966 11250 26968
rect 10225 26963 10291 26966
rect 11130 26936 11250 26966
rect 1117 26890 1183 26893
rect 1117 26888 2744 26890
rect 1117 26832 1122 26888
rect 1178 26832 2744 26888
rect 1117 26830 2744 26832
rect 1117 26827 1183 26830
rect 2684 26754 2744 26830
rect 2865 26888 2931 26893
rect 2865 26832 2870 26888
rect 2926 26832 2931 26888
rect 2865 26827 2931 26832
rect 3550 26828 3556 26892
rect 3620 26890 3626 26892
rect 4102 26890 4108 26892
rect 3620 26830 4108 26890
rect 3620 26828 3626 26830
rect 4102 26828 4108 26830
rect 4172 26828 4178 26892
rect 8385 26890 8451 26893
rect 8702 26890 8708 26892
rect 8385 26888 8708 26890
rect 8385 26832 8390 26888
rect 8446 26832 8708 26888
rect 8385 26830 8708 26832
rect 8385 26827 8451 26830
rect 8702 26828 8708 26830
rect 8772 26828 8778 26892
rect 4429 26754 4495 26757
rect 2684 26752 4495 26754
rect 2684 26696 4434 26752
rect 4490 26696 4495 26752
rect 2684 26694 4495 26696
rect 4429 26691 4495 26694
rect 9305 26754 9371 26757
rect 11130 26754 11250 26784
rect 9305 26752 11250 26754
rect 9305 26696 9310 26752
rect 9366 26696 11250 26752
rect 9305 26694 11250 26696
rect 9305 26691 9371 26694
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 7946 26688 8262 26689
rect 7946 26624 7952 26688
rect 8016 26624 8032 26688
rect 8096 26624 8112 26688
rect 8176 26624 8192 26688
rect 8256 26624 8262 26688
rect 11130 26664 11250 26694
rect 7946 26623 8262 26624
rect 5625 26618 5691 26621
rect 6085 26618 6151 26621
rect 8477 26618 8543 26621
rect 8661 26618 8727 26621
rect 5625 26616 6010 26618
rect 5625 26560 5630 26616
rect 5686 26560 6010 26616
rect 5625 26558 6010 26560
rect 5625 26555 5691 26558
rect 422 26420 428 26484
rect 492 26482 498 26484
rect 657 26482 723 26485
rect 492 26480 723 26482
rect 492 26424 662 26480
rect 718 26424 723 26480
rect 492 26422 723 26424
rect 492 26420 498 26422
rect 657 26419 723 26422
rect 4889 26482 4955 26485
rect 5257 26482 5323 26485
rect 4889 26480 5323 26482
rect 4889 26424 4894 26480
rect 4950 26424 5262 26480
rect 5318 26424 5323 26480
rect 4889 26422 5323 26424
rect 4889 26419 4955 26422
rect 5257 26419 5323 26422
rect 1117 26346 1183 26349
rect 3877 26346 3943 26349
rect 1117 26344 3943 26346
rect 1117 26288 1122 26344
rect 1178 26288 3882 26344
rect 3938 26288 3943 26344
rect 1117 26286 3943 26288
rect 1117 26283 1183 26286
rect 3877 26283 3943 26286
rect 4429 26346 4495 26349
rect 5809 26346 5875 26349
rect 4429 26344 5875 26346
rect 4429 26288 4434 26344
rect 4490 26288 5814 26344
rect 5870 26288 5875 26344
rect 4429 26286 5875 26288
rect 4429 26283 4495 26286
rect 5809 26283 5875 26286
rect 0 26210 120 26240
rect 657 26210 723 26213
rect 0 26208 723 26210
rect 0 26152 662 26208
rect 718 26152 723 26208
rect 0 26150 723 26152
rect 0 26120 120 26150
rect 657 26147 723 26150
rect 5625 26210 5691 26213
rect 5950 26210 6010 26558
rect 6085 26616 6194 26618
rect 6085 26560 6090 26616
rect 6146 26560 6194 26616
rect 6085 26555 6194 26560
rect 8477 26616 8727 26618
rect 8477 26560 8482 26616
rect 8538 26560 8666 26616
rect 8722 26560 8727 26616
rect 8477 26558 8727 26560
rect 8477 26555 8543 26558
rect 8661 26555 8727 26558
rect 5625 26208 6010 26210
rect 5625 26152 5630 26208
rect 5686 26152 6010 26208
rect 5625 26150 6010 26152
rect 6134 26213 6194 26555
rect 10777 26482 10843 26485
rect 11130 26482 11250 26512
rect 10777 26480 11250 26482
rect 10777 26424 10782 26480
rect 10838 26424 11250 26480
rect 10777 26422 11250 26424
rect 10777 26419 10843 26422
rect 11130 26392 11250 26422
rect 8334 26284 8340 26348
rect 8404 26346 8410 26348
rect 9489 26346 9555 26349
rect 8404 26344 9555 26346
rect 8404 26288 9494 26344
rect 9550 26288 9555 26344
rect 8404 26286 9555 26288
rect 8404 26284 8410 26286
rect 9489 26283 9555 26286
rect 6134 26208 6243 26213
rect 6134 26152 6182 26208
rect 6238 26152 6243 26208
rect 6134 26150 6243 26152
rect 5625 26147 5691 26150
rect 6177 26147 6243 26150
rect 8201 26210 8267 26213
rect 9949 26212 10015 26213
rect 9949 26210 9996 26212
rect 8201 26208 8540 26210
rect 8201 26152 8206 26208
rect 8262 26152 8540 26208
rect 8201 26150 8540 26152
rect 9904 26208 9996 26210
rect 9904 26152 9954 26208
rect 9904 26150 9996 26152
rect 8201 26147 8267 26150
rect 3006 26144 3322 26145
rect 3006 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3322 26144
rect 3006 26079 3322 26080
rect 3601 26074 3667 26077
rect 3734 26074 3740 26076
rect 3601 26072 3740 26074
rect 3601 26016 3606 26072
rect 3662 26016 3740 26072
rect 3601 26014 3740 26016
rect 3601 26011 3667 26014
rect 3734 26012 3740 26014
rect 3804 26012 3810 26076
rect 4337 26074 4403 26077
rect 4337 26072 8172 26074
rect 4337 26016 4342 26072
rect 4398 26016 8172 26072
rect 4337 26014 8172 26016
rect 4337 26011 4403 26014
rect 2681 25940 2747 25941
rect 2630 25938 2636 25940
rect 2590 25878 2636 25938
rect 2700 25936 2747 25940
rect 7097 25938 7163 25941
rect 2742 25880 2747 25936
rect 2630 25876 2636 25878
rect 2700 25876 2747 25880
rect 2681 25875 2747 25876
rect 2822 25936 7163 25938
rect 2822 25880 7102 25936
rect 7158 25880 7163 25936
rect 2822 25878 7163 25880
rect 197 25802 263 25805
rect 2822 25802 2882 25878
rect 7097 25875 7163 25878
rect 197 25800 2882 25802
rect 197 25744 202 25800
rect 258 25744 2882 25800
rect 197 25742 2882 25744
rect 197 25739 263 25742
rect 7046 25740 7052 25804
rect 7116 25802 7122 25804
rect 7925 25802 7991 25805
rect 7116 25800 7991 25802
rect 7116 25744 7930 25800
rect 7986 25744 7991 25800
rect 7116 25742 7991 25744
rect 8112 25802 8172 26014
rect 8480 25938 8540 26150
rect 9949 26148 9996 26150
rect 10060 26148 10066 26212
rect 10317 26210 10383 26213
rect 11130 26210 11250 26240
rect 10317 26208 11250 26210
rect 10317 26152 10322 26208
rect 10378 26152 11250 26208
rect 10317 26150 11250 26152
rect 9949 26147 10015 26148
rect 10317 26147 10383 26150
rect 9006 26144 9322 26145
rect 9006 26080 9012 26144
rect 9076 26080 9092 26144
rect 9156 26080 9172 26144
rect 9236 26080 9252 26144
rect 9316 26080 9322 26144
rect 11130 26120 11250 26150
rect 9006 26079 9322 26080
rect 9622 26012 9628 26076
rect 9692 26074 9698 26076
rect 10041 26074 10107 26077
rect 9692 26072 10107 26074
rect 9692 26016 10046 26072
rect 10102 26016 10107 26072
rect 9692 26014 10107 26016
rect 9692 26012 9698 26014
rect 10041 26011 10107 26014
rect 8845 25938 8911 25941
rect 8480 25936 8911 25938
rect 8480 25880 8850 25936
rect 8906 25880 8911 25936
rect 8480 25878 8911 25880
rect 8845 25875 8911 25878
rect 9673 25938 9739 25941
rect 11130 25938 11250 25968
rect 9673 25936 11250 25938
rect 9673 25880 9678 25936
rect 9734 25880 11250 25936
rect 9673 25878 11250 25880
rect 9673 25875 9739 25878
rect 11130 25848 11250 25878
rect 10726 25802 10732 25804
rect 8112 25742 10732 25802
rect 7116 25740 7122 25742
rect 7925 25739 7991 25742
rect 10726 25740 10732 25742
rect 10796 25740 10802 25804
rect 10225 25666 10291 25669
rect 11130 25666 11250 25696
rect 10225 25664 11250 25666
rect 10225 25608 10230 25664
rect 10286 25608 11250 25664
rect 10225 25606 11250 25608
rect 10225 25603 10291 25606
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 7946 25600 8262 25601
rect 7946 25536 7952 25600
rect 8016 25536 8032 25600
rect 8096 25536 8112 25600
rect 8176 25536 8192 25600
rect 8256 25536 8262 25600
rect 11130 25576 11250 25606
rect 7946 25535 8262 25536
rect 2497 25530 2563 25533
rect 4102 25530 4108 25532
rect 2497 25528 4108 25530
rect 2497 25472 2502 25528
rect 2558 25472 4108 25528
rect 2497 25470 4108 25472
rect 2497 25467 2563 25470
rect 4102 25468 4108 25470
rect 4172 25468 4178 25532
rect 0 25394 120 25424
rect 1393 25394 1459 25397
rect 0 25392 1459 25394
rect 0 25336 1398 25392
rect 1454 25336 1459 25392
rect 0 25334 1459 25336
rect 0 25304 120 25334
rect 1393 25331 1459 25334
rect 2630 25332 2636 25396
rect 2700 25394 2706 25396
rect 5533 25394 5599 25397
rect 2700 25392 5599 25394
rect 2700 25336 5538 25392
rect 5594 25336 5599 25392
rect 2700 25334 5599 25336
rect 2700 25332 2706 25334
rect 5533 25331 5599 25334
rect 6269 25394 6335 25397
rect 6494 25394 6500 25396
rect 6269 25392 6500 25394
rect 6269 25336 6274 25392
rect 6330 25336 6500 25392
rect 6269 25334 6500 25336
rect 6269 25331 6335 25334
rect 6494 25332 6500 25334
rect 6564 25394 6570 25396
rect 8017 25394 8083 25397
rect 6564 25392 8083 25394
rect 6564 25336 8022 25392
rect 8078 25336 8083 25392
rect 6564 25334 8083 25336
rect 6564 25332 6570 25334
rect 8017 25331 8083 25334
rect 9581 25394 9647 25397
rect 11130 25394 11250 25424
rect 9581 25392 11250 25394
rect 9581 25336 9586 25392
rect 9642 25336 11250 25392
rect 9581 25334 11250 25336
rect 9581 25331 9647 25334
rect 11130 25304 11250 25334
rect 5257 25122 5323 25125
rect 7414 25122 7420 25124
rect 5257 25120 7420 25122
rect 5257 25064 5262 25120
rect 5318 25064 7420 25120
rect 5257 25062 7420 25064
rect 5257 25059 5323 25062
rect 7414 25060 7420 25062
rect 7484 25060 7490 25124
rect 9673 25122 9739 25125
rect 11130 25122 11250 25152
rect 9673 25120 11250 25122
rect 9673 25064 9678 25120
rect 9734 25064 11250 25120
rect 9673 25062 11250 25064
rect 9673 25059 9739 25062
rect 3006 25056 3322 25057
rect 3006 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3322 25056
rect 3006 24991 3322 24992
rect 9006 25056 9322 25057
rect 9006 24992 9012 25056
rect 9076 24992 9092 25056
rect 9156 24992 9172 25056
rect 9236 24992 9252 25056
rect 9316 24992 9322 25056
rect 11130 25032 11250 25062
rect 9006 24991 9322 24992
rect 238 24924 244 24988
rect 308 24986 314 24988
rect 381 24986 447 24989
rect 308 24984 447 24986
rect 308 24928 386 24984
rect 442 24928 447 24984
rect 308 24926 447 24928
rect 308 24924 314 24926
rect 381 24923 447 24926
rect 5022 24924 5028 24988
rect 5092 24986 5098 24988
rect 5901 24986 5967 24989
rect 7097 24986 7163 24989
rect 5092 24984 5967 24986
rect 5092 24928 5906 24984
rect 5962 24928 5967 24984
rect 5092 24926 5967 24928
rect 5092 24924 5098 24926
rect 5901 24923 5967 24926
rect 7054 24984 7163 24986
rect 7054 24928 7102 24984
rect 7158 24928 7163 24984
rect 7054 24923 7163 24928
rect 7782 24924 7788 24988
rect 7852 24986 7858 24988
rect 7852 24926 8816 24986
rect 7852 24924 7858 24926
rect 5022 24788 5028 24852
rect 5092 24850 5098 24852
rect 6862 24850 6868 24852
rect 5092 24790 6868 24850
rect 5092 24788 5098 24790
rect 6862 24788 6868 24790
rect 6932 24788 6938 24852
rect 1526 24652 1532 24716
rect 1596 24714 1602 24716
rect 2129 24714 2195 24717
rect 1596 24712 2195 24714
rect 1596 24656 2134 24712
rect 2190 24656 2195 24712
rect 1596 24654 2195 24656
rect 1596 24652 1602 24654
rect 2129 24651 2195 24654
rect 6862 24652 6868 24716
rect 6932 24714 6938 24716
rect 7054 24714 7114 24923
rect 7414 24788 7420 24852
rect 7484 24850 7490 24852
rect 8201 24850 8267 24853
rect 7484 24848 8267 24850
rect 7484 24792 8206 24848
rect 8262 24792 8267 24848
rect 7484 24790 8267 24792
rect 8756 24850 8816 24926
rect 9305 24850 9371 24853
rect 8756 24848 9371 24850
rect 8756 24792 9310 24848
rect 9366 24792 9371 24848
rect 8756 24790 9371 24792
rect 7484 24788 7490 24790
rect 8201 24787 8267 24790
rect 9305 24787 9371 24790
rect 10225 24850 10291 24853
rect 11130 24850 11250 24880
rect 10225 24848 11250 24850
rect 10225 24792 10230 24848
rect 10286 24792 11250 24848
rect 10225 24790 11250 24792
rect 10225 24787 10291 24790
rect 11130 24760 11250 24790
rect 6932 24654 7114 24714
rect 7189 24714 7255 24717
rect 7782 24714 7788 24716
rect 7189 24712 7788 24714
rect 7189 24656 7194 24712
rect 7250 24656 7788 24712
rect 7189 24654 7788 24656
rect 6932 24652 6938 24654
rect 7189 24651 7255 24654
rect 7782 24652 7788 24654
rect 7852 24652 7858 24716
rect 0 24578 120 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 120 24518
rect 1393 24515 1459 24518
rect 9765 24578 9831 24581
rect 11130 24578 11250 24608
rect 9765 24576 11250 24578
rect 9765 24520 9770 24576
rect 9826 24520 11250 24576
rect 9765 24518 11250 24520
rect 9765 24515 9831 24518
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 7946 24512 8262 24513
rect 7946 24448 7952 24512
rect 8016 24448 8032 24512
rect 8096 24448 8112 24512
rect 8176 24448 8192 24512
rect 8256 24448 8262 24512
rect 11130 24488 11250 24518
rect 7946 24447 8262 24448
rect 2446 24380 2452 24444
rect 2516 24442 2522 24444
rect 2516 24382 7482 24442
rect 2516 24380 2522 24382
rect 7281 24306 7347 24309
rect 6916 24304 7347 24306
rect 6916 24248 7286 24304
rect 7342 24248 7347 24304
rect 6916 24246 7347 24248
rect 7422 24306 7482 24382
rect 9121 24306 9187 24309
rect 7422 24304 9187 24306
rect 7422 24248 9126 24304
rect 9182 24248 9187 24304
rect 7422 24246 9187 24248
rect 6916 24173 6976 24246
rect 7281 24243 7347 24246
rect 9121 24243 9187 24246
rect 9673 24306 9739 24309
rect 11130 24306 11250 24336
rect 9673 24304 11250 24306
rect 9673 24248 9678 24304
rect 9734 24248 11250 24304
rect 9673 24246 11250 24248
rect 9673 24243 9739 24246
rect 11130 24216 11250 24246
rect 2957 24170 3023 24173
rect 2822 24168 3023 24170
rect 2822 24112 2962 24168
rect 3018 24112 3023 24168
rect 2822 24110 3023 24112
rect 0 23762 120 23792
rect 1393 23762 1459 23765
rect 0 23760 1459 23762
rect 0 23704 1398 23760
rect 1454 23704 1459 23760
rect 0 23702 1459 23704
rect 2822 23762 2882 24110
rect 2957 24107 3023 24110
rect 3141 24170 3207 24173
rect 4429 24170 4495 24173
rect 3141 24168 3618 24170
rect 3141 24112 3146 24168
rect 3202 24112 3618 24168
rect 3141 24110 3618 24112
rect 3141 24107 3207 24110
rect 3006 23968 3322 23969
rect 3006 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3322 23968
rect 3006 23903 3322 23904
rect 2957 23762 3023 23765
rect 2822 23760 3023 23762
rect 2822 23704 2962 23760
rect 3018 23704 3023 23760
rect 2822 23702 3023 23704
rect 0 23672 120 23702
rect 1393 23699 1459 23702
rect 2957 23699 3023 23702
rect 3233 23762 3299 23765
rect 3558 23762 3618 24110
rect 4156 24168 4495 24170
rect 4156 24112 4434 24168
rect 4490 24112 4495 24168
rect 4156 24110 4495 24112
rect 4156 24037 4216 24110
rect 4429 24107 4495 24110
rect 6913 24168 6979 24173
rect 6913 24112 6918 24168
rect 6974 24112 6979 24168
rect 6913 24107 6979 24112
rect 4153 24032 4219 24037
rect 4153 23976 4158 24032
rect 4214 23976 4219 24032
rect 4153 23971 4219 23976
rect 10225 24034 10291 24037
rect 11130 24034 11250 24064
rect 10225 24032 11250 24034
rect 10225 23976 10230 24032
rect 10286 23976 11250 24032
rect 10225 23974 11250 23976
rect 10225 23971 10291 23974
rect 9006 23968 9322 23969
rect 9006 23904 9012 23968
rect 9076 23904 9092 23968
rect 9156 23904 9172 23968
rect 9236 23904 9252 23968
rect 9316 23904 9322 23968
rect 11130 23944 11250 23974
rect 9006 23903 9322 23904
rect 5390 23836 5396 23900
rect 5460 23898 5466 23900
rect 5901 23898 5967 23901
rect 5460 23896 5967 23898
rect 5460 23840 5906 23896
rect 5962 23840 5967 23896
rect 5460 23838 5967 23840
rect 5460 23836 5466 23838
rect 5901 23835 5967 23838
rect 8293 23898 8359 23901
rect 8518 23898 8524 23900
rect 8293 23896 8524 23898
rect 8293 23840 8298 23896
rect 8354 23840 8524 23896
rect 8293 23838 8524 23840
rect 8293 23835 8359 23838
rect 8518 23836 8524 23838
rect 8588 23836 8594 23900
rect 7925 23762 7991 23765
rect 8518 23762 8524 23764
rect 3233 23760 8524 23762
rect 3233 23704 3238 23760
rect 3294 23704 7930 23760
rect 7986 23704 8524 23760
rect 3233 23702 8524 23704
rect 3233 23699 3299 23702
rect 7925 23699 7991 23702
rect 8518 23700 8524 23702
rect 8588 23700 8594 23764
rect 9673 23762 9739 23765
rect 11130 23762 11250 23792
rect 9673 23760 11250 23762
rect 9673 23704 9678 23760
rect 9734 23704 11250 23760
rect 9673 23702 11250 23704
rect 9673 23699 9739 23702
rect 11130 23672 11250 23702
rect 8017 23626 8083 23629
rect 7468 23624 8083 23626
rect 7468 23568 8022 23624
rect 8078 23568 8083 23624
rect 7468 23566 8083 23568
rect 3877 23490 3943 23493
rect 4838 23490 4844 23492
rect 3877 23488 4844 23490
rect 3877 23432 3882 23488
rect 3938 23432 4844 23488
rect 3877 23430 4844 23432
rect 3877 23427 3943 23430
rect 4838 23428 4844 23430
rect 4908 23428 4914 23492
rect 7230 23428 7236 23492
rect 7300 23428 7306 23492
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 4286 23292 4292 23356
rect 4356 23354 4362 23356
rect 4521 23354 4587 23357
rect 4356 23352 4587 23354
rect 4356 23296 4526 23352
rect 4582 23296 4587 23352
rect 4356 23294 4587 23296
rect 4356 23292 4362 23294
rect 4521 23291 4587 23294
rect 13 23218 79 23221
rect 422 23218 428 23220
rect 13 23216 428 23218
rect 13 23160 18 23216
rect 74 23160 428 23216
rect 13 23158 428 23160
rect 13 23155 79 23158
rect 422 23156 428 23158
rect 492 23156 498 23220
rect 1945 23218 2011 23221
rect 2446 23218 2452 23220
rect 1945 23216 2452 23218
rect 1945 23160 1950 23216
rect 2006 23160 2452 23216
rect 1945 23158 2452 23160
rect 1945 23155 2011 23158
rect 2446 23156 2452 23158
rect 2516 23218 2522 23220
rect 2681 23218 2747 23221
rect 2516 23216 2747 23218
rect 2516 23160 2686 23216
rect 2742 23160 2747 23216
rect 2516 23158 2747 23160
rect 2516 23156 2522 23158
rect 2681 23155 2747 23158
rect 5390 23020 5396 23084
rect 5460 23082 5466 23084
rect 5993 23082 6059 23085
rect 5460 23080 6059 23082
rect 5460 23024 5998 23080
rect 6054 23024 6059 23080
rect 5460 23022 6059 23024
rect 5460 23020 5466 23022
rect 5993 23019 6059 23022
rect 6269 23080 6335 23085
rect 6269 23024 6274 23080
rect 6330 23024 6335 23080
rect 6269 23019 6335 23024
rect 7005 23082 7071 23085
rect 7238 23082 7298 23428
rect 7005 23080 7298 23082
rect 7005 23024 7010 23080
rect 7066 23024 7298 23080
rect 7005 23022 7298 23024
rect 7005 23019 7071 23022
rect 0 22946 120 22976
rect 1393 22946 1459 22949
rect 0 22944 1459 22946
rect 0 22888 1398 22944
rect 1454 22888 1459 22944
rect 0 22886 1459 22888
rect 6272 22946 6332 23019
rect 7281 22946 7347 22949
rect 6272 22944 7347 22946
rect 6272 22888 7286 22944
rect 7342 22888 7347 22944
rect 6272 22886 7347 22888
rect 0 22856 120 22886
rect 1393 22883 1459 22886
rect 7281 22883 7347 22886
rect 3006 22880 3322 22881
rect 3006 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3322 22880
rect 3006 22815 3322 22816
rect 4337 22810 4403 22813
rect 6269 22810 6335 22813
rect 4337 22808 6335 22810
rect 4337 22752 4342 22808
rect 4398 22752 6274 22808
rect 6330 22752 6335 22808
rect 4337 22750 6335 22752
rect 4337 22747 4403 22750
rect 6269 22747 6335 22750
rect 6494 22748 6500 22812
rect 6564 22810 6570 22812
rect 7005 22810 7071 22813
rect 6564 22808 7071 22810
rect 6564 22752 7010 22808
rect 7066 22752 7071 22808
rect 6564 22750 7071 22752
rect 6564 22748 6570 22750
rect 7005 22747 7071 22750
rect 3233 22674 3299 22677
rect 5574 22674 5580 22676
rect 3233 22672 5580 22674
rect 3233 22616 3238 22672
rect 3294 22616 5580 22672
rect 3233 22614 5580 22616
rect 3233 22611 3299 22614
rect 5574 22612 5580 22614
rect 5644 22612 5650 22676
rect 6729 22674 6795 22677
rect 7046 22674 7052 22676
rect 6729 22672 7052 22674
rect 6729 22616 6734 22672
rect 6790 22616 7052 22672
rect 6729 22614 7052 22616
rect 6729 22611 6795 22614
rect 7046 22612 7052 22614
rect 7116 22612 7122 22676
rect 2814 22476 2820 22540
rect 2884 22538 2890 22540
rect 7005 22538 7071 22541
rect 2884 22536 7071 22538
rect 2884 22480 7010 22536
rect 7066 22480 7071 22536
rect 2884 22478 7071 22480
rect 2884 22476 2890 22478
rect 7005 22475 7071 22478
rect 3325 22402 3391 22405
rect 3734 22402 3740 22404
rect 3325 22400 3740 22402
rect 3325 22344 3330 22400
rect 3386 22344 3740 22400
rect 3325 22342 3740 22344
rect 3325 22339 3391 22342
rect 3734 22340 3740 22342
rect 3804 22340 3810 22404
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 3509 22266 3575 22269
rect 3734 22266 3740 22268
rect 3509 22264 3740 22266
rect 3509 22208 3514 22264
rect 3570 22208 3740 22264
rect 3509 22206 3740 22208
rect 3509 22203 3575 22206
rect 3734 22204 3740 22206
rect 3804 22204 3810 22268
rect 4061 22266 4127 22269
rect 4286 22266 4292 22268
rect 4061 22264 4292 22266
rect 4061 22208 4066 22264
rect 4122 22208 4292 22264
rect 4061 22206 4292 22208
rect 4061 22203 4127 22206
rect 4286 22204 4292 22206
rect 4356 22204 4362 22268
rect 6678 22204 6684 22268
rect 6748 22266 6754 22268
rect 6913 22266 6979 22269
rect 7189 22268 7255 22269
rect 7189 22266 7236 22268
rect 6748 22264 6979 22266
rect 6748 22208 6918 22264
rect 6974 22208 6979 22264
rect 6748 22206 6979 22208
rect 7144 22264 7236 22266
rect 7144 22208 7194 22264
rect 7144 22206 7236 22208
rect 6748 22204 6754 22206
rect 6913 22203 6979 22206
rect 7189 22204 7236 22206
rect 7300 22204 7306 22268
rect 7189 22203 7255 22204
rect 0 22130 120 22160
rect 7468 22133 7528 23566
rect 8017 23563 8083 23566
rect 8201 23626 8267 23629
rect 8201 23624 8402 23626
rect 8201 23568 8206 23624
rect 8262 23568 8402 23624
rect 8201 23566 8402 23568
rect 8201 23563 8267 23566
rect 7946 23424 8262 23425
rect 7946 23360 7952 23424
rect 8016 23360 8032 23424
rect 8096 23360 8112 23424
rect 8176 23360 8192 23424
rect 8256 23360 8262 23424
rect 7946 23359 8262 23360
rect 8017 23218 8083 23221
rect 8342 23218 8402 23566
rect 10225 23490 10291 23493
rect 11130 23490 11250 23520
rect 10225 23488 11250 23490
rect 10225 23432 10230 23488
rect 10286 23432 11250 23488
rect 10225 23430 11250 23432
rect 10225 23427 10291 23430
rect 11130 23400 11250 23430
rect 8017 23216 8402 23218
rect 8017 23160 8022 23216
rect 8078 23160 8402 23216
rect 8017 23158 8402 23160
rect 9673 23218 9739 23221
rect 11130 23218 11250 23248
rect 9673 23216 11250 23218
rect 9673 23160 9678 23216
rect 9734 23160 11250 23216
rect 9673 23158 11250 23160
rect 8017 23155 8083 23158
rect 9673 23155 9739 23158
rect 11130 23128 11250 23158
rect 10225 22946 10291 22949
rect 11130 22946 11250 22976
rect 10225 22944 11250 22946
rect 10225 22888 10230 22944
rect 10286 22888 11250 22944
rect 10225 22886 11250 22888
rect 10225 22883 10291 22886
rect 9006 22880 9322 22881
rect 9006 22816 9012 22880
rect 9076 22816 9092 22880
rect 9156 22816 9172 22880
rect 9236 22816 9252 22880
rect 9316 22816 9322 22880
rect 11130 22856 11250 22886
rect 9006 22815 9322 22816
rect 9765 22674 9831 22677
rect 11130 22674 11250 22704
rect 9765 22672 11250 22674
rect 9765 22616 9770 22672
rect 9826 22616 11250 22672
rect 9765 22614 11250 22616
rect 9765 22611 9831 22614
rect 11130 22584 11250 22614
rect 8017 22538 8083 22541
rect 9990 22538 9996 22540
rect 8017 22536 9996 22538
rect 8017 22480 8022 22536
rect 8078 22480 9996 22536
rect 8017 22478 9996 22480
rect 8017 22475 8083 22478
rect 9990 22476 9996 22478
rect 10060 22476 10066 22540
rect 9673 22402 9739 22405
rect 11130 22402 11250 22432
rect 9673 22400 11250 22402
rect 9673 22344 9678 22400
rect 9734 22344 11250 22400
rect 9673 22342 11250 22344
rect 9673 22339 9739 22342
rect 7946 22336 8262 22337
rect 7946 22272 7952 22336
rect 8016 22272 8032 22336
rect 8096 22272 8112 22336
rect 8176 22272 8192 22336
rect 8256 22272 8262 22336
rect 11130 22312 11250 22342
rect 7946 22271 8262 22272
rect 1393 22130 1459 22133
rect 0 22128 1459 22130
rect 0 22072 1398 22128
rect 1454 22072 1459 22128
rect 0 22070 1459 22072
rect 0 22040 120 22070
rect 1393 22067 1459 22070
rect 1526 22068 1532 22132
rect 1596 22068 1602 22132
rect 3693 22130 3759 22133
rect 3693 22128 7344 22130
rect 3693 22072 3698 22128
rect 3754 22072 7344 22128
rect 3693 22070 7344 22072
rect 1534 21997 1594 22068
rect 3693 22067 3759 22070
rect 1485 21992 1594 21997
rect 1485 21936 1490 21992
rect 1546 21936 1594 21992
rect 1485 21934 1594 21936
rect 2681 21994 2747 21997
rect 4889 21994 4955 21997
rect 2681 21992 4955 21994
rect 2681 21936 2686 21992
rect 2742 21936 4894 21992
rect 4950 21936 4955 21992
rect 2681 21934 4955 21936
rect 1485 21931 1551 21934
rect 2681 21931 2747 21934
rect 4889 21931 4955 21934
rect 6913 21994 6979 21997
rect 7097 21994 7163 21997
rect 6913 21992 7163 21994
rect 6913 21936 6918 21992
rect 6974 21936 7102 21992
rect 7158 21936 7163 21992
rect 6913 21934 7163 21936
rect 6913 21931 6979 21934
rect 7097 21931 7163 21934
rect 3969 21858 4035 21861
rect 4797 21860 4863 21861
rect 4797 21858 4844 21860
rect 3604 21856 4035 21858
rect 3604 21800 3974 21856
rect 4030 21800 4035 21856
rect 3604 21798 4035 21800
rect 4752 21856 4844 21858
rect 4752 21800 4802 21856
rect 4752 21798 4844 21800
rect 3006 21792 3322 21793
rect 3006 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3322 21792
rect 3006 21727 3322 21728
rect 1526 21524 1532 21588
rect 1596 21586 1602 21588
rect 2446 21586 2452 21588
rect 1596 21526 2452 21586
rect 1596 21524 1602 21526
rect 2446 21524 2452 21526
rect 2516 21524 2522 21588
rect 2221 21450 2287 21453
rect 2221 21448 2468 21450
rect 2221 21392 2226 21448
rect 2282 21392 2468 21448
rect 2221 21390 2468 21392
rect 2221 21387 2287 21390
rect 0 21314 120 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 120 21254
rect 1393 21251 1459 21254
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 2037 21042 2103 21045
rect 2408 21042 2468 21390
rect 3604 21178 3664 21798
rect 3969 21795 4035 21798
rect 4797 21796 4844 21798
rect 4908 21796 4914 21860
rect 5809 21858 5875 21861
rect 7097 21860 7163 21861
rect 7046 21858 7052 21860
rect 5398 21856 5875 21858
rect 5398 21800 5814 21856
rect 5870 21800 5875 21856
rect 5398 21798 5875 21800
rect 7006 21798 7052 21858
rect 7116 21856 7163 21860
rect 7158 21800 7163 21856
rect 4797 21795 4863 21796
rect 5398 21725 5458 21798
rect 5809 21795 5875 21798
rect 7046 21796 7052 21798
rect 7116 21796 7163 21800
rect 7284 21858 7344 22070
rect 7465 22128 7531 22133
rect 7465 22072 7470 22128
rect 7526 22072 7531 22128
rect 7465 22067 7531 22072
rect 9857 22130 9923 22133
rect 11130 22130 11250 22160
rect 9857 22128 11250 22130
rect 9857 22072 9862 22128
rect 9918 22072 11250 22128
rect 9857 22070 11250 22072
rect 9857 22067 9923 22070
rect 11130 22040 11250 22070
rect 8702 21932 8708 21996
rect 8772 21994 8778 21996
rect 9397 21994 9463 21997
rect 8772 21992 9463 21994
rect 8772 21936 9402 21992
rect 9458 21936 9463 21992
rect 8772 21934 9463 21936
rect 8772 21932 8778 21934
rect 9397 21931 9463 21934
rect 8477 21858 8543 21861
rect 7284 21856 8543 21858
rect 7284 21800 8482 21856
rect 8538 21800 8543 21856
rect 7284 21798 8543 21800
rect 7097 21795 7163 21796
rect 8477 21795 8543 21798
rect 9673 21858 9739 21861
rect 11130 21858 11250 21888
rect 9673 21856 11250 21858
rect 9673 21800 9678 21856
rect 9734 21800 11250 21856
rect 9673 21798 11250 21800
rect 9673 21795 9739 21798
rect 9006 21792 9322 21793
rect 9006 21728 9012 21792
rect 9076 21728 9092 21792
rect 9156 21728 9172 21792
rect 9236 21728 9252 21792
rect 9316 21728 9322 21792
rect 11130 21768 11250 21798
rect 9006 21727 9322 21728
rect 3785 21724 3851 21725
rect 3734 21660 3740 21724
rect 3804 21722 3851 21724
rect 4061 21722 4127 21725
rect 4981 21722 5047 21725
rect 3804 21720 3896 21722
rect 3846 21664 3896 21720
rect 3804 21662 3896 21664
rect 4061 21720 5047 21722
rect 4061 21664 4066 21720
rect 4122 21664 4986 21720
rect 5042 21664 5047 21720
rect 4061 21662 5047 21664
rect 5398 21720 5507 21725
rect 5398 21664 5446 21720
rect 5502 21664 5507 21720
rect 5398 21662 5507 21664
rect 3804 21660 3851 21662
rect 3785 21659 3851 21660
rect 4061 21659 4127 21662
rect 4981 21659 5047 21662
rect 5441 21659 5507 21662
rect 5574 21660 5580 21724
rect 5644 21722 5650 21724
rect 7741 21722 7807 21725
rect 5644 21720 7807 21722
rect 5644 21664 7746 21720
rect 7802 21664 7807 21720
rect 5644 21662 7807 21664
rect 5644 21660 5650 21662
rect 7741 21659 7807 21662
rect 7925 21722 7991 21725
rect 8702 21722 8708 21724
rect 7925 21720 8708 21722
rect 7925 21664 7930 21720
rect 7986 21664 8708 21720
rect 7925 21662 8708 21664
rect 7925 21659 7991 21662
rect 8702 21660 8708 21662
rect 8772 21660 8778 21724
rect 10685 21722 10751 21725
rect 10910 21722 10916 21724
rect 10685 21720 10916 21722
rect 10685 21664 10690 21720
rect 10746 21664 10916 21720
rect 10685 21662 10916 21664
rect 10685 21659 10751 21662
rect 10910 21660 10916 21662
rect 10980 21660 10986 21724
rect 3734 21524 3740 21588
rect 3804 21586 3810 21588
rect 6494 21586 6500 21588
rect 3804 21526 6500 21586
rect 3804 21524 3810 21526
rect 6494 21524 6500 21526
rect 6564 21524 6570 21588
rect 9857 21586 9923 21589
rect 11130 21586 11250 21616
rect 9857 21584 11250 21586
rect 9857 21528 9862 21584
rect 9918 21528 11250 21584
rect 9857 21526 11250 21528
rect 9857 21523 9923 21526
rect 11130 21496 11250 21526
rect 4061 21450 4127 21453
rect 4245 21450 4311 21453
rect 5390 21450 5396 21452
rect 4061 21448 4170 21450
rect 4061 21392 4066 21448
rect 4122 21392 4170 21448
rect 4061 21387 4170 21392
rect 4245 21448 5396 21450
rect 4245 21392 4250 21448
rect 4306 21392 5396 21448
rect 4245 21390 5396 21392
rect 4245 21387 4311 21390
rect 5390 21388 5396 21390
rect 5460 21388 5466 21452
rect 5809 21450 5875 21453
rect 9029 21450 9095 21453
rect 5809 21448 9095 21450
rect 5809 21392 5814 21448
rect 5870 21392 9034 21448
rect 9090 21392 9095 21448
rect 5809 21390 9095 21392
rect 5809 21387 5875 21390
rect 9029 21387 9095 21390
rect 4110 21314 4170 21387
rect 4705 21314 4771 21317
rect 4110 21312 4771 21314
rect 4110 21256 4710 21312
rect 4766 21256 4771 21312
rect 4110 21254 4771 21256
rect 4705 21251 4771 21254
rect 6637 21314 6703 21317
rect 6862 21314 6868 21316
rect 6637 21312 6868 21314
rect 6637 21256 6642 21312
rect 6698 21256 6868 21312
rect 6637 21254 6868 21256
rect 6637 21251 6703 21254
rect 6862 21252 6868 21254
rect 6932 21252 6938 21316
rect 7189 21314 7255 21317
rect 9673 21314 9739 21317
rect 11130 21314 11250 21344
rect 7189 21312 7850 21314
rect 7189 21256 7194 21312
rect 7250 21256 7850 21312
rect 7189 21254 7850 21256
rect 7189 21251 7255 21254
rect 3785 21178 3851 21181
rect 3604 21176 3851 21178
rect 3604 21120 3790 21176
rect 3846 21120 3851 21176
rect 3604 21118 3851 21120
rect 3785 21115 3851 21118
rect 5073 21178 5139 21181
rect 5206 21178 5212 21180
rect 5073 21176 5212 21178
rect 5073 21120 5078 21176
rect 5134 21120 5212 21176
rect 5073 21118 5212 21120
rect 5073 21115 5139 21118
rect 5206 21116 5212 21118
rect 5276 21116 5282 21180
rect 7649 21178 7715 21181
rect 7606 21176 7715 21178
rect 7606 21120 7654 21176
rect 7710 21120 7715 21176
rect 7606 21115 7715 21120
rect 2037 21040 2468 21042
rect 2037 20984 2042 21040
rect 2098 20984 2468 21040
rect 2037 20982 2468 20984
rect 2037 20979 2103 20982
rect 2630 20844 2636 20908
rect 2700 20906 2706 20908
rect 4797 20906 4863 20909
rect 2700 20904 4863 20906
rect 2700 20848 4802 20904
rect 4858 20848 4863 20904
rect 2700 20846 4863 20848
rect 2700 20844 2706 20846
rect 4797 20843 4863 20846
rect 3785 20768 3851 20773
rect 3785 20712 3790 20768
rect 3846 20712 3851 20768
rect 3785 20707 3851 20712
rect 3969 20770 4035 20773
rect 4102 20770 4108 20772
rect 3969 20768 4108 20770
rect 3969 20712 3974 20768
rect 4030 20712 4108 20768
rect 3969 20710 4108 20712
rect 3969 20707 4035 20710
rect 4102 20708 4108 20710
rect 4172 20708 4178 20772
rect 3006 20704 3322 20705
rect 3006 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3322 20704
rect 3006 20639 3322 20640
rect 1393 20636 1459 20637
rect 1342 20572 1348 20636
rect 1412 20634 1459 20636
rect 3788 20634 3848 20707
rect 4102 20634 4108 20636
rect 1412 20632 1504 20634
rect 1454 20576 1504 20632
rect 1412 20574 1504 20576
rect 3788 20574 4108 20634
rect 1412 20572 1459 20574
rect 4102 20572 4108 20574
rect 4172 20572 4178 20636
rect 6361 20634 6427 20637
rect 7230 20634 7236 20636
rect 6361 20632 7236 20634
rect 6361 20576 6366 20632
rect 6422 20576 7236 20632
rect 6361 20574 7236 20576
rect 1393 20571 1459 20572
rect 6361 20571 6427 20574
rect 7230 20572 7236 20574
rect 7300 20572 7306 20636
rect 0 20498 120 20528
rect 841 20498 907 20501
rect 0 20496 907 20498
rect 0 20440 846 20496
rect 902 20440 907 20496
rect 0 20438 907 20440
rect 0 20408 120 20438
rect 841 20435 907 20438
rect 2313 20362 2379 20365
rect 7189 20362 7255 20365
rect 7606 20362 7666 21115
rect 7790 21042 7850 21254
rect 9673 21312 11250 21314
rect 9673 21256 9678 21312
rect 9734 21256 11250 21312
rect 9673 21254 11250 21256
rect 9673 21251 9739 21254
rect 7946 21248 8262 21249
rect 7946 21184 7952 21248
rect 8016 21184 8032 21248
rect 8096 21184 8112 21248
rect 8176 21184 8192 21248
rect 8256 21184 8262 21248
rect 11130 21224 11250 21254
rect 7946 21183 8262 21184
rect 7925 21042 7991 21045
rect 7790 21040 7991 21042
rect 7790 20984 7930 21040
rect 7986 20984 7991 21040
rect 7790 20982 7991 20984
rect 7925 20979 7991 20982
rect 8477 21042 8543 21045
rect 10225 21042 10291 21045
rect 11130 21042 11250 21072
rect 8477 21040 8724 21042
rect 8477 20984 8482 21040
rect 8538 20984 8724 21040
rect 8477 20982 8724 20984
rect 8477 20979 8543 20982
rect 8664 20501 8724 20982
rect 10225 21040 11250 21042
rect 10225 20984 10230 21040
rect 10286 20984 11250 21040
rect 10225 20982 11250 20984
rect 10225 20979 10291 20982
rect 11130 20952 11250 20982
rect 9673 20770 9739 20773
rect 11130 20770 11250 20800
rect 9673 20768 11250 20770
rect 9673 20712 9678 20768
rect 9734 20712 11250 20768
rect 9673 20710 11250 20712
rect 9673 20707 9739 20710
rect 9006 20704 9322 20705
rect 9006 20640 9012 20704
rect 9076 20640 9092 20704
rect 9156 20640 9172 20704
rect 9236 20640 9252 20704
rect 9316 20640 9322 20704
rect 11130 20680 11250 20710
rect 9006 20639 9322 20640
rect 8661 20496 8727 20501
rect 8661 20440 8666 20496
rect 8722 20440 8727 20496
rect 8661 20435 8727 20440
rect 9121 20498 9187 20501
rect 9622 20498 9628 20500
rect 9121 20496 9628 20498
rect 9121 20440 9126 20496
rect 9182 20440 9628 20496
rect 9121 20438 9628 20440
rect 9121 20435 9187 20438
rect 9622 20436 9628 20438
rect 9692 20436 9698 20500
rect 10225 20498 10291 20501
rect 11130 20498 11250 20528
rect 10225 20496 11250 20498
rect 10225 20440 10230 20496
rect 10286 20440 11250 20496
rect 10225 20438 11250 20440
rect 10225 20435 10291 20438
rect 11130 20408 11250 20438
rect 2313 20360 2514 20362
rect 2313 20304 2318 20360
rect 2374 20304 2514 20360
rect 2313 20302 2514 20304
rect 2313 20299 2379 20302
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 2313 19818 2379 19821
rect 2454 19818 2514 20302
rect 7189 20360 7666 20362
rect 7189 20304 7194 20360
rect 7250 20304 7666 20360
rect 7189 20302 7666 20304
rect 7189 20299 7255 20302
rect 8702 20300 8708 20364
rect 8772 20362 8778 20364
rect 8937 20362 9003 20365
rect 8772 20360 9003 20362
rect 8772 20304 8942 20360
rect 8998 20304 9003 20360
rect 8772 20302 9003 20304
rect 8772 20300 8778 20302
rect 8937 20299 9003 20302
rect 9673 20226 9739 20229
rect 11130 20226 11250 20256
rect 9673 20224 11250 20226
rect 9673 20168 9678 20224
rect 9734 20168 11250 20224
rect 9673 20166 11250 20168
rect 9673 20163 9739 20166
rect 7946 20160 8262 20161
rect 7946 20096 7952 20160
rect 8016 20096 8032 20160
rect 8096 20096 8112 20160
rect 8176 20096 8192 20160
rect 8256 20096 8262 20160
rect 11130 20136 11250 20166
rect 7946 20095 8262 20096
rect 2865 19954 2931 19957
rect 2313 19816 2514 19818
rect 2313 19760 2318 19816
rect 2374 19760 2514 19816
rect 2313 19758 2514 19760
rect 2822 19952 2931 19954
rect 2822 19896 2870 19952
rect 2926 19896 2931 19952
rect 2822 19891 2931 19896
rect 6637 19952 6703 19957
rect 6637 19896 6642 19952
rect 6698 19896 6703 19952
rect 6637 19891 6703 19896
rect 10041 19954 10107 19957
rect 11130 19954 11250 19984
rect 10041 19952 11250 19954
rect 10041 19896 10046 19952
rect 10102 19896 11250 19952
rect 10041 19894 11250 19896
rect 10041 19891 10107 19894
rect 2313 19755 2379 19758
rect 0 19682 120 19712
rect 1393 19682 1459 19685
rect 0 19680 1459 19682
rect 0 19624 1398 19680
rect 1454 19624 1459 19680
rect 0 19622 1459 19624
rect 0 19592 120 19622
rect 1393 19619 1459 19622
rect 2822 19410 2882 19891
rect 6361 19818 6427 19821
rect 6640 19818 6700 19891
rect 11130 19864 11250 19894
rect 9029 19818 9095 19821
rect 6361 19816 6700 19818
rect 6361 19760 6366 19816
rect 6422 19760 6700 19816
rect 6361 19758 6700 19760
rect 8756 19816 9095 19818
rect 8756 19760 9034 19816
rect 9090 19760 9095 19816
rect 8756 19758 9095 19760
rect 6361 19755 6427 19758
rect 3877 19682 3943 19685
rect 6678 19682 6684 19684
rect 3877 19680 6684 19682
rect 3877 19624 3882 19680
rect 3938 19624 6684 19680
rect 3877 19622 6684 19624
rect 3877 19619 3943 19622
rect 6678 19620 6684 19622
rect 6748 19682 6754 19684
rect 7557 19682 7623 19685
rect 6748 19680 7623 19682
rect 6748 19624 7562 19680
rect 7618 19624 7623 19680
rect 6748 19622 7623 19624
rect 6748 19620 6754 19622
rect 7557 19619 7623 19622
rect 3006 19616 3322 19617
rect 3006 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3322 19616
rect 3006 19551 3322 19552
rect 2957 19410 3023 19413
rect 2822 19408 3023 19410
rect 2822 19352 2962 19408
rect 3018 19352 3023 19408
rect 2822 19350 3023 19352
rect 2957 19347 3023 19350
rect 7782 19348 7788 19412
rect 7852 19410 7858 19412
rect 8756 19410 8816 19758
rect 9029 19755 9095 19758
rect 10225 19682 10291 19685
rect 11130 19682 11250 19712
rect 10225 19680 11250 19682
rect 10225 19624 10230 19680
rect 10286 19624 11250 19680
rect 10225 19622 11250 19624
rect 10225 19619 10291 19622
rect 9006 19616 9322 19617
rect 9006 19552 9012 19616
rect 9076 19552 9092 19616
rect 9156 19552 9172 19616
rect 9236 19552 9252 19616
rect 9316 19552 9322 19616
rect 11130 19592 11250 19622
rect 9006 19551 9322 19552
rect 10409 19546 10475 19549
rect 10726 19546 10732 19548
rect 10409 19544 10732 19546
rect 10409 19488 10414 19544
rect 10470 19488 10732 19544
rect 10409 19486 10732 19488
rect 10409 19483 10475 19486
rect 10726 19484 10732 19486
rect 10796 19484 10802 19548
rect 8937 19410 9003 19413
rect 7852 19350 8402 19410
rect 8756 19408 9003 19410
rect 8756 19352 8942 19408
rect 8998 19352 9003 19408
rect 8756 19350 9003 19352
rect 7852 19348 7858 19350
rect 7925 19274 7991 19277
rect 7790 19272 7991 19274
rect 7790 19216 7930 19272
rect 7986 19216 7991 19272
rect 7790 19214 7991 19216
rect 8342 19274 8402 19350
rect 8937 19347 9003 19350
rect 9673 19410 9739 19413
rect 11130 19410 11250 19440
rect 9673 19408 11250 19410
rect 9673 19352 9678 19408
rect 9734 19352 11250 19408
rect 9673 19350 11250 19352
rect 9673 19347 9739 19350
rect 11130 19320 11250 19350
rect 10685 19274 10751 19277
rect 8342 19272 10751 19274
rect 8342 19216 10690 19272
rect 10746 19216 10751 19272
rect 8342 19214 10751 19216
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 5901 19004 5967 19005
rect 5901 19002 5948 19004
rect 5856 19000 5948 19002
rect 5856 18944 5906 19000
rect 5856 18942 5948 18944
rect 5901 18940 5948 18942
rect 6012 18940 6018 19004
rect 5901 18939 5967 18940
rect 0 18866 120 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 120 18806
rect 1393 18803 1459 18806
rect 3877 18866 3943 18869
rect 5165 18866 5231 18869
rect 3877 18864 5231 18866
rect 3877 18808 3882 18864
rect 3938 18808 5170 18864
rect 5226 18808 5231 18864
rect 3877 18806 5231 18808
rect 3877 18803 3943 18806
rect 5165 18803 5231 18806
rect 6361 18866 6427 18869
rect 6678 18866 6684 18868
rect 6361 18864 6684 18866
rect 6361 18808 6366 18864
rect 6422 18808 6684 18864
rect 6361 18806 6684 18808
rect 6361 18803 6427 18806
rect 6678 18804 6684 18806
rect 6748 18804 6754 18868
rect 7790 18866 7850 19214
rect 7925 19211 7991 19214
rect 10685 19211 10751 19214
rect 9673 19138 9739 19141
rect 11130 19138 11250 19168
rect 9673 19136 11250 19138
rect 9673 19080 9678 19136
rect 9734 19080 11250 19136
rect 9673 19078 11250 19080
rect 9673 19075 9739 19078
rect 7946 19072 8262 19073
rect 7946 19008 7952 19072
rect 8016 19008 8032 19072
rect 8096 19008 8112 19072
rect 8176 19008 8192 19072
rect 8256 19008 8262 19072
rect 11130 19048 11250 19078
rect 7946 19007 8262 19008
rect 8702 18866 8708 18868
rect 7790 18806 8708 18866
rect 8702 18804 8708 18806
rect 8772 18804 8778 18868
rect 10225 18866 10291 18869
rect 11130 18866 11250 18896
rect 10225 18864 11250 18866
rect 10225 18808 10230 18864
rect 10286 18808 11250 18864
rect 10225 18806 11250 18808
rect 10225 18803 10291 18806
rect 11130 18776 11250 18806
rect 3693 18730 3759 18733
rect 5349 18730 5415 18733
rect 3693 18728 5415 18730
rect 3693 18672 3698 18728
rect 3754 18672 5354 18728
rect 5410 18672 5415 18728
rect 3693 18670 5415 18672
rect 3693 18667 3759 18670
rect 5349 18667 5415 18670
rect 5942 18668 5948 18732
rect 6012 18730 6018 18732
rect 9305 18730 9371 18733
rect 6012 18728 9371 18730
rect 6012 18672 9310 18728
rect 9366 18672 9371 18728
rect 6012 18670 9371 18672
rect 6012 18668 6018 18670
rect 9305 18667 9371 18670
rect 9673 18730 9739 18733
rect 10910 18730 10916 18732
rect 9673 18728 10916 18730
rect 9673 18672 9678 18728
rect 9734 18672 10916 18728
rect 9673 18670 10916 18672
rect 9673 18667 9739 18670
rect 10910 18668 10916 18670
rect 10980 18668 10986 18732
rect 3877 18594 3943 18597
rect 4102 18594 4108 18596
rect 3877 18592 4108 18594
rect 3877 18536 3882 18592
rect 3938 18536 4108 18592
rect 3877 18534 4108 18536
rect 3877 18531 3943 18534
rect 4102 18532 4108 18534
rect 4172 18532 4178 18596
rect 9673 18594 9739 18597
rect 11130 18594 11250 18624
rect 9673 18592 11250 18594
rect 9673 18536 9678 18592
rect 9734 18536 11250 18592
rect 9673 18534 11250 18536
rect 9673 18531 9739 18534
rect 3006 18528 3322 18529
rect 3006 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3322 18528
rect 3006 18463 3322 18464
rect 9006 18528 9322 18529
rect 9006 18464 9012 18528
rect 9076 18464 9092 18528
rect 9156 18464 9172 18528
rect 9236 18464 9252 18528
rect 9316 18464 9322 18528
rect 11130 18504 11250 18534
rect 9006 18463 9322 18464
rect 4286 18260 4292 18324
rect 4356 18322 4362 18324
rect 9029 18322 9095 18325
rect 4356 18320 9095 18322
rect 4356 18264 9034 18320
rect 9090 18264 9095 18320
rect 4356 18262 9095 18264
rect 4356 18260 4362 18262
rect 9029 18259 9095 18262
rect 9949 18322 10015 18325
rect 11130 18322 11250 18352
rect 9949 18320 11250 18322
rect 9949 18264 9954 18320
rect 10010 18264 11250 18320
rect 9949 18262 11250 18264
rect 9949 18259 10015 18262
rect 11130 18232 11250 18262
rect 197 18186 263 18189
rect 5574 18186 5580 18188
rect 197 18184 5580 18186
rect 197 18128 202 18184
rect 258 18128 5580 18184
rect 197 18126 5580 18128
rect 197 18123 263 18126
rect 5574 18124 5580 18126
rect 5644 18124 5650 18188
rect 6862 18124 6868 18188
rect 6932 18186 6938 18188
rect 7782 18186 7788 18188
rect 6932 18126 7788 18186
rect 6932 18124 6938 18126
rect 7782 18124 7788 18126
rect 7852 18186 7858 18188
rect 8109 18186 8175 18189
rect 7852 18184 8175 18186
rect 7852 18128 8114 18184
rect 8170 18128 8175 18184
rect 7852 18126 8175 18128
rect 7852 18124 7858 18126
rect 8109 18123 8175 18126
rect 0 18050 120 18080
rect 1393 18050 1459 18053
rect 0 18048 1459 18050
rect 0 17992 1398 18048
rect 1454 17992 1459 18048
rect 0 17990 1459 17992
rect 0 17960 120 17990
rect 1393 17987 1459 17990
rect 2814 17988 2820 18052
rect 2884 18050 2890 18052
rect 3325 18050 3391 18053
rect 3969 18050 4035 18053
rect 2884 18048 3391 18050
rect 2884 17992 3330 18048
rect 3386 17992 3391 18048
rect 2884 17990 3391 17992
rect 2884 17988 2890 17990
rect 3325 17987 3391 17990
rect 3926 18048 4035 18050
rect 3926 17992 3974 18048
rect 4030 17992 4035 18048
rect 3926 17987 4035 17992
rect 4654 17988 4660 18052
rect 4724 18050 4730 18052
rect 9857 18050 9923 18053
rect 11130 18050 11250 18080
rect 4724 17990 4906 18050
rect 4724 17988 4730 17990
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 2446 17852 2452 17916
rect 2516 17914 2522 17916
rect 2681 17914 2747 17917
rect 2516 17912 2747 17914
rect 2516 17856 2686 17912
rect 2742 17856 2747 17912
rect 2516 17854 2747 17856
rect 2516 17852 2522 17854
rect 2681 17851 2747 17854
rect 2814 17852 2820 17916
rect 2884 17914 2890 17916
rect 3509 17914 3575 17917
rect 2884 17912 3575 17914
rect 2884 17856 3514 17912
rect 3570 17856 3575 17912
rect 2884 17854 3575 17856
rect 3926 17914 3986 17987
rect 4654 17914 4660 17916
rect 3926 17854 4660 17914
rect 2884 17852 2890 17854
rect 3509 17851 3575 17854
rect 4654 17852 4660 17854
rect 4724 17852 4730 17916
rect 4846 17914 4906 17990
rect 9857 18048 11250 18050
rect 9857 17992 9862 18048
rect 9918 17992 11250 18048
rect 9857 17990 11250 17992
rect 9857 17987 9923 17990
rect 7946 17984 8262 17985
rect 7946 17920 7952 17984
rect 8016 17920 8032 17984
rect 8096 17920 8112 17984
rect 8176 17920 8192 17984
rect 8256 17920 8262 17984
rect 11130 17960 11250 17990
rect 7946 17919 8262 17920
rect 5533 17914 5599 17917
rect 6269 17916 6335 17917
rect 6269 17914 6316 17916
rect 4846 17912 5599 17914
rect 4846 17856 5538 17912
rect 5594 17856 5599 17912
rect 4846 17854 5599 17856
rect 6224 17912 6316 17914
rect 6224 17856 6274 17912
rect 6224 17854 6316 17856
rect 5533 17851 5599 17854
rect 6269 17852 6316 17854
rect 6380 17852 6386 17916
rect 9622 17914 9628 17916
rect 8342 17854 9628 17914
rect 6269 17851 6335 17852
rect 7649 17778 7715 17781
rect 8342 17778 8402 17854
rect 9622 17852 9628 17854
rect 9692 17914 9698 17916
rect 9990 17914 9996 17916
rect 9692 17854 9996 17914
rect 9692 17852 9698 17854
rect 9990 17852 9996 17854
rect 10060 17852 10066 17916
rect 7649 17776 8402 17778
rect 7649 17720 7654 17776
rect 7710 17720 8402 17776
rect 7649 17718 8402 17720
rect 9765 17778 9831 17781
rect 11130 17778 11250 17808
rect 9765 17776 11250 17778
rect 9765 17720 9770 17776
rect 9826 17720 11250 17776
rect 9765 17718 11250 17720
rect 7649 17715 7715 17718
rect 9765 17715 9831 17718
rect 11130 17688 11250 17718
rect 9673 17506 9739 17509
rect 11130 17506 11250 17536
rect 9673 17504 11250 17506
rect 9673 17448 9678 17504
rect 9734 17448 11250 17504
rect 9673 17446 11250 17448
rect 9673 17443 9739 17446
rect 3006 17440 3322 17441
rect 3006 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3322 17440
rect 3006 17375 3322 17376
rect 9006 17440 9322 17441
rect 9006 17376 9012 17440
rect 9076 17376 9092 17440
rect 9156 17376 9172 17440
rect 9236 17376 9252 17440
rect 9316 17376 9322 17440
rect 11130 17416 11250 17446
rect 9006 17375 9322 17376
rect 2405 17370 2471 17373
rect 9581 17370 9647 17373
rect 2405 17368 2698 17370
rect 2405 17312 2410 17368
rect 2466 17312 2698 17368
rect 2405 17310 2698 17312
rect 2405 17307 2471 17310
rect 0 17234 120 17264
rect 657 17234 723 17237
rect 0 17232 723 17234
rect 0 17176 662 17232
rect 718 17176 723 17232
rect 0 17174 723 17176
rect 0 17144 120 17174
rect 657 17171 723 17174
rect 2313 17098 2379 17101
rect 2446 17098 2452 17100
rect 2313 17096 2452 17098
rect 2313 17040 2318 17096
rect 2374 17040 2452 17096
rect 2313 17038 2452 17040
rect 2313 17035 2379 17038
rect 2446 17036 2452 17038
rect 2516 17036 2522 17100
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 2638 16690 2698 17310
rect 9446 17368 9647 17370
rect 9446 17312 9586 17368
rect 9642 17312 9647 17368
rect 9446 17310 9647 17312
rect 9305 17234 9371 17237
rect 9446 17234 9506 17310
rect 9581 17307 9647 17310
rect 9305 17232 9506 17234
rect 9305 17176 9310 17232
rect 9366 17176 9506 17232
rect 9305 17174 9506 17176
rect 9765 17234 9831 17237
rect 11130 17234 11250 17264
rect 9765 17232 11250 17234
rect 9765 17176 9770 17232
rect 9826 17176 11250 17232
rect 9765 17174 11250 17176
rect 9305 17171 9371 17174
rect 9765 17171 9831 17174
rect 11130 17144 11250 17174
rect 3233 17098 3299 17101
rect 3509 17098 3575 17101
rect 5073 17100 5139 17101
rect 3734 17098 3740 17100
rect 3233 17096 3740 17098
rect 3233 17040 3238 17096
rect 3294 17040 3514 17096
rect 3570 17040 3740 17096
rect 3233 17038 3740 17040
rect 3233 17035 3299 17038
rect 3509 17035 3575 17038
rect 3734 17036 3740 17038
rect 3804 17036 3810 17100
rect 5022 17036 5028 17100
rect 5092 17098 5139 17100
rect 5092 17096 5184 17098
rect 5134 17040 5184 17096
rect 5092 17038 5184 17040
rect 5092 17036 5139 17038
rect 7782 17036 7788 17100
rect 7852 17098 7858 17100
rect 8109 17098 8175 17101
rect 7852 17096 8175 17098
rect 7852 17040 8114 17096
rect 8170 17040 8175 17096
rect 7852 17038 8175 17040
rect 7852 17036 7858 17038
rect 5073 17035 5139 17036
rect 8109 17035 8175 17038
rect 2957 16962 3023 16965
rect 3734 16962 3740 16964
rect 2957 16960 3740 16962
rect 2957 16904 2962 16960
rect 3018 16904 3740 16960
rect 2957 16902 3740 16904
rect 2957 16899 3023 16902
rect 3734 16900 3740 16902
rect 3804 16900 3810 16964
rect 4470 16900 4476 16964
rect 4540 16962 4546 16964
rect 5441 16962 5507 16965
rect 4540 16960 5507 16962
rect 4540 16904 5446 16960
rect 5502 16904 5507 16960
rect 4540 16902 5507 16904
rect 4540 16900 4546 16902
rect 5441 16899 5507 16902
rect 9673 16962 9739 16965
rect 11130 16962 11250 16992
rect 9673 16960 11250 16962
rect 9673 16904 9678 16960
rect 9734 16904 11250 16960
rect 9673 16902 11250 16904
rect 9673 16899 9739 16902
rect 7946 16896 8262 16897
rect 7946 16832 7952 16896
rect 8016 16832 8032 16896
rect 8096 16832 8112 16896
rect 8176 16832 8192 16896
rect 8256 16832 8262 16896
rect 11130 16872 11250 16902
rect 7946 16831 8262 16832
rect 2773 16690 2839 16693
rect 2638 16688 2839 16690
rect 2638 16632 2778 16688
rect 2834 16632 2839 16688
rect 2638 16630 2839 16632
rect 2773 16627 2839 16630
rect 4286 16628 4292 16692
rect 4356 16690 4362 16692
rect 4889 16690 4955 16693
rect 4356 16688 4955 16690
rect 4356 16632 4894 16688
rect 4950 16632 4955 16688
rect 4356 16630 4955 16632
rect 4356 16628 4362 16630
rect 4889 16627 4955 16630
rect 9673 16690 9739 16693
rect 11130 16690 11250 16720
rect 9673 16688 11250 16690
rect 9673 16632 9678 16688
rect 9734 16632 11250 16688
rect 9673 16630 11250 16632
rect 9673 16627 9739 16630
rect 11130 16600 11250 16630
rect 6085 16554 6151 16557
rect 6494 16554 6500 16556
rect 6085 16552 6500 16554
rect 6085 16496 6090 16552
rect 6146 16496 6500 16552
rect 6085 16494 6500 16496
rect 6085 16491 6151 16494
rect 6494 16492 6500 16494
rect 6564 16492 6570 16556
rect 0 16418 120 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 120 16358
rect 1393 16355 1459 16358
rect 9765 16418 9831 16421
rect 11130 16418 11250 16448
rect 9765 16416 11250 16418
rect 9765 16360 9770 16416
rect 9826 16360 11250 16416
rect 9765 16358 11250 16360
rect 9765 16355 9831 16358
rect 3006 16352 3322 16353
rect 3006 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3322 16352
rect 3006 16287 3322 16288
rect 9006 16352 9322 16353
rect 9006 16288 9012 16352
rect 9076 16288 9092 16352
rect 9156 16288 9172 16352
rect 9236 16288 9252 16352
rect 9316 16288 9322 16352
rect 11130 16328 11250 16358
rect 9006 16287 9322 16288
rect 3601 16280 3667 16285
rect 3601 16224 3606 16280
rect 3662 16224 3667 16280
rect 3601 16219 3667 16224
rect 3325 15874 3391 15877
rect 3604 15874 3664 16219
rect 5758 16084 5764 16148
rect 5828 16146 5834 16148
rect 6269 16146 6335 16149
rect 7557 16148 7623 16149
rect 7557 16146 7604 16148
rect 5828 16144 6335 16146
rect 5828 16088 6274 16144
rect 6330 16088 6335 16144
rect 5828 16086 6335 16088
rect 7512 16144 7604 16146
rect 7512 16088 7562 16144
rect 7512 16086 7604 16088
rect 5828 16084 5834 16086
rect 6269 16083 6335 16086
rect 7557 16084 7604 16086
rect 7668 16084 7674 16148
rect 8017 16146 8083 16149
rect 8569 16146 8635 16149
rect 8017 16144 8635 16146
rect 8017 16088 8022 16144
rect 8078 16088 8574 16144
rect 8630 16088 8635 16144
rect 8017 16086 8635 16088
rect 7557 16083 7623 16084
rect 8017 16083 8083 16086
rect 8569 16083 8635 16086
rect 9857 16146 9923 16149
rect 11130 16146 11250 16176
rect 9857 16144 11250 16146
rect 9857 16088 9862 16144
rect 9918 16088 11250 16144
rect 9857 16086 11250 16088
rect 9857 16083 9923 16086
rect 11130 16056 11250 16086
rect 5533 16008 5599 16013
rect 5533 15952 5538 16008
rect 5594 15952 5599 16008
rect 5533 15947 5599 15952
rect 5758 15948 5764 16012
rect 5828 16010 5834 16012
rect 10358 16010 10364 16012
rect 5828 15950 10364 16010
rect 5828 15948 5834 15950
rect 10358 15948 10364 15950
rect 10428 15948 10434 16012
rect 4981 15874 5047 15877
rect 3325 15872 5047 15874
rect 3325 15816 3330 15872
rect 3386 15816 4986 15872
rect 5042 15816 5047 15872
rect 3325 15814 5047 15816
rect 5536 15874 5596 15947
rect 5993 15874 6059 15877
rect 5536 15872 6059 15874
rect 5536 15816 5998 15872
rect 6054 15816 6059 15872
rect 5536 15814 6059 15816
rect 3325 15811 3391 15814
rect 4981 15811 5047 15814
rect 5993 15811 6059 15814
rect 9673 15874 9739 15877
rect 11130 15874 11250 15904
rect 9673 15872 11250 15874
rect 9673 15816 9678 15872
rect 9734 15816 11250 15872
rect 9673 15814 11250 15816
rect 9673 15811 9739 15814
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 7946 15808 8262 15809
rect 7946 15744 7952 15808
rect 8016 15744 8032 15808
rect 8096 15744 8112 15808
rect 8176 15744 8192 15808
rect 8256 15744 8262 15808
rect 11130 15784 11250 15814
rect 7946 15743 8262 15744
rect 4245 15738 4311 15741
rect 5717 15738 5783 15741
rect 4245 15736 6056 15738
rect 4245 15680 4250 15736
rect 4306 15680 5722 15736
rect 5778 15680 6056 15736
rect 4245 15678 6056 15680
rect 4245 15675 4311 15678
rect 5717 15675 5783 15678
rect 0 15602 120 15632
rect 1209 15602 1275 15605
rect 0 15600 1275 15602
rect 0 15544 1214 15600
rect 1270 15544 1275 15600
rect 0 15542 1275 15544
rect 0 15512 120 15542
rect 1209 15539 1275 15542
rect 5996 15469 6056 15678
rect 7230 15676 7236 15740
rect 7300 15738 7306 15740
rect 7373 15738 7439 15741
rect 7300 15736 7439 15738
rect 7300 15680 7378 15736
rect 7434 15680 7439 15736
rect 7300 15678 7439 15680
rect 7300 15676 7306 15678
rect 7373 15675 7439 15678
rect 7649 15602 7715 15605
rect 9438 15602 9444 15604
rect 7649 15600 9444 15602
rect 7649 15544 7654 15600
rect 7710 15544 9444 15600
rect 7649 15542 9444 15544
rect 7649 15539 7715 15542
rect 9438 15540 9444 15542
rect 9508 15540 9514 15604
rect 9765 15602 9831 15605
rect 11130 15602 11250 15632
rect 9765 15600 11250 15602
rect 9765 15544 9770 15600
rect 9826 15544 11250 15600
rect 9765 15542 11250 15544
rect 9765 15539 9831 15542
rect 11130 15512 11250 15542
rect 5993 15464 6059 15469
rect 5993 15408 5998 15464
rect 6054 15408 6059 15464
rect 5993 15403 6059 15408
rect 7598 15404 7604 15468
rect 7668 15466 7674 15468
rect 10317 15466 10383 15469
rect 7668 15464 10383 15466
rect 7668 15408 10322 15464
rect 10378 15408 10383 15464
rect 7668 15406 10383 15408
rect 7668 15404 7674 15406
rect 10317 15403 10383 15406
rect 10501 15330 10567 15333
rect 11130 15330 11250 15360
rect 10501 15328 11250 15330
rect 10501 15272 10506 15328
rect 10562 15272 11250 15328
rect 10501 15270 11250 15272
rect 10501 15267 10567 15270
rect 3006 15264 3322 15265
rect 3006 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3322 15264
rect 3006 15199 3322 15200
rect 9006 15264 9322 15265
rect 9006 15200 9012 15264
rect 9076 15200 9092 15264
rect 9156 15200 9172 15264
rect 9236 15200 9252 15264
rect 9316 15200 9322 15264
rect 11130 15240 11250 15270
rect 9006 15199 9322 15200
rect 4153 15194 4219 15197
rect 8385 15194 8451 15197
rect 8661 15194 8727 15197
rect 4153 15192 8727 15194
rect 4153 15136 4158 15192
rect 4214 15136 8390 15192
rect 8446 15136 8666 15192
rect 8722 15136 8727 15192
rect 4153 15134 8727 15136
rect 4153 15131 4219 15134
rect 8385 15131 8451 15134
rect 8661 15131 8727 15134
rect 2630 14996 2636 15060
rect 2700 15058 2706 15060
rect 5349 15058 5415 15061
rect 2700 15056 5415 15058
rect 2700 15000 5354 15056
rect 5410 15000 5415 15056
rect 2700 14998 5415 15000
rect 2700 14996 2706 14998
rect 5349 14995 5415 14998
rect 8753 15058 8819 15061
rect 11130 15058 11250 15088
rect 8753 15056 11250 15058
rect 8753 15000 8758 15056
rect 8814 15000 11250 15056
rect 8753 14998 11250 15000
rect 8753 14995 8819 14998
rect 11130 14968 11250 14998
rect 1209 14922 1275 14925
rect 4286 14922 4292 14924
rect 1209 14920 4292 14922
rect 1209 14864 1214 14920
rect 1270 14864 4292 14920
rect 1209 14862 4292 14864
rect 1209 14859 1275 14862
rect 4286 14860 4292 14862
rect 4356 14860 4362 14924
rect 5022 14860 5028 14924
rect 5092 14922 5098 14924
rect 5390 14922 5396 14924
rect 5092 14862 5396 14922
rect 5092 14860 5098 14862
rect 5390 14860 5396 14862
rect 5460 14860 5466 14924
rect 9489 14922 9555 14925
rect 5536 14920 9555 14922
rect 5536 14864 9494 14920
rect 9550 14864 9555 14920
rect 5536 14862 9555 14864
rect 0 14786 120 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 120 14726
rect 1485 14723 1551 14726
rect 3785 14786 3851 14789
rect 5536 14786 5596 14862
rect 9489 14859 9555 14862
rect 3785 14784 5596 14786
rect 3785 14728 3790 14784
rect 3846 14728 5596 14784
rect 3785 14726 5596 14728
rect 9765 14786 9831 14789
rect 11130 14786 11250 14816
rect 9765 14784 11250 14786
rect 9765 14728 9770 14784
rect 9826 14728 11250 14784
rect 9765 14726 11250 14728
rect 3785 14723 3851 14726
rect 9765 14723 9831 14726
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 7946 14720 8262 14721
rect 7946 14656 7952 14720
rect 8016 14656 8032 14720
rect 8096 14656 8112 14720
rect 8176 14656 8192 14720
rect 8256 14656 8262 14720
rect 11130 14696 11250 14726
rect 7946 14655 8262 14656
rect 6678 14588 6684 14652
rect 6748 14650 6754 14652
rect 6748 14590 7850 14650
rect 6748 14588 6754 14590
rect 6729 14516 6795 14517
rect 6678 14514 6684 14516
rect 6638 14454 6684 14514
rect 6748 14512 6795 14516
rect 6790 14456 6795 14512
rect 6678 14452 6684 14454
rect 6748 14452 6795 14456
rect 7790 14514 7850 14590
rect 8334 14588 8340 14652
rect 8404 14650 8410 14652
rect 9305 14650 9371 14653
rect 8404 14648 9371 14650
rect 8404 14592 9310 14648
rect 9366 14592 9371 14648
rect 8404 14590 9371 14592
rect 8404 14588 8410 14590
rect 9305 14587 9371 14590
rect 8661 14514 8727 14517
rect 7790 14512 8727 14514
rect 7790 14456 8666 14512
rect 8722 14456 8727 14512
rect 7790 14454 8727 14456
rect 6729 14451 6795 14452
rect 8661 14451 8727 14454
rect 8845 14514 8911 14517
rect 11130 14514 11250 14544
rect 8845 14512 11250 14514
rect 8845 14456 8850 14512
rect 8906 14456 11250 14512
rect 8845 14454 11250 14456
rect 8845 14451 8911 14454
rect 11130 14424 11250 14454
rect 1526 14316 1532 14380
rect 1596 14378 1602 14380
rect 4153 14378 4219 14381
rect 1596 14376 4219 14378
rect 1596 14320 4158 14376
rect 4214 14320 4219 14376
rect 1596 14318 4219 14320
rect 1596 14316 1602 14318
rect 4153 14315 4219 14318
rect 10685 14242 10751 14245
rect 11130 14242 11250 14272
rect 10685 14240 11250 14242
rect 10685 14184 10690 14240
rect 10746 14184 11250 14240
rect 10685 14182 11250 14184
rect 10685 14179 10751 14182
rect 3006 14176 3322 14177
rect 3006 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3322 14176
rect 3006 14111 3322 14112
rect 9006 14176 9322 14177
rect 9006 14112 9012 14176
rect 9076 14112 9092 14176
rect 9156 14112 9172 14176
rect 9236 14112 9252 14176
rect 9316 14112 9322 14176
rect 11130 14152 11250 14182
rect 9006 14111 9322 14112
rect 0 13970 120 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 120 13910
rect 1485 13907 1551 13910
rect 10317 13970 10383 13973
rect 11130 13970 11250 14000
rect 10317 13968 11250 13970
rect 10317 13912 10322 13968
rect 10378 13912 11250 13968
rect 10317 13910 11250 13912
rect 10317 13907 10383 13910
rect 11130 13880 11250 13910
rect 7598 13834 7604 13836
rect 5766 13774 7604 13834
rect 4981 13698 5047 13701
rect 5574 13698 5580 13700
rect 4981 13696 5580 13698
rect 4981 13640 4986 13696
rect 5042 13640 5580 13696
rect 4981 13638 5580 13640
rect 4981 13635 5047 13638
rect 5574 13636 5580 13638
rect 5644 13636 5650 13700
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 5022 13500 5028 13564
rect 5092 13562 5098 13564
rect 5766 13562 5826 13774
rect 7598 13772 7604 13774
rect 7668 13772 7674 13836
rect 8109 13834 8175 13837
rect 8334 13834 8340 13836
rect 8109 13832 8340 13834
rect 8109 13776 8114 13832
rect 8170 13776 8340 13832
rect 8109 13774 8340 13776
rect 8109 13771 8175 13774
rect 8334 13772 8340 13774
rect 8404 13772 8410 13836
rect 9949 13698 10015 13701
rect 11130 13698 11250 13728
rect 9949 13696 11250 13698
rect 9949 13640 9954 13696
rect 10010 13640 11250 13696
rect 9949 13638 11250 13640
rect 9949 13635 10015 13638
rect 7946 13632 8262 13633
rect 7946 13568 7952 13632
rect 8016 13568 8032 13632
rect 8096 13568 8112 13632
rect 8176 13568 8192 13632
rect 8256 13568 8262 13632
rect 11130 13608 11250 13638
rect 7946 13567 8262 13568
rect 5092 13502 5826 13562
rect 5092 13500 5098 13502
rect 7414 13500 7420 13564
rect 7484 13562 7490 13564
rect 7741 13562 7807 13565
rect 7484 13560 7807 13562
rect 7484 13504 7746 13560
rect 7802 13504 7807 13560
rect 7484 13502 7807 13504
rect 7484 13500 7490 13502
rect 7741 13499 7807 13502
rect 8385 13562 8451 13565
rect 9397 13562 9463 13565
rect 8385 13560 9463 13562
rect 8385 13504 8390 13560
rect 8446 13504 9402 13560
rect 9458 13504 9463 13560
rect 8385 13502 9463 13504
rect 8385 13499 8451 13502
rect 9397 13499 9463 13502
rect 10961 13426 11027 13429
rect 11130 13426 11250 13456
rect 10961 13424 11250 13426
rect 10961 13368 10966 13424
rect 11022 13368 11250 13424
rect 10961 13366 11250 13368
rect 10961 13363 11027 13366
rect 11130 13336 11250 13366
rect 6269 13290 6335 13293
rect 9581 13290 9647 13293
rect 6269 13288 9647 13290
rect 6269 13232 6274 13288
rect 6330 13232 9586 13288
rect 9642 13232 9647 13288
rect 6269 13230 9647 13232
rect 6269 13227 6335 13230
rect 9581 13227 9647 13230
rect 9949 13290 10015 13293
rect 10409 13290 10475 13293
rect 9949 13288 10475 13290
rect 9949 13232 9954 13288
rect 10010 13232 10414 13288
rect 10470 13232 10475 13288
rect 9949 13230 10475 13232
rect 9949 13227 10015 13230
rect 10409 13227 10475 13230
rect 0 13154 120 13184
rect 1485 13154 1551 13157
rect 0 13152 1551 13154
rect 0 13096 1490 13152
rect 1546 13096 1551 13152
rect 0 13094 1551 13096
rect 0 13064 120 13094
rect 1485 13091 1551 13094
rect 9673 13154 9739 13157
rect 11130 13154 11250 13184
rect 9673 13152 11250 13154
rect 9673 13096 9678 13152
rect 9734 13096 11250 13152
rect 9673 13094 11250 13096
rect 9673 13091 9739 13094
rect 3006 13088 3322 13089
rect 3006 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3322 13088
rect 3006 13023 3322 13024
rect 9006 13088 9322 13089
rect 9006 13024 9012 13088
rect 9076 13024 9092 13088
rect 9156 13024 9172 13088
rect 9236 13024 9252 13088
rect 9316 13024 9322 13088
rect 11130 13064 11250 13094
rect 9006 13023 9322 13024
rect 7782 12956 7788 13020
rect 7852 13018 7858 13020
rect 8293 13018 8359 13021
rect 7852 13016 8359 13018
rect 7852 12960 8298 13016
rect 8354 12960 8359 13016
rect 7852 12958 8359 12960
rect 7852 12956 7858 12958
rect 8293 12955 8359 12958
rect 7925 12882 7991 12885
rect 8845 12882 8911 12885
rect 7925 12880 8911 12882
rect 7925 12824 7930 12880
rect 7986 12824 8850 12880
rect 8906 12824 8911 12880
rect 7925 12822 8911 12824
rect 7925 12819 7991 12822
rect 8845 12819 8911 12822
rect 9765 12882 9831 12885
rect 11130 12882 11250 12912
rect 9765 12880 11250 12882
rect 9765 12824 9770 12880
rect 9826 12824 11250 12880
rect 9765 12822 11250 12824
rect 9765 12819 9831 12822
rect 11130 12792 11250 12822
rect 2957 12746 3023 12749
rect 4061 12746 4127 12749
rect 4838 12746 4844 12748
rect 2957 12744 4844 12746
rect 2957 12688 2962 12744
rect 3018 12688 4066 12744
rect 4122 12688 4844 12744
rect 2957 12686 4844 12688
rect 2957 12683 3023 12686
rect 4061 12683 4127 12686
rect 4838 12684 4844 12686
rect 4908 12684 4914 12748
rect 5809 12746 5875 12749
rect 7373 12746 7439 12749
rect 7833 12746 7899 12749
rect 5809 12744 7899 12746
rect 5809 12688 5814 12744
rect 5870 12688 7378 12744
rect 7434 12688 7838 12744
rect 7894 12688 7899 12744
rect 5809 12686 7899 12688
rect 5809 12683 5875 12686
rect 7373 12683 7439 12686
rect 7833 12683 7899 12686
rect 8109 12746 8175 12749
rect 8569 12746 8635 12749
rect 8109 12744 8635 12746
rect 8109 12688 8114 12744
rect 8170 12688 8574 12744
rect 8630 12688 8635 12744
rect 8109 12686 8635 12688
rect 8109 12683 8175 12686
rect 8569 12683 8635 12686
rect 10225 12610 10291 12613
rect 11130 12610 11250 12640
rect 10225 12608 11250 12610
rect 10225 12552 10230 12608
rect 10286 12552 11250 12608
rect 10225 12550 11250 12552
rect 10225 12547 10291 12550
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 7946 12544 8262 12545
rect 7946 12480 7952 12544
rect 8016 12480 8032 12544
rect 8096 12480 8112 12544
rect 8176 12480 8192 12544
rect 8256 12480 8262 12544
rect 11130 12520 11250 12550
rect 7946 12479 8262 12480
rect 5441 12474 5507 12477
rect 5441 12472 7850 12474
rect 5441 12416 5446 12472
rect 5502 12416 7850 12472
rect 5441 12414 7850 12416
rect 5441 12411 5507 12414
rect 0 12338 120 12368
rect 1025 12338 1091 12341
rect 0 12336 1091 12338
rect 0 12280 1030 12336
rect 1086 12280 1091 12336
rect 0 12278 1091 12280
rect 7790 12338 7850 12414
rect 8201 12338 8267 12341
rect 7790 12336 8267 12338
rect 7790 12280 8206 12336
rect 8262 12280 8267 12336
rect 7790 12278 8267 12280
rect 0 12248 120 12278
rect 1025 12275 1091 12278
rect 8201 12275 8267 12278
rect 8518 12276 8524 12340
rect 8588 12338 8594 12340
rect 9121 12338 9187 12341
rect 8588 12336 9187 12338
rect 8588 12280 9126 12336
rect 9182 12280 9187 12336
rect 8588 12278 9187 12280
rect 8588 12276 8594 12278
rect 9121 12275 9187 12278
rect 9857 12338 9923 12341
rect 11130 12338 11250 12368
rect 9857 12336 11250 12338
rect 9857 12280 9862 12336
rect 9918 12280 11250 12336
rect 9857 12278 11250 12280
rect 9857 12275 9923 12278
rect 11130 12248 11250 12278
rect 3049 12202 3115 12205
rect 2822 12200 3115 12202
rect 2822 12144 3054 12200
rect 3110 12144 3115 12200
rect 2822 12142 3115 12144
rect 2822 11794 2882 12142
rect 3049 12139 3115 12142
rect 6269 12202 6335 12205
rect 6729 12202 6795 12205
rect 6269 12200 6795 12202
rect 6269 12144 6274 12200
rect 6330 12144 6734 12200
rect 6790 12144 6795 12200
rect 6269 12142 6795 12144
rect 6269 12139 6335 12142
rect 6729 12139 6795 12142
rect 9673 12066 9739 12069
rect 11130 12066 11250 12096
rect 9673 12064 11250 12066
rect 9673 12008 9678 12064
rect 9734 12008 11250 12064
rect 9673 12006 11250 12008
rect 9673 12003 9739 12006
rect 3006 12000 3322 12001
rect 3006 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3322 12000
rect 3006 11935 3322 11936
rect 9006 12000 9322 12001
rect 9006 11936 9012 12000
rect 9076 11936 9092 12000
rect 9156 11936 9172 12000
rect 9236 11936 9252 12000
rect 9316 11936 9322 12000
rect 11130 11976 11250 12006
rect 9006 11935 9322 11936
rect 4102 11868 4108 11932
rect 4172 11930 4178 11932
rect 4521 11930 4587 11933
rect 4172 11928 4587 11930
rect 4172 11872 4526 11928
rect 4582 11872 4587 11928
rect 4172 11870 4587 11872
rect 4172 11868 4178 11870
rect 4521 11867 4587 11870
rect 5257 11930 5323 11933
rect 5942 11930 5948 11932
rect 5257 11928 5948 11930
rect 5257 11872 5262 11928
rect 5318 11872 5948 11928
rect 5257 11870 5948 11872
rect 5257 11867 5323 11870
rect 5942 11868 5948 11870
rect 6012 11868 6018 11932
rect 3049 11794 3115 11797
rect 2822 11792 3115 11794
rect 2822 11736 3054 11792
rect 3110 11736 3115 11792
rect 2822 11734 3115 11736
rect 3049 11731 3115 11734
rect 7833 11794 7899 11797
rect 9622 11794 9628 11796
rect 7833 11792 9628 11794
rect 7833 11736 7838 11792
rect 7894 11736 9628 11792
rect 7833 11734 9628 11736
rect 7833 11731 7899 11734
rect 9622 11732 9628 11734
rect 9692 11732 9698 11796
rect 9765 11794 9831 11797
rect 11130 11794 11250 11824
rect 9765 11792 11250 11794
rect 9765 11736 9770 11792
rect 9826 11736 11250 11792
rect 9765 11734 11250 11736
rect 9765 11731 9831 11734
rect 11130 11704 11250 11734
rect 5993 11658 6059 11661
rect 6126 11658 6132 11660
rect 5993 11656 6132 11658
rect 5993 11600 5998 11656
rect 6054 11600 6132 11656
rect 5993 11598 6132 11600
rect 5993 11595 6059 11598
rect 6126 11596 6132 11598
rect 6196 11658 6202 11660
rect 9121 11658 9187 11661
rect 6196 11656 9187 11658
rect 6196 11600 9126 11656
rect 9182 11600 9187 11656
rect 6196 11598 9187 11600
rect 6196 11596 6202 11598
rect 9121 11595 9187 11598
rect 0 11522 120 11552
rect 1485 11522 1551 11525
rect 0 11520 1551 11522
rect 0 11464 1490 11520
rect 1546 11464 1551 11520
rect 0 11462 1551 11464
rect 0 11432 120 11462
rect 1485 11459 1551 11462
rect 8334 11460 8340 11524
rect 8404 11522 8410 11524
rect 8937 11522 9003 11525
rect 8404 11520 9003 11522
rect 8404 11464 8942 11520
rect 8998 11464 9003 11520
rect 8404 11462 9003 11464
rect 8404 11460 8410 11462
rect 8937 11459 9003 11462
rect 9765 11522 9831 11525
rect 11130 11522 11250 11552
rect 9765 11520 11250 11522
rect 9765 11464 9770 11520
rect 9826 11464 11250 11520
rect 9765 11462 11250 11464
rect 9765 11459 9831 11462
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 7946 11456 8262 11457
rect 7946 11392 7952 11456
rect 8016 11392 8032 11456
rect 8096 11392 8112 11456
rect 8176 11392 8192 11456
rect 8256 11392 8262 11456
rect 11130 11432 11250 11462
rect 7946 11391 8262 11392
rect 3734 11324 3740 11388
rect 3804 11386 3810 11388
rect 4245 11386 4311 11389
rect 3804 11384 4311 11386
rect 3804 11328 4250 11384
rect 4306 11328 4311 11384
rect 3804 11326 4311 11328
rect 3804 11324 3810 11326
rect 4245 11323 4311 11326
rect 3049 11250 3115 11253
rect 9489 11250 9555 11253
rect 3049 11248 9555 11250
rect 3049 11192 3054 11248
rect 3110 11192 9494 11248
rect 9550 11192 9555 11248
rect 3049 11190 9555 11192
rect 3049 11187 3115 11190
rect 9489 11187 9555 11190
rect 9949 11250 10015 11253
rect 11130 11250 11250 11280
rect 9949 11248 11250 11250
rect 9949 11192 9954 11248
rect 10010 11192 11250 11248
rect 9949 11190 11250 11192
rect 9949 11187 10015 11190
rect 11130 11160 11250 11190
rect 1945 11114 2011 11117
rect 3550 11114 3556 11116
rect 1945 11112 3556 11114
rect 1945 11056 1950 11112
rect 2006 11056 3556 11112
rect 1945 11054 3556 11056
rect 1945 11051 2011 11054
rect 3550 11052 3556 11054
rect 3620 11052 3626 11116
rect 790 10916 796 10980
rect 860 10978 866 10980
rect 1485 10978 1551 10981
rect 860 10976 1551 10978
rect 860 10920 1490 10976
rect 1546 10920 1551 10976
rect 860 10918 1551 10920
rect 860 10916 866 10918
rect 1485 10915 1551 10918
rect 9857 10978 9923 10981
rect 11130 10978 11250 11008
rect 9857 10976 11250 10978
rect 9857 10920 9862 10976
rect 9918 10920 11250 10976
rect 9857 10918 11250 10920
rect 9857 10915 9923 10918
rect 3006 10912 3322 10913
rect 3006 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3322 10912
rect 3006 10847 3322 10848
rect 9006 10912 9322 10913
rect 9006 10848 9012 10912
rect 9076 10848 9092 10912
rect 9156 10848 9172 10912
rect 9236 10848 9252 10912
rect 9316 10848 9322 10912
rect 11130 10888 11250 10918
rect 9006 10847 9322 10848
rect 0 10706 120 10736
rect 841 10706 907 10709
rect 0 10704 907 10706
rect 0 10648 846 10704
rect 902 10648 907 10704
rect 0 10646 907 10648
rect 0 10616 120 10646
rect 841 10643 907 10646
rect 8845 10706 8911 10709
rect 11130 10706 11250 10736
rect 8845 10704 11250 10706
rect 8845 10648 8850 10704
rect 8906 10648 11250 10704
rect 8845 10646 11250 10648
rect 8845 10643 8911 10646
rect 11130 10616 11250 10646
rect 2037 10570 2103 10573
rect 6821 10570 6887 10573
rect 2037 10568 6887 10570
rect 2037 10512 2042 10568
rect 2098 10512 6826 10568
rect 6882 10512 6887 10568
rect 2037 10510 6887 10512
rect 2037 10507 2103 10510
rect 6821 10507 6887 10510
rect 7046 10508 7052 10572
rect 7116 10570 7122 10572
rect 8477 10570 8543 10573
rect 7116 10568 8543 10570
rect 7116 10512 8482 10568
rect 8538 10512 8543 10568
rect 7116 10510 8543 10512
rect 7116 10508 7122 10510
rect 8477 10507 8543 10510
rect 9765 10434 9831 10437
rect 11130 10434 11250 10464
rect 9765 10432 11250 10434
rect 9765 10376 9770 10432
rect 9826 10376 11250 10432
rect 9765 10374 11250 10376
rect 9765 10371 9831 10374
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 7946 10368 8262 10369
rect 7946 10304 7952 10368
rect 8016 10304 8032 10368
rect 8096 10304 8112 10368
rect 8176 10304 8192 10368
rect 8256 10304 8262 10368
rect 11130 10344 11250 10374
rect 7946 10303 8262 10304
rect 1710 10100 1716 10164
rect 1780 10162 1786 10164
rect 1945 10162 2011 10165
rect 1780 10160 2011 10162
rect 1780 10104 1950 10160
rect 2006 10104 2011 10160
rect 1780 10102 2011 10104
rect 1780 10100 1786 10102
rect 1945 10099 2011 10102
rect 6678 10100 6684 10164
rect 6748 10162 6754 10164
rect 7005 10162 7071 10165
rect 6748 10160 7071 10162
rect 6748 10104 7010 10160
rect 7066 10104 7071 10160
rect 6748 10102 7071 10104
rect 6748 10100 6754 10102
rect 7005 10099 7071 10102
rect 8334 10100 8340 10164
rect 8404 10162 8410 10164
rect 8845 10162 8911 10165
rect 8404 10160 8911 10162
rect 8404 10104 8850 10160
rect 8906 10104 8911 10160
rect 8404 10102 8911 10104
rect 8404 10100 8410 10102
rect 8845 10099 8911 10102
rect 10777 10162 10843 10165
rect 11130 10162 11250 10192
rect 10777 10160 11250 10162
rect 10777 10104 10782 10160
rect 10838 10104 11250 10160
rect 10777 10102 11250 10104
rect 10777 10099 10843 10102
rect 11130 10072 11250 10102
rect 0 9890 120 9920
rect 1485 9890 1551 9893
rect 0 9888 1551 9890
rect 0 9832 1490 9888
rect 1546 9832 1551 9888
rect 0 9830 1551 9832
rect 0 9800 120 9830
rect 1485 9827 1551 9830
rect 4797 9890 4863 9893
rect 8017 9890 8083 9893
rect 4797 9888 8083 9890
rect 4797 9832 4802 9888
rect 4858 9832 8022 9888
rect 8078 9832 8083 9888
rect 4797 9830 8083 9832
rect 4797 9827 4863 9830
rect 8017 9827 8083 9830
rect 9673 9890 9739 9893
rect 11130 9890 11250 9920
rect 9673 9888 11250 9890
rect 9673 9832 9678 9888
rect 9734 9832 11250 9888
rect 9673 9830 11250 9832
rect 9673 9827 9739 9830
rect 3006 9824 3322 9825
rect 3006 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3322 9824
rect 3006 9759 3322 9760
rect 9006 9824 9322 9825
rect 9006 9760 9012 9824
rect 9076 9760 9092 9824
rect 9156 9760 9172 9824
rect 9236 9760 9252 9824
rect 9316 9760 9322 9824
rect 11130 9800 11250 9830
rect 9006 9759 9322 9760
rect 1025 9754 1091 9757
rect 2814 9754 2820 9756
rect 1025 9752 2820 9754
rect 1025 9696 1030 9752
rect 1086 9696 2820 9752
rect 1025 9694 2820 9696
rect 1025 9691 1091 9694
rect 2814 9692 2820 9694
rect 2884 9692 2890 9756
rect 3693 9754 3759 9757
rect 4654 9754 4660 9756
rect 3693 9752 4660 9754
rect 3693 9696 3698 9752
rect 3754 9696 4660 9752
rect 3693 9694 4660 9696
rect 3693 9691 3759 9694
rect 4654 9692 4660 9694
rect 4724 9692 4730 9756
rect 5349 9618 5415 9621
rect 8661 9618 8727 9621
rect 5349 9616 8727 9618
rect 5349 9560 5354 9616
rect 5410 9560 8666 9616
rect 8722 9560 8727 9616
rect 5349 9558 8727 9560
rect 5349 9555 5415 9558
rect 8661 9555 8727 9558
rect 10041 9618 10107 9621
rect 11130 9618 11250 9648
rect 10041 9616 11250 9618
rect 10041 9560 10046 9616
rect 10102 9560 11250 9616
rect 10041 9558 11250 9560
rect 10041 9555 10107 9558
rect 11130 9528 11250 9558
rect 4613 9482 4679 9485
rect 4889 9482 4955 9485
rect 6085 9482 6151 9485
rect 4613 9480 6151 9482
rect 4613 9424 4618 9480
rect 4674 9424 4894 9480
rect 4950 9424 6090 9480
rect 6146 9424 6151 9480
rect 4613 9422 6151 9424
rect 4613 9419 4679 9422
rect 4889 9419 4955 9422
rect 6085 9419 6151 9422
rect 6729 9482 6795 9485
rect 7465 9482 7531 9485
rect 9489 9484 9555 9485
rect 6729 9480 7531 9482
rect 6729 9424 6734 9480
rect 6790 9424 7470 9480
rect 7526 9424 7531 9480
rect 6729 9422 7531 9424
rect 6729 9419 6795 9422
rect 7465 9419 7531 9422
rect 9438 9420 9444 9484
rect 9508 9482 9555 9484
rect 9508 9480 9600 9482
rect 9550 9424 9600 9480
rect 9508 9422 9600 9424
rect 9508 9420 9555 9422
rect 9489 9419 9555 9420
rect 5073 9346 5139 9349
rect 6269 9346 6335 9349
rect 5073 9344 6335 9346
rect 5073 9288 5078 9344
rect 5134 9288 6274 9344
rect 6330 9288 6335 9344
rect 5073 9286 6335 9288
rect 5073 9283 5139 9286
rect 6269 9283 6335 9286
rect 10961 9346 11027 9349
rect 11130 9346 11250 9376
rect 10961 9344 11250 9346
rect 10961 9288 10966 9344
rect 11022 9288 11250 9344
rect 10961 9286 11250 9288
rect 10961 9283 11027 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 7946 9280 8262 9281
rect 7946 9216 7952 9280
rect 8016 9216 8032 9280
rect 8096 9216 8112 9280
rect 8176 9216 8192 9280
rect 8256 9216 8262 9280
rect 11130 9256 11250 9286
rect 7946 9215 8262 9216
rect 0 9074 120 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 120 9014
rect 1485 9011 1551 9014
rect 9765 9074 9831 9077
rect 11130 9074 11250 9104
rect 9765 9072 11250 9074
rect 9765 9016 9770 9072
rect 9826 9016 11250 9072
rect 9765 9014 11250 9016
rect 9765 9011 9831 9014
rect 11130 8984 11250 9014
rect 9305 8938 9371 8941
rect 9305 8936 9506 8938
rect 9305 8880 9310 8936
rect 9366 8880 9506 8936
rect 9305 8878 9506 8880
rect 9305 8875 9371 8878
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 6269 8666 6335 8669
rect 8477 8666 8543 8669
rect 6269 8664 8543 8666
rect 6269 8608 6274 8664
rect 6330 8608 8482 8664
rect 8538 8608 8543 8664
rect 6269 8606 8543 8608
rect 6269 8603 6335 8606
rect 8477 8603 8543 8606
rect 7373 8530 7439 8533
rect 8201 8530 8267 8533
rect 7373 8528 8267 8530
rect 7373 8472 7378 8528
rect 7434 8472 8206 8528
rect 8262 8472 8267 8528
rect 7373 8470 8267 8472
rect 7373 8467 7439 8470
rect 8201 8467 8267 8470
rect 9305 8530 9371 8533
rect 9446 8530 9506 8878
rect 9857 8802 9923 8805
rect 11130 8802 11250 8832
rect 9857 8800 11250 8802
rect 9857 8744 9862 8800
rect 9918 8744 11250 8800
rect 9857 8742 11250 8744
rect 9857 8739 9923 8742
rect 11130 8712 11250 8742
rect 9305 8528 9506 8530
rect 9305 8472 9310 8528
rect 9366 8472 9506 8528
rect 9305 8470 9506 8472
rect 9673 8530 9739 8533
rect 11130 8530 11250 8560
rect 9673 8528 11250 8530
rect 9673 8472 9678 8528
rect 9734 8472 11250 8528
rect 9673 8470 11250 8472
rect 9305 8467 9371 8470
rect 9673 8467 9739 8470
rect 11130 8440 11250 8470
rect 6821 8394 6887 8397
rect 8569 8394 8635 8397
rect 6821 8392 8635 8394
rect 6821 8336 6826 8392
rect 6882 8336 8574 8392
rect 8630 8336 8635 8392
rect 6821 8334 8635 8336
rect 6821 8331 6887 8334
rect 8569 8331 8635 8334
rect 0 8258 120 8288
rect 841 8258 907 8261
rect 0 8256 907 8258
rect 0 8200 846 8256
rect 902 8200 907 8256
rect 0 8198 907 8200
rect 0 8168 120 8198
rect 841 8195 907 8198
rect 2405 8260 2471 8261
rect 2405 8256 2452 8260
rect 2516 8258 2522 8260
rect 9949 8258 10015 8261
rect 11130 8258 11250 8288
rect 2405 8200 2410 8256
rect 2405 8196 2452 8200
rect 2516 8198 2562 8258
rect 9949 8256 11250 8258
rect 9949 8200 9954 8256
rect 10010 8200 11250 8256
rect 9949 8198 11250 8200
rect 2516 8196 2522 8198
rect 2405 8195 2471 8196
rect 9949 8195 10015 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 11130 8168 11250 8198
rect 7946 8127 8262 8128
rect 1158 7924 1164 7988
rect 1228 7986 1234 7988
rect 2037 7986 2103 7989
rect 1228 7984 2103 7986
rect 1228 7928 2042 7984
rect 2098 7928 2103 7984
rect 1228 7926 2103 7928
rect 1228 7924 1234 7926
rect 2037 7923 2103 7926
rect 7373 7986 7439 7989
rect 9305 7986 9371 7989
rect 7373 7984 9371 7986
rect 7373 7928 7378 7984
rect 7434 7928 9310 7984
rect 9366 7928 9371 7984
rect 7373 7926 9371 7928
rect 7373 7923 7439 7926
rect 9305 7923 9371 7926
rect 9673 7986 9739 7989
rect 11130 7986 11250 8016
rect 9673 7984 11250 7986
rect 9673 7928 9678 7984
rect 9734 7928 11250 7984
rect 9673 7926 11250 7928
rect 9673 7923 9739 7926
rect 11130 7896 11250 7926
rect 2773 7850 2839 7853
rect 8937 7850 9003 7853
rect 2773 7848 9003 7850
rect 2773 7792 2778 7848
rect 2834 7792 8942 7848
rect 8998 7792 9003 7848
rect 2773 7790 9003 7792
rect 2773 7787 2839 7790
rect 8937 7787 9003 7790
rect 9489 7716 9555 7717
rect 9438 7652 9444 7716
rect 9508 7714 9555 7716
rect 9765 7714 9831 7717
rect 11130 7714 11250 7744
rect 9508 7712 9600 7714
rect 9550 7656 9600 7712
rect 9508 7654 9600 7656
rect 9765 7712 11250 7714
rect 9765 7656 9770 7712
rect 9826 7656 11250 7712
rect 9765 7654 11250 7656
rect 9508 7652 9555 7654
rect 9489 7651 9555 7652
rect 9765 7651 9831 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 11130 7624 11250 7654
rect 9006 7583 9322 7584
rect 5390 7516 5396 7580
rect 5460 7578 5466 7580
rect 6913 7578 6979 7581
rect 5460 7576 6979 7578
rect 5460 7520 6918 7576
rect 6974 7520 6979 7576
rect 5460 7518 6979 7520
rect 5460 7516 5466 7518
rect 6913 7515 6979 7518
rect 7281 7578 7347 7581
rect 8569 7578 8635 7581
rect 7281 7576 8635 7578
rect 7281 7520 7286 7576
rect 7342 7520 8574 7576
rect 8630 7520 8635 7576
rect 7281 7518 8635 7520
rect 7281 7515 7347 7518
rect 8569 7515 8635 7518
rect 0 7442 120 7472
rect 1485 7442 1551 7445
rect 0 7440 1551 7442
rect 0 7384 1490 7440
rect 1546 7384 1551 7440
rect 0 7382 1551 7384
rect 0 7352 120 7382
rect 1485 7379 1551 7382
rect 4613 7442 4679 7445
rect 5625 7442 5691 7445
rect 4613 7440 5691 7442
rect 4613 7384 4618 7440
rect 4674 7384 5630 7440
rect 5686 7384 5691 7440
rect 4613 7382 5691 7384
rect 4613 7379 4679 7382
rect 5625 7379 5691 7382
rect 7373 7442 7439 7445
rect 8845 7442 8911 7445
rect 7373 7440 8911 7442
rect 7373 7384 7378 7440
rect 7434 7384 8850 7440
rect 8906 7384 8911 7440
rect 7373 7382 8911 7384
rect 7373 7379 7439 7382
rect 8845 7379 8911 7382
rect 9857 7442 9923 7445
rect 11130 7442 11250 7472
rect 9857 7440 11250 7442
rect 9857 7384 9862 7440
rect 9918 7384 11250 7440
rect 9857 7382 11250 7384
rect 9857 7379 9923 7382
rect 11130 7352 11250 7382
rect 8293 7306 8359 7309
rect 9489 7306 9555 7309
rect 8293 7304 9555 7306
rect 8293 7248 8298 7304
rect 8354 7248 9494 7304
rect 9550 7248 9555 7304
rect 8293 7246 9555 7248
rect 8293 7243 8359 7246
rect 9489 7243 9555 7246
rect 5717 7170 5783 7173
rect 5993 7170 6059 7173
rect 5717 7168 6059 7170
rect 5717 7112 5722 7168
rect 5778 7112 5998 7168
rect 6054 7112 6059 7168
rect 5717 7110 6059 7112
rect 5717 7107 5783 7110
rect 5993 7107 6059 7110
rect 9673 7170 9739 7173
rect 11130 7170 11250 7200
rect 9673 7168 11250 7170
rect 9673 7112 9678 7168
rect 9734 7112 11250 7168
rect 9673 7110 11250 7112
rect 9673 7107 9739 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 11130 7080 11250 7110
rect 7946 7039 8262 7040
rect 8702 6836 8708 6900
rect 8772 6898 8778 6900
rect 9397 6898 9463 6901
rect 8772 6896 9463 6898
rect 8772 6840 9402 6896
rect 9458 6840 9463 6896
rect 8772 6838 9463 6840
rect 8772 6836 8778 6838
rect 9397 6835 9463 6838
rect 9949 6898 10015 6901
rect 11130 6898 11250 6928
rect 9949 6896 11250 6898
rect 9949 6840 9954 6896
rect 10010 6840 11250 6896
rect 9949 6838 11250 6840
rect 9949 6835 10015 6838
rect 11130 6808 11250 6838
rect 9489 6762 9555 6765
rect 10910 6762 10916 6764
rect 9489 6760 10916 6762
rect 9489 6704 9494 6760
rect 9550 6704 10916 6760
rect 9489 6702 10916 6704
rect 9489 6699 9555 6702
rect 10910 6700 10916 6702
rect 10980 6700 10986 6764
rect 0 6626 120 6656
rect 1393 6626 1459 6629
rect 0 6624 1459 6626
rect 0 6568 1398 6624
rect 1454 6568 1459 6624
rect 0 6566 1459 6568
rect 0 6536 120 6566
rect 1393 6563 1459 6566
rect 9673 6626 9739 6629
rect 11130 6626 11250 6656
rect 9673 6624 11250 6626
rect 9673 6568 9678 6624
rect 9734 6568 11250 6624
rect 9673 6566 11250 6568
rect 9673 6563 9739 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 11130 6536 11250 6566
rect 9006 6495 9322 6496
rect 9765 6354 9831 6357
rect 11130 6354 11250 6384
rect 9765 6352 11250 6354
rect 9765 6296 9770 6352
rect 9826 6296 11250 6352
rect 9765 6294 11250 6296
rect 9765 6291 9831 6294
rect 11130 6264 11250 6294
rect 9765 6082 9831 6085
rect 11130 6082 11250 6112
rect 9765 6080 11250 6082
rect 9765 6024 9770 6080
rect 9826 6024 11250 6080
rect 9765 6022 11250 6024
rect 9765 6019 9831 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 11130 5992 11250 6022
rect 7946 5951 8262 5952
rect 5717 5948 5783 5949
rect 6453 5948 6519 5949
rect 5717 5946 5764 5948
rect 5672 5944 5764 5946
rect 5672 5888 5722 5944
rect 5672 5886 5764 5888
rect 5717 5884 5764 5886
rect 5828 5884 5834 5948
rect 6453 5946 6500 5948
rect 6408 5944 6500 5946
rect 6408 5888 6458 5944
rect 6408 5886 6500 5888
rect 6453 5884 6500 5886
rect 6564 5884 6570 5948
rect 5717 5883 5783 5884
rect 6453 5883 6519 5884
rect 0 5810 120 5840
rect 1853 5810 1919 5813
rect 5533 5812 5599 5813
rect 5533 5810 5580 5812
rect 0 5808 1919 5810
rect 0 5752 1858 5808
rect 1914 5752 1919 5808
rect 0 5750 1919 5752
rect 5488 5808 5580 5810
rect 5488 5752 5538 5808
rect 5488 5750 5580 5752
rect 0 5720 120 5750
rect 1853 5747 1919 5750
rect 5533 5748 5580 5750
rect 5644 5748 5650 5812
rect 10685 5810 10751 5813
rect 11130 5810 11250 5840
rect 10685 5808 11250 5810
rect 10685 5752 10690 5808
rect 10746 5752 11250 5808
rect 10685 5750 11250 5752
rect 5533 5747 5599 5748
rect 10685 5747 10751 5750
rect 11130 5720 11250 5750
rect 9673 5538 9739 5541
rect 11130 5538 11250 5568
rect 9673 5536 11250 5538
rect 9673 5480 9678 5536
rect 9734 5480 11250 5536
rect 9673 5478 11250 5480
rect 9673 5475 9739 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 11130 5448 11250 5478
rect 9006 5407 9322 5408
rect 9765 5266 9831 5269
rect 11130 5266 11250 5296
rect 9765 5264 11250 5266
rect 9765 5208 9770 5264
rect 9826 5208 11250 5264
rect 9765 5206 11250 5208
rect 9765 5203 9831 5206
rect 11130 5176 11250 5206
rect 8293 5130 8359 5133
rect 9806 5130 9812 5132
rect 8293 5128 9812 5130
rect 8293 5072 8298 5128
rect 8354 5072 9812 5128
rect 8293 5070 9812 5072
rect 8293 5067 8359 5070
rect 9806 5068 9812 5070
rect 9876 5068 9882 5132
rect 0 4994 120 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 120 4934
rect 1485 4931 1551 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 0 4178 120 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 120 4118
rect 1485 4115 1551 4118
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 3918 2620 3924 2684
rect 3988 2682 3994 2684
rect 6913 2682 6979 2685
rect 3988 2680 6979 2682
rect 3988 2624 6918 2680
rect 6974 2624 6979 2680
rect 3988 2622 6979 2624
rect 3988 2620 3994 2622
rect 6913 2619 6979 2622
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 974 1260 980 1324
rect 1044 1322 1050 1324
rect 3693 1322 3759 1325
rect 1044 1320 3759 1322
rect 1044 1264 3698 1320
rect 3754 1264 3759 1320
rect 1044 1262 3759 1264
rect 1044 1260 1050 1262
rect 3693 1259 3759 1262
rect 5073 1322 5139 1325
rect 10133 1324 10199 1325
rect 5206 1322 5212 1324
rect 5073 1320 5212 1322
rect 5073 1264 5078 1320
rect 5134 1264 5212 1320
rect 5073 1262 5212 1264
rect 5073 1259 5139 1262
rect 5206 1260 5212 1262
rect 5276 1260 5282 1324
rect 10133 1322 10180 1324
rect 10088 1320 10180 1322
rect 10088 1264 10138 1320
rect 10088 1262 10180 1264
rect 10133 1260 10180 1262
rect 10244 1260 10250 1324
rect 10133 1259 10199 1260
rect 606 1124 612 1188
rect 676 1186 682 1188
rect 4613 1186 4679 1189
rect 676 1184 4679 1186
rect 676 1128 4618 1184
rect 4674 1128 4679 1184
rect 676 1126 4679 1128
rect 676 1124 682 1126
rect 4613 1123 4679 1126
rect 4838 1124 4844 1188
rect 4908 1186 4914 1188
rect 6453 1186 6519 1189
rect 4908 1184 6519 1186
rect 4908 1128 6458 1184
rect 6514 1128 6519 1184
rect 4908 1126 6519 1128
rect 4908 1124 4914 1126
rect 6453 1123 6519 1126
rect 9213 1186 9279 1189
rect 10542 1186 10548 1188
rect 9213 1184 10548 1186
rect 9213 1128 9218 1184
rect 9274 1128 10548 1184
rect 9213 1126 10548 1128
rect 9213 1123 9279 1126
rect 10542 1124 10548 1126
rect 10612 1124 10618 1188
<< via3 >>
rect 3012 42460 3076 42464
rect 3012 42404 3016 42460
rect 3016 42404 3072 42460
rect 3072 42404 3076 42460
rect 3012 42400 3076 42404
rect 3092 42460 3156 42464
rect 3092 42404 3096 42460
rect 3096 42404 3152 42460
rect 3152 42404 3156 42460
rect 3092 42400 3156 42404
rect 3172 42460 3236 42464
rect 3172 42404 3176 42460
rect 3176 42404 3232 42460
rect 3232 42404 3236 42460
rect 3172 42400 3236 42404
rect 3252 42460 3316 42464
rect 3252 42404 3256 42460
rect 3256 42404 3312 42460
rect 3312 42404 3316 42460
rect 3252 42400 3316 42404
rect 9012 42460 9076 42464
rect 9012 42404 9016 42460
rect 9016 42404 9072 42460
rect 9072 42404 9076 42460
rect 9012 42400 9076 42404
rect 9092 42460 9156 42464
rect 9092 42404 9096 42460
rect 9096 42404 9152 42460
rect 9152 42404 9156 42460
rect 9092 42400 9156 42404
rect 9172 42460 9236 42464
rect 9172 42404 9176 42460
rect 9176 42404 9232 42460
rect 9232 42404 9236 42460
rect 9172 42400 9236 42404
rect 9252 42460 9316 42464
rect 9252 42404 9256 42460
rect 9256 42404 9312 42460
rect 9312 42404 9316 42460
rect 9252 42400 9316 42404
rect 1952 41916 2016 41920
rect 1952 41860 1956 41916
rect 1956 41860 2012 41916
rect 2012 41860 2016 41916
rect 1952 41856 2016 41860
rect 2032 41916 2096 41920
rect 2032 41860 2036 41916
rect 2036 41860 2092 41916
rect 2092 41860 2096 41916
rect 2032 41856 2096 41860
rect 2112 41916 2176 41920
rect 2112 41860 2116 41916
rect 2116 41860 2172 41916
rect 2172 41860 2176 41916
rect 2112 41856 2176 41860
rect 2192 41916 2256 41920
rect 2192 41860 2196 41916
rect 2196 41860 2252 41916
rect 2252 41860 2256 41916
rect 2192 41856 2256 41860
rect 7952 41916 8016 41920
rect 7952 41860 7956 41916
rect 7956 41860 8012 41916
rect 8012 41860 8016 41916
rect 7952 41856 8016 41860
rect 8032 41916 8096 41920
rect 8032 41860 8036 41916
rect 8036 41860 8092 41916
rect 8092 41860 8096 41916
rect 8032 41856 8096 41860
rect 8112 41916 8176 41920
rect 8112 41860 8116 41916
rect 8116 41860 8172 41916
rect 8172 41860 8176 41916
rect 8112 41856 8176 41860
rect 8192 41916 8256 41920
rect 8192 41860 8196 41916
rect 8196 41860 8252 41916
rect 8252 41860 8256 41916
rect 8192 41856 8256 41860
rect 796 41516 860 41580
rect 3012 41372 3076 41376
rect 3012 41316 3016 41372
rect 3016 41316 3072 41372
rect 3072 41316 3076 41372
rect 3012 41312 3076 41316
rect 3092 41372 3156 41376
rect 3092 41316 3096 41372
rect 3096 41316 3152 41372
rect 3152 41316 3156 41372
rect 3092 41312 3156 41316
rect 3172 41372 3236 41376
rect 3172 41316 3176 41372
rect 3176 41316 3232 41372
rect 3232 41316 3236 41372
rect 3172 41312 3236 41316
rect 3252 41372 3316 41376
rect 3252 41316 3256 41372
rect 3256 41316 3312 41372
rect 3312 41316 3316 41372
rect 3252 41312 3316 41316
rect 9012 41372 9076 41376
rect 9012 41316 9016 41372
rect 9016 41316 9072 41372
rect 9072 41316 9076 41372
rect 9012 41312 9076 41316
rect 9092 41372 9156 41376
rect 9092 41316 9096 41372
rect 9096 41316 9152 41372
rect 9152 41316 9156 41372
rect 9092 41312 9156 41316
rect 9172 41372 9236 41376
rect 9172 41316 9176 41372
rect 9176 41316 9232 41372
rect 9232 41316 9236 41372
rect 9172 41312 9236 41316
rect 9252 41372 9316 41376
rect 9252 41316 9256 41372
rect 9256 41316 9312 41372
rect 9312 41316 9316 41372
rect 9252 41312 9316 41316
rect 612 40972 676 41036
rect 1952 40828 2016 40832
rect 1952 40772 1956 40828
rect 1956 40772 2012 40828
rect 2012 40772 2016 40828
rect 1952 40768 2016 40772
rect 2032 40828 2096 40832
rect 2032 40772 2036 40828
rect 2036 40772 2092 40828
rect 2092 40772 2096 40828
rect 2032 40768 2096 40772
rect 2112 40828 2176 40832
rect 2112 40772 2116 40828
rect 2116 40772 2172 40828
rect 2172 40772 2176 40828
rect 2112 40768 2176 40772
rect 2192 40828 2256 40832
rect 2192 40772 2196 40828
rect 2196 40772 2252 40828
rect 2252 40772 2256 40828
rect 2192 40768 2256 40772
rect 7952 40828 8016 40832
rect 7952 40772 7956 40828
rect 7956 40772 8012 40828
rect 8012 40772 8016 40828
rect 7952 40768 8016 40772
rect 8032 40828 8096 40832
rect 8032 40772 8036 40828
rect 8036 40772 8092 40828
rect 8092 40772 8096 40828
rect 8032 40768 8096 40772
rect 8112 40828 8176 40832
rect 8112 40772 8116 40828
rect 8116 40772 8172 40828
rect 8172 40772 8176 40828
rect 8112 40768 8176 40772
rect 8192 40828 8256 40832
rect 8192 40772 8196 40828
rect 8196 40772 8252 40828
rect 8252 40772 8256 40828
rect 8192 40768 8256 40772
rect 7788 40352 7852 40356
rect 7788 40296 7802 40352
rect 7802 40296 7852 40352
rect 7788 40292 7852 40296
rect 9812 40352 9876 40356
rect 9812 40296 9826 40352
rect 9826 40296 9876 40352
rect 9812 40292 9876 40296
rect 3012 40284 3076 40288
rect 3012 40228 3016 40284
rect 3016 40228 3072 40284
rect 3072 40228 3076 40284
rect 3012 40224 3076 40228
rect 3092 40284 3156 40288
rect 3092 40228 3096 40284
rect 3096 40228 3152 40284
rect 3152 40228 3156 40284
rect 3092 40224 3156 40228
rect 3172 40284 3236 40288
rect 3172 40228 3176 40284
rect 3176 40228 3232 40284
rect 3232 40228 3236 40284
rect 3172 40224 3236 40228
rect 3252 40284 3316 40288
rect 3252 40228 3256 40284
rect 3256 40228 3312 40284
rect 3312 40228 3316 40284
rect 3252 40224 3316 40228
rect 9012 40284 9076 40288
rect 9012 40228 9016 40284
rect 9016 40228 9072 40284
rect 9072 40228 9076 40284
rect 9012 40224 9076 40228
rect 9092 40284 9156 40288
rect 9092 40228 9096 40284
rect 9096 40228 9152 40284
rect 9152 40228 9156 40284
rect 9092 40224 9156 40228
rect 9172 40284 9236 40288
rect 9172 40228 9176 40284
rect 9176 40228 9232 40284
rect 9232 40228 9236 40284
rect 9172 40224 9236 40228
rect 9252 40284 9316 40288
rect 9252 40228 9256 40284
rect 9256 40228 9312 40284
rect 9312 40228 9316 40284
rect 9252 40224 9316 40228
rect 10180 40156 10244 40220
rect 5212 40020 5276 40084
rect 1952 39740 2016 39744
rect 1952 39684 1956 39740
rect 1956 39684 2012 39740
rect 2012 39684 2016 39740
rect 1952 39680 2016 39684
rect 2032 39740 2096 39744
rect 2032 39684 2036 39740
rect 2036 39684 2092 39740
rect 2092 39684 2096 39740
rect 2032 39680 2096 39684
rect 2112 39740 2176 39744
rect 2112 39684 2116 39740
rect 2116 39684 2172 39740
rect 2172 39684 2176 39740
rect 2112 39680 2176 39684
rect 2192 39740 2256 39744
rect 2192 39684 2196 39740
rect 2196 39684 2252 39740
rect 2252 39684 2256 39740
rect 2192 39680 2256 39684
rect 7952 39740 8016 39744
rect 7952 39684 7956 39740
rect 7956 39684 8012 39740
rect 8012 39684 8016 39740
rect 7952 39680 8016 39684
rect 8032 39740 8096 39744
rect 8032 39684 8036 39740
rect 8036 39684 8092 39740
rect 8092 39684 8096 39740
rect 8032 39680 8096 39684
rect 8112 39740 8176 39744
rect 8112 39684 8116 39740
rect 8116 39684 8172 39740
rect 8172 39684 8176 39740
rect 8112 39680 8176 39684
rect 8192 39740 8256 39744
rect 8192 39684 8196 39740
rect 8196 39684 8252 39740
rect 8252 39684 8256 39740
rect 8192 39680 8256 39684
rect 10548 39612 10612 39676
rect 980 39476 1044 39540
rect 8708 39340 8772 39404
rect 3012 39196 3076 39200
rect 3012 39140 3016 39196
rect 3016 39140 3072 39196
rect 3072 39140 3076 39196
rect 3012 39136 3076 39140
rect 3092 39196 3156 39200
rect 3092 39140 3096 39196
rect 3096 39140 3152 39196
rect 3152 39140 3156 39196
rect 3092 39136 3156 39140
rect 3172 39196 3236 39200
rect 3172 39140 3176 39196
rect 3176 39140 3232 39196
rect 3232 39140 3236 39196
rect 3172 39136 3236 39140
rect 3252 39196 3316 39200
rect 3252 39140 3256 39196
rect 3256 39140 3312 39196
rect 3312 39140 3316 39196
rect 3252 39136 3316 39140
rect 9012 39196 9076 39200
rect 9012 39140 9016 39196
rect 9016 39140 9072 39196
rect 9072 39140 9076 39196
rect 9012 39136 9076 39140
rect 9092 39196 9156 39200
rect 9092 39140 9096 39196
rect 9096 39140 9152 39196
rect 9152 39140 9156 39196
rect 9092 39136 9156 39140
rect 9172 39196 9236 39200
rect 9172 39140 9176 39196
rect 9176 39140 9232 39196
rect 9232 39140 9236 39196
rect 9172 39136 9236 39140
rect 9252 39196 9316 39200
rect 9252 39140 9256 39196
rect 9256 39140 9312 39196
rect 9312 39140 9316 39196
rect 9252 39136 9316 39140
rect 5948 38796 6012 38860
rect 8340 38660 8404 38724
rect 1952 38652 2016 38656
rect 1952 38596 1956 38652
rect 1956 38596 2012 38652
rect 2012 38596 2016 38652
rect 1952 38592 2016 38596
rect 2032 38652 2096 38656
rect 2032 38596 2036 38652
rect 2036 38596 2092 38652
rect 2092 38596 2096 38652
rect 2032 38592 2096 38596
rect 2112 38652 2176 38656
rect 2112 38596 2116 38652
rect 2116 38596 2172 38652
rect 2172 38596 2176 38652
rect 2112 38592 2176 38596
rect 2192 38652 2256 38656
rect 2192 38596 2196 38652
rect 2196 38596 2252 38652
rect 2252 38596 2256 38652
rect 2192 38592 2256 38596
rect 7952 38652 8016 38656
rect 7952 38596 7956 38652
rect 7956 38596 8012 38652
rect 8012 38596 8016 38652
rect 7952 38592 8016 38596
rect 8032 38652 8096 38656
rect 8032 38596 8036 38652
rect 8036 38596 8092 38652
rect 8092 38596 8096 38652
rect 8032 38592 8096 38596
rect 8112 38652 8176 38656
rect 8112 38596 8116 38652
rect 8116 38596 8172 38652
rect 8172 38596 8176 38652
rect 8112 38592 8176 38596
rect 8192 38652 8256 38656
rect 8192 38596 8196 38652
rect 8196 38596 8252 38652
rect 8252 38596 8256 38652
rect 8192 38592 8256 38596
rect 10364 38252 10428 38316
rect 3012 38108 3076 38112
rect 3012 38052 3016 38108
rect 3016 38052 3072 38108
rect 3072 38052 3076 38108
rect 3012 38048 3076 38052
rect 3092 38108 3156 38112
rect 3092 38052 3096 38108
rect 3096 38052 3152 38108
rect 3152 38052 3156 38108
rect 3092 38048 3156 38052
rect 3172 38108 3236 38112
rect 3172 38052 3176 38108
rect 3176 38052 3232 38108
rect 3232 38052 3236 38108
rect 3172 38048 3236 38052
rect 3252 38108 3316 38112
rect 3252 38052 3256 38108
rect 3256 38052 3312 38108
rect 3312 38052 3316 38108
rect 3252 38048 3316 38052
rect 9012 38108 9076 38112
rect 9012 38052 9016 38108
rect 9016 38052 9072 38108
rect 9072 38052 9076 38108
rect 9012 38048 9076 38052
rect 9092 38108 9156 38112
rect 9092 38052 9096 38108
rect 9096 38052 9152 38108
rect 9152 38052 9156 38108
rect 9092 38048 9156 38052
rect 9172 38108 9236 38112
rect 9172 38052 9176 38108
rect 9176 38052 9232 38108
rect 9232 38052 9236 38108
rect 9172 38048 9236 38052
rect 9252 38108 9316 38112
rect 9252 38052 9256 38108
rect 9256 38052 9312 38108
rect 9312 38052 9316 38108
rect 9252 38048 9316 38052
rect 4476 37708 4540 37772
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 7952 37564 8016 37568
rect 7952 37508 7956 37564
rect 7956 37508 8012 37564
rect 8012 37508 8016 37564
rect 7952 37504 8016 37508
rect 8032 37564 8096 37568
rect 8032 37508 8036 37564
rect 8036 37508 8092 37564
rect 8092 37508 8096 37564
rect 8032 37504 8096 37508
rect 8112 37564 8176 37568
rect 8112 37508 8116 37564
rect 8116 37508 8172 37564
rect 8172 37508 8176 37564
rect 8112 37504 8176 37508
rect 8192 37564 8256 37568
rect 8192 37508 8196 37564
rect 8196 37508 8252 37564
rect 8252 37508 8256 37564
rect 8192 37504 8256 37508
rect 6500 37300 6564 37364
rect 5028 37224 5092 37228
rect 5028 37168 5042 37224
rect 5042 37168 5092 37224
rect 5028 37164 5092 37168
rect 6868 37164 6932 37228
rect 3012 37020 3076 37024
rect 3012 36964 3016 37020
rect 3016 36964 3072 37020
rect 3072 36964 3076 37020
rect 3012 36960 3076 36964
rect 3092 37020 3156 37024
rect 3092 36964 3096 37020
rect 3096 36964 3152 37020
rect 3152 36964 3156 37020
rect 3092 36960 3156 36964
rect 3172 37020 3236 37024
rect 3172 36964 3176 37020
rect 3176 36964 3232 37020
rect 3232 36964 3236 37020
rect 3172 36960 3236 36964
rect 3252 37020 3316 37024
rect 3252 36964 3256 37020
rect 3256 36964 3312 37020
rect 3312 36964 3316 37020
rect 3252 36960 3316 36964
rect 9012 37020 9076 37024
rect 9012 36964 9016 37020
rect 9016 36964 9072 37020
rect 9072 36964 9076 37020
rect 9012 36960 9076 36964
rect 9092 37020 9156 37024
rect 9092 36964 9096 37020
rect 9096 36964 9152 37020
rect 9152 36964 9156 37020
rect 9092 36960 9156 36964
rect 9172 37020 9236 37024
rect 9172 36964 9176 37020
rect 9176 36964 9232 37020
rect 9232 36964 9236 37020
rect 9172 36960 9236 36964
rect 9252 37020 9316 37024
rect 9252 36964 9256 37020
rect 9256 36964 9312 37020
rect 9312 36964 9316 37020
rect 9252 36960 9316 36964
rect 4660 36756 4724 36820
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 7952 36476 8016 36480
rect 7952 36420 7956 36476
rect 7956 36420 8012 36476
rect 8012 36420 8016 36476
rect 7952 36416 8016 36420
rect 8032 36476 8096 36480
rect 8032 36420 8036 36476
rect 8036 36420 8092 36476
rect 8092 36420 8096 36476
rect 8032 36416 8096 36420
rect 8112 36476 8176 36480
rect 8112 36420 8116 36476
rect 8116 36420 8172 36476
rect 8172 36420 8176 36476
rect 8112 36416 8176 36420
rect 8192 36476 8256 36480
rect 8192 36420 8196 36476
rect 8196 36420 8252 36476
rect 8252 36420 8256 36476
rect 8192 36416 8256 36420
rect 3740 36076 3804 36140
rect 1532 35804 1596 35868
rect 3012 35932 3076 35936
rect 3012 35876 3016 35932
rect 3016 35876 3072 35932
rect 3072 35876 3076 35932
rect 3012 35872 3076 35876
rect 3092 35932 3156 35936
rect 3092 35876 3096 35932
rect 3096 35876 3152 35932
rect 3152 35876 3156 35932
rect 3092 35872 3156 35876
rect 3172 35932 3236 35936
rect 3172 35876 3176 35932
rect 3176 35876 3232 35932
rect 3232 35876 3236 35932
rect 3172 35872 3236 35876
rect 3252 35932 3316 35936
rect 3252 35876 3256 35932
rect 3256 35876 3312 35932
rect 3312 35876 3316 35932
rect 3252 35872 3316 35876
rect 9012 35932 9076 35936
rect 9012 35876 9016 35932
rect 9016 35876 9072 35932
rect 9072 35876 9076 35932
rect 9012 35872 9076 35876
rect 9092 35932 9156 35936
rect 9092 35876 9096 35932
rect 9096 35876 9152 35932
rect 9152 35876 9156 35932
rect 9092 35872 9156 35876
rect 9172 35932 9236 35936
rect 9172 35876 9176 35932
rect 9176 35876 9232 35932
rect 9232 35876 9236 35932
rect 9172 35872 9236 35876
rect 9252 35932 9316 35936
rect 9252 35876 9256 35932
rect 9256 35876 9312 35932
rect 9312 35876 9316 35932
rect 9252 35872 9316 35876
rect 7420 35804 7484 35868
rect 8524 35864 8588 35868
rect 8524 35808 8574 35864
rect 8574 35808 8588 35864
rect 8524 35804 8588 35808
rect 2636 35668 2700 35732
rect 7788 35668 7852 35732
rect 9996 35668 10060 35732
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 7952 35388 8016 35392
rect 7952 35332 7956 35388
rect 7956 35332 8012 35388
rect 8012 35332 8016 35388
rect 7952 35328 8016 35332
rect 8032 35388 8096 35392
rect 8032 35332 8036 35388
rect 8036 35332 8092 35388
rect 8092 35332 8096 35388
rect 8032 35328 8096 35332
rect 8112 35388 8176 35392
rect 8112 35332 8116 35388
rect 8116 35332 8172 35388
rect 8172 35332 8176 35388
rect 8112 35328 8176 35332
rect 8192 35388 8256 35392
rect 8192 35332 8196 35388
rect 8196 35332 8252 35388
rect 8252 35332 8256 35388
rect 8192 35328 8256 35332
rect 5396 35124 5460 35188
rect 9444 35124 9508 35188
rect 3012 34844 3076 34848
rect 3012 34788 3016 34844
rect 3016 34788 3072 34844
rect 3072 34788 3076 34844
rect 3012 34784 3076 34788
rect 3092 34844 3156 34848
rect 3092 34788 3096 34844
rect 3096 34788 3152 34844
rect 3152 34788 3156 34844
rect 3092 34784 3156 34788
rect 3172 34844 3236 34848
rect 3172 34788 3176 34844
rect 3176 34788 3232 34844
rect 3232 34788 3236 34844
rect 3172 34784 3236 34788
rect 3252 34844 3316 34848
rect 3252 34788 3256 34844
rect 3256 34788 3312 34844
rect 3312 34788 3316 34844
rect 3252 34784 3316 34788
rect 9012 34844 9076 34848
rect 9012 34788 9016 34844
rect 9016 34788 9072 34844
rect 9072 34788 9076 34844
rect 9012 34784 9076 34788
rect 9092 34844 9156 34848
rect 9092 34788 9096 34844
rect 9096 34788 9152 34844
rect 9152 34788 9156 34844
rect 9092 34784 9156 34788
rect 9172 34844 9236 34848
rect 9172 34788 9176 34844
rect 9176 34788 9232 34844
rect 9232 34788 9236 34844
rect 9172 34784 9236 34788
rect 9252 34844 9316 34848
rect 9252 34788 9256 34844
rect 9256 34788 9312 34844
rect 9312 34788 9316 34844
rect 9252 34784 9316 34788
rect 3556 34580 3620 34644
rect 2452 34444 2516 34508
rect 7052 34444 7116 34508
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 7952 34300 8016 34304
rect 7952 34244 7956 34300
rect 7956 34244 8012 34300
rect 8012 34244 8016 34300
rect 7952 34240 8016 34244
rect 8032 34300 8096 34304
rect 8032 34244 8036 34300
rect 8036 34244 8092 34300
rect 8092 34244 8096 34300
rect 8032 34240 8096 34244
rect 8112 34300 8176 34304
rect 8112 34244 8116 34300
rect 8116 34244 8172 34300
rect 8172 34244 8176 34300
rect 8112 34240 8176 34244
rect 8192 34300 8256 34304
rect 8192 34244 8196 34300
rect 8196 34244 8252 34300
rect 8252 34244 8256 34300
rect 8192 34240 8256 34244
rect 6868 34232 6932 34236
rect 6868 34176 6882 34232
rect 6882 34176 6932 34232
rect 6868 34172 6932 34176
rect 6316 33900 6380 33964
rect 3012 33756 3076 33760
rect 3012 33700 3016 33756
rect 3016 33700 3072 33756
rect 3072 33700 3076 33756
rect 3012 33696 3076 33700
rect 3092 33756 3156 33760
rect 3092 33700 3096 33756
rect 3096 33700 3152 33756
rect 3152 33700 3156 33756
rect 3092 33696 3156 33700
rect 3172 33756 3236 33760
rect 3172 33700 3176 33756
rect 3176 33700 3232 33756
rect 3232 33700 3236 33756
rect 3172 33696 3236 33700
rect 3252 33756 3316 33760
rect 3252 33700 3256 33756
rect 3256 33700 3312 33756
rect 3312 33700 3316 33756
rect 3252 33696 3316 33700
rect 9012 33756 9076 33760
rect 9012 33700 9016 33756
rect 9016 33700 9072 33756
rect 9072 33700 9076 33756
rect 9012 33696 9076 33700
rect 9092 33756 9156 33760
rect 9092 33700 9096 33756
rect 9096 33700 9152 33756
rect 9152 33700 9156 33756
rect 9092 33696 9156 33700
rect 9172 33756 9236 33760
rect 9172 33700 9176 33756
rect 9176 33700 9232 33756
rect 9232 33700 9236 33756
rect 9172 33696 9236 33700
rect 9252 33756 9316 33760
rect 9252 33700 9256 33756
rect 9256 33700 9312 33756
rect 9312 33700 9316 33756
rect 9252 33696 9316 33700
rect 4292 33356 4356 33420
rect 5580 33356 5644 33420
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 2820 33084 2884 33148
rect 7952 33212 8016 33216
rect 7952 33156 7956 33212
rect 7956 33156 8012 33212
rect 8012 33156 8016 33212
rect 7952 33152 8016 33156
rect 8032 33212 8096 33216
rect 8032 33156 8036 33212
rect 8036 33156 8092 33212
rect 8092 33156 8096 33212
rect 8032 33152 8096 33156
rect 8112 33212 8176 33216
rect 8112 33156 8116 33212
rect 8116 33156 8172 33212
rect 8172 33156 8176 33212
rect 8112 33152 8176 33156
rect 8192 33212 8256 33216
rect 8192 33156 8196 33212
rect 8196 33156 8252 33212
rect 8252 33156 8256 33212
rect 8192 33152 8256 33156
rect 3924 32948 3988 33012
rect 8524 32948 8588 33012
rect 1716 32872 1780 32876
rect 1716 32816 1730 32872
rect 1730 32816 1780 32872
rect 1716 32812 1780 32816
rect 5764 32812 5828 32876
rect 7788 32676 7852 32740
rect 3012 32668 3076 32672
rect 3012 32612 3016 32668
rect 3016 32612 3072 32668
rect 3072 32612 3076 32668
rect 3012 32608 3076 32612
rect 3092 32668 3156 32672
rect 3092 32612 3096 32668
rect 3096 32612 3152 32668
rect 3152 32612 3156 32668
rect 3092 32608 3156 32612
rect 3172 32668 3236 32672
rect 3172 32612 3176 32668
rect 3176 32612 3232 32668
rect 3232 32612 3236 32668
rect 3172 32608 3236 32612
rect 3252 32668 3316 32672
rect 3252 32612 3256 32668
rect 3256 32612 3312 32668
rect 3312 32612 3316 32668
rect 3252 32608 3316 32612
rect 9012 32668 9076 32672
rect 9012 32612 9016 32668
rect 9016 32612 9072 32668
rect 9072 32612 9076 32668
rect 9012 32608 9076 32612
rect 9092 32668 9156 32672
rect 9092 32612 9096 32668
rect 9096 32612 9152 32668
rect 9152 32612 9156 32668
rect 9092 32608 9156 32612
rect 9172 32668 9236 32672
rect 9172 32612 9176 32668
rect 9176 32612 9232 32668
rect 9232 32612 9236 32668
rect 9172 32608 9236 32612
rect 9252 32668 9316 32672
rect 9252 32612 9256 32668
rect 9256 32612 9312 32668
rect 9312 32612 9316 32668
rect 9252 32608 9316 32612
rect 7604 32268 7668 32332
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 7952 32124 8016 32128
rect 7952 32068 7956 32124
rect 7956 32068 8012 32124
rect 8012 32068 8016 32124
rect 7952 32064 8016 32068
rect 8032 32124 8096 32128
rect 8032 32068 8036 32124
rect 8036 32068 8092 32124
rect 8092 32068 8096 32124
rect 8032 32064 8096 32068
rect 8112 32124 8176 32128
rect 8112 32068 8116 32124
rect 8116 32068 8172 32124
rect 8172 32068 8176 32124
rect 8112 32064 8176 32068
rect 8192 32124 8256 32128
rect 8192 32068 8196 32124
rect 8196 32068 8252 32124
rect 8252 32068 8256 32124
rect 8192 32064 8256 32068
rect 2636 31860 2700 31924
rect 6132 31724 6196 31788
rect 7236 31784 7300 31788
rect 7236 31728 7250 31784
rect 7250 31728 7300 31784
rect 7236 31724 7300 31728
rect 244 31588 308 31652
rect 3012 31580 3076 31584
rect 3012 31524 3016 31580
rect 3016 31524 3072 31580
rect 3072 31524 3076 31580
rect 3012 31520 3076 31524
rect 3092 31580 3156 31584
rect 3092 31524 3096 31580
rect 3096 31524 3152 31580
rect 3152 31524 3156 31580
rect 3092 31520 3156 31524
rect 3172 31580 3236 31584
rect 3172 31524 3176 31580
rect 3176 31524 3232 31580
rect 3232 31524 3236 31580
rect 3172 31520 3236 31524
rect 3252 31580 3316 31584
rect 3252 31524 3256 31580
rect 3256 31524 3312 31580
rect 3312 31524 3316 31580
rect 3252 31520 3316 31524
rect 9012 31580 9076 31584
rect 9012 31524 9016 31580
rect 9016 31524 9072 31580
rect 9072 31524 9076 31580
rect 9012 31520 9076 31524
rect 9092 31580 9156 31584
rect 9092 31524 9096 31580
rect 9096 31524 9152 31580
rect 9152 31524 9156 31580
rect 9092 31520 9156 31524
rect 9172 31580 9236 31584
rect 9172 31524 9176 31580
rect 9176 31524 9232 31580
rect 9232 31524 9236 31580
rect 9172 31520 9236 31524
rect 9252 31580 9316 31584
rect 9252 31524 9256 31580
rect 9256 31524 9312 31580
rect 9312 31524 9316 31580
rect 9252 31520 9316 31524
rect 4292 31452 4356 31516
rect 7236 31452 7300 31516
rect 8524 31452 8588 31516
rect 4844 31316 4908 31380
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 7952 31036 8016 31040
rect 7952 30980 7956 31036
rect 7956 30980 8012 31036
rect 8012 30980 8016 31036
rect 7952 30976 8016 30980
rect 8032 31036 8096 31040
rect 8032 30980 8036 31036
rect 8036 30980 8092 31036
rect 8092 30980 8096 31036
rect 8032 30976 8096 30980
rect 8112 31036 8176 31040
rect 8112 30980 8116 31036
rect 8116 30980 8172 31036
rect 8172 30980 8176 31036
rect 8112 30976 8176 30980
rect 8192 31036 8256 31040
rect 8192 30980 8196 31036
rect 8196 30980 8252 31036
rect 8252 30980 8256 31036
rect 8192 30976 8256 30980
rect 9628 30908 9692 30972
rect 5580 30500 5644 30564
rect 3012 30492 3076 30496
rect 3012 30436 3016 30492
rect 3016 30436 3072 30492
rect 3072 30436 3076 30492
rect 3012 30432 3076 30436
rect 3092 30492 3156 30496
rect 3092 30436 3096 30492
rect 3096 30436 3152 30492
rect 3152 30436 3156 30492
rect 3092 30432 3156 30436
rect 3172 30492 3236 30496
rect 3172 30436 3176 30492
rect 3176 30436 3232 30492
rect 3232 30436 3236 30492
rect 3172 30432 3236 30436
rect 3252 30492 3316 30496
rect 3252 30436 3256 30492
rect 3256 30436 3312 30492
rect 3312 30436 3316 30492
rect 3252 30432 3316 30436
rect 9012 30492 9076 30496
rect 9012 30436 9016 30492
rect 9016 30436 9072 30492
rect 9072 30436 9076 30492
rect 9012 30432 9076 30436
rect 9092 30492 9156 30496
rect 9092 30436 9096 30492
rect 9096 30436 9152 30492
rect 9152 30436 9156 30492
rect 9092 30432 9156 30436
rect 9172 30492 9236 30496
rect 9172 30436 9176 30492
rect 9176 30436 9232 30492
rect 9232 30436 9236 30492
rect 9172 30432 9236 30436
rect 9252 30492 9316 30496
rect 9252 30436 9256 30492
rect 9256 30436 9312 30492
rect 9312 30436 9316 30492
rect 9252 30432 9316 30436
rect 2820 30364 2884 30428
rect 4108 30424 4172 30428
rect 4108 30368 4122 30424
rect 4122 30368 4172 30424
rect 4108 30364 4172 30368
rect 6500 30364 6564 30428
rect 8340 30364 8404 30428
rect 2452 30228 2516 30292
rect 4292 30228 4356 30292
rect 7052 30228 7116 30292
rect 3924 30092 3988 30156
rect 7052 30092 7116 30156
rect 4660 29956 4724 30020
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 7952 29948 8016 29952
rect 7952 29892 7956 29948
rect 7956 29892 8012 29948
rect 8012 29892 8016 29948
rect 7952 29888 8016 29892
rect 8032 29948 8096 29952
rect 8032 29892 8036 29948
rect 8036 29892 8092 29948
rect 8092 29892 8096 29948
rect 8032 29888 8096 29892
rect 8112 29948 8176 29952
rect 8112 29892 8116 29948
rect 8116 29892 8172 29948
rect 8172 29892 8176 29948
rect 8112 29888 8176 29892
rect 8192 29948 8256 29952
rect 8192 29892 8196 29948
rect 8196 29892 8252 29948
rect 8252 29892 8256 29948
rect 8192 29888 8256 29892
rect 7788 29684 7852 29748
rect 4660 29608 4724 29612
rect 4660 29552 4710 29608
rect 4710 29552 4724 29608
rect 4660 29548 4724 29552
rect 5028 29412 5092 29476
rect 3012 29404 3076 29408
rect 3012 29348 3016 29404
rect 3016 29348 3072 29404
rect 3072 29348 3076 29404
rect 3012 29344 3076 29348
rect 3092 29404 3156 29408
rect 3092 29348 3096 29404
rect 3096 29348 3152 29404
rect 3152 29348 3156 29404
rect 3092 29344 3156 29348
rect 3172 29404 3236 29408
rect 3172 29348 3176 29404
rect 3176 29348 3232 29404
rect 3232 29348 3236 29404
rect 3172 29344 3236 29348
rect 3252 29404 3316 29408
rect 3252 29348 3256 29404
rect 3256 29348 3312 29404
rect 3312 29348 3316 29404
rect 3252 29344 3316 29348
rect 9012 29404 9076 29408
rect 9012 29348 9016 29404
rect 9016 29348 9072 29404
rect 9072 29348 9076 29404
rect 9012 29344 9076 29348
rect 9092 29404 9156 29408
rect 9092 29348 9096 29404
rect 9096 29348 9152 29404
rect 9152 29348 9156 29404
rect 9092 29344 9156 29348
rect 9172 29404 9236 29408
rect 9172 29348 9176 29404
rect 9176 29348 9232 29404
rect 9232 29348 9236 29404
rect 9172 29344 9236 29348
rect 9252 29404 9316 29408
rect 9252 29348 9256 29404
rect 9256 29348 9312 29404
rect 9312 29348 9316 29404
rect 9252 29344 9316 29348
rect 1716 29140 1780 29204
rect 6868 29276 6932 29340
rect 1716 28928 1780 28932
rect 1716 28872 1730 28928
rect 1730 28872 1780 28928
rect 1716 28868 1780 28872
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 1164 28596 1228 28660
rect 1348 28460 1412 28524
rect 3012 28316 3076 28320
rect 3012 28260 3016 28316
rect 3016 28260 3072 28316
rect 3072 28260 3076 28316
rect 3012 28256 3076 28260
rect 3092 28316 3156 28320
rect 3092 28260 3096 28316
rect 3096 28260 3152 28316
rect 3152 28260 3156 28316
rect 3092 28256 3156 28260
rect 3172 28316 3236 28320
rect 3172 28260 3176 28316
rect 3176 28260 3232 28316
rect 3232 28260 3236 28316
rect 3172 28256 3236 28260
rect 3252 28316 3316 28320
rect 3252 28260 3256 28316
rect 3256 28260 3312 28316
rect 3312 28260 3316 28316
rect 3252 28256 3316 28260
rect 2636 28052 2700 28116
rect 2636 27916 2700 27980
rect 7952 28860 8016 28864
rect 7952 28804 7956 28860
rect 7956 28804 8012 28860
rect 8012 28804 8016 28860
rect 7952 28800 8016 28804
rect 8032 28860 8096 28864
rect 8032 28804 8036 28860
rect 8036 28804 8092 28860
rect 8092 28804 8096 28860
rect 8032 28800 8096 28804
rect 8112 28860 8176 28864
rect 8112 28804 8116 28860
rect 8116 28804 8172 28860
rect 8172 28804 8176 28860
rect 8112 28800 8176 28804
rect 8192 28860 8256 28864
rect 8192 28804 8196 28860
rect 8196 28804 8252 28860
rect 8252 28804 8256 28860
rect 8192 28800 8256 28804
rect 10916 28732 10980 28796
rect 6500 28656 6564 28660
rect 6500 28600 6550 28656
rect 6550 28600 6564 28656
rect 6500 28596 6564 28600
rect 7236 28656 7300 28660
rect 7236 28600 7250 28656
rect 7250 28600 7300 28656
rect 7236 28596 7300 28600
rect 8340 28596 8404 28660
rect 6684 28460 6748 28524
rect 9012 28316 9076 28320
rect 9012 28260 9016 28316
rect 9016 28260 9072 28316
rect 9072 28260 9076 28316
rect 9012 28256 9076 28260
rect 9092 28316 9156 28320
rect 9092 28260 9096 28316
rect 9096 28260 9152 28316
rect 9152 28260 9156 28316
rect 9092 28256 9156 28260
rect 9172 28316 9236 28320
rect 9172 28260 9176 28316
rect 9176 28260 9232 28316
rect 9232 28260 9236 28316
rect 9172 28256 9236 28260
rect 9252 28316 9316 28320
rect 9252 28260 9256 28316
rect 9256 28260 9312 28316
rect 9312 28260 9316 28316
rect 9252 28256 9316 28260
rect 7420 28188 7484 28252
rect 9444 28112 9508 28116
rect 9444 28056 9494 28112
rect 9494 28056 9508 28112
rect 9444 28052 9508 28056
rect 5580 27976 5644 27980
rect 5580 27920 5594 27976
rect 5594 27920 5644 27976
rect 5580 27916 5644 27920
rect 7788 27916 7852 27980
rect 9628 27916 9692 27980
rect 7236 27780 7300 27844
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 7952 27772 8016 27776
rect 7952 27716 7956 27772
rect 7956 27716 8012 27772
rect 8012 27716 8016 27772
rect 7952 27712 8016 27716
rect 8032 27772 8096 27776
rect 8032 27716 8036 27772
rect 8036 27716 8092 27772
rect 8092 27716 8096 27772
rect 8032 27712 8096 27716
rect 8112 27772 8176 27776
rect 8112 27716 8116 27772
rect 8116 27716 8172 27772
rect 8172 27716 8176 27772
rect 8112 27712 8176 27716
rect 8192 27772 8256 27776
rect 8192 27716 8196 27772
rect 8196 27716 8252 27772
rect 8252 27716 8256 27772
rect 8192 27712 8256 27716
rect 3924 27644 3988 27708
rect 9444 27704 9508 27708
rect 9444 27648 9458 27704
rect 9458 27648 9508 27704
rect 9444 27644 9508 27648
rect 3740 27508 3804 27572
rect 8708 27568 8772 27572
rect 8708 27512 8758 27568
rect 8758 27512 8772 27568
rect 8708 27508 8772 27512
rect 2820 27372 2884 27436
rect 5028 27372 5092 27436
rect 8524 27372 8588 27436
rect 3012 27228 3076 27232
rect 3012 27172 3016 27228
rect 3016 27172 3072 27228
rect 3072 27172 3076 27228
rect 3012 27168 3076 27172
rect 3092 27228 3156 27232
rect 3092 27172 3096 27228
rect 3096 27172 3152 27228
rect 3152 27172 3156 27228
rect 3092 27168 3156 27172
rect 3172 27228 3236 27232
rect 3172 27172 3176 27228
rect 3176 27172 3232 27228
rect 3232 27172 3236 27228
rect 3172 27168 3236 27172
rect 3252 27228 3316 27232
rect 3252 27172 3256 27228
rect 3256 27172 3312 27228
rect 3312 27172 3316 27228
rect 3252 27168 3316 27172
rect 9012 27228 9076 27232
rect 9012 27172 9016 27228
rect 9016 27172 9072 27228
rect 9072 27172 9076 27228
rect 9012 27168 9076 27172
rect 9092 27228 9156 27232
rect 9092 27172 9096 27228
rect 9096 27172 9152 27228
rect 9152 27172 9156 27228
rect 9092 27168 9156 27172
rect 9172 27228 9236 27232
rect 9172 27172 9176 27228
rect 9176 27172 9232 27228
rect 9232 27172 9236 27228
rect 9172 27168 9236 27172
rect 9252 27228 9316 27232
rect 9252 27172 9256 27228
rect 9256 27172 9312 27228
rect 9312 27172 9316 27228
rect 9252 27168 9316 27172
rect 3556 26964 3620 27028
rect 3556 26828 3620 26892
rect 4108 26828 4172 26892
rect 8708 26828 8772 26892
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 7952 26684 8016 26688
rect 7952 26628 7956 26684
rect 7956 26628 8012 26684
rect 8012 26628 8016 26684
rect 7952 26624 8016 26628
rect 8032 26684 8096 26688
rect 8032 26628 8036 26684
rect 8036 26628 8092 26684
rect 8092 26628 8096 26684
rect 8032 26624 8096 26628
rect 8112 26684 8176 26688
rect 8112 26628 8116 26684
rect 8116 26628 8172 26684
rect 8172 26628 8176 26684
rect 8112 26624 8176 26628
rect 8192 26684 8256 26688
rect 8192 26628 8196 26684
rect 8196 26628 8252 26684
rect 8252 26628 8256 26684
rect 8192 26624 8256 26628
rect 428 26420 492 26484
rect 8340 26284 8404 26348
rect 9996 26208 10060 26212
rect 9996 26152 10010 26208
rect 10010 26152 10060 26208
rect 3012 26140 3076 26144
rect 3012 26084 3016 26140
rect 3016 26084 3072 26140
rect 3072 26084 3076 26140
rect 3012 26080 3076 26084
rect 3092 26140 3156 26144
rect 3092 26084 3096 26140
rect 3096 26084 3152 26140
rect 3152 26084 3156 26140
rect 3092 26080 3156 26084
rect 3172 26140 3236 26144
rect 3172 26084 3176 26140
rect 3176 26084 3232 26140
rect 3232 26084 3236 26140
rect 3172 26080 3236 26084
rect 3252 26140 3316 26144
rect 3252 26084 3256 26140
rect 3256 26084 3312 26140
rect 3312 26084 3316 26140
rect 3252 26080 3316 26084
rect 3740 26012 3804 26076
rect 2636 25936 2700 25940
rect 2636 25880 2686 25936
rect 2686 25880 2700 25936
rect 2636 25876 2700 25880
rect 7052 25740 7116 25804
rect 9996 26148 10060 26152
rect 9012 26140 9076 26144
rect 9012 26084 9016 26140
rect 9016 26084 9072 26140
rect 9072 26084 9076 26140
rect 9012 26080 9076 26084
rect 9092 26140 9156 26144
rect 9092 26084 9096 26140
rect 9096 26084 9152 26140
rect 9152 26084 9156 26140
rect 9092 26080 9156 26084
rect 9172 26140 9236 26144
rect 9172 26084 9176 26140
rect 9176 26084 9232 26140
rect 9232 26084 9236 26140
rect 9172 26080 9236 26084
rect 9252 26140 9316 26144
rect 9252 26084 9256 26140
rect 9256 26084 9312 26140
rect 9312 26084 9316 26140
rect 9252 26080 9316 26084
rect 9628 26012 9692 26076
rect 10732 25740 10796 25804
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 7952 25596 8016 25600
rect 7952 25540 7956 25596
rect 7956 25540 8012 25596
rect 8012 25540 8016 25596
rect 7952 25536 8016 25540
rect 8032 25596 8096 25600
rect 8032 25540 8036 25596
rect 8036 25540 8092 25596
rect 8092 25540 8096 25596
rect 8032 25536 8096 25540
rect 8112 25596 8176 25600
rect 8112 25540 8116 25596
rect 8116 25540 8172 25596
rect 8172 25540 8176 25596
rect 8112 25536 8176 25540
rect 8192 25596 8256 25600
rect 8192 25540 8196 25596
rect 8196 25540 8252 25596
rect 8252 25540 8256 25596
rect 8192 25536 8256 25540
rect 4108 25468 4172 25532
rect 2636 25332 2700 25396
rect 6500 25332 6564 25396
rect 7420 25060 7484 25124
rect 3012 25052 3076 25056
rect 3012 24996 3016 25052
rect 3016 24996 3072 25052
rect 3072 24996 3076 25052
rect 3012 24992 3076 24996
rect 3092 25052 3156 25056
rect 3092 24996 3096 25052
rect 3096 24996 3152 25052
rect 3152 24996 3156 25052
rect 3092 24992 3156 24996
rect 3172 25052 3236 25056
rect 3172 24996 3176 25052
rect 3176 24996 3232 25052
rect 3232 24996 3236 25052
rect 3172 24992 3236 24996
rect 3252 25052 3316 25056
rect 3252 24996 3256 25052
rect 3256 24996 3312 25052
rect 3312 24996 3316 25052
rect 3252 24992 3316 24996
rect 9012 25052 9076 25056
rect 9012 24996 9016 25052
rect 9016 24996 9072 25052
rect 9072 24996 9076 25052
rect 9012 24992 9076 24996
rect 9092 25052 9156 25056
rect 9092 24996 9096 25052
rect 9096 24996 9152 25052
rect 9152 24996 9156 25052
rect 9092 24992 9156 24996
rect 9172 25052 9236 25056
rect 9172 24996 9176 25052
rect 9176 24996 9232 25052
rect 9232 24996 9236 25052
rect 9172 24992 9236 24996
rect 9252 25052 9316 25056
rect 9252 24996 9256 25052
rect 9256 24996 9312 25052
rect 9312 24996 9316 25052
rect 9252 24992 9316 24996
rect 244 24924 308 24988
rect 5028 24924 5092 24988
rect 7788 24924 7852 24988
rect 5028 24788 5092 24852
rect 6868 24788 6932 24852
rect 1532 24652 1596 24716
rect 6868 24652 6932 24716
rect 7420 24788 7484 24852
rect 7788 24652 7852 24716
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 7952 24508 8016 24512
rect 7952 24452 7956 24508
rect 7956 24452 8012 24508
rect 8012 24452 8016 24508
rect 7952 24448 8016 24452
rect 8032 24508 8096 24512
rect 8032 24452 8036 24508
rect 8036 24452 8092 24508
rect 8092 24452 8096 24508
rect 8032 24448 8096 24452
rect 8112 24508 8176 24512
rect 8112 24452 8116 24508
rect 8116 24452 8172 24508
rect 8172 24452 8176 24508
rect 8112 24448 8176 24452
rect 8192 24508 8256 24512
rect 8192 24452 8196 24508
rect 8196 24452 8252 24508
rect 8252 24452 8256 24508
rect 8192 24448 8256 24452
rect 2452 24380 2516 24444
rect 3012 23964 3076 23968
rect 3012 23908 3016 23964
rect 3016 23908 3072 23964
rect 3072 23908 3076 23964
rect 3012 23904 3076 23908
rect 3092 23964 3156 23968
rect 3092 23908 3096 23964
rect 3096 23908 3152 23964
rect 3152 23908 3156 23964
rect 3092 23904 3156 23908
rect 3172 23964 3236 23968
rect 3172 23908 3176 23964
rect 3176 23908 3232 23964
rect 3232 23908 3236 23964
rect 3172 23904 3236 23908
rect 3252 23964 3316 23968
rect 3252 23908 3256 23964
rect 3256 23908 3312 23964
rect 3312 23908 3316 23964
rect 3252 23904 3316 23908
rect 9012 23964 9076 23968
rect 9012 23908 9016 23964
rect 9016 23908 9072 23964
rect 9072 23908 9076 23964
rect 9012 23904 9076 23908
rect 9092 23964 9156 23968
rect 9092 23908 9096 23964
rect 9096 23908 9152 23964
rect 9152 23908 9156 23964
rect 9092 23904 9156 23908
rect 9172 23964 9236 23968
rect 9172 23908 9176 23964
rect 9176 23908 9232 23964
rect 9232 23908 9236 23964
rect 9172 23904 9236 23908
rect 9252 23964 9316 23968
rect 9252 23908 9256 23964
rect 9256 23908 9312 23964
rect 9312 23908 9316 23964
rect 9252 23904 9316 23908
rect 5396 23836 5460 23900
rect 8524 23836 8588 23900
rect 8524 23700 8588 23764
rect 4844 23428 4908 23492
rect 7236 23428 7300 23492
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 4292 23292 4356 23356
rect 428 23156 492 23220
rect 2452 23156 2516 23220
rect 5396 23020 5460 23084
rect 3012 22876 3076 22880
rect 3012 22820 3016 22876
rect 3016 22820 3072 22876
rect 3072 22820 3076 22876
rect 3012 22816 3076 22820
rect 3092 22876 3156 22880
rect 3092 22820 3096 22876
rect 3096 22820 3152 22876
rect 3152 22820 3156 22876
rect 3092 22816 3156 22820
rect 3172 22876 3236 22880
rect 3172 22820 3176 22876
rect 3176 22820 3232 22876
rect 3232 22820 3236 22876
rect 3172 22816 3236 22820
rect 3252 22876 3316 22880
rect 3252 22820 3256 22876
rect 3256 22820 3312 22876
rect 3312 22820 3316 22876
rect 3252 22816 3316 22820
rect 6500 22748 6564 22812
rect 5580 22612 5644 22676
rect 7052 22612 7116 22676
rect 2820 22476 2884 22540
rect 3740 22340 3804 22404
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 3740 22204 3804 22268
rect 4292 22204 4356 22268
rect 6684 22204 6748 22268
rect 7236 22264 7300 22268
rect 7236 22208 7250 22264
rect 7250 22208 7300 22264
rect 7236 22204 7300 22208
rect 7952 23420 8016 23424
rect 7952 23364 7956 23420
rect 7956 23364 8012 23420
rect 8012 23364 8016 23420
rect 7952 23360 8016 23364
rect 8032 23420 8096 23424
rect 8032 23364 8036 23420
rect 8036 23364 8092 23420
rect 8092 23364 8096 23420
rect 8032 23360 8096 23364
rect 8112 23420 8176 23424
rect 8112 23364 8116 23420
rect 8116 23364 8172 23420
rect 8172 23364 8176 23420
rect 8112 23360 8176 23364
rect 8192 23420 8256 23424
rect 8192 23364 8196 23420
rect 8196 23364 8252 23420
rect 8252 23364 8256 23420
rect 8192 23360 8256 23364
rect 9012 22876 9076 22880
rect 9012 22820 9016 22876
rect 9016 22820 9072 22876
rect 9072 22820 9076 22876
rect 9012 22816 9076 22820
rect 9092 22876 9156 22880
rect 9092 22820 9096 22876
rect 9096 22820 9152 22876
rect 9152 22820 9156 22876
rect 9092 22816 9156 22820
rect 9172 22876 9236 22880
rect 9172 22820 9176 22876
rect 9176 22820 9232 22876
rect 9232 22820 9236 22876
rect 9172 22816 9236 22820
rect 9252 22876 9316 22880
rect 9252 22820 9256 22876
rect 9256 22820 9312 22876
rect 9312 22820 9316 22876
rect 9252 22816 9316 22820
rect 9996 22476 10060 22540
rect 7952 22332 8016 22336
rect 7952 22276 7956 22332
rect 7956 22276 8012 22332
rect 8012 22276 8016 22332
rect 7952 22272 8016 22276
rect 8032 22332 8096 22336
rect 8032 22276 8036 22332
rect 8036 22276 8092 22332
rect 8092 22276 8096 22332
rect 8032 22272 8096 22276
rect 8112 22332 8176 22336
rect 8112 22276 8116 22332
rect 8116 22276 8172 22332
rect 8172 22276 8176 22332
rect 8112 22272 8176 22276
rect 8192 22332 8256 22336
rect 8192 22276 8196 22332
rect 8196 22276 8252 22332
rect 8252 22276 8256 22332
rect 8192 22272 8256 22276
rect 1532 22068 1596 22132
rect 4844 21856 4908 21860
rect 4844 21800 4858 21856
rect 4858 21800 4908 21856
rect 3012 21788 3076 21792
rect 3012 21732 3016 21788
rect 3016 21732 3072 21788
rect 3072 21732 3076 21788
rect 3012 21728 3076 21732
rect 3092 21788 3156 21792
rect 3092 21732 3096 21788
rect 3096 21732 3152 21788
rect 3152 21732 3156 21788
rect 3092 21728 3156 21732
rect 3172 21788 3236 21792
rect 3172 21732 3176 21788
rect 3176 21732 3232 21788
rect 3232 21732 3236 21788
rect 3172 21728 3236 21732
rect 3252 21788 3316 21792
rect 3252 21732 3256 21788
rect 3256 21732 3312 21788
rect 3312 21732 3316 21788
rect 3252 21728 3316 21732
rect 1532 21524 1596 21588
rect 2452 21524 2516 21588
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 4844 21796 4908 21800
rect 7052 21856 7116 21860
rect 7052 21800 7102 21856
rect 7102 21800 7116 21856
rect 7052 21796 7116 21800
rect 8708 21932 8772 21996
rect 9012 21788 9076 21792
rect 9012 21732 9016 21788
rect 9016 21732 9072 21788
rect 9072 21732 9076 21788
rect 9012 21728 9076 21732
rect 9092 21788 9156 21792
rect 9092 21732 9096 21788
rect 9096 21732 9152 21788
rect 9152 21732 9156 21788
rect 9092 21728 9156 21732
rect 9172 21788 9236 21792
rect 9172 21732 9176 21788
rect 9176 21732 9232 21788
rect 9232 21732 9236 21788
rect 9172 21728 9236 21732
rect 9252 21788 9316 21792
rect 9252 21732 9256 21788
rect 9256 21732 9312 21788
rect 9312 21732 9316 21788
rect 9252 21728 9316 21732
rect 3740 21720 3804 21724
rect 3740 21664 3790 21720
rect 3790 21664 3804 21720
rect 3740 21660 3804 21664
rect 5580 21660 5644 21724
rect 8708 21660 8772 21724
rect 10916 21660 10980 21724
rect 3740 21524 3804 21588
rect 6500 21524 6564 21588
rect 5396 21388 5460 21452
rect 6868 21252 6932 21316
rect 5212 21116 5276 21180
rect 2636 20844 2700 20908
rect 4108 20708 4172 20772
rect 3012 20700 3076 20704
rect 3012 20644 3016 20700
rect 3016 20644 3072 20700
rect 3072 20644 3076 20700
rect 3012 20640 3076 20644
rect 3092 20700 3156 20704
rect 3092 20644 3096 20700
rect 3096 20644 3152 20700
rect 3152 20644 3156 20700
rect 3092 20640 3156 20644
rect 3172 20700 3236 20704
rect 3172 20644 3176 20700
rect 3176 20644 3232 20700
rect 3232 20644 3236 20700
rect 3172 20640 3236 20644
rect 3252 20700 3316 20704
rect 3252 20644 3256 20700
rect 3256 20644 3312 20700
rect 3312 20644 3316 20700
rect 3252 20640 3316 20644
rect 1348 20632 1412 20636
rect 1348 20576 1398 20632
rect 1398 20576 1412 20632
rect 1348 20572 1412 20576
rect 4108 20572 4172 20636
rect 7236 20572 7300 20636
rect 7952 21244 8016 21248
rect 7952 21188 7956 21244
rect 7956 21188 8012 21244
rect 8012 21188 8016 21244
rect 7952 21184 8016 21188
rect 8032 21244 8096 21248
rect 8032 21188 8036 21244
rect 8036 21188 8092 21244
rect 8092 21188 8096 21244
rect 8032 21184 8096 21188
rect 8112 21244 8176 21248
rect 8112 21188 8116 21244
rect 8116 21188 8172 21244
rect 8172 21188 8176 21244
rect 8112 21184 8176 21188
rect 8192 21244 8256 21248
rect 8192 21188 8196 21244
rect 8196 21188 8252 21244
rect 8252 21188 8256 21244
rect 8192 21184 8256 21188
rect 9012 20700 9076 20704
rect 9012 20644 9016 20700
rect 9016 20644 9072 20700
rect 9072 20644 9076 20700
rect 9012 20640 9076 20644
rect 9092 20700 9156 20704
rect 9092 20644 9096 20700
rect 9096 20644 9152 20700
rect 9152 20644 9156 20700
rect 9092 20640 9156 20644
rect 9172 20700 9236 20704
rect 9172 20644 9176 20700
rect 9176 20644 9232 20700
rect 9232 20644 9236 20700
rect 9172 20640 9236 20644
rect 9252 20700 9316 20704
rect 9252 20644 9256 20700
rect 9256 20644 9312 20700
rect 9312 20644 9316 20700
rect 9252 20640 9316 20644
rect 9628 20436 9692 20500
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 8708 20300 8772 20364
rect 7952 20156 8016 20160
rect 7952 20100 7956 20156
rect 7956 20100 8012 20156
rect 8012 20100 8016 20156
rect 7952 20096 8016 20100
rect 8032 20156 8096 20160
rect 8032 20100 8036 20156
rect 8036 20100 8092 20156
rect 8092 20100 8096 20156
rect 8032 20096 8096 20100
rect 8112 20156 8176 20160
rect 8112 20100 8116 20156
rect 8116 20100 8172 20156
rect 8172 20100 8176 20156
rect 8112 20096 8176 20100
rect 8192 20156 8256 20160
rect 8192 20100 8196 20156
rect 8196 20100 8252 20156
rect 8252 20100 8256 20156
rect 8192 20096 8256 20100
rect 6684 19620 6748 19684
rect 3012 19612 3076 19616
rect 3012 19556 3016 19612
rect 3016 19556 3072 19612
rect 3072 19556 3076 19612
rect 3012 19552 3076 19556
rect 3092 19612 3156 19616
rect 3092 19556 3096 19612
rect 3096 19556 3152 19612
rect 3152 19556 3156 19612
rect 3092 19552 3156 19556
rect 3172 19612 3236 19616
rect 3172 19556 3176 19612
rect 3176 19556 3232 19612
rect 3232 19556 3236 19612
rect 3172 19552 3236 19556
rect 3252 19612 3316 19616
rect 3252 19556 3256 19612
rect 3256 19556 3312 19612
rect 3312 19556 3316 19612
rect 3252 19552 3316 19556
rect 7788 19348 7852 19412
rect 9012 19612 9076 19616
rect 9012 19556 9016 19612
rect 9016 19556 9072 19612
rect 9072 19556 9076 19612
rect 9012 19552 9076 19556
rect 9092 19612 9156 19616
rect 9092 19556 9096 19612
rect 9096 19556 9152 19612
rect 9152 19556 9156 19612
rect 9092 19552 9156 19556
rect 9172 19612 9236 19616
rect 9172 19556 9176 19612
rect 9176 19556 9232 19612
rect 9232 19556 9236 19612
rect 9172 19552 9236 19556
rect 9252 19612 9316 19616
rect 9252 19556 9256 19612
rect 9256 19556 9312 19612
rect 9312 19556 9316 19612
rect 9252 19552 9316 19556
rect 10732 19484 10796 19548
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 5948 19000 6012 19004
rect 5948 18944 5962 19000
rect 5962 18944 6012 19000
rect 5948 18940 6012 18944
rect 6684 18804 6748 18868
rect 7952 19068 8016 19072
rect 7952 19012 7956 19068
rect 7956 19012 8012 19068
rect 8012 19012 8016 19068
rect 7952 19008 8016 19012
rect 8032 19068 8096 19072
rect 8032 19012 8036 19068
rect 8036 19012 8092 19068
rect 8092 19012 8096 19068
rect 8032 19008 8096 19012
rect 8112 19068 8176 19072
rect 8112 19012 8116 19068
rect 8116 19012 8172 19068
rect 8172 19012 8176 19068
rect 8112 19008 8176 19012
rect 8192 19068 8256 19072
rect 8192 19012 8196 19068
rect 8196 19012 8252 19068
rect 8252 19012 8256 19068
rect 8192 19008 8256 19012
rect 8708 18804 8772 18868
rect 5948 18668 6012 18732
rect 10916 18668 10980 18732
rect 4108 18532 4172 18596
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 3172 18524 3236 18528
rect 3172 18468 3176 18524
rect 3176 18468 3232 18524
rect 3232 18468 3236 18524
rect 3172 18464 3236 18468
rect 3252 18524 3316 18528
rect 3252 18468 3256 18524
rect 3256 18468 3312 18524
rect 3312 18468 3316 18524
rect 3252 18464 3316 18468
rect 9012 18524 9076 18528
rect 9012 18468 9016 18524
rect 9016 18468 9072 18524
rect 9072 18468 9076 18524
rect 9012 18464 9076 18468
rect 9092 18524 9156 18528
rect 9092 18468 9096 18524
rect 9096 18468 9152 18524
rect 9152 18468 9156 18524
rect 9092 18464 9156 18468
rect 9172 18524 9236 18528
rect 9172 18468 9176 18524
rect 9176 18468 9232 18524
rect 9232 18468 9236 18524
rect 9172 18464 9236 18468
rect 9252 18524 9316 18528
rect 9252 18468 9256 18524
rect 9256 18468 9312 18524
rect 9312 18468 9316 18524
rect 9252 18464 9316 18468
rect 4292 18260 4356 18324
rect 5580 18124 5644 18188
rect 6868 18124 6932 18188
rect 7788 18124 7852 18188
rect 2820 17988 2884 18052
rect 4660 17988 4724 18052
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 2452 17852 2516 17916
rect 2820 17852 2884 17916
rect 4660 17852 4724 17916
rect 7952 17980 8016 17984
rect 7952 17924 7956 17980
rect 7956 17924 8012 17980
rect 8012 17924 8016 17980
rect 7952 17920 8016 17924
rect 8032 17980 8096 17984
rect 8032 17924 8036 17980
rect 8036 17924 8092 17980
rect 8092 17924 8096 17980
rect 8032 17920 8096 17924
rect 8112 17980 8176 17984
rect 8112 17924 8116 17980
rect 8116 17924 8172 17980
rect 8172 17924 8176 17980
rect 8112 17920 8176 17924
rect 8192 17980 8256 17984
rect 8192 17924 8196 17980
rect 8196 17924 8252 17980
rect 8252 17924 8256 17980
rect 8192 17920 8256 17924
rect 6316 17912 6380 17916
rect 6316 17856 6330 17912
rect 6330 17856 6380 17912
rect 6316 17852 6380 17856
rect 9628 17852 9692 17916
rect 9996 17852 10060 17916
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 3172 17436 3236 17440
rect 3172 17380 3176 17436
rect 3176 17380 3232 17436
rect 3232 17380 3236 17436
rect 3172 17376 3236 17380
rect 3252 17436 3316 17440
rect 3252 17380 3256 17436
rect 3256 17380 3312 17436
rect 3312 17380 3316 17436
rect 3252 17376 3316 17380
rect 9012 17436 9076 17440
rect 9012 17380 9016 17436
rect 9016 17380 9072 17436
rect 9072 17380 9076 17436
rect 9012 17376 9076 17380
rect 9092 17436 9156 17440
rect 9092 17380 9096 17436
rect 9096 17380 9152 17436
rect 9152 17380 9156 17436
rect 9092 17376 9156 17380
rect 9172 17436 9236 17440
rect 9172 17380 9176 17436
rect 9176 17380 9232 17436
rect 9232 17380 9236 17436
rect 9172 17376 9236 17380
rect 9252 17436 9316 17440
rect 9252 17380 9256 17436
rect 9256 17380 9312 17436
rect 9312 17380 9316 17436
rect 9252 17376 9316 17380
rect 2452 17036 2516 17100
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 3740 17036 3804 17100
rect 5028 17096 5092 17100
rect 5028 17040 5078 17096
rect 5078 17040 5092 17096
rect 5028 17036 5092 17040
rect 7788 17036 7852 17100
rect 3740 16900 3804 16964
rect 4476 16900 4540 16964
rect 7952 16892 8016 16896
rect 7952 16836 7956 16892
rect 7956 16836 8012 16892
rect 8012 16836 8016 16892
rect 7952 16832 8016 16836
rect 8032 16892 8096 16896
rect 8032 16836 8036 16892
rect 8036 16836 8092 16892
rect 8092 16836 8096 16892
rect 8032 16832 8096 16836
rect 8112 16892 8176 16896
rect 8112 16836 8116 16892
rect 8116 16836 8172 16892
rect 8172 16836 8176 16892
rect 8112 16832 8176 16836
rect 8192 16892 8256 16896
rect 8192 16836 8196 16892
rect 8196 16836 8252 16892
rect 8252 16836 8256 16892
rect 8192 16832 8256 16836
rect 4292 16628 4356 16692
rect 6500 16492 6564 16556
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 3172 16348 3236 16352
rect 3172 16292 3176 16348
rect 3176 16292 3232 16348
rect 3232 16292 3236 16348
rect 3172 16288 3236 16292
rect 3252 16348 3316 16352
rect 3252 16292 3256 16348
rect 3256 16292 3312 16348
rect 3312 16292 3316 16348
rect 3252 16288 3316 16292
rect 9012 16348 9076 16352
rect 9012 16292 9016 16348
rect 9016 16292 9072 16348
rect 9072 16292 9076 16348
rect 9012 16288 9076 16292
rect 9092 16348 9156 16352
rect 9092 16292 9096 16348
rect 9096 16292 9152 16348
rect 9152 16292 9156 16348
rect 9092 16288 9156 16292
rect 9172 16348 9236 16352
rect 9172 16292 9176 16348
rect 9176 16292 9232 16348
rect 9232 16292 9236 16348
rect 9172 16288 9236 16292
rect 9252 16348 9316 16352
rect 9252 16292 9256 16348
rect 9256 16292 9312 16348
rect 9312 16292 9316 16348
rect 9252 16288 9316 16292
rect 5764 16084 5828 16148
rect 7604 16144 7668 16148
rect 7604 16088 7618 16144
rect 7618 16088 7668 16144
rect 7604 16084 7668 16088
rect 5764 15948 5828 16012
rect 10364 15948 10428 16012
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 7952 15804 8016 15808
rect 7952 15748 7956 15804
rect 7956 15748 8012 15804
rect 8012 15748 8016 15804
rect 7952 15744 8016 15748
rect 8032 15804 8096 15808
rect 8032 15748 8036 15804
rect 8036 15748 8092 15804
rect 8092 15748 8096 15804
rect 8032 15744 8096 15748
rect 8112 15804 8176 15808
rect 8112 15748 8116 15804
rect 8116 15748 8172 15804
rect 8172 15748 8176 15804
rect 8112 15744 8176 15748
rect 8192 15804 8256 15808
rect 8192 15748 8196 15804
rect 8196 15748 8252 15804
rect 8252 15748 8256 15804
rect 8192 15744 8256 15748
rect 7236 15676 7300 15740
rect 9444 15540 9508 15604
rect 7604 15404 7668 15468
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 3172 15260 3236 15264
rect 3172 15204 3176 15260
rect 3176 15204 3232 15260
rect 3232 15204 3236 15260
rect 3172 15200 3236 15204
rect 3252 15260 3316 15264
rect 3252 15204 3256 15260
rect 3256 15204 3312 15260
rect 3312 15204 3316 15260
rect 3252 15200 3316 15204
rect 9012 15260 9076 15264
rect 9012 15204 9016 15260
rect 9016 15204 9072 15260
rect 9072 15204 9076 15260
rect 9012 15200 9076 15204
rect 9092 15260 9156 15264
rect 9092 15204 9096 15260
rect 9096 15204 9152 15260
rect 9152 15204 9156 15260
rect 9092 15200 9156 15204
rect 9172 15260 9236 15264
rect 9172 15204 9176 15260
rect 9176 15204 9232 15260
rect 9232 15204 9236 15260
rect 9172 15200 9236 15204
rect 9252 15260 9316 15264
rect 9252 15204 9256 15260
rect 9256 15204 9312 15260
rect 9312 15204 9316 15260
rect 9252 15200 9316 15204
rect 2636 14996 2700 15060
rect 4292 14860 4356 14924
rect 5028 14860 5092 14924
rect 5396 14860 5460 14924
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 7952 14716 8016 14720
rect 7952 14660 7956 14716
rect 7956 14660 8012 14716
rect 8012 14660 8016 14716
rect 7952 14656 8016 14660
rect 8032 14716 8096 14720
rect 8032 14660 8036 14716
rect 8036 14660 8092 14716
rect 8092 14660 8096 14716
rect 8032 14656 8096 14660
rect 8112 14716 8176 14720
rect 8112 14660 8116 14716
rect 8116 14660 8172 14716
rect 8172 14660 8176 14716
rect 8112 14656 8176 14660
rect 8192 14716 8256 14720
rect 8192 14660 8196 14716
rect 8196 14660 8252 14716
rect 8252 14660 8256 14716
rect 8192 14656 8256 14660
rect 6684 14588 6748 14652
rect 6684 14512 6748 14516
rect 6684 14456 6734 14512
rect 6734 14456 6748 14512
rect 6684 14452 6748 14456
rect 8340 14588 8404 14652
rect 1532 14316 1596 14380
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 3172 14172 3236 14176
rect 3172 14116 3176 14172
rect 3176 14116 3232 14172
rect 3232 14116 3236 14172
rect 3172 14112 3236 14116
rect 3252 14172 3316 14176
rect 3252 14116 3256 14172
rect 3256 14116 3312 14172
rect 3312 14116 3316 14172
rect 3252 14112 3316 14116
rect 9012 14172 9076 14176
rect 9012 14116 9016 14172
rect 9016 14116 9072 14172
rect 9072 14116 9076 14172
rect 9012 14112 9076 14116
rect 9092 14172 9156 14176
rect 9092 14116 9096 14172
rect 9096 14116 9152 14172
rect 9152 14116 9156 14172
rect 9092 14112 9156 14116
rect 9172 14172 9236 14176
rect 9172 14116 9176 14172
rect 9176 14116 9232 14172
rect 9232 14116 9236 14172
rect 9172 14112 9236 14116
rect 9252 14172 9316 14176
rect 9252 14116 9256 14172
rect 9256 14116 9312 14172
rect 9312 14116 9316 14172
rect 9252 14112 9316 14116
rect 5580 13636 5644 13700
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 5028 13500 5092 13564
rect 7604 13772 7668 13836
rect 8340 13772 8404 13836
rect 7952 13628 8016 13632
rect 7952 13572 7956 13628
rect 7956 13572 8012 13628
rect 8012 13572 8016 13628
rect 7952 13568 8016 13572
rect 8032 13628 8096 13632
rect 8032 13572 8036 13628
rect 8036 13572 8092 13628
rect 8092 13572 8096 13628
rect 8032 13568 8096 13572
rect 8112 13628 8176 13632
rect 8112 13572 8116 13628
rect 8116 13572 8172 13628
rect 8172 13572 8176 13628
rect 8112 13568 8176 13572
rect 8192 13628 8256 13632
rect 8192 13572 8196 13628
rect 8196 13572 8252 13628
rect 8252 13572 8256 13628
rect 8192 13568 8256 13572
rect 7420 13500 7484 13564
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 3172 13084 3236 13088
rect 3172 13028 3176 13084
rect 3176 13028 3232 13084
rect 3232 13028 3236 13084
rect 3172 13024 3236 13028
rect 3252 13084 3316 13088
rect 3252 13028 3256 13084
rect 3256 13028 3312 13084
rect 3312 13028 3316 13084
rect 3252 13024 3316 13028
rect 9012 13084 9076 13088
rect 9012 13028 9016 13084
rect 9016 13028 9072 13084
rect 9072 13028 9076 13084
rect 9012 13024 9076 13028
rect 9092 13084 9156 13088
rect 9092 13028 9096 13084
rect 9096 13028 9152 13084
rect 9152 13028 9156 13084
rect 9092 13024 9156 13028
rect 9172 13084 9236 13088
rect 9172 13028 9176 13084
rect 9176 13028 9232 13084
rect 9232 13028 9236 13084
rect 9172 13024 9236 13028
rect 9252 13084 9316 13088
rect 9252 13028 9256 13084
rect 9256 13028 9312 13084
rect 9312 13028 9316 13084
rect 9252 13024 9316 13028
rect 7788 12956 7852 13020
rect 4844 12684 4908 12748
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 7952 12540 8016 12544
rect 7952 12484 7956 12540
rect 7956 12484 8012 12540
rect 8012 12484 8016 12540
rect 7952 12480 8016 12484
rect 8032 12540 8096 12544
rect 8032 12484 8036 12540
rect 8036 12484 8092 12540
rect 8092 12484 8096 12540
rect 8032 12480 8096 12484
rect 8112 12540 8176 12544
rect 8112 12484 8116 12540
rect 8116 12484 8172 12540
rect 8172 12484 8176 12540
rect 8112 12480 8176 12484
rect 8192 12540 8256 12544
rect 8192 12484 8196 12540
rect 8196 12484 8252 12540
rect 8252 12484 8256 12540
rect 8192 12480 8256 12484
rect 8524 12276 8588 12340
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 3172 11996 3236 12000
rect 3172 11940 3176 11996
rect 3176 11940 3232 11996
rect 3232 11940 3236 11996
rect 3172 11936 3236 11940
rect 3252 11996 3316 12000
rect 3252 11940 3256 11996
rect 3256 11940 3312 11996
rect 3312 11940 3316 11996
rect 3252 11936 3316 11940
rect 9012 11996 9076 12000
rect 9012 11940 9016 11996
rect 9016 11940 9072 11996
rect 9072 11940 9076 11996
rect 9012 11936 9076 11940
rect 9092 11996 9156 12000
rect 9092 11940 9096 11996
rect 9096 11940 9152 11996
rect 9152 11940 9156 11996
rect 9092 11936 9156 11940
rect 9172 11996 9236 12000
rect 9172 11940 9176 11996
rect 9176 11940 9232 11996
rect 9232 11940 9236 11996
rect 9172 11936 9236 11940
rect 9252 11996 9316 12000
rect 9252 11940 9256 11996
rect 9256 11940 9312 11996
rect 9312 11940 9316 11996
rect 9252 11936 9316 11940
rect 4108 11868 4172 11932
rect 5948 11868 6012 11932
rect 9628 11732 9692 11796
rect 6132 11596 6196 11660
rect 8340 11460 8404 11524
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 7952 11452 8016 11456
rect 7952 11396 7956 11452
rect 7956 11396 8012 11452
rect 8012 11396 8016 11452
rect 7952 11392 8016 11396
rect 8032 11452 8096 11456
rect 8032 11396 8036 11452
rect 8036 11396 8092 11452
rect 8092 11396 8096 11452
rect 8032 11392 8096 11396
rect 8112 11452 8176 11456
rect 8112 11396 8116 11452
rect 8116 11396 8172 11452
rect 8172 11396 8176 11452
rect 8112 11392 8176 11396
rect 8192 11452 8256 11456
rect 8192 11396 8196 11452
rect 8196 11396 8252 11452
rect 8252 11396 8256 11452
rect 8192 11392 8256 11396
rect 3740 11324 3804 11388
rect 3556 11052 3620 11116
rect 796 10916 860 10980
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 3172 10908 3236 10912
rect 3172 10852 3176 10908
rect 3176 10852 3232 10908
rect 3232 10852 3236 10908
rect 3172 10848 3236 10852
rect 3252 10908 3316 10912
rect 3252 10852 3256 10908
rect 3256 10852 3312 10908
rect 3312 10852 3316 10908
rect 3252 10848 3316 10852
rect 9012 10908 9076 10912
rect 9012 10852 9016 10908
rect 9016 10852 9072 10908
rect 9072 10852 9076 10908
rect 9012 10848 9076 10852
rect 9092 10908 9156 10912
rect 9092 10852 9096 10908
rect 9096 10852 9152 10908
rect 9152 10852 9156 10908
rect 9092 10848 9156 10852
rect 9172 10908 9236 10912
rect 9172 10852 9176 10908
rect 9176 10852 9232 10908
rect 9232 10852 9236 10908
rect 9172 10848 9236 10852
rect 9252 10908 9316 10912
rect 9252 10852 9256 10908
rect 9256 10852 9312 10908
rect 9312 10852 9316 10908
rect 9252 10848 9316 10852
rect 7052 10508 7116 10572
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 7952 10364 8016 10368
rect 7952 10308 7956 10364
rect 7956 10308 8012 10364
rect 8012 10308 8016 10364
rect 7952 10304 8016 10308
rect 8032 10364 8096 10368
rect 8032 10308 8036 10364
rect 8036 10308 8092 10364
rect 8092 10308 8096 10364
rect 8032 10304 8096 10308
rect 8112 10364 8176 10368
rect 8112 10308 8116 10364
rect 8116 10308 8172 10364
rect 8172 10308 8176 10364
rect 8112 10304 8176 10308
rect 8192 10364 8256 10368
rect 8192 10308 8196 10364
rect 8196 10308 8252 10364
rect 8252 10308 8256 10364
rect 8192 10304 8256 10308
rect 1716 10100 1780 10164
rect 6684 10100 6748 10164
rect 8340 10100 8404 10164
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 3172 9820 3236 9824
rect 3172 9764 3176 9820
rect 3176 9764 3232 9820
rect 3232 9764 3236 9820
rect 3172 9760 3236 9764
rect 3252 9820 3316 9824
rect 3252 9764 3256 9820
rect 3256 9764 3312 9820
rect 3312 9764 3316 9820
rect 3252 9760 3316 9764
rect 9012 9820 9076 9824
rect 9012 9764 9016 9820
rect 9016 9764 9072 9820
rect 9072 9764 9076 9820
rect 9012 9760 9076 9764
rect 9092 9820 9156 9824
rect 9092 9764 9096 9820
rect 9096 9764 9152 9820
rect 9152 9764 9156 9820
rect 9092 9760 9156 9764
rect 9172 9820 9236 9824
rect 9172 9764 9176 9820
rect 9176 9764 9232 9820
rect 9232 9764 9236 9820
rect 9172 9760 9236 9764
rect 9252 9820 9316 9824
rect 9252 9764 9256 9820
rect 9256 9764 9312 9820
rect 9312 9764 9316 9820
rect 9252 9760 9316 9764
rect 2820 9692 2884 9756
rect 4660 9692 4724 9756
rect 9444 9480 9508 9484
rect 9444 9424 9494 9480
rect 9494 9424 9508 9480
rect 9444 9420 9508 9424
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 7952 9276 8016 9280
rect 7952 9220 7956 9276
rect 7956 9220 8012 9276
rect 8012 9220 8016 9276
rect 7952 9216 8016 9220
rect 8032 9276 8096 9280
rect 8032 9220 8036 9276
rect 8036 9220 8092 9276
rect 8092 9220 8096 9276
rect 8032 9216 8096 9220
rect 8112 9276 8176 9280
rect 8112 9220 8116 9276
rect 8116 9220 8172 9276
rect 8172 9220 8176 9276
rect 8112 9216 8176 9220
rect 8192 9276 8256 9280
rect 8192 9220 8196 9276
rect 8196 9220 8252 9276
rect 8252 9220 8256 9276
rect 8192 9216 8256 9220
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 2452 8256 2516 8260
rect 2452 8200 2466 8256
rect 2466 8200 2516 8256
rect 2452 8196 2516 8200
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 1164 7924 1228 7988
rect 9444 7712 9508 7716
rect 9444 7656 9494 7712
rect 9494 7656 9508 7712
rect 9444 7652 9508 7656
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 5396 7516 5460 7580
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 8708 6836 8772 6900
rect 10916 6700 10980 6764
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 5764 5944 5828 5948
rect 5764 5888 5778 5944
rect 5778 5888 5828 5944
rect 5764 5884 5828 5888
rect 6500 5944 6564 5948
rect 6500 5888 6514 5944
rect 6514 5888 6564 5944
rect 6500 5884 6564 5888
rect 5580 5808 5644 5812
rect 5580 5752 5594 5808
rect 5594 5752 5644 5808
rect 5580 5748 5644 5752
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 9812 5068 9876 5132
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 3924 2620 3988 2684
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 980 1260 1044 1324
rect 5212 1260 5276 1324
rect 10180 1320 10244 1324
rect 10180 1264 10194 1320
rect 10194 1264 10244 1320
rect 10180 1260 10244 1264
rect 612 1124 676 1188
rect 4844 1124 4908 1188
rect 10548 1124 10612 1188
<< metal4 >>
rect 1944 41920 2264 45000
rect 1944 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2264 41920
rect 795 41580 861 41581
rect 795 41516 796 41580
rect 860 41516 861 41580
rect 795 41515 861 41516
rect 611 41036 677 41037
rect 611 40972 612 41036
rect 676 40972 677 41036
rect 611 40971 677 40972
rect 243 31652 309 31653
rect 243 31588 244 31652
rect 308 31588 309 31652
rect 243 31587 309 31588
rect 246 24989 306 31587
rect 427 26484 493 26485
rect 427 26420 428 26484
rect 492 26420 493 26484
rect 427 26419 493 26420
rect 243 24988 309 24989
rect 243 24924 244 24988
rect 308 24924 309 24988
rect 243 24923 309 24924
rect 430 23221 490 26419
rect 427 23220 493 23221
rect 427 23156 428 23220
rect 492 23156 493 23220
rect 427 23155 493 23156
rect 614 1189 674 40971
rect 798 10981 858 41515
rect 1944 40832 2264 41856
rect 1944 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2264 40832
rect 1944 39744 2264 40768
rect 1944 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2264 39744
rect 979 39540 1045 39541
rect 979 39476 980 39540
rect 1044 39476 1045 39540
rect 979 39475 1045 39476
rect 795 10980 861 10981
rect 795 10916 796 10980
rect 860 10916 861 10980
rect 795 10915 861 10916
rect 982 1325 1042 39475
rect 1944 38656 2264 39680
rect 1944 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2264 38656
rect 1944 37568 2264 38592
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1531 35868 1597 35869
rect 1531 35804 1532 35868
rect 1596 35804 1597 35868
rect 1531 35803 1597 35804
rect 1163 28660 1229 28661
rect 1163 28596 1164 28660
rect 1228 28596 1229 28660
rect 1163 28595 1229 28596
rect 1166 7989 1226 28595
rect 1347 28524 1413 28525
rect 1347 28460 1348 28524
rect 1412 28460 1413 28524
rect 1347 28459 1413 28460
rect 1350 20637 1410 28459
rect 1534 24717 1594 35803
rect 1944 35392 2264 36416
rect 3004 42464 3324 45000
rect 3004 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3324 42464
rect 3004 41376 3324 42400
rect 3004 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3324 41376
rect 3004 40288 3324 41312
rect 7944 41920 8264 45000
rect 7944 41856 7952 41920
rect 8016 41856 8032 41920
rect 8096 41856 8112 41920
rect 8176 41856 8192 41920
rect 8256 41856 8264 41920
rect 7944 40832 8264 41856
rect 7944 40768 7952 40832
rect 8016 40768 8032 40832
rect 8096 40768 8112 40832
rect 8176 40768 8192 40832
rect 8256 40768 8264 40832
rect 7787 40356 7853 40357
rect 7787 40292 7788 40356
rect 7852 40292 7853 40356
rect 7787 40291 7853 40292
rect 3004 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3324 40288
rect 3004 39200 3324 40224
rect 5211 40084 5277 40085
rect 5211 40020 5212 40084
rect 5276 40020 5277 40084
rect 5211 40019 5277 40020
rect 3004 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3324 39200
rect 3004 38112 3324 39136
rect 3004 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3324 38112
rect 3004 37024 3324 38048
rect 4475 37772 4541 37773
rect 4475 37708 4476 37772
rect 4540 37708 4541 37772
rect 4475 37707 4541 37708
rect 3004 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3324 37024
rect 3004 35936 3324 36960
rect 3739 36140 3805 36141
rect 3739 36076 3740 36140
rect 3804 36076 3805 36140
rect 3739 36075 3805 36076
rect 3004 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3324 35936
rect 2635 35732 2701 35733
rect 2635 35668 2636 35732
rect 2700 35668 2701 35732
rect 2635 35667 2701 35668
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 2451 34508 2517 34509
rect 2451 34444 2452 34508
rect 2516 34444 2517 34508
rect 2451 34443 2517 34444
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33216 2264 34240
rect 1944 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2264 33216
rect 1715 32876 1781 32877
rect 1715 32812 1716 32876
rect 1780 32812 1781 32876
rect 1715 32811 1781 32812
rect 1718 29205 1778 32811
rect 1944 32128 2264 33152
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 2454 31770 2514 34443
rect 2638 31925 2698 35667
rect 3004 34848 3324 35872
rect 3004 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3324 34848
rect 3004 33760 3324 34784
rect 3555 34644 3621 34645
rect 3555 34580 3556 34644
rect 3620 34580 3621 34644
rect 3555 34579 3621 34580
rect 3004 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3324 33760
rect 2819 33148 2885 33149
rect 2819 33084 2820 33148
rect 2884 33084 2885 33148
rect 2819 33083 2885 33084
rect 2635 31924 2701 31925
rect 2635 31860 2636 31924
rect 2700 31860 2701 31924
rect 2635 31859 2701 31860
rect 2454 31710 2698 31770
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 2451 30292 2517 30293
rect 2451 30228 2452 30292
rect 2516 30228 2517 30292
rect 2451 30227 2517 30228
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1715 29204 1781 29205
rect 1715 29140 1716 29204
rect 1780 29140 1781 29204
rect 1715 29139 1781 29140
rect 1715 28932 1781 28933
rect 1715 28868 1716 28932
rect 1780 28868 1781 28932
rect 1715 28867 1781 28868
rect 1531 24716 1597 24717
rect 1531 24652 1532 24716
rect 1596 24652 1597 24716
rect 1531 24651 1597 24652
rect 1534 22133 1594 24651
rect 1531 22132 1597 22133
rect 1531 22068 1532 22132
rect 1596 22068 1597 22132
rect 1531 22067 1597 22068
rect 1531 21588 1597 21589
rect 1531 21524 1532 21588
rect 1596 21524 1597 21588
rect 1531 21523 1597 21524
rect 1347 20636 1413 20637
rect 1347 20572 1348 20636
rect 1412 20572 1413 20636
rect 1347 20571 1413 20572
rect 1534 14381 1594 21523
rect 1531 14380 1597 14381
rect 1531 14316 1532 14380
rect 1596 14316 1597 14380
rect 1531 14315 1597 14316
rect 1718 10165 1778 28867
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 27776 2264 28800
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 2454 24445 2514 30227
rect 2638 28117 2698 31710
rect 2822 30429 2882 33083
rect 3004 32672 3324 33696
rect 3004 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3324 32672
rect 3004 31584 3324 32608
rect 3004 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3324 31584
rect 3004 30496 3324 31520
rect 3004 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3324 30496
rect 2819 30428 2885 30429
rect 2819 30364 2820 30428
rect 2884 30364 2885 30428
rect 2819 30363 2885 30364
rect 3004 29408 3324 30432
rect 3004 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3324 29408
rect 3004 28320 3324 29344
rect 3004 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3324 28320
rect 2635 28116 2701 28117
rect 2635 28052 2636 28116
rect 2700 28052 2701 28116
rect 2635 28051 2701 28052
rect 2635 27980 2701 27981
rect 2635 27916 2636 27980
rect 2700 27916 2701 27980
rect 2635 27915 2701 27916
rect 2638 25941 2698 27915
rect 2819 27436 2885 27437
rect 2819 27372 2820 27436
rect 2884 27372 2885 27436
rect 2819 27371 2885 27372
rect 2635 25940 2701 25941
rect 2635 25876 2636 25940
rect 2700 25876 2701 25940
rect 2635 25875 2701 25876
rect 2635 25396 2701 25397
rect 2635 25332 2636 25396
rect 2700 25332 2701 25396
rect 2635 25331 2701 25332
rect 2451 24444 2517 24445
rect 2451 24380 2452 24444
rect 2516 24380 2517 24444
rect 2451 24379 2517 24380
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 22336 2264 23360
rect 2451 23220 2517 23221
rect 2451 23156 2452 23220
rect 2516 23156 2517 23220
rect 2451 23155 2517 23156
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 2454 21589 2514 23155
rect 2451 21588 2517 21589
rect 2451 21524 2452 21588
rect 2516 21524 2517 21588
rect 2451 21523 2517 21524
rect 2638 21450 2698 25331
rect 2822 22541 2882 27371
rect 3004 27232 3324 28256
rect 3004 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3324 27232
rect 3004 26144 3324 27168
rect 3558 27029 3618 34579
rect 3742 27573 3802 36075
rect 4291 33420 4357 33421
rect 4291 33356 4292 33420
rect 4356 33356 4357 33420
rect 4291 33355 4357 33356
rect 3923 33012 3989 33013
rect 3923 32948 3924 33012
rect 3988 32948 3989 33012
rect 3923 32947 3989 32948
rect 3926 30157 3986 32947
rect 4294 31517 4354 33355
rect 4291 31516 4357 31517
rect 4291 31452 4292 31516
rect 4356 31452 4357 31516
rect 4291 31451 4357 31452
rect 4107 30428 4173 30429
rect 4107 30364 4108 30428
rect 4172 30364 4173 30428
rect 4107 30363 4173 30364
rect 3923 30156 3989 30157
rect 3923 30092 3924 30156
rect 3988 30092 3989 30156
rect 3923 30091 3989 30092
rect 3923 27708 3989 27709
rect 3923 27644 3924 27708
rect 3988 27644 3989 27708
rect 3923 27643 3989 27644
rect 3739 27572 3805 27573
rect 3739 27508 3740 27572
rect 3804 27508 3805 27572
rect 3739 27507 3805 27508
rect 3555 27028 3621 27029
rect 3555 26964 3556 27028
rect 3620 26964 3621 27028
rect 3555 26963 3621 26964
rect 3555 26892 3621 26893
rect 3555 26828 3556 26892
rect 3620 26828 3621 26892
rect 3555 26827 3621 26828
rect 3004 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3324 26144
rect 3004 25056 3324 26080
rect 3004 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3324 25056
rect 3004 23968 3324 24992
rect 3004 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3324 23968
rect 3004 22880 3324 23904
rect 3004 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3324 22880
rect 2819 22540 2885 22541
rect 2819 22476 2820 22540
rect 2884 22476 2885 22540
rect 2819 22475 2885 22476
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 17984 2264 19008
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 2454 21390 2698 21450
rect 2454 17917 2514 21390
rect 2635 20908 2701 20909
rect 2635 20844 2636 20908
rect 2700 20844 2701 20908
rect 2635 20843 2701 20844
rect 2451 17916 2517 17917
rect 2451 17852 2452 17916
rect 2516 17852 2517 17916
rect 2451 17851 2517 17852
rect 2451 17100 2517 17101
rect 2451 17036 2452 17100
rect 2516 17036 2517 17100
rect 2451 17035 2517 17036
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 12544 2264 13568
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1715 10164 1781 10165
rect 1715 10100 1716 10164
rect 1780 10100 1781 10164
rect 1715 10099 1781 10100
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 2454 8261 2514 17035
rect 2638 15061 2698 20843
rect 2822 18053 2882 22475
rect 3004 21792 3324 22816
rect 3004 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3324 21792
rect 3004 20704 3324 21728
rect 3004 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3324 20704
rect 3004 19616 3324 20640
rect 3004 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3324 19616
rect 3004 18528 3324 19552
rect 3004 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3324 18528
rect 2819 18052 2885 18053
rect 2819 17988 2820 18052
rect 2884 17988 2885 18052
rect 2819 17987 2885 17988
rect 2819 17916 2885 17917
rect 2819 17852 2820 17916
rect 2884 17852 2885 17916
rect 2819 17851 2885 17852
rect 2635 15060 2701 15061
rect 2635 14996 2636 15060
rect 2700 14996 2701 15060
rect 2635 14995 2701 14996
rect 2822 9757 2882 17851
rect 3004 17440 3324 18464
rect 3004 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3324 17440
rect 3004 16352 3324 17376
rect 3004 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3324 16352
rect 3004 15264 3324 16288
rect 3004 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3324 15264
rect 3004 14176 3324 15200
rect 3004 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3324 14176
rect 3004 13088 3324 14112
rect 3004 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3324 13088
rect 3004 12000 3324 13024
rect 3004 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3324 12000
rect 3004 10912 3324 11936
rect 3558 11117 3618 26827
rect 3739 26076 3805 26077
rect 3739 26012 3740 26076
rect 3804 26012 3805 26076
rect 3739 26011 3805 26012
rect 3742 22405 3802 26011
rect 3739 22404 3805 22405
rect 3739 22340 3740 22404
rect 3804 22340 3805 22404
rect 3739 22339 3805 22340
rect 3739 22268 3805 22269
rect 3739 22204 3740 22268
rect 3804 22204 3805 22268
rect 3739 22203 3805 22204
rect 3742 21725 3802 22203
rect 3739 21724 3805 21725
rect 3739 21660 3740 21724
rect 3804 21660 3805 21724
rect 3739 21659 3805 21660
rect 3739 21588 3805 21589
rect 3739 21524 3740 21588
rect 3804 21524 3805 21588
rect 3739 21523 3805 21524
rect 3742 17101 3802 21523
rect 3739 17100 3805 17101
rect 3739 17036 3740 17100
rect 3804 17036 3805 17100
rect 3739 17035 3805 17036
rect 3739 16964 3805 16965
rect 3739 16900 3740 16964
rect 3804 16900 3805 16964
rect 3739 16899 3805 16900
rect 3742 16690 3802 16899
rect 3926 16690 3986 27643
rect 4110 26893 4170 30363
rect 4291 30292 4357 30293
rect 4291 30228 4292 30292
rect 4356 30228 4357 30292
rect 4291 30227 4357 30228
rect 4107 26892 4173 26893
rect 4107 26828 4108 26892
rect 4172 26828 4173 26892
rect 4107 26827 4173 26828
rect 4107 25532 4173 25533
rect 4107 25468 4108 25532
rect 4172 25468 4173 25532
rect 4107 25467 4173 25468
rect 4110 20773 4170 25467
rect 4294 23357 4354 30227
rect 4291 23356 4357 23357
rect 4291 23292 4292 23356
rect 4356 23292 4357 23356
rect 4291 23291 4357 23292
rect 4291 22268 4357 22269
rect 4291 22204 4292 22268
rect 4356 22204 4357 22268
rect 4291 22203 4357 22204
rect 4107 20772 4173 20773
rect 4107 20708 4108 20772
rect 4172 20708 4173 20772
rect 4107 20707 4173 20708
rect 4107 20636 4173 20637
rect 4107 20572 4108 20636
rect 4172 20572 4173 20636
rect 4107 20571 4173 20572
rect 4110 18597 4170 20571
rect 4107 18596 4173 18597
rect 4107 18532 4108 18596
rect 4172 18532 4173 18596
rect 4107 18531 4173 18532
rect 4294 18325 4354 22203
rect 4291 18324 4357 18325
rect 4291 18260 4292 18324
rect 4356 18260 4357 18324
rect 4291 18259 4357 18260
rect 4478 17370 4538 37707
rect 5027 37228 5093 37229
rect 5027 37164 5028 37228
rect 5092 37164 5093 37228
rect 5027 37163 5093 37164
rect 4659 36820 4725 36821
rect 4659 36756 4660 36820
rect 4724 36756 4725 36820
rect 4659 36755 4725 36756
rect 4662 30021 4722 36755
rect 4843 31380 4909 31381
rect 4843 31316 4844 31380
rect 4908 31316 4909 31380
rect 4843 31315 4909 31316
rect 4659 30020 4725 30021
rect 4659 29956 4660 30020
rect 4724 29956 4725 30020
rect 4659 29955 4725 29956
rect 4659 29612 4725 29613
rect 4659 29548 4660 29612
rect 4724 29548 4725 29612
rect 4659 29547 4725 29548
rect 4662 18053 4722 29547
rect 4846 23493 4906 31315
rect 5030 29477 5090 37163
rect 5027 29476 5093 29477
rect 5027 29412 5028 29476
rect 5092 29412 5093 29476
rect 5027 29411 5093 29412
rect 5027 27436 5093 27437
rect 5027 27372 5028 27436
rect 5092 27372 5093 27436
rect 5027 27371 5093 27372
rect 5030 24989 5090 27371
rect 5027 24988 5093 24989
rect 5027 24924 5028 24988
rect 5092 24924 5093 24988
rect 5027 24923 5093 24924
rect 5027 24852 5093 24853
rect 5027 24788 5028 24852
rect 5092 24788 5093 24852
rect 5027 24787 5093 24788
rect 4843 23492 4909 23493
rect 4843 23428 4844 23492
rect 4908 23428 4909 23492
rect 4843 23427 4909 23428
rect 4843 21860 4909 21861
rect 4843 21796 4844 21860
rect 4908 21796 4909 21860
rect 4843 21795 4909 21796
rect 4659 18052 4725 18053
rect 4659 17988 4660 18052
rect 4724 17988 4725 18052
rect 4659 17987 4725 17988
rect 4659 17916 4725 17917
rect 4659 17852 4660 17916
rect 4724 17852 4725 17916
rect 4659 17851 4725 17852
rect 3742 16630 3986 16690
rect 4110 17310 4538 17370
rect 3742 11389 3802 16630
rect 4110 11933 4170 17310
rect 4475 16964 4541 16965
rect 4475 16900 4476 16964
rect 4540 16900 4541 16964
rect 4475 16899 4541 16900
rect 4291 16692 4357 16693
rect 4291 16628 4292 16692
rect 4356 16628 4357 16692
rect 4291 16627 4357 16628
rect 4294 14925 4354 16627
rect 4291 14924 4357 14925
rect 4291 14860 4292 14924
rect 4356 14860 4357 14924
rect 4291 14859 4357 14860
rect 4107 11932 4173 11933
rect 4107 11868 4108 11932
rect 4172 11868 4173 11932
rect 4107 11867 4173 11868
rect 3739 11388 3805 11389
rect 3739 11324 3740 11388
rect 3804 11324 3805 11388
rect 3739 11323 3805 11324
rect 3555 11116 3621 11117
rect 3555 11052 3556 11116
rect 3620 11052 3621 11116
rect 3555 11051 3621 11052
rect 3004 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3324 10912
rect 3004 9824 3324 10848
rect 3004 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3324 9824
rect 2819 9756 2885 9757
rect 2819 9692 2820 9756
rect 2884 9692 2885 9756
rect 2819 9691 2885 9692
rect 3004 8736 3324 9760
rect 4478 9690 4538 16899
rect 4662 9757 4722 17851
rect 4846 12749 4906 21795
rect 5030 17101 5090 24787
rect 5214 21181 5274 40019
rect 5947 38860 6013 38861
rect 5947 38796 5948 38860
rect 6012 38796 6013 38860
rect 5947 38795 6013 38796
rect 5395 35188 5461 35189
rect 5395 35124 5396 35188
rect 5460 35124 5461 35188
rect 5395 35123 5461 35124
rect 5398 23901 5458 35123
rect 5579 33420 5645 33421
rect 5579 33356 5580 33420
rect 5644 33356 5645 33420
rect 5579 33355 5645 33356
rect 5582 30565 5642 33355
rect 5763 32876 5829 32877
rect 5763 32812 5764 32876
rect 5828 32812 5829 32876
rect 5763 32811 5829 32812
rect 5579 30564 5645 30565
rect 5579 30500 5580 30564
rect 5644 30500 5645 30564
rect 5579 30499 5645 30500
rect 5579 27980 5645 27981
rect 5579 27916 5580 27980
rect 5644 27916 5645 27980
rect 5579 27915 5645 27916
rect 5395 23900 5461 23901
rect 5395 23836 5396 23900
rect 5460 23836 5461 23900
rect 5395 23835 5461 23836
rect 5395 23084 5461 23085
rect 5395 23020 5396 23084
rect 5460 23020 5461 23084
rect 5395 23019 5461 23020
rect 5398 21453 5458 23019
rect 5582 22677 5642 27915
rect 5579 22676 5645 22677
rect 5579 22612 5580 22676
rect 5644 22612 5645 22676
rect 5579 22611 5645 22612
rect 5579 21724 5645 21725
rect 5579 21660 5580 21724
rect 5644 21660 5645 21724
rect 5579 21659 5645 21660
rect 5395 21452 5461 21453
rect 5395 21388 5396 21452
rect 5460 21388 5461 21452
rect 5395 21387 5461 21388
rect 5211 21180 5277 21181
rect 5211 21116 5212 21180
rect 5276 21116 5277 21180
rect 5211 21115 5277 21116
rect 5582 18730 5642 21659
rect 5214 18670 5642 18730
rect 5027 17100 5093 17101
rect 5027 17036 5028 17100
rect 5092 17036 5093 17100
rect 5027 17035 5093 17036
rect 5214 15330 5274 18670
rect 5579 18188 5645 18189
rect 5579 18124 5580 18188
rect 5644 18124 5645 18188
rect 5579 18123 5645 18124
rect 5582 15330 5642 18123
rect 5766 16149 5826 32811
rect 5950 19005 6010 38795
rect 6499 37364 6565 37365
rect 6499 37300 6500 37364
rect 6564 37300 6565 37364
rect 6499 37299 6565 37300
rect 6315 33964 6381 33965
rect 6315 33900 6316 33964
rect 6380 33900 6381 33964
rect 6315 33899 6381 33900
rect 6131 31788 6197 31789
rect 6131 31724 6132 31788
rect 6196 31724 6197 31788
rect 6131 31723 6197 31724
rect 5947 19004 6013 19005
rect 5947 18940 5948 19004
rect 6012 18940 6013 19004
rect 5947 18939 6013 18940
rect 5947 18732 6013 18733
rect 5947 18668 5948 18732
rect 6012 18668 6013 18732
rect 5947 18667 6013 18668
rect 5763 16148 5829 16149
rect 5763 16084 5764 16148
rect 5828 16084 5829 16148
rect 5763 16083 5829 16084
rect 5763 16012 5829 16013
rect 5763 15948 5764 16012
rect 5828 15948 5829 16012
rect 5763 15947 5829 15948
rect 5030 15270 5274 15330
rect 5398 15270 5642 15330
rect 5030 14925 5090 15270
rect 5398 15058 5458 15270
rect 5214 14998 5458 15058
rect 5027 14924 5093 14925
rect 5027 14860 5028 14924
rect 5092 14860 5093 14924
rect 5027 14859 5093 14860
rect 5027 13564 5093 13565
rect 5027 13500 5028 13564
rect 5092 13500 5093 13564
rect 5027 13499 5093 13500
rect 4843 12748 4909 12749
rect 4843 12684 4844 12748
rect 4908 12684 4909 12748
rect 4843 12683 4909 12684
rect 4659 9756 4725 9757
rect 4659 9692 4660 9756
rect 4724 9692 4725 9756
rect 4659 9691 4725 9692
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 2451 8260 2517 8261
rect 2451 8196 2452 8260
rect 2516 8196 2517 8260
rect 2451 8195 2517 8196
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1163 7988 1229 7989
rect 1163 7924 1164 7988
rect 1228 7924 1229 7988
rect 1163 7923 1229 7924
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 979 1324 1045 1325
rect 979 1260 980 1324
rect 1044 1260 1045 1324
rect 979 1259 1045 1260
rect 611 1188 677 1189
rect 611 1124 612 1188
rect 676 1124 677 1188
rect 611 1123 677 1124
rect 1944 0 2264 2688
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3926 9630 4538 9690
rect 3926 2685 3986 9630
rect 5030 2790 5090 13499
rect 4846 2730 5090 2790
rect 3923 2684 3989 2685
rect 3923 2620 3924 2684
rect 3988 2620 3989 2684
rect 3923 2619 3989 2620
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 4846 1189 4906 2730
rect 5214 1325 5274 14998
rect 5395 14924 5461 14925
rect 5395 14860 5396 14924
rect 5460 14860 5461 14924
rect 5395 14859 5461 14860
rect 5398 7581 5458 14859
rect 5579 13700 5645 13701
rect 5579 13636 5580 13700
rect 5644 13636 5645 13700
rect 5579 13635 5645 13636
rect 5395 7580 5461 7581
rect 5395 7516 5396 7580
rect 5460 7516 5461 7580
rect 5395 7515 5461 7516
rect 5582 5813 5642 13635
rect 5766 5949 5826 15947
rect 5950 11933 6010 18667
rect 5947 11932 6013 11933
rect 5947 11868 5948 11932
rect 6012 11868 6013 11932
rect 5947 11867 6013 11868
rect 6134 11661 6194 31723
rect 6318 17917 6378 33899
rect 6502 30429 6562 37299
rect 6867 37228 6933 37229
rect 6867 37164 6868 37228
rect 6932 37164 6933 37228
rect 6867 37163 6933 37164
rect 6870 34237 6930 37163
rect 7419 35868 7485 35869
rect 7419 35804 7420 35868
rect 7484 35804 7485 35868
rect 7419 35803 7485 35804
rect 7051 34508 7117 34509
rect 7051 34444 7052 34508
rect 7116 34444 7117 34508
rect 7051 34443 7117 34444
rect 6867 34236 6933 34237
rect 6867 34172 6868 34236
rect 6932 34172 6933 34236
rect 6867 34171 6933 34172
rect 6499 30428 6565 30429
rect 6499 30364 6500 30428
rect 6564 30364 6565 30428
rect 6499 30363 6565 30364
rect 7054 30293 7114 34443
rect 7235 31788 7301 31789
rect 7235 31724 7236 31788
rect 7300 31724 7301 31788
rect 7235 31723 7301 31724
rect 7238 31517 7298 31723
rect 7235 31516 7301 31517
rect 7235 31452 7236 31516
rect 7300 31452 7301 31516
rect 7235 31451 7301 31452
rect 7051 30292 7117 30293
rect 7051 30228 7052 30292
rect 7116 30228 7117 30292
rect 7051 30227 7117 30228
rect 7051 30156 7117 30157
rect 7051 30092 7052 30156
rect 7116 30092 7117 30156
rect 7051 30091 7117 30092
rect 6867 29340 6933 29341
rect 6867 29276 6868 29340
rect 6932 29276 6933 29340
rect 6867 29275 6933 29276
rect 6499 28660 6565 28661
rect 6499 28596 6500 28660
rect 6564 28596 6565 28660
rect 6499 28595 6565 28596
rect 6502 25397 6562 28595
rect 6683 28524 6749 28525
rect 6683 28460 6684 28524
rect 6748 28460 6749 28524
rect 6683 28459 6749 28460
rect 6499 25396 6565 25397
rect 6499 25332 6500 25396
rect 6564 25332 6565 25396
rect 6499 25331 6565 25332
rect 6499 22812 6565 22813
rect 6499 22748 6500 22812
rect 6564 22748 6565 22812
rect 6499 22747 6565 22748
rect 6502 21589 6562 22747
rect 6686 22269 6746 28459
rect 6870 24853 6930 29275
rect 7054 25805 7114 30091
rect 7235 28660 7301 28661
rect 7235 28596 7236 28660
rect 7300 28596 7301 28660
rect 7235 28595 7301 28596
rect 7238 27978 7298 28595
rect 7422 28253 7482 35803
rect 7790 35733 7850 40291
rect 7944 39744 8264 40768
rect 7944 39680 7952 39744
rect 8016 39680 8032 39744
rect 8096 39680 8112 39744
rect 8176 39680 8192 39744
rect 8256 39680 8264 39744
rect 7944 38656 8264 39680
rect 9004 42464 9324 45000
rect 9004 42400 9012 42464
rect 9076 42400 9092 42464
rect 9156 42400 9172 42464
rect 9236 42400 9252 42464
rect 9316 42400 9324 42464
rect 9004 41376 9324 42400
rect 9004 41312 9012 41376
rect 9076 41312 9092 41376
rect 9156 41312 9172 41376
rect 9236 41312 9252 41376
rect 9316 41312 9324 41376
rect 9004 40288 9324 41312
rect 9811 40356 9877 40357
rect 9811 40292 9812 40356
rect 9876 40292 9877 40356
rect 9811 40291 9877 40292
rect 9004 40224 9012 40288
rect 9076 40224 9092 40288
rect 9156 40224 9172 40288
rect 9236 40224 9252 40288
rect 9316 40224 9324 40288
rect 8707 39404 8773 39405
rect 8707 39340 8708 39404
rect 8772 39340 8773 39404
rect 8707 39339 8773 39340
rect 8339 38724 8405 38725
rect 8339 38660 8340 38724
rect 8404 38660 8405 38724
rect 8339 38659 8405 38660
rect 7944 38592 7952 38656
rect 8016 38592 8032 38656
rect 8096 38592 8112 38656
rect 8176 38592 8192 38656
rect 8256 38592 8264 38656
rect 7944 37568 8264 38592
rect 7944 37504 7952 37568
rect 8016 37504 8032 37568
rect 8096 37504 8112 37568
rect 8176 37504 8192 37568
rect 8256 37504 8264 37568
rect 7944 36480 8264 37504
rect 7944 36416 7952 36480
rect 8016 36416 8032 36480
rect 8096 36416 8112 36480
rect 8176 36416 8192 36480
rect 8256 36416 8264 36480
rect 7787 35732 7853 35733
rect 7787 35668 7788 35732
rect 7852 35668 7853 35732
rect 7787 35667 7853 35668
rect 7944 35392 8264 36416
rect 7944 35328 7952 35392
rect 8016 35328 8032 35392
rect 8096 35328 8112 35392
rect 8176 35328 8192 35392
rect 8256 35328 8264 35392
rect 7944 34304 8264 35328
rect 7944 34240 7952 34304
rect 8016 34240 8032 34304
rect 8096 34240 8112 34304
rect 8176 34240 8192 34304
rect 8256 34240 8264 34304
rect 7944 33216 8264 34240
rect 7944 33152 7952 33216
rect 8016 33152 8032 33216
rect 8096 33152 8112 33216
rect 8176 33152 8192 33216
rect 8256 33152 8264 33216
rect 7787 32740 7853 32741
rect 7787 32676 7788 32740
rect 7852 32676 7853 32740
rect 7787 32675 7853 32676
rect 7603 32332 7669 32333
rect 7603 32268 7604 32332
rect 7668 32268 7669 32332
rect 7603 32267 7669 32268
rect 7419 28252 7485 28253
rect 7419 28188 7420 28252
rect 7484 28188 7485 28252
rect 7419 28187 7485 28188
rect 7238 27918 7482 27978
rect 7235 27844 7301 27845
rect 7235 27780 7236 27844
rect 7300 27780 7301 27844
rect 7235 27779 7301 27780
rect 7051 25804 7117 25805
rect 7051 25740 7052 25804
rect 7116 25740 7117 25804
rect 7051 25739 7117 25740
rect 6867 24852 6933 24853
rect 6867 24788 6868 24852
rect 6932 24788 6933 24852
rect 6867 24787 6933 24788
rect 6867 24716 6933 24717
rect 6867 24652 6868 24716
rect 6932 24652 6933 24716
rect 6867 24651 6933 24652
rect 6683 22268 6749 22269
rect 6683 22204 6684 22268
rect 6748 22204 6749 22268
rect 6683 22203 6749 22204
rect 6870 22130 6930 24651
rect 7054 22677 7114 25739
rect 7238 23493 7298 27779
rect 7422 25125 7482 27918
rect 7419 25124 7485 25125
rect 7419 25060 7420 25124
rect 7484 25060 7485 25124
rect 7419 25059 7485 25060
rect 7419 24852 7485 24853
rect 7419 24788 7420 24852
rect 7484 24788 7485 24852
rect 7419 24787 7485 24788
rect 7235 23492 7301 23493
rect 7235 23428 7236 23492
rect 7300 23428 7301 23492
rect 7235 23427 7301 23428
rect 7051 22676 7117 22677
rect 7051 22612 7052 22676
rect 7116 22612 7117 22676
rect 7051 22611 7117 22612
rect 6686 22070 6930 22130
rect 6499 21588 6565 21589
rect 6499 21524 6500 21588
rect 6564 21524 6565 21588
rect 6499 21523 6565 21524
rect 6686 19685 6746 22070
rect 7054 21861 7114 22611
rect 7235 22268 7301 22269
rect 7235 22204 7236 22268
rect 7300 22204 7301 22268
rect 7235 22203 7301 22204
rect 7051 21860 7117 21861
rect 7051 21796 7052 21860
rect 7116 21796 7117 21860
rect 7051 21795 7117 21796
rect 6867 21316 6933 21317
rect 6867 21252 6868 21316
rect 6932 21252 6933 21316
rect 6867 21251 6933 21252
rect 6683 19684 6749 19685
rect 6683 19620 6684 19684
rect 6748 19620 6749 19684
rect 6683 19619 6749 19620
rect 6683 18868 6749 18869
rect 6683 18804 6684 18868
rect 6748 18804 6749 18868
rect 6683 18803 6749 18804
rect 6315 17916 6381 17917
rect 6315 17852 6316 17916
rect 6380 17852 6381 17916
rect 6315 17851 6381 17852
rect 6499 16556 6565 16557
rect 6499 16492 6500 16556
rect 6564 16492 6565 16556
rect 6499 16491 6565 16492
rect 6131 11660 6197 11661
rect 6131 11596 6132 11660
rect 6196 11596 6197 11660
rect 6131 11595 6197 11596
rect 6502 5949 6562 16491
rect 6686 14653 6746 18803
rect 6870 18189 6930 21251
rect 7238 20770 7298 22203
rect 7054 20710 7298 20770
rect 6867 18188 6933 18189
rect 6867 18124 6868 18188
rect 6932 18124 6933 18188
rect 6867 18123 6933 18124
rect 6683 14652 6749 14653
rect 6683 14588 6684 14652
rect 6748 14588 6749 14652
rect 6683 14587 6749 14588
rect 6683 14516 6749 14517
rect 6683 14452 6684 14516
rect 6748 14452 6749 14516
rect 6683 14451 6749 14452
rect 6686 10165 6746 14451
rect 7054 10573 7114 20710
rect 7235 20636 7301 20637
rect 7235 20572 7236 20636
rect 7300 20572 7301 20636
rect 7235 20571 7301 20572
rect 7238 15741 7298 20571
rect 7235 15740 7301 15741
rect 7235 15676 7236 15740
rect 7300 15676 7301 15740
rect 7235 15675 7301 15676
rect 7422 13565 7482 24787
rect 7606 16149 7666 32267
rect 7790 29749 7850 32675
rect 7944 32128 8264 33152
rect 7944 32064 7952 32128
rect 8016 32064 8032 32128
rect 8096 32064 8112 32128
rect 8176 32064 8192 32128
rect 8256 32064 8264 32128
rect 7944 31040 8264 32064
rect 7944 30976 7952 31040
rect 8016 30976 8032 31040
rect 8096 30976 8112 31040
rect 8176 30976 8192 31040
rect 8256 30976 8264 31040
rect 7944 29952 8264 30976
rect 8342 30429 8402 38659
rect 8523 35868 8589 35869
rect 8523 35804 8524 35868
rect 8588 35804 8589 35868
rect 8523 35803 8589 35804
rect 8526 33013 8586 35803
rect 8523 33012 8589 33013
rect 8523 32948 8524 33012
rect 8588 32948 8589 33012
rect 8523 32947 8589 32948
rect 8523 31516 8589 31517
rect 8523 31452 8524 31516
rect 8588 31452 8589 31516
rect 8523 31451 8589 31452
rect 8339 30428 8405 30429
rect 8339 30364 8340 30428
rect 8404 30364 8405 30428
rect 8339 30363 8405 30364
rect 7944 29888 7952 29952
rect 8016 29888 8032 29952
rect 8096 29888 8112 29952
rect 8176 29888 8192 29952
rect 8256 29888 8264 29952
rect 7787 29748 7853 29749
rect 7787 29684 7788 29748
rect 7852 29684 7853 29748
rect 7787 29683 7853 29684
rect 7944 28864 8264 29888
rect 7944 28800 7952 28864
rect 8016 28800 8032 28864
rect 8096 28800 8112 28864
rect 8176 28800 8192 28864
rect 8256 28800 8264 28864
rect 7787 27980 7853 27981
rect 7787 27916 7788 27980
rect 7852 27916 7853 27980
rect 7787 27915 7853 27916
rect 7790 24989 7850 27915
rect 7944 27776 8264 28800
rect 8339 28660 8405 28661
rect 8339 28596 8340 28660
rect 8404 28596 8405 28660
rect 8339 28595 8405 28596
rect 7944 27712 7952 27776
rect 8016 27712 8032 27776
rect 8096 27712 8112 27776
rect 8176 27712 8192 27776
rect 8256 27712 8264 27776
rect 7944 26688 8264 27712
rect 7944 26624 7952 26688
rect 8016 26624 8032 26688
rect 8096 26624 8112 26688
rect 8176 26624 8192 26688
rect 8256 26624 8264 26688
rect 7944 25600 8264 26624
rect 8342 26482 8402 28595
rect 8526 27437 8586 31451
rect 8710 27573 8770 39339
rect 9004 39200 9324 40224
rect 9004 39136 9012 39200
rect 9076 39136 9092 39200
rect 9156 39136 9172 39200
rect 9236 39136 9252 39200
rect 9316 39136 9324 39200
rect 9004 38112 9324 39136
rect 9004 38048 9012 38112
rect 9076 38048 9092 38112
rect 9156 38048 9172 38112
rect 9236 38048 9252 38112
rect 9316 38048 9324 38112
rect 9004 37024 9324 38048
rect 9004 36960 9012 37024
rect 9076 36960 9092 37024
rect 9156 36960 9172 37024
rect 9236 36960 9252 37024
rect 9316 36960 9324 37024
rect 9004 35936 9324 36960
rect 9004 35872 9012 35936
rect 9076 35872 9092 35936
rect 9156 35872 9172 35936
rect 9236 35872 9252 35936
rect 9316 35872 9324 35936
rect 9004 34848 9324 35872
rect 9443 35188 9509 35189
rect 9443 35124 9444 35188
rect 9508 35124 9509 35188
rect 9443 35123 9509 35124
rect 9004 34784 9012 34848
rect 9076 34784 9092 34848
rect 9156 34784 9172 34848
rect 9236 34784 9252 34848
rect 9316 34784 9324 34848
rect 9004 33760 9324 34784
rect 9004 33696 9012 33760
rect 9076 33696 9092 33760
rect 9156 33696 9172 33760
rect 9236 33696 9252 33760
rect 9316 33696 9324 33760
rect 9004 32672 9324 33696
rect 9004 32608 9012 32672
rect 9076 32608 9092 32672
rect 9156 32608 9172 32672
rect 9236 32608 9252 32672
rect 9316 32608 9324 32672
rect 9004 31584 9324 32608
rect 9004 31520 9012 31584
rect 9076 31520 9092 31584
rect 9156 31520 9172 31584
rect 9236 31520 9252 31584
rect 9316 31520 9324 31584
rect 9004 30496 9324 31520
rect 9004 30432 9012 30496
rect 9076 30432 9092 30496
rect 9156 30432 9172 30496
rect 9236 30432 9252 30496
rect 9316 30432 9324 30496
rect 9004 29408 9324 30432
rect 9004 29344 9012 29408
rect 9076 29344 9092 29408
rect 9156 29344 9172 29408
rect 9236 29344 9252 29408
rect 9316 29344 9324 29408
rect 9004 28320 9324 29344
rect 9004 28256 9012 28320
rect 9076 28256 9092 28320
rect 9156 28256 9172 28320
rect 9236 28256 9252 28320
rect 9316 28256 9324 28320
rect 8707 27572 8773 27573
rect 8707 27508 8708 27572
rect 8772 27508 8773 27572
rect 8707 27507 8773 27508
rect 8523 27436 8589 27437
rect 8523 27372 8524 27436
rect 8588 27372 8589 27436
rect 8523 27371 8589 27372
rect 9004 27232 9324 28256
rect 9446 28117 9506 35123
rect 9627 30972 9693 30973
rect 9627 30908 9628 30972
rect 9692 30908 9693 30972
rect 9627 30907 9693 30908
rect 9443 28116 9509 28117
rect 9443 28052 9444 28116
rect 9508 28052 9509 28116
rect 9443 28051 9509 28052
rect 9630 27981 9690 30907
rect 9627 27980 9693 27981
rect 9627 27916 9628 27980
rect 9692 27916 9693 27980
rect 9627 27915 9693 27916
rect 9443 27708 9509 27709
rect 9443 27644 9444 27708
rect 9508 27644 9509 27708
rect 9443 27643 9509 27644
rect 9004 27168 9012 27232
rect 9076 27168 9092 27232
rect 9156 27168 9172 27232
rect 9236 27168 9252 27232
rect 9316 27168 9324 27232
rect 8707 26892 8773 26893
rect 8707 26828 8708 26892
rect 8772 26828 8773 26892
rect 8707 26827 8773 26828
rect 8342 26422 8586 26482
rect 8339 26348 8405 26349
rect 8339 26284 8340 26348
rect 8404 26284 8405 26348
rect 8339 26283 8405 26284
rect 7944 25536 7952 25600
rect 8016 25536 8032 25600
rect 8096 25536 8112 25600
rect 8176 25536 8192 25600
rect 8256 25536 8264 25600
rect 7787 24988 7853 24989
rect 7787 24924 7788 24988
rect 7852 24924 7853 24988
rect 7787 24923 7853 24924
rect 7787 24716 7853 24717
rect 7787 24652 7788 24716
rect 7852 24652 7853 24716
rect 7787 24651 7853 24652
rect 7790 19413 7850 24651
rect 7944 24512 8264 25536
rect 7944 24448 7952 24512
rect 8016 24448 8032 24512
rect 8096 24448 8112 24512
rect 8176 24448 8192 24512
rect 8256 24448 8264 24512
rect 7944 23424 8264 24448
rect 7944 23360 7952 23424
rect 8016 23360 8032 23424
rect 8096 23360 8112 23424
rect 8176 23360 8192 23424
rect 8256 23360 8264 23424
rect 7944 22336 8264 23360
rect 7944 22272 7952 22336
rect 8016 22272 8032 22336
rect 8096 22272 8112 22336
rect 8176 22272 8192 22336
rect 8256 22272 8264 22336
rect 7944 21248 8264 22272
rect 7944 21184 7952 21248
rect 8016 21184 8032 21248
rect 8096 21184 8112 21248
rect 8176 21184 8192 21248
rect 8256 21184 8264 21248
rect 7944 20160 8264 21184
rect 7944 20096 7952 20160
rect 8016 20096 8032 20160
rect 8096 20096 8112 20160
rect 8176 20096 8192 20160
rect 8256 20096 8264 20160
rect 7787 19412 7853 19413
rect 7787 19348 7788 19412
rect 7852 19348 7853 19412
rect 7787 19347 7853 19348
rect 7944 19072 8264 20096
rect 7944 19008 7952 19072
rect 8016 19008 8032 19072
rect 8096 19008 8112 19072
rect 8176 19008 8192 19072
rect 8256 19008 8264 19072
rect 7787 18188 7853 18189
rect 7787 18124 7788 18188
rect 7852 18124 7853 18188
rect 7787 18123 7853 18124
rect 7790 17101 7850 18123
rect 7944 17984 8264 19008
rect 7944 17920 7952 17984
rect 8016 17920 8032 17984
rect 8096 17920 8112 17984
rect 8176 17920 8192 17984
rect 8256 17920 8264 17984
rect 7787 17100 7853 17101
rect 7787 17036 7788 17100
rect 7852 17036 7853 17100
rect 7787 17035 7853 17036
rect 7603 16148 7669 16149
rect 7603 16084 7604 16148
rect 7668 16084 7669 16148
rect 7603 16083 7669 16084
rect 7603 15468 7669 15469
rect 7603 15404 7604 15468
rect 7668 15404 7669 15468
rect 7603 15403 7669 15404
rect 7606 13837 7666 15403
rect 7603 13836 7669 13837
rect 7603 13772 7604 13836
rect 7668 13772 7669 13836
rect 7603 13771 7669 13772
rect 7419 13564 7485 13565
rect 7419 13500 7420 13564
rect 7484 13500 7485 13564
rect 7419 13499 7485 13500
rect 7790 13021 7850 17035
rect 7944 16896 8264 17920
rect 7944 16832 7952 16896
rect 8016 16832 8032 16896
rect 8096 16832 8112 16896
rect 8176 16832 8192 16896
rect 8256 16832 8264 16896
rect 7944 15808 8264 16832
rect 7944 15744 7952 15808
rect 8016 15744 8032 15808
rect 8096 15744 8112 15808
rect 8176 15744 8192 15808
rect 8256 15744 8264 15808
rect 7944 14720 8264 15744
rect 7944 14656 7952 14720
rect 8016 14656 8032 14720
rect 8096 14656 8112 14720
rect 8176 14656 8192 14720
rect 8256 14656 8264 14720
rect 7944 13632 8264 14656
rect 8342 14653 8402 26283
rect 8526 23901 8586 26422
rect 8523 23900 8589 23901
rect 8523 23836 8524 23900
rect 8588 23836 8589 23900
rect 8523 23835 8589 23836
rect 8523 23764 8589 23765
rect 8523 23700 8524 23764
rect 8588 23700 8589 23764
rect 8523 23699 8589 23700
rect 8339 14652 8405 14653
rect 8339 14588 8340 14652
rect 8404 14588 8405 14652
rect 8339 14587 8405 14588
rect 8339 13836 8405 13837
rect 8339 13772 8340 13836
rect 8404 13772 8405 13836
rect 8339 13771 8405 13772
rect 7944 13568 7952 13632
rect 8016 13568 8032 13632
rect 8096 13568 8112 13632
rect 8176 13568 8192 13632
rect 8256 13568 8264 13632
rect 7787 13020 7853 13021
rect 7787 12956 7788 13020
rect 7852 12956 7853 13020
rect 7787 12955 7853 12956
rect 7944 12544 8264 13568
rect 7944 12480 7952 12544
rect 8016 12480 8032 12544
rect 8096 12480 8112 12544
rect 8176 12480 8192 12544
rect 8256 12480 8264 12544
rect 7944 11456 8264 12480
rect 8342 11525 8402 13771
rect 8526 12341 8586 23699
rect 8710 21997 8770 26827
rect 9004 26144 9324 27168
rect 9004 26080 9012 26144
rect 9076 26080 9092 26144
rect 9156 26080 9172 26144
rect 9236 26080 9252 26144
rect 9316 26080 9324 26144
rect 9004 25056 9324 26080
rect 9004 24992 9012 25056
rect 9076 24992 9092 25056
rect 9156 24992 9172 25056
rect 9236 24992 9252 25056
rect 9316 24992 9324 25056
rect 9004 23968 9324 24992
rect 9004 23904 9012 23968
rect 9076 23904 9092 23968
rect 9156 23904 9172 23968
rect 9236 23904 9252 23968
rect 9316 23904 9324 23968
rect 9004 22880 9324 23904
rect 9004 22816 9012 22880
rect 9076 22816 9092 22880
rect 9156 22816 9172 22880
rect 9236 22816 9252 22880
rect 9316 22816 9324 22880
rect 8707 21996 8773 21997
rect 8707 21932 8708 21996
rect 8772 21932 8773 21996
rect 8707 21931 8773 21932
rect 9004 21792 9324 22816
rect 9004 21728 9012 21792
rect 9076 21728 9092 21792
rect 9156 21728 9172 21792
rect 9236 21728 9252 21792
rect 9316 21728 9324 21792
rect 8707 21724 8773 21725
rect 8707 21660 8708 21724
rect 8772 21660 8773 21724
rect 8707 21659 8773 21660
rect 8710 20365 8770 21659
rect 9004 20704 9324 21728
rect 9004 20640 9012 20704
rect 9076 20640 9092 20704
rect 9156 20640 9172 20704
rect 9236 20640 9252 20704
rect 9316 20640 9324 20704
rect 8707 20364 8773 20365
rect 8707 20300 8708 20364
rect 8772 20300 8773 20364
rect 8707 20299 8773 20300
rect 9004 19616 9324 20640
rect 9004 19552 9012 19616
rect 9076 19552 9092 19616
rect 9156 19552 9172 19616
rect 9236 19552 9252 19616
rect 9316 19552 9324 19616
rect 8707 18868 8773 18869
rect 8707 18804 8708 18868
rect 8772 18804 8773 18868
rect 8707 18803 8773 18804
rect 8523 12340 8589 12341
rect 8523 12276 8524 12340
rect 8588 12276 8589 12340
rect 8523 12275 8589 12276
rect 8339 11524 8405 11525
rect 8339 11460 8340 11524
rect 8404 11460 8405 11524
rect 8339 11459 8405 11460
rect 7944 11392 7952 11456
rect 8016 11392 8032 11456
rect 8096 11392 8112 11456
rect 8176 11392 8192 11456
rect 8256 11392 8264 11456
rect 7051 10572 7117 10573
rect 7051 10508 7052 10572
rect 7116 10508 7117 10572
rect 7051 10507 7117 10508
rect 7944 10368 8264 11392
rect 7944 10304 7952 10368
rect 8016 10304 8032 10368
rect 8096 10304 8112 10368
rect 8176 10304 8192 10368
rect 8256 10304 8264 10368
rect 6683 10164 6749 10165
rect 6683 10100 6684 10164
rect 6748 10100 6749 10164
rect 6683 10099 6749 10100
rect 7944 9280 8264 10304
rect 8342 10165 8402 11459
rect 8339 10164 8405 10165
rect 8339 10100 8340 10164
rect 8404 10100 8405 10164
rect 8339 10099 8405 10100
rect 7944 9216 7952 9280
rect 8016 9216 8032 9280
rect 8096 9216 8112 9280
rect 8176 9216 8192 9280
rect 8256 9216 8264 9280
rect 7944 8192 8264 9216
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 8710 6901 8770 18803
rect 9004 18528 9324 19552
rect 9004 18464 9012 18528
rect 9076 18464 9092 18528
rect 9156 18464 9172 18528
rect 9236 18464 9252 18528
rect 9316 18464 9324 18528
rect 9004 17440 9324 18464
rect 9004 17376 9012 17440
rect 9076 17376 9092 17440
rect 9156 17376 9172 17440
rect 9236 17376 9252 17440
rect 9316 17376 9324 17440
rect 9004 16352 9324 17376
rect 9004 16288 9012 16352
rect 9076 16288 9092 16352
rect 9156 16288 9172 16352
rect 9236 16288 9252 16352
rect 9316 16288 9324 16352
rect 9004 15264 9324 16288
rect 9446 15605 9506 27643
rect 9627 26076 9693 26077
rect 9627 26012 9628 26076
rect 9692 26012 9693 26076
rect 9627 26011 9693 26012
rect 9630 20501 9690 26011
rect 9627 20500 9693 20501
rect 9627 20436 9628 20500
rect 9692 20436 9693 20500
rect 9627 20435 9693 20436
rect 9627 17916 9693 17917
rect 9627 17852 9628 17916
rect 9692 17852 9693 17916
rect 9627 17851 9693 17852
rect 9443 15604 9509 15605
rect 9443 15540 9444 15604
rect 9508 15540 9509 15604
rect 9443 15539 9509 15540
rect 9004 15200 9012 15264
rect 9076 15200 9092 15264
rect 9156 15200 9172 15264
rect 9236 15200 9252 15264
rect 9316 15200 9324 15264
rect 9004 14176 9324 15200
rect 9004 14112 9012 14176
rect 9076 14112 9092 14176
rect 9156 14112 9172 14176
rect 9236 14112 9252 14176
rect 9316 14112 9324 14176
rect 9004 13088 9324 14112
rect 9004 13024 9012 13088
rect 9076 13024 9092 13088
rect 9156 13024 9172 13088
rect 9236 13024 9252 13088
rect 9316 13024 9324 13088
rect 9004 12000 9324 13024
rect 9004 11936 9012 12000
rect 9076 11936 9092 12000
rect 9156 11936 9172 12000
rect 9236 11936 9252 12000
rect 9316 11936 9324 12000
rect 9004 10912 9324 11936
rect 9630 11797 9690 17851
rect 9627 11796 9693 11797
rect 9627 11732 9628 11796
rect 9692 11732 9693 11796
rect 9627 11731 9693 11732
rect 9004 10848 9012 10912
rect 9076 10848 9092 10912
rect 9156 10848 9172 10912
rect 9236 10848 9252 10912
rect 9316 10848 9324 10912
rect 9004 9824 9324 10848
rect 9004 9760 9012 9824
rect 9076 9760 9092 9824
rect 9156 9760 9172 9824
rect 9236 9760 9252 9824
rect 9316 9760 9324 9824
rect 9004 8736 9324 9760
rect 9443 9484 9509 9485
rect 9443 9420 9444 9484
rect 9508 9420 9509 9484
rect 9443 9419 9509 9420
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9446 7717 9506 9419
rect 9443 7716 9509 7717
rect 9443 7652 9444 7716
rect 9508 7652 9509 7716
rect 9443 7651 9509 7652
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 8707 6900 8773 6901
rect 8707 6836 8708 6900
rect 8772 6836 8773 6900
rect 8707 6835 8773 6836
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 5763 5948 5829 5949
rect 5763 5884 5764 5948
rect 5828 5884 5829 5948
rect 5763 5883 5829 5884
rect 6499 5948 6565 5949
rect 6499 5884 6500 5948
rect 6564 5884 6565 5948
rect 6499 5883 6565 5884
rect 5579 5812 5645 5813
rect 5579 5748 5580 5812
rect 5644 5748 5645 5812
rect 5579 5747 5645 5748
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 5211 1324 5277 1325
rect 5211 1260 5212 1324
rect 5276 1260 5277 1324
rect 5211 1259 5277 1260
rect 4843 1188 4909 1189
rect 4843 1124 4844 1188
rect 4908 1124 4909 1188
rect 4843 1123 4909 1124
rect 7944 0 8264 2688
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9814 5133 9874 40291
rect 10179 40220 10245 40221
rect 10179 40156 10180 40220
rect 10244 40156 10245 40220
rect 10179 40155 10245 40156
rect 9995 35732 10061 35733
rect 9995 35668 9996 35732
rect 10060 35668 10061 35732
rect 9995 35667 10061 35668
rect 9998 26213 10058 35667
rect 9995 26212 10061 26213
rect 9995 26148 9996 26212
rect 10060 26148 10061 26212
rect 9995 26147 10061 26148
rect 9995 22540 10061 22541
rect 9995 22476 9996 22540
rect 10060 22476 10061 22540
rect 9995 22475 10061 22476
rect 9998 17917 10058 22475
rect 9995 17916 10061 17917
rect 9995 17852 9996 17916
rect 10060 17852 10061 17916
rect 9995 17851 10061 17852
rect 9811 5132 9877 5133
rect 9811 5068 9812 5132
rect 9876 5068 9877 5132
rect 9811 5067 9877 5068
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 10182 1325 10242 40155
rect 10547 39676 10613 39677
rect 10547 39612 10548 39676
rect 10612 39612 10613 39676
rect 10547 39611 10613 39612
rect 10363 38316 10429 38317
rect 10363 38252 10364 38316
rect 10428 38252 10429 38316
rect 10363 38251 10429 38252
rect 10366 16013 10426 38251
rect 10363 16012 10429 16013
rect 10363 15948 10364 16012
rect 10428 15948 10429 16012
rect 10363 15947 10429 15948
rect 10179 1324 10245 1325
rect 10179 1260 10180 1324
rect 10244 1260 10245 1324
rect 10179 1259 10245 1260
rect 10550 1189 10610 39611
rect 10915 28796 10981 28797
rect 10915 28732 10916 28796
rect 10980 28732 10981 28796
rect 10915 28731 10981 28732
rect 10731 25804 10797 25805
rect 10731 25740 10732 25804
rect 10796 25740 10797 25804
rect 10731 25739 10797 25740
rect 10734 19549 10794 25739
rect 10918 22110 10978 28731
rect 10918 22050 11162 22110
rect 10915 21724 10981 21725
rect 10915 21660 10916 21724
rect 10980 21660 10981 21724
rect 10915 21659 10981 21660
rect 10731 19548 10797 19549
rect 10731 19484 10732 19548
rect 10796 19484 10797 19548
rect 10731 19483 10797 19484
rect 10918 18733 10978 21659
rect 10915 18732 10981 18733
rect 10915 18668 10916 18732
rect 10980 18668 10981 18732
rect 10915 18667 10981 18668
rect 11102 12450 11162 22050
rect 10918 12390 11162 12450
rect 10918 6765 10978 12390
rect 10915 6764 10981 6765
rect 10915 6700 10916 6764
rect 10980 6700 10981 6764
rect 10915 6699 10981 6700
rect 10547 1188 10613 1189
rect 10547 1124 10548 1188
rect 10612 1124 10613 1188
rect 10547 1123 10613 1124
use sky130_fd_sc_hd__inv_1  _032_
timestamp -3599
transform 1 0 6624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp -3599
transform 1 0 6440 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _034_
timestamp -3599
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _035_
timestamp -3599
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _036_
timestamp -3599
transform -1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _037_
timestamp -3599
transform -1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _038_
timestamp -3599
transform 1 0 5428 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _039_
timestamp -3599
transform -1 0 7360 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _040_
timestamp -3599
transform 1 0 4968 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _041_
timestamp -3599
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _042_
timestamp -3599
transform 1 0 7452 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _043_
timestamp -3599
transform 1 0 7360 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _044_
timestamp -3599
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _045_
timestamp -3599
transform -1 0 7544 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _046_
timestamp -3599
transform 1 0 7084 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _047_
timestamp -3599
transform 1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _048_
timestamp -3599
transform 1 0 5060 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _049_
timestamp -3599
transform -1 0 8740 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _050_
timestamp -3599
transform 1 0 6900 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _051_
timestamp -3599
transform 1 0 7544 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _052_
timestamp -3599
transform -1 0 9752 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _053_
timestamp -3599
transform -1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _054_
timestamp -3599
transform 1 0 7544 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _055_
timestamp -3599
transform 1 0 7452 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _056_
timestamp -3599
transform -1 0 9108 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _057_
timestamp -3599
transform -1 0 4416 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _058_
timestamp -3599
transform 1 0 7636 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _059_
timestamp -3599
transform 1 0 6900 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _060_
timestamp -3599
transform 1 0 2484 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _061_
timestamp -3599
transform 1 0 2760 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _062_
timestamp -3599
transform -1 0 5612 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _063_
timestamp -3599
transform 1 0 3220 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _064_
timestamp -3599
transform -1 0 4324 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _065_
timestamp -3599
transform 1 0 4600 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _066_
timestamp -3599
transform 1 0 7544 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _067_
timestamp -3599
transform -1 0 9476 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _068_
timestamp -3599
transform 1 0 7176 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _069_
timestamp -3599
transform 1 0 2484 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _070_
timestamp -3599
transform 1 0 3772 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _071_
timestamp -3599
transform -1 0 4876 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _072_
timestamp -3599
transform 1 0 4140 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _073_
timestamp -3599
transform -1 0 4324 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _074_
timestamp -3599
transform 1 0 7544 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _075_
timestamp -3599
transform 1 0 7544 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _076_
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _077_
timestamp -3599
transform 1 0 4968 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _078_
timestamp -3599
transform 1 0 7176 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _079_
timestamp -3599
transform 1 0 2484 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _080_
timestamp -3599
transform -1 0 3680 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _081_
timestamp -3599
transform 1 0 5060 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _082_
timestamp -3599
transform 1 0 7176 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _083_
timestamp -3599
transform 1 0 7636 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _084_
timestamp -3599
transform 1 0 4324 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _085_
timestamp -3599
transform 1 0 3036 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _086_
timestamp -3599
transform -1 0 9568 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _087_
timestamp -3599
transform -1 0 4784 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _088_
timestamp -3599
transform -1 0 6256 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _089_
timestamp -3599
transform 1 0 3496 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _090_
timestamp -3599
transform 1 0 7820 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _091_
timestamp -3599
transform 1 0 7544 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _092_
timestamp -3599
transform 1 0 2392 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _093_
timestamp -3599
transform 1 0 2852 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _094_
timestamp -3599
transform 1 0 6900 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _095_
timestamp -3599
transform -1 0 5704 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _096_
timestamp -3599
transform 1 0 4600 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _097_
timestamp -3599
transform -1 0 7084 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _098_
timestamp -3599
transform 1 0 8924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp -3599
transform -1 0 9568 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _100_
timestamp -3599
transform 1 0 6164 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp -3599
transform 1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _103_
timestamp -3599
transform 1 0 7452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _104_
timestamp -3599
transform -1 0 8556 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _105_
timestamp -3599
transform -1 0 9200 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _106_
timestamp -3599
transform -1 0 9568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _107_
timestamp -3599
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _108_
timestamp -3599
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _109_
timestamp -3599
transform 1 0 5888 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _110_
timestamp -3599
transform 1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _111_
timestamp -3599
transform -1 0 5612 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _112_
timestamp -3599
transform -1 0 6992 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _113_
timestamp -3599
transform -1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _114_
timestamp -3599
transform -1 0 5796 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _115_
timestamp -3599
transform 1 0 4784 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlxtp_1  _116_
timestamp -3599
transform -1 0 2668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _117_
timestamp -3599
transform -1 0 2668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _118_
timestamp -3599
transform -1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _119_
timestamp -3599
transform -1 0 6256 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _120_
timestamp -3599
transform -1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _121_
timestamp -3599
transform -1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _122_
timestamp -3599
transform -1 0 6164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _123_
timestamp -3599
transform -1 0 6072 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _124_
timestamp -3599
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _125_
timestamp -3599
transform -1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _126_
timestamp -3599
transform 1 0 7728 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _127_
timestamp -3599
transform 1 0 8372 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _128_
timestamp -3599
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _129_
timestamp -3599
transform 1 0 4784 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _130_
timestamp -3599
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _131_
timestamp -3599
transform 1 0 3956 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _132_
timestamp -3599
transform 1 0 1932 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _133_
timestamp -3599
transform 1 0 2024 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _134_
timestamp -3599
transform 1 0 5796 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _135_
timestamp -3599
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _136_
timestamp -3599
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _137_
timestamp -3599
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _138_
timestamp -3599
transform 1 0 2024 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _139_
timestamp -3599
transform 1 0 1932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _140_
timestamp -3599
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _141_
timestamp -3599
transform 1 0 7452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _142_
timestamp -3599
transform 1 0 7176 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _143_
timestamp -3599
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _144_
timestamp -3599
transform 1 0 2024 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _145_
timestamp -3599
transform 1 0 1932 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _146_
timestamp -3599
transform 1 0 4232 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _147_
timestamp -3599
transform 1 0 4416 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _148_
timestamp -3599
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _149_
timestamp -3599
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _150_
timestamp -3599
transform 1 0 7544 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _151_
timestamp -3599
transform 1 0 7176 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _152_
timestamp -3599
transform 1 0 1840 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _153_
timestamp -3599
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _154_
timestamp -3599
transform -1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _155_
timestamp -3599
transform 1 0 4600 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _156_
timestamp -3599
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _157_
timestamp -3599
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _158_
timestamp -3599
transform 1 0 7268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _159_
timestamp -3599
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _160_
timestamp -3599
transform 1 0 4508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _161_
timestamp -3599
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _162_
timestamp -3599
transform 1 0 1472 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _163_
timestamp -3599
transform 1 0 1472 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _164_
timestamp -3599
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _165_
timestamp -3599
transform 1 0 1932 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _166_
timestamp -3599
transform 1 0 6256 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _167_
timestamp -3599
transform 1 0 6532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _168_
timestamp -3599
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _169_
timestamp -3599
transform 1 0 1472 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _170_
timestamp -3599
transform 1 0 2576 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _171_
timestamp -3599
transform 1 0 2668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _172_
timestamp -3599
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _173_
timestamp -3599
transform 1 0 6716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _174_
timestamp -3599
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _175_
timestamp -3599
transform 1 0 6532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _176_
timestamp -3599
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _177_
timestamp -3599
transform 1 0 1656 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _178_
timestamp -3599
transform 1 0 4416 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _179_
timestamp -3599
transform -1 0 5520 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _180_
timestamp -3599
transform 1 0 2208 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _181_
timestamp -3599
transform 1 0 1840 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _182_
timestamp -3599
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _183_
timestamp -3599
transform -1 0 5704 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _184_
timestamp -3599
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _185_
timestamp -3599
transform 1 0 2024 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _186_
timestamp -3599
transform 1 0 6440 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _187_
timestamp -3599
transform 1 0 6440 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _188_
timestamp -3599
transform 1 0 6532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _189_
timestamp -3599
transform 1 0 6440 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _190_
timestamp -3599
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _191_
timestamp -3599
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _192_
timestamp -3599
transform 1 0 4232 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _193_
timestamp -3599
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _194_
timestamp -3599
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _195_
timestamp -3599
transform 1 0 1748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _196_
timestamp -3599
transform 1 0 2392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _197_
timestamp -3599
transform 1 0 2392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _198_
timestamp -3599
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _199_
timestamp -3599
transform 1 0 2576 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _200_
timestamp -3599
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _201_
timestamp -3599
transform 1 0 1656 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _202_
timestamp -3599
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _203_
timestamp -3599
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _204_
timestamp -3599
transform 1 0 6348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _205_
timestamp -3599
transform 1 0 6624 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _206_
timestamp -3599
transform 1 0 7268 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _207_
timestamp -3599
transform 1 0 6808 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _208_
timestamp -3599
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _209_
timestamp -3599
transform 1 0 1656 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _210_
timestamp -3599
transform 1 0 7544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _211_
timestamp -3599
transform 1 0 6440 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _212_
timestamp -3599
transform 1 0 2208 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _213_
timestamp -3599
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _214_
timestamp -3599
transform 1 0 6900 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _215_
timestamp -3599
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _216_
timestamp -3599
transform 1 0 2024 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _217_
timestamp -3599
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _218_
timestamp -3599
transform 1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _219_
timestamp -3599
transform 1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _220_
timestamp -3599
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _221_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _222_
timestamp -3599
transform 1 0 7544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _223_
timestamp -3599
transform -1 0 6808 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _224_
timestamp -3599
transform 1 0 4600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _225_
timestamp -3599
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _226_
timestamp -3599
transform 1 0 3864 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _227_
timestamp -3599
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _228_
timestamp -3599
transform 1 0 2668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _229_
timestamp -3599
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp -3599
transform 1 0 4232 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp -3599
transform 1 0 5704 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  _232_
timestamp -3599
transform 1 0 4416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp -3599
transform -1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp -3599
transform -1 0 8832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _235_
timestamp -3599
transform 1 0 4048 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp -3599
transform 1 0 8464 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp -3599
transform -1 0 8464 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp -3599
transform -1 0 8464 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp -3599
transform -1 0 6992 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _240_
timestamp -3599
transform 1 0 3404 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _241_
timestamp -3599
transform 1 0 3864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp -3599
transform 1 0 9568 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _243_
timestamp -3599
transform 1 0 6440 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _244_
timestamp -3599
transform 1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp -3599
transform -1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp -3599
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _247_
timestamp -3599
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _248_
timestamp -3599
transform 1 0 5704 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp -3599
transform -1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp -3599
transform -1 0 5980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _251_
timestamp -3599
transform 1 0 3956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp -3599
transform -1 0 8832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp -3599
transform -1 0 7912 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp -3599
transform -1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp -3599
transform -1 0 3588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp -3599
transform -1 0 4048 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _257_
timestamp -3599
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _258_
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _259_
timestamp -3599
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _260_
timestamp -3599
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _261_
timestamp -3599
transform 1 0 6072 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _262_
timestamp -3599
transform 1 0 6532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp -3599
transform -1 0 7728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp -3599
transform -1 0 6808 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp -3599
transform -1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp -3599
transform -1 0 1656 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _267_
timestamp -3599
transform -1 0 6624 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp -3599
transform -1 0 6440 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _269_
timestamp -3599
transform 1 0 1748 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _270_
timestamp -3599
transform 1 0 1748 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp -3599
transform -1 0 6624 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp -3599
transform -1 0 6624 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _273_
timestamp -3599
transform -1 0 2024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp -3599
transform -1 0 2484 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _275_
timestamp -3599
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _276_
timestamp -3599
transform 1 0 5428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _277_
timestamp -3599
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _278_
timestamp -3599
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _279_
timestamp -3599
transform 1 0 8372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp -3599
transform -1 0 8832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _281_
timestamp -3599
transform 1 0 5704 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _282_
timestamp -3599
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _283_
timestamp -3599
transform 1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _284_
timestamp -3599
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp -3599
transform -1 0 2392 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp -3599
transform -1 0 2668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _287_
timestamp -3599
transform -1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp -3599
transform -1 0 2024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp -3599
transform -1 0 2024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _290_
timestamp -3599
transform -1 0 8372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp -3599
transform 1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp -3599
transform 1 0 7360 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp -3599
transform 1 0 7360 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp -3599
transform 1 0 6992 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp -3599
transform 1 0 8096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp -3599
transform 1 0 8740 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp -3599
transform 1 0 6716 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp -3599
transform -1 0 6624 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp -3599
transform -1 0 7544 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp -3599
transform 1 0 8556 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp -3599
transform 1 0 8924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp -3599
transform 1 0 9476 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp -3599
transform -1 0 7912 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp -3599
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp -3599
transform 1 0 8188 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp -3599
transform 1 0 9200 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _307_
timestamp -3599
transform -1 0 6072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _308_
timestamp -3599
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp -3599
transform -1 0 6256 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp -3599
transform 1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _311_
timestamp -3599
transform -1 0 8096 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp -3599
transform -1 0 8740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _313_
timestamp -3599
transform 1 0 6348 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp -3599
transform -1 0 5060 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp -3599
transform 1 0 8188 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp -3599
transform -1 0 4508 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp -3599
transform -1 0 4600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp -3599
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp -3599
transform -1 0 8832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp -3599
transform -1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp -3599
transform 1 0 4876 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp -3599
transform -1 0 4600 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp -3599
transform -1 0 8740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _324_
timestamp -3599
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp -3599
transform -1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _326_
timestamp -3599
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp -3599
transform -1 0 8832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp -3599
transform -1 0 6808 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp -3599
transform -1 0 3680 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp -3599
transform -1 0 5704 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp -3599
transform -1 0 5888 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _332_
timestamp -3599
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 9292 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 9108 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 9660 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 6348 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 7728 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform 1 0 8556 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 9476 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 7820 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 8740 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 8372 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform -1 0 9384 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform 1 0 5520 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform 1 0 7912 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform 1 0 6992 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 7176 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform -1 0 8280 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 6716 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp -3599
transform 1 0 7360 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK
timestamp -3599
transform 1 0 5704 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp -3599
transform 1 0 5704 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp -3599
transform 1 0 6348 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp -3599
transform -1 0 5612 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp -3599
transform 1 0 8004 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp -3599
transform 1 0 3404 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp -3599
transform -1 0 5612 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout45
timestamp -3599
transform -1 0 5060 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp -3599
transform 1 0 8004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp -3599
transform -1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp -3599
transform 1 0 1840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout49
timestamp -3599
transform -1 0 3588 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp -3599
transform 1 0 4416 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout51
timestamp -3599
transform 1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp -3599
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp -3599
transform 1 0 5612 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp -3599
transform 1 0 5520 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp -3599
transform 1 0 3496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout56
timestamp -3599
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp -3599
transform 1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp -3599
transform -1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp -3599
transform 1 0 2116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17
timestamp -3599
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25
timestamp -3599
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp -3599
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp -3599
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp -3599
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636964856
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp -3599
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_7
timestamp 1636964856
transform 1 0 1748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp -3599
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_51
timestamp 1636964856
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_63
timestamp 1636964856
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp -3599
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp -3599
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1636964856
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_19
timestamp -3599
transform 1 0 2852 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp -3599
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_29
timestamp -3599
transform 1 0 3772 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_38
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_46
timestamp -3599
transform 1 0 5336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp -3599
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_23
timestamp -3599
transform 1 0 3220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp -3599
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1636964856
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_63
timestamp -3599
transform 1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp -3599
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_16
timestamp -3599
transform 1 0 2576 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp -3599
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp -3599
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_64
timestamp -3599
transform 1 0 6992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_71
timestamp -3599
transform 1 0 7636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636964856
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_64
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp -3599
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_25
timestamp 1636964856
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_37
timestamp 1636964856
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp -3599
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_7
timestamp 1636964856
transform 1 0 1748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp -3599
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -3599
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636964856
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636964856
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636964856
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp -3599
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -3599
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_90
timestamp -3599
transform 1 0 9384 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_7
timestamp -3599
transform 1 0 1748 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp -3599
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_29
timestamp -3599
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp -3599
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_64
timestamp -3599
transform 1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_79
timestamp -3599
transform 1 0 8372 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_84
timestamp -3599
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp -3599
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp -3599
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp -3599
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_49
timestamp -3599
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_61
timestamp -3599
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_74
timestamp -3599
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_5
timestamp -3599
transform 1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp -3599
transform 1 0 3128 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 1636964856
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_42
timestamp -3599
transform 1 0 4968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp -3599
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp -3599
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp -3599
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp -3599
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp -3599
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636964856
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp -3599
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp -3599
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_94
timestamp -3599
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp -3599
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp -3599
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp -3599
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp -3599
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_61
timestamp -3599
transform 1 0 6716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_69
timestamp -3599
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_5
timestamp -3599
transform 1 0 1564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_22
timestamp -3599
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp -3599
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp -3599
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp -3599
transform 1 0 7912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp -3599
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_42
timestamp 1636964856
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp -3599
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1636964856
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp -3599
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp -3599
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636964856
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636964856
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp -3599
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_59
timestamp -3599
transform 1 0 6532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_63
timestamp -3599
transform 1 0 6900 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_71
timestamp -3599
transform 1 0 7636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_94
timestamp -3599
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_40
timestamp -3599
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp -3599
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636964856
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp -3599
transform 1 0 9384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp -3599
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp -3599
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp -3599
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_37
timestamp -3599
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_62
timestamp -3599
transform 1 0 6808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp -3599
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_90
timestamp -3599
transform 1 0 9384 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp -3599
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1636964856
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1636964856
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp -3599
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp -3599
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp -3599
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp -3599
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_9
timestamp -3599
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_22
timestamp -3599
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp -3599
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_50
timestamp -3599
transform 1 0 5704 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_54
timestamp 1636964856
transform 1 0 6072 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp -3599
transform 1 0 7176 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_13
timestamp -3599
transform 1 0 2300 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_69
timestamp -3599
transform 1 0 7452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp -3599
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp -3599
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp -3599
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp -3599
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_49
timestamp 1636964856
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_73
timestamp -3599
transform 1 0 7820 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636964856
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp -3599
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp -3599
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636964856
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_69
timestamp -3599
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_17
timestamp -3599
transform 1 0 2668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp -3599
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636964856
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636964856
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_53
timestamp -3599
transform 1 0 5980 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_57
timestamp -3599
transform 1 0 6348 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_77
timestamp -3599
transform 1 0 8188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp -3599
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_22
timestamp -3599
transform 1 0 3128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_49
timestamp -3599
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp -3599
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp -3599
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp -3599
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp -3599
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -3599
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp -3599
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp -3599
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_75
timestamp -3599
transform 1 0 8004 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp -3599
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_6
timestamp -3599
transform 1 0 1656 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1636964856
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp -3599
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_69
timestamp -3599
transform 1 0 7452 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_6
timestamp -3599
transform 1 0 1656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_19
timestamp -3599
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp -3599
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp -3599
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_38
timestamp 1636964856
transform 1 0 4600 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_50
timestamp -3599
transform 1 0 5704 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_56
timestamp -3599
transform 1 0 6256 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp -3599
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp -3599
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp -3599
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_12
timestamp 1636964856
transform 1 0 2208 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_24
timestamp 1636964856
transform 1 0 3312 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_36
timestamp 1636964856
transform 1 0 4416 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp -3599
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp -3599
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_72
timestamp -3599
transform 1 0 7728 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_9
timestamp -3599
transform 1 0 1932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp -3599
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp -3599
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_35
timestamp -3599
transform 1 0 4324 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_44
timestamp 1636964856
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_56
timestamp -3599
transform 1 0 6256 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp -3599
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp -3599
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp -3599
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636964856
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_90
timestamp -3599
transform 1 0 9384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp -3599
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp -3599
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -3599
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp -3599
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp -3599
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_62
timestamp 1636964856
transform 1 0 6808 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_74
timestamp -3599
transform 1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp -3599
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_18
timestamp 1636964856
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp -3599
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_46
timestamp -3599
transform 1 0 5336 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_52
timestamp -3599
transform 1 0 5888 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_69
timestamp -3599
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_77
timestamp -3599
transform 1 0 8188 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp -3599
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp -3599
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636964856
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636964856
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_53
timestamp -3599
transform 1 0 5980 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_64
timestamp -3599
transform 1 0 6992 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp -3599
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp -3599
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_9
timestamp -3599
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_22
timestamp -3599
transform 1 0 3128 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp -3599
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -3599
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp -3599
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_65
timestamp -3599
transform 1 0 7084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp -3599
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_86
timestamp -3599
transform 1 0 9016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_6
timestamp -3599
transform 1 0 1656 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp -3599
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636964856
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_41
timestamp -3599
transform 1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_77
timestamp -3599
transform 1 0 8188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp -3599
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_6
timestamp -3599
transform 1 0 1656 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp -3599
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp -3599
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_65
timestamp -3599
transform 1 0 7084 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_89
timestamp -3599
transform 1 0 9292 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_6
timestamp -3599
transform 1 0 1656 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_10
timestamp 1636964856
transform 1 0 2024 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp -3599
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_29
timestamp -3599
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_37
timestamp -3599
transform 1 0 4508 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_52
timestamp -3599
transform 1 0 5888 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_56
timestamp -3599
transform 1 0 6256 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp -3599
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp -3599
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636964856
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636964856
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp -3599
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp -3599
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp -3599
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_71
timestamp -3599
transform 1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_94
timestamp -3599
transform 1 0 9752 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_6
timestamp -3599
transform 1 0 1656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_10
timestamp -3599
transform 1 0 2024 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp -3599
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_29
timestamp -3599
transform 1 0 3772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_35
timestamp -3599
transform 1 0 4324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_64
timestamp -3599
transform 1 0 6992 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_78
timestamp -3599
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp -3599
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_6
timestamp -3599
transform 1 0 1656 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp -3599
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp -3599
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_64
timestamp 1636964856
transform 1 0 6992 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_76
timestamp -3599
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp -3599
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_17
timestamp -3599
transform 1 0 2668 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp -3599
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp -3599
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_33
timestamp -3599
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_49
timestamp 1636964856
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_61
timestamp 1636964856
transform 1 0 6716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_73
timestamp -3599
transform 1 0 7820 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_79
timestamp -3599
transform 1 0 8372 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp -3599
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_6
timestamp -3599
transform 1 0 1656 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_35
timestamp -3599
transform 1 0 4324 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_41
timestamp -3599
transform 1 0 4876 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp -3599
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_57
timestamp -3599
transform 1 0 6348 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_70
timestamp -3599
transform 1 0 7544 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_19
timestamp -3599
transform 1 0 2852 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp -3599
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_43
timestamp -3599
transform 1 0 5060 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_53
timestamp -3599
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_57
timestamp -3599
transform 1 0 6348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_70
timestamp -3599
transform 1 0 7544 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_78
timestamp -3599
transform 1 0 8280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp -3599
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_6
timestamp -3599
transform 1 0 1656 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_19
timestamp 1636964856
transform 1 0 2852 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_31
timestamp -3599
transform 1 0 3956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp -3599
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp -3599
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp -3599
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_65
timestamp -3599
transform 1 0 7084 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_6
timestamp -3599
transform 1 0 1656 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_10
timestamp 1636964856
transform 1 0 2024 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_22
timestamp -3599
transform 1 0 3128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp -3599
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_37
timestamp -3599
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_71
timestamp -3599
transform 1 0 7636 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_94
timestamp -3599
transform 1 0 9752 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_7
timestamp 1636964856
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1636964856
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1636964856
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp -3599
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_60
timestamp -3599
transform 1 0 6624 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_3
timestamp -3599
transform 1 0 1380 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_32
timestamp 1636964856
transform 1 0 4048 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_44
timestamp 1636964856
transform 1 0 5152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_68
timestamp -3599
transform 1 0 7360 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_72
timestamp -3599
transform 1 0 7728 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp -3599
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_3
timestamp -3599
transform 1 0 1380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_16
timestamp -3599
transform 1 0 2576 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_27
timestamp -3599
transform 1 0 3588 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp -3599
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636964856
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_69
timestamp -3599
transform 1 0 7452 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_29
timestamp -3599
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_56
timestamp -3599
transform 1 0 6256 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_64
timestamp -3599
transform 1 0 6992 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_79
timestamp -3599
transform 1 0 8372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp -3599
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1636964856
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_19
timestamp -3599
transform 1 0 2852 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1636964856
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_40
timestamp -3599
transform 1 0 4784 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp -3599
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_74
timestamp -3599
transform 1 0 7912 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp -3599
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp -3599
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636964856
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp -3599
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_49
timestamp -3599
transform 1 0 5612 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_7
timestamp -3599
transform 1 0 1748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_12
timestamp -3599
transform 1 0 2208 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_35
timestamp 1636964856
transform 1 0 4324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp -3599
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp -3599
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636964856
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_69
timestamp -3599
transform 1 0 7452 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_93
timestamp -3599
transform 1 0 9660 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_18
timestamp -3599
transform 1 0 2760 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_24
timestamp -3599
transform 1 0 3312 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636964856
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp -3599
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_11
timestamp -3599
transform 1 0 2116 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_19
timestamp -3599
transform 1 0 2852 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_60
timestamp -3599
transform 1 0 6624 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp -3599
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_10
timestamp 1636964856
transform 1 0 2024 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_22
timestamp -3599
transform 1 0 3128 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_29
timestamp -3599
transform 1 0 3772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_37
timestamp -3599
transform 1 0 4508 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_78
timestamp -3599
transform 1 0 8280 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp -3599
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_10
timestamp -3599
transform 1 0 2024 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_36
timestamp 1636964856
transform 1 0 4416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_48
timestamp -3599
transform 1 0 5520 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_60
timestamp -3599
transform 1 0 6624 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_68
timestamp -3599
transform 1 0 7360 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_92
timestamp -3599
transform 1 0 9568 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_7
timestamp -3599
transform 1 0 1748 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_22
timestamp -3599
transform 1 0 3128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_49
timestamp -3599
transform 1 0 5612 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp -3599
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp -3599
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp -3599
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_19
timestamp 1636964856
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp -3599
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp -3599
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_65
timestamp -3599
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_10
timestamp -3599
transform 1 0 2024 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_17
timestamp -3599
transform 1 0 2668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp -3599
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp -3599
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_33
timestamp -3599
transform 1 0 4140 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_46
timestamp -3599
transform 1 0 5336 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp -3599
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp -3599
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_52
timestamp -3599
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_77
timestamp -3599
transform 1 0 8188 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_7
timestamp -3599
transform 1 0 1748 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp -3599
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp -3599
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp -3599
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_54
timestamp -3599
transform 1 0 6072 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_70
timestamp -3599
transform 1 0 7544 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_78
timestamp -3599
transform 1 0 8280 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_85
timestamp -3599
transform 1 0 8924 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_7
timestamp 1636964856
transform 1 0 1748 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_19
timestamp -3599
transform 1 0 2852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp -3599
transform 1 0 3588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_33
timestamp -3599
transform 1 0 4140 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_48
timestamp -3599
transform 1 0 5520 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp -3599
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_60
timestamp 1636964856
transform 1 0 6624 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_72
timestamp -3599
transform 1 0 7728 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_80
timestamp -3599
transform 1 0 8464 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_7
timestamp 1636964856
transform 1 0 1748 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_19
timestamp -3599
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp -3599
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_29
timestamp -3599
transform 1 0 3772 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_35
timestamp -3599
transform 1 0 4324 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_48
timestamp 1636964856
transform 1 0 5520 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_60
timestamp 1636964856
transform 1 0 6624 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_72
timestamp 1636964856
transform 1 0 7728 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp -3599
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636964856
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636964856
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636964856
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636964856
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp -3599
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp -3599
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_57
timestamp -3599
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_65
timestamp -3599
transform 1 0 7084 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_70
timestamp -3599
transform 1 0 7544 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_78
timestamp -3599
transform 1 0 8280 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_86
timestamp -3599
transform 1 0 9016 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_7
timestamp 1636964856
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp -3599
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp -3599
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636964856
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636964856
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_53
timestamp -3599
transform 1 0 5980 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_63
timestamp -3599
transform 1 0 6900 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_67
timestamp -3599
transform 1 0 7268 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_73
timestamp -3599
transform 1 0 7820 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_76
timestamp -3599
transform 1 0 8096 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_79
timestamp -3599
transform 1 0 8372 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_90
timestamp -3599
transform 1 0 9384 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_93
timestamp -3599
transform 1 0 9660 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_7
timestamp 1636964856
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_19
timestamp 1636964856
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_31
timestamp 1636964856
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_43
timestamp 1636964856
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp -3599
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_57
timestamp -3599
transform 1 0 6348 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_66
timestamp -3599
transform 1 0 7176 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_80
timestamp -3599
transform 1 0 8464 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_83
timestamp -3599
transform 1 0 8740 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_94
timestamp -3599
transform 1 0 9752 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_6
timestamp 1636964856
transform 1 0 1656 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_18
timestamp -3599
transform 1 0 2760 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp -3599
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636964856
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636964856
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_53
timestamp -3599
transform 1 0 5980 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_79
timestamp -3599
transform 1 0 8372 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_85
timestamp -3599
transform 1 0 8924 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_3
timestamp -3599
transform 1 0 1380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_8
timestamp -3599
transform 1 0 1840 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_13
timestamp -3599
transform 1 0 2300 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_18
timestamp -3599
transform 1 0 2760 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_23
timestamp -3599
transform 1 0 3220 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_33
timestamp -3599
transform 1 0 4140 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_38
timestamp -3599
transform 1 0 4600 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_43
timestamp -3599
transform 1 0 5060 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_57
timestamp -3599
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_63
timestamp -3599
transform 1 0 6900 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_74
timestamp -3599
transform 1 0 7912 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_82
timestamp -3599
transform 1 0 8648 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_93
timestamp -3599
transform 1 0 9660 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp -3599
transform 1 0 1380 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input4
timestamp -3599
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -3599
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -3599
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3599
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3599
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -3599
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -3599
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -3599
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp -3599
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp -3599
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp -3599
transform 1 0 1380 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -3599
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp -3599
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp -3599
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp -3599
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp -3599
transform 1 0 1380 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp -3599
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -3599
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -3599
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp -3599
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp -3599
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp -3599
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp -3599
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp -3599
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -3599
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -3599
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -3599
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform 1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp -3599
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp -3599
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -3599
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp -3599
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp -3599
transform -1 0 9844 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input37
timestamp -3599
transform -1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -3599
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp -3599
transform -1 0 9844 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp -3599
transform -1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input41
timestamp -3599
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp -3599
transform -1 0 9844 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input43
timestamp -3599
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp -3599
transform -1 0 8832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input45
timestamp -3599
transform -1 0 8464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp -3599
transform -1 0 9844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp -3599
transform -1 0 9844 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp -3599
transform -1 0 9844 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input49
timestamp -3599
transform -1 0 7452 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp -3599
transform -1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp -3599
transform -1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp -3599
transform -1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input53
timestamp -3599
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp -3599
transform -1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp -3599
transform -1 0 8832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp -3599
transform -1 0 8832 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp -3599
transform -1 0 9844 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input58
timestamp -3599
transform -1 0 8464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp -3599
transform -1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp -3599
transform -1 0 9844 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp -3599
transform -1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp -3599
transform -1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp -3599
transform -1 0 8832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp -3599
transform -1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp -3599
transform -1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp -3599
transform -1 0 9844 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input67
timestamp -3599
transform 1 0 6808 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp -3599
transform -1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp -3599
transform -1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp -3599
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp -3599
transform -1 0 9568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp -3599
transform -1 0 9844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp -3599
transform -1 0 7636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp -3599
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp -3599
transform -1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp -3599
transform -1 0 8832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp -3599
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp -3599
transform -1 0 9844 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input79
timestamp -3599
transform -1 0 8280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp -3599
transform -1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp -3599
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp -3599
transform -1 0 8004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp -3599
transform -1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform -1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 9476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 9108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 8740 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 9476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 9108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform 1 0 8372 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform 1 0 9108 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform 1 0 9476 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform 1 0 9108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform 1 0 9476 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform 1 0 9476 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform 1 0 9108 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform 1 0 9108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 9476 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform 1 0 9108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform 1 0 8096 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform 1 0 9108 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform -1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform 1 0 9476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform 1 0 9476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 8740 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform 1 0 9108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform 1 0 9476 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform 1 0 9476 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform 1 0 9108 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform 1 0 9108 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform 1 0 9476 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform 1 0 9476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform 1 0 9108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform 1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform 1 0 9108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform 1 0 9476 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform 1 0 9108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform 1 0 9476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform 1 0 9476 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform 1 0 9108 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform 1 0 9476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform 1 0 9108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform 1 0 9476 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform 1 0 9108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform 1 0 9476 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform 1 0 9108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform 1 0 9108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform 1 0 9476 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform 1 0 9108 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform 1 0 8740 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform 1 0 9108 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform 1 0 9476 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform 1 0 8740 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp -3599
transform 1 0 9476 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp -3599
transform 1 0 9108 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp -3599
transform 1 0 9476 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp -3599
transform 1 0 9476 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp -3599
transform 1 0 9108 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp -3599
transform 1 0 8832 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp -3599
transform 1 0 8740 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp -3599
transform 1 0 9108 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp -3599
transform 1 0 9476 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp -3599
transform 1 0 9108 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp -3599
transform 1 0 9476 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp -3599
transform 1 0 9292 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp -3599
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp -3599
transform -1 0 1840 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp -3599
transform -1 0 6256 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp -3599
transform 1 0 6532 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp -3599
transform -1 0 7544 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp -3599
transform -1 0 7912 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp -3599
transform -1 0 8648 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp -3599
transform -1 0 9292 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp -3599
transform 1 0 9292 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp -3599
transform -1 0 6992 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp -3599
transform -1 0 8096 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp -3599
transform 1 0 9108 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp -3599
transform 1 0 1932 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp -3599
transform 1 0 2392 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp -3599
transform -1 0 3220 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp -3599
transform -1 0 3680 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp -3599
transform -1 0 4140 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp -3599
transform -1 0 4600 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp -3599
transform -1 0 5060 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp -3599
transform -1 0 5520 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp -3599
transform -1 0 5888 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output196
timestamp -3599
transform -1 0 1656 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_74
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_75
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_76
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_77
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_78
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_79
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_80
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_81
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_82
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_83
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_84
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_85
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_86
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_87
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_88
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_89
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_90
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 10120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_91
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_92
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 10120 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_93
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_94
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 10120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_95
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 10120 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_96
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 10120 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_97
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 10120 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_98
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 10120 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_99
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 10120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_100
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_101
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_102
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 10120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_103
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_104
timestamp -3599
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3599
transform -1 0 10120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_105
timestamp -3599
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3599
transform -1 0 10120 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_106
timestamp -3599
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3599
transform -1 0 10120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_107
timestamp -3599
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -3599
transform -1 0 10120 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_108
timestamp -3599
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -3599
transform -1 0 10120 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_109
timestamp -3599
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -3599
transform -1 0 10120 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_110
timestamp -3599
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -3599
transform -1 0 10120 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_111
timestamp -3599
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -3599
transform -1 0 10120 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_112
timestamp -3599
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -3599
transform -1 0 10120 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_113
timestamp -3599
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -3599
transform -1 0 10120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_114
timestamp -3599
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -3599
transform -1 0 10120 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_115
timestamp -3599
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -3599
transform -1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_116
timestamp -3599
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -3599
transform -1 0 10120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_117
timestamp -3599
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -3599
transform -1 0 10120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_118
timestamp -3599
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -3599
transform -1 0 10120 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_119
timestamp -3599
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -3599
transform -1 0 10120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_120
timestamp -3599
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -3599
transform -1 0 10120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_121
timestamp -3599
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp -3599
transform -1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_122
timestamp -3599
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp -3599
transform -1 0 10120 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_123
timestamp -3599
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp -3599
transform -1 0 10120 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_124
timestamp -3599
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp -3599
transform -1 0 10120 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_125
timestamp -3599
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp -3599
transform -1 0 10120 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_126
timestamp -3599
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp -3599
transform -1 0 10120 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_127
timestamp -3599
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp -3599
transform -1 0 10120 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_128
timestamp -3599
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp -3599
transform -1 0 10120 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_129
timestamp -3599
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp -3599
transform -1 0 10120 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_130
timestamp -3599
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp -3599
transform -1 0 10120 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_131
timestamp -3599
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp -3599
transform -1 0 10120 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_132
timestamp -3599
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp -3599
transform -1 0 10120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_133
timestamp -3599
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp -3599
transform -1 0 10120 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_134
timestamp -3599
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp -3599
transform -1 0 10120 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_135
timestamp -3599
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp -3599
transform -1 0 10120 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_136
timestamp -3599
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp -3599
transform -1 0 10120 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_137
timestamp -3599
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp -3599
transform -1 0 10120 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_138
timestamp -3599
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp -3599
transform -1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_139
timestamp -3599
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp -3599
transform -1 0 10120 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_140
timestamp -3599
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp -3599
transform -1 0 10120 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_141
timestamp -3599
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp -3599
transform -1 0 10120 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_142
timestamp -3599
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp -3599
transform -1 0 10120 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_143
timestamp -3599
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp -3599
transform -1 0 10120 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_144
timestamp -3599
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp -3599
transform -1 0 10120 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_145
timestamp -3599
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp -3599
transform -1 0 10120 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_146
timestamp -3599
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp -3599
transform -1 0 10120 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_147
timestamp -3599
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp -3599
transform -1 0 10120 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_150
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_151
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_154
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_155
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_156
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_157
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_158
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_159
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_160
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_161
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_162
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_163
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_164
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_165
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_166
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_167
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_168
timestamp -3599
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_169
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_170
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_171
timestamp -3599
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_172
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp -3599
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_175
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp -3599
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp -3599
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_179
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_180
timestamp -3599
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_181
timestamp -3599
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_182
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_183
timestamp -3599
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_184
timestamp -3599
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp -3599
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_187
timestamp -3599
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_188
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_189
timestamp -3599
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_190
timestamp -3599
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_191
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_192
timestamp -3599
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_193
timestamp -3599
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_194
timestamp -3599
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_195
timestamp -3599
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_196
timestamp -3599
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_197
timestamp -3599
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_198
timestamp -3599
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_199
timestamp -3599
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_200
timestamp -3599
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_201
timestamp -3599
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_202
timestamp -3599
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_203
timestamp -3599
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_204
timestamp -3599
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_205
timestamp -3599
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_206
timestamp -3599
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_207
timestamp -3599
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_208
timestamp -3599
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_209
timestamp -3599
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_210
timestamp -3599
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_211
timestamp -3599
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_212
timestamp -3599
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_213
timestamp -3599
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_214
timestamp -3599
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_215
timestamp -3599
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_216
timestamp -3599
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_217
timestamp -3599
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_218
timestamp -3599
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_219
timestamp -3599
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_220
timestamp -3599
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_221
timestamp -3599
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_222
timestamp -3599
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_223
timestamp -3599
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_224
timestamp -3599
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_225
timestamp -3599
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_226
timestamp -3599
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_227
timestamp -3599
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_228
timestamp -3599
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_229
timestamp -3599
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_230
timestamp -3599
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_231
timestamp -3599
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_232
timestamp -3599
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_233
timestamp -3599
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_234
timestamp -3599
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_235
timestamp -3599
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_236
timestamp -3599
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_237
timestamp -3599
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_238
timestamp -3599
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_239
timestamp -3599
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_240
timestamp -3599
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_241
timestamp -3599
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_242
timestamp -3599
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_243
timestamp -3599
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_244
timestamp -3599
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_245
timestamp -3599
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_246
timestamp -3599
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_247
timestamp -3599
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_248
timestamp -3599
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_249
timestamp -3599
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_250
timestamp -3599
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_251
timestamp -3599
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_252
timestamp -3599
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_253
timestamp -3599
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_254
timestamp -3599
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_255
timestamp -3599
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_256
timestamp -3599
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_257
timestamp -3599
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_258
timestamp -3599
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_259
timestamp -3599
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_260
timestamp -3599
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_261
timestamp -3599
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 A_I_top
port 0 nsew signal output
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 A_T_top
port 2 nsew signal output
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal3 s 0 10616 120 10736 0 FreeSans 480 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal3 s 0 11432 120 11552 0 FreeSans 480 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 B_I_top
port 7 nsew signal output
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 B_T_top
port 9 nsew signal output
flabel metal3 s 0 12248 120 12368 0 FreeSans 480 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal3 s 0 13064 120 13184 0 FreeSans 480 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal3 s 0 13880 120 14000 0 FreeSans 480 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal3 s 0 14696 120 14816 0 FreeSans 480 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal3 s 11130 18232 11250 18352 0 FreeSans 480 0 0 0 E1BEG[0]
port 14 nsew signal output
flabel metal3 s 11130 18504 11250 18624 0 FreeSans 480 0 0 0 E1BEG[1]
port 15 nsew signal output
flabel metal3 s 11130 18776 11250 18896 0 FreeSans 480 0 0 0 E1BEG[2]
port 16 nsew signal output
flabel metal3 s 11130 19048 11250 19168 0 FreeSans 480 0 0 0 E1BEG[3]
port 17 nsew signal output
flabel metal3 s 11130 19320 11250 19440 0 FreeSans 480 0 0 0 E2BEG[0]
port 18 nsew signal output
flabel metal3 s 11130 19592 11250 19712 0 FreeSans 480 0 0 0 E2BEG[1]
port 19 nsew signal output
flabel metal3 s 11130 19864 11250 19984 0 FreeSans 480 0 0 0 E2BEG[2]
port 20 nsew signal output
flabel metal3 s 11130 20136 11250 20256 0 FreeSans 480 0 0 0 E2BEG[3]
port 21 nsew signal output
flabel metal3 s 11130 20408 11250 20528 0 FreeSans 480 0 0 0 E2BEG[4]
port 22 nsew signal output
flabel metal3 s 11130 20680 11250 20800 0 FreeSans 480 0 0 0 E2BEG[5]
port 23 nsew signal output
flabel metal3 s 11130 20952 11250 21072 0 FreeSans 480 0 0 0 E2BEG[6]
port 24 nsew signal output
flabel metal3 s 11130 21224 11250 21344 0 FreeSans 480 0 0 0 E2BEG[7]
port 25 nsew signal output
flabel metal3 s 11130 21496 11250 21616 0 FreeSans 480 0 0 0 E2BEGb[0]
port 26 nsew signal output
flabel metal3 s 11130 21768 11250 21888 0 FreeSans 480 0 0 0 E2BEGb[1]
port 27 nsew signal output
flabel metal3 s 11130 22040 11250 22160 0 FreeSans 480 0 0 0 E2BEGb[2]
port 28 nsew signal output
flabel metal3 s 11130 22312 11250 22432 0 FreeSans 480 0 0 0 E2BEGb[3]
port 29 nsew signal output
flabel metal3 s 11130 22584 11250 22704 0 FreeSans 480 0 0 0 E2BEGb[4]
port 30 nsew signal output
flabel metal3 s 11130 22856 11250 22976 0 FreeSans 480 0 0 0 E2BEGb[5]
port 31 nsew signal output
flabel metal3 s 11130 23128 11250 23248 0 FreeSans 480 0 0 0 E2BEGb[6]
port 32 nsew signal output
flabel metal3 s 11130 23400 11250 23520 0 FreeSans 480 0 0 0 E2BEGb[7]
port 33 nsew signal output
flabel metal3 s 11130 28024 11250 28144 0 FreeSans 480 0 0 0 E6BEG[0]
port 34 nsew signal output
flabel metal3 s 11130 30744 11250 30864 0 FreeSans 480 0 0 0 E6BEG[10]
port 35 nsew signal output
flabel metal3 s 11130 31016 11250 31136 0 FreeSans 480 0 0 0 E6BEG[11]
port 36 nsew signal output
flabel metal3 s 11130 28296 11250 28416 0 FreeSans 480 0 0 0 E6BEG[1]
port 37 nsew signal output
flabel metal3 s 11130 28568 11250 28688 0 FreeSans 480 0 0 0 E6BEG[2]
port 38 nsew signal output
flabel metal3 s 11130 28840 11250 28960 0 FreeSans 480 0 0 0 E6BEG[3]
port 39 nsew signal output
flabel metal3 s 11130 29112 11250 29232 0 FreeSans 480 0 0 0 E6BEG[4]
port 40 nsew signal output
flabel metal3 s 11130 29384 11250 29504 0 FreeSans 480 0 0 0 E6BEG[5]
port 41 nsew signal output
flabel metal3 s 11130 29656 11250 29776 0 FreeSans 480 0 0 0 E6BEG[6]
port 42 nsew signal output
flabel metal3 s 11130 29928 11250 30048 0 FreeSans 480 0 0 0 E6BEG[7]
port 43 nsew signal output
flabel metal3 s 11130 30200 11250 30320 0 FreeSans 480 0 0 0 E6BEG[8]
port 44 nsew signal output
flabel metal3 s 11130 30472 11250 30592 0 FreeSans 480 0 0 0 E6BEG[9]
port 45 nsew signal output
flabel metal3 s 11130 23672 11250 23792 0 FreeSans 480 0 0 0 EE4BEG[0]
port 46 nsew signal output
flabel metal3 s 11130 26392 11250 26512 0 FreeSans 480 0 0 0 EE4BEG[10]
port 47 nsew signal output
flabel metal3 s 11130 26664 11250 26784 0 FreeSans 480 0 0 0 EE4BEG[11]
port 48 nsew signal output
flabel metal3 s 11130 26936 11250 27056 0 FreeSans 480 0 0 0 EE4BEG[12]
port 49 nsew signal output
flabel metal3 s 11130 27208 11250 27328 0 FreeSans 480 0 0 0 EE4BEG[13]
port 50 nsew signal output
flabel metal3 s 11130 27480 11250 27600 0 FreeSans 480 0 0 0 EE4BEG[14]
port 51 nsew signal output
flabel metal3 s 11130 27752 11250 27872 0 FreeSans 480 0 0 0 EE4BEG[15]
port 52 nsew signal output
flabel metal3 s 11130 23944 11250 24064 0 FreeSans 480 0 0 0 EE4BEG[1]
port 53 nsew signal output
flabel metal3 s 11130 24216 11250 24336 0 FreeSans 480 0 0 0 EE4BEG[2]
port 54 nsew signal output
flabel metal3 s 11130 24488 11250 24608 0 FreeSans 480 0 0 0 EE4BEG[3]
port 55 nsew signal output
flabel metal3 s 11130 24760 11250 24880 0 FreeSans 480 0 0 0 EE4BEG[4]
port 56 nsew signal output
flabel metal3 s 11130 25032 11250 25152 0 FreeSans 480 0 0 0 EE4BEG[5]
port 57 nsew signal output
flabel metal3 s 11130 25304 11250 25424 0 FreeSans 480 0 0 0 EE4BEG[6]
port 58 nsew signal output
flabel metal3 s 11130 25576 11250 25696 0 FreeSans 480 0 0 0 EE4BEG[7]
port 59 nsew signal output
flabel metal3 s 11130 25848 11250 25968 0 FreeSans 480 0 0 0 EE4BEG[8]
port 60 nsew signal output
flabel metal3 s 11130 26120 11250 26240 0 FreeSans 480 0 0 0 EE4BEG[9]
port 61 nsew signal output
flabel metal3 s 0 15512 120 15632 0 FreeSans 480 0 0 0 FrameData[0]
port 62 nsew signal input
flabel metal3 s 0 23672 120 23792 0 FreeSans 480 0 0 0 FrameData[10]
port 63 nsew signal input
flabel metal3 s 0 24488 120 24608 0 FreeSans 480 0 0 0 FrameData[11]
port 64 nsew signal input
flabel metal3 s 0 25304 120 25424 0 FreeSans 480 0 0 0 FrameData[12]
port 65 nsew signal input
flabel metal3 s 0 26120 120 26240 0 FreeSans 480 0 0 0 FrameData[13]
port 66 nsew signal input
flabel metal3 s 0 26936 120 27056 0 FreeSans 480 0 0 0 FrameData[14]
port 67 nsew signal input
flabel metal3 s 0 27752 120 27872 0 FreeSans 480 0 0 0 FrameData[15]
port 68 nsew signal input
flabel metal3 s 0 28568 120 28688 0 FreeSans 480 0 0 0 FrameData[16]
port 69 nsew signal input
flabel metal3 s 0 29384 120 29504 0 FreeSans 480 0 0 0 FrameData[17]
port 70 nsew signal input
flabel metal3 s 0 30200 120 30320 0 FreeSans 480 0 0 0 FrameData[18]
port 71 nsew signal input
flabel metal3 s 0 31016 120 31136 0 FreeSans 480 0 0 0 FrameData[19]
port 72 nsew signal input
flabel metal3 s 0 16328 120 16448 0 FreeSans 480 0 0 0 FrameData[1]
port 73 nsew signal input
flabel metal3 s 0 31832 120 31952 0 FreeSans 480 0 0 0 FrameData[20]
port 74 nsew signal input
flabel metal3 s 0 32648 120 32768 0 FreeSans 480 0 0 0 FrameData[21]
port 75 nsew signal input
flabel metal3 s 0 33464 120 33584 0 FreeSans 480 0 0 0 FrameData[22]
port 76 nsew signal input
flabel metal3 s 0 34280 120 34400 0 FreeSans 480 0 0 0 FrameData[23]
port 77 nsew signal input
flabel metal3 s 0 35096 120 35216 0 FreeSans 480 0 0 0 FrameData[24]
port 78 nsew signal input
flabel metal3 s 0 35912 120 36032 0 FreeSans 480 0 0 0 FrameData[25]
port 79 nsew signal input
flabel metal3 s 0 36728 120 36848 0 FreeSans 480 0 0 0 FrameData[26]
port 80 nsew signal input
flabel metal3 s 0 37544 120 37664 0 FreeSans 480 0 0 0 FrameData[27]
port 81 nsew signal input
flabel metal3 s 0 38360 120 38480 0 FreeSans 480 0 0 0 FrameData[28]
port 82 nsew signal input
flabel metal3 s 0 39176 120 39296 0 FreeSans 480 0 0 0 FrameData[29]
port 83 nsew signal input
flabel metal3 s 0 17144 120 17264 0 FreeSans 480 0 0 0 FrameData[2]
port 84 nsew signal input
flabel metal3 s 0 39992 120 40112 0 FreeSans 480 0 0 0 FrameData[30]
port 85 nsew signal input
flabel metal3 s 0 40808 120 40928 0 FreeSans 480 0 0 0 FrameData[31]
port 86 nsew signal input
flabel metal3 s 0 17960 120 18080 0 FreeSans 480 0 0 0 FrameData[3]
port 87 nsew signal input
flabel metal3 s 0 18776 120 18896 0 FreeSans 480 0 0 0 FrameData[4]
port 88 nsew signal input
flabel metal3 s 0 19592 120 19712 0 FreeSans 480 0 0 0 FrameData[5]
port 89 nsew signal input
flabel metal3 s 0 20408 120 20528 0 FreeSans 480 0 0 0 FrameData[6]
port 90 nsew signal input
flabel metal3 s 0 21224 120 21344 0 FreeSans 480 0 0 0 FrameData[7]
port 91 nsew signal input
flabel metal3 s 0 22040 120 22160 0 FreeSans 480 0 0 0 FrameData[8]
port 92 nsew signal input
flabel metal3 s 0 22856 120 22976 0 FreeSans 480 0 0 0 FrameData[9]
port 93 nsew signal input
flabel metal3 s 11130 31288 11250 31408 0 FreeSans 480 0 0 0 FrameData_O[0]
port 94 nsew signal output
flabel metal3 s 11130 34008 11250 34128 0 FreeSans 480 0 0 0 FrameData_O[10]
port 95 nsew signal output
flabel metal3 s 11130 34280 11250 34400 0 FreeSans 480 0 0 0 FrameData_O[11]
port 96 nsew signal output
flabel metal3 s 11130 34552 11250 34672 0 FreeSans 480 0 0 0 FrameData_O[12]
port 97 nsew signal output
flabel metal3 s 11130 34824 11250 34944 0 FreeSans 480 0 0 0 FrameData_O[13]
port 98 nsew signal output
flabel metal3 s 11130 35096 11250 35216 0 FreeSans 480 0 0 0 FrameData_O[14]
port 99 nsew signal output
flabel metal3 s 11130 35368 11250 35488 0 FreeSans 480 0 0 0 FrameData_O[15]
port 100 nsew signal output
flabel metal3 s 11130 35640 11250 35760 0 FreeSans 480 0 0 0 FrameData_O[16]
port 101 nsew signal output
flabel metal3 s 11130 35912 11250 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 102 nsew signal output
flabel metal3 s 11130 36184 11250 36304 0 FreeSans 480 0 0 0 FrameData_O[18]
port 103 nsew signal output
flabel metal3 s 11130 36456 11250 36576 0 FreeSans 480 0 0 0 FrameData_O[19]
port 104 nsew signal output
flabel metal3 s 11130 31560 11250 31680 0 FreeSans 480 0 0 0 FrameData_O[1]
port 105 nsew signal output
flabel metal3 s 11130 36728 11250 36848 0 FreeSans 480 0 0 0 FrameData_O[20]
port 106 nsew signal output
flabel metal3 s 11130 37000 11250 37120 0 FreeSans 480 0 0 0 FrameData_O[21]
port 107 nsew signal output
flabel metal3 s 11130 37272 11250 37392 0 FreeSans 480 0 0 0 FrameData_O[22]
port 108 nsew signal output
flabel metal3 s 11130 37544 11250 37664 0 FreeSans 480 0 0 0 FrameData_O[23]
port 109 nsew signal output
flabel metal3 s 11130 37816 11250 37936 0 FreeSans 480 0 0 0 FrameData_O[24]
port 110 nsew signal output
flabel metal3 s 11130 38088 11250 38208 0 FreeSans 480 0 0 0 FrameData_O[25]
port 111 nsew signal output
flabel metal3 s 11130 38360 11250 38480 0 FreeSans 480 0 0 0 FrameData_O[26]
port 112 nsew signal output
flabel metal3 s 11130 38632 11250 38752 0 FreeSans 480 0 0 0 FrameData_O[27]
port 113 nsew signal output
flabel metal3 s 11130 38904 11250 39024 0 FreeSans 480 0 0 0 FrameData_O[28]
port 114 nsew signal output
flabel metal3 s 11130 39176 11250 39296 0 FreeSans 480 0 0 0 FrameData_O[29]
port 115 nsew signal output
flabel metal3 s 11130 31832 11250 31952 0 FreeSans 480 0 0 0 FrameData_O[2]
port 116 nsew signal output
flabel metal3 s 11130 39448 11250 39568 0 FreeSans 480 0 0 0 FrameData_O[30]
port 117 nsew signal output
flabel metal3 s 11130 39720 11250 39840 0 FreeSans 480 0 0 0 FrameData_O[31]
port 118 nsew signal output
flabel metal3 s 11130 32104 11250 32224 0 FreeSans 480 0 0 0 FrameData_O[3]
port 119 nsew signal output
flabel metal3 s 11130 32376 11250 32496 0 FreeSans 480 0 0 0 FrameData_O[4]
port 120 nsew signal output
flabel metal3 s 11130 32648 11250 32768 0 FreeSans 480 0 0 0 FrameData_O[5]
port 121 nsew signal output
flabel metal3 s 11130 32920 11250 33040 0 FreeSans 480 0 0 0 FrameData_O[6]
port 122 nsew signal output
flabel metal3 s 11130 33192 11250 33312 0 FreeSans 480 0 0 0 FrameData_O[7]
port 123 nsew signal output
flabel metal3 s 11130 33464 11250 33584 0 FreeSans 480 0 0 0 FrameData_O[8]
port 124 nsew signal output
flabel metal3 s 11130 33736 11250 33856 0 FreeSans 480 0 0 0 FrameData_O[9]
port 125 nsew signal output
flabel metal2 s 1398 0 1454 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 126 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 127 nsew signal input
flabel metal2 s 6458 0 6514 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 128 nsew signal input
flabel metal2 s 6918 0 6974 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 129 nsew signal input
flabel metal2 s 7378 0 7434 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 130 nsew signal input
flabel metal2 s 7838 0 7894 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 131 nsew signal input
flabel metal2 s 8298 0 8354 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 132 nsew signal input
flabel metal2 s 8758 0 8814 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 133 nsew signal input
flabel metal2 s 9218 0 9274 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 134 nsew signal input
flabel metal2 s 9678 0 9734 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 135 nsew signal input
flabel metal2 s 10138 0 10194 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 136 nsew signal input
flabel metal2 s 1858 0 1914 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 137 nsew signal input
flabel metal2 s 2318 0 2374 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 138 nsew signal input
flabel metal2 s 2778 0 2834 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 139 nsew signal input
flabel metal2 s 3238 0 3294 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 140 nsew signal input
flabel metal2 s 3698 0 3754 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 141 nsew signal input
flabel metal2 s 4158 0 4214 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 142 nsew signal input
flabel metal2 s 4618 0 4674 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 143 nsew signal input
flabel metal2 s 5078 0 5134 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 144 nsew signal input
flabel metal2 s 5538 0 5594 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 145 nsew signal input
flabel metal2 s 1398 44944 1454 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 146 nsew signal output
flabel metal2 s 5998 44944 6054 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 147 nsew signal output
flabel metal2 s 6458 44944 6514 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 148 nsew signal output
flabel metal2 s 6918 44944 6974 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 149 nsew signal output
flabel metal2 s 7378 44944 7434 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 150 nsew signal output
flabel metal2 s 7838 44944 7894 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 151 nsew signal output
flabel metal2 s 8298 44944 8354 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 152 nsew signal output
flabel metal2 s 8758 44944 8814 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 153 nsew signal output
flabel metal2 s 9218 44944 9274 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 154 nsew signal output
flabel metal2 s 9678 44944 9734 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 155 nsew signal output
flabel metal2 s 10138 44944 10194 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 156 nsew signal output
flabel metal2 s 1858 44944 1914 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 157 nsew signal output
flabel metal2 s 2318 44944 2374 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 158 nsew signal output
flabel metal2 s 2778 44944 2834 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 159 nsew signal output
flabel metal2 s 3238 44944 3294 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 160 nsew signal output
flabel metal2 s 3698 44944 3754 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 161 nsew signal output
flabel metal2 s 4158 44944 4214 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 162 nsew signal output
flabel metal2 s 4618 44944 4674 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 163 nsew signal output
flabel metal2 s 5078 44944 5134 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 164 nsew signal output
flabel metal2 s 5538 44944 5594 45000 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 165 nsew signal output
flabel metal2 s 938 0 994 56 0 FreeSans 224 0 0 0 UserCLK
port 166 nsew signal input
flabel metal2 s 938 44944 994 45000 0 FreeSans 224 0 0 0 UserCLKo
port 167 nsew signal output
flabel metal4 s 3004 0 3324 45000 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 3004 44940 3324 45000 0 FreeSans 480 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 9004 0 9324 45000 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 9004 44940 9324 45000 0 FreeSans 480 0 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 1944 0 2264 45000 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 1944 44940 2264 45000 0 FreeSans 480 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 7944 0 8264 45000 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 7944 44940 8264 45000 0 FreeSans 480 0 0 0 VPWR
port 169 nsew power bidirectional
flabel metal3 s 11130 5176 11250 5296 0 FreeSans 480 0 0 0 W1END[0]
port 170 nsew signal input
flabel metal3 s 11130 5448 11250 5568 0 FreeSans 480 0 0 0 W1END[1]
port 171 nsew signal input
flabel metal3 s 11130 5720 11250 5840 0 FreeSans 480 0 0 0 W1END[2]
port 172 nsew signal input
flabel metal3 s 11130 5992 11250 6112 0 FreeSans 480 0 0 0 W1END[3]
port 173 nsew signal input
flabel metal3 s 11130 8440 11250 8560 0 FreeSans 480 0 0 0 W2END[0]
port 174 nsew signal input
flabel metal3 s 11130 8712 11250 8832 0 FreeSans 480 0 0 0 W2END[1]
port 175 nsew signal input
flabel metal3 s 11130 8984 11250 9104 0 FreeSans 480 0 0 0 W2END[2]
port 176 nsew signal input
flabel metal3 s 11130 9256 11250 9376 0 FreeSans 480 0 0 0 W2END[3]
port 177 nsew signal input
flabel metal3 s 11130 9528 11250 9648 0 FreeSans 480 0 0 0 W2END[4]
port 178 nsew signal input
flabel metal3 s 11130 9800 11250 9920 0 FreeSans 480 0 0 0 W2END[5]
port 179 nsew signal input
flabel metal3 s 11130 10072 11250 10192 0 FreeSans 480 0 0 0 W2END[6]
port 180 nsew signal input
flabel metal3 s 11130 10344 11250 10464 0 FreeSans 480 0 0 0 W2END[7]
port 181 nsew signal input
flabel metal3 s 11130 6264 11250 6384 0 FreeSans 480 0 0 0 W2MID[0]
port 182 nsew signal input
flabel metal3 s 11130 6536 11250 6656 0 FreeSans 480 0 0 0 W2MID[1]
port 183 nsew signal input
flabel metal3 s 11130 6808 11250 6928 0 FreeSans 480 0 0 0 W2MID[2]
port 184 nsew signal input
flabel metal3 s 11130 7080 11250 7200 0 FreeSans 480 0 0 0 W2MID[3]
port 185 nsew signal input
flabel metal3 s 11130 7352 11250 7472 0 FreeSans 480 0 0 0 W2MID[4]
port 186 nsew signal input
flabel metal3 s 11130 7624 11250 7744 0 FreeSans 480 0 0 0 W2MID[5]
port 187 nsew signal input
flabel metal3 s 11130 7896 11250 8016 0 FreeSans 480 0 0 0 W2MID[6]
port 188 nsew signal input
flabel metal3 s 11130 8168 11250 8288 0 FreeSans 480 0 0 0 W2MID[7]
port 189 nsew signal input
flabel metal3 s 11130 14968 11250 15088 0 FreeSans 480 0 0 0 W6END[0]
port 190 nsew signal input
flabel metal3 s 11130 17688 11250 17808 0 FreeSans 480 0 0 0 W6END[10]
port 191 nsew signal input
flabel metal3 s 11130 17960 11250 18080 0 FreeSans 480 0 0 0 W6END[11]
port 192 nsew signal input
flabel metal3 s 11130 15240 11250 15360 0 FreeSans 480 0 0 0 W6END[1]
port 193 nsew signal input
flabel metal3 s 11130 15512 11250 15632 0 FreeSans 480 0 0 0 W6END[2]
port 194 nsew signal input
flabel metal3 s 11130 15784 11250 15904 0 FreeSans 480 0 0 0 W6END[3]
port 195 nsew signal input
flabel metal3 s 11130 16056 11250 16176 0 FreeSans 480 0 0 0 W6END[4]
port 196 nsew signal input
flabel metal3 s 11130 16328 11250 16448 0 FreeSans 480 0 0 0 W6END[5]
port 197 nsew signal input
flabel metal3 s 11130 16600 11250 16720 0 FreeSans 480 0 0 0 W6END[6]
port 198 nsew signal input
flabel metal3 s 11130 16872 11250 16992 0 FreeSans 480 0 0 0 W6END[7]
port 199 nsew signal input
flabel metal3 s 11130 17144 11250 17264 0 FreeSans 480 0 0 0 W6END[8]
port 200 nsew signal input
flabel metal3 s 11130 17416 11250 17536 0 FreeSans 480 0 0 0 W6END[9]
port 201 nsew signal input
flabel metal3 s 11130 10616 11250 10736 0 FreeSans 480 0 0 0 WW4END[0]
port 202 nsew signal input
flabel metal3 s 11130 13336 11250 13456 0 FreeSans 480 0 0 0 WW4END[10]
port 203 nsew signal input
flabel metal3 s 11130 13608 11250 13728 0 FreeSans 480 0 0 0 WW4END[11]
port 204 nsew signal input
flabel metal3 s 11130 13880 11250 14000 0 FreeSans 480 0 0 0 WW4END[12]
port 205 nsew signal input
flabel metal3 s 11130 14152 11250 14272 0 FreeSans 480 0 0 0 WW4END[13]
port 206 nsew signal input
flabel metal3 s 11130 14424 11250 14544 0 FreeSans 480 0 0 0 WW4END[14]
port 207 nsew signal input
flabel metal3 s 11130 14696 11250 14816 0 FreeSans 480 0 0 0 WW4END[15]
port 208 nsew signal input
flabel metal3 s 11130 10888 11250 11008 0 FreeSans 480 0 0 0 WW4END[1]
port 209 nsew signal input
flabel metal3 s 11130 11160 11250 11280 0 FreeSans 480 0 0 0 WW4END[2]
port 210 nsew signal input
flabel metal3 s 11130 11432 11250 11552 0 FreeSans 480 0 0 0 WW4END[3]
port 211 nsew signal input
flabel metal3 s 11130 11704 11250 11824 0 FreeSans 480 0 0 0 WW4END[4]
port 212 nsew signal input
flabel metal3 s 11130 11976 11250 12096 0 FreeSans 480 0 0 0 WW4END[5]
port 213 nsew signal input
flabel metal3 s 11130 12248 11250 12368 0 FreeSans 480 0 0 0 WW4END[6]
port 214 nsew signal input
flabel metal3 s 11130 12520 11250 12640 0 FreeSans 480 0 0 0 WW4END[7]
port 215 nsew signal input
flabel metal3 s 11130 12792 11250 12912 0 FreeSans 480 0 0 0 WW4END[8]
port 216 nsew signal input
flabel metal3 s 11130 13064 11250 13184 0 FreeSans 480 0 0 0 WW4END[9]
port 217 nsew signal input
rlabel metal1 5612 42432 5612 42432 0 VGND
rlabel metal1 5612 41888 5612 41888 0 VPWR
rlabel metal3 804 4964 804 4964 0 A_I_top
rlabel metal3 804 4148 804 4148 0 A_O_top
rlabel metal3 988 5780 988 5780 0 A_T_top
rlabel metal3 804 9044 804 9044 0 A_config_C_bit0
rlabel metal3 804 9860 804 9860 0 A_config_C_bit1
rlabel metal3 482 10676 482 10676 0 A_config_C_bit2
rlabel metal3 804 11492 804 11492 0 A_config_C_bit3
rlabel metal3 804 7412 804 7412 0 B_I_top
rlabel metal3 758 6596 758 6596 0 B_O_top
rlabel metal3 482 8228 482 8228 0 B_T_top
rlabel metal3 574 12308 574 12308 0 B_config_C_bit0
rlabel metal3 804 13124 804 13124 0 B_config_C_bit1
rlabel metal3 804 13940 804 13940 0 B_config_C_bit2
rlabel metal3 804 14756 804 14756 0 B_config_C_bit3
rlabel metal3 10571 18292 10571 18292 0 E1BEG[0]
rlabel metal2 9706 18479 9706 18479 0 E1BEG[1]
rlabel metal3 10709 18836 10709 18836 0 E1BEG[2]
rlabel metal2 9706 19023 9706 19023 0 E1BEG[3]
rlabel metal3 10433 19380 10433 19380 0 E2BEG[0]
rlabel metal3 10709 19652 10709 19652 0 E2BEG[1]
rlabel metal3 10617 19924 10617 19924 0 E2BEG[2]
rlabel metal2 9706 20111 9706 20111 0 E2BEG[3]
rlabel metal3 10709 20468 10709 20468 0 E2BEG[4]
rlabel metal2 9706 20655 9706 20655 0 E2BEG[5]
rlabel metal3 10709 21012 10709 21012 0 E2BEG[6]
rlabel metal2 9706 21199 9706 21199 0 E2BEG[7]
rlabel metal2 9890 21743 9890 21743 0 E2BEGb[0]
rlabel metal2 9706 21743 9706 21743 0 E2BEGb[1]
rlabel metal3 10525 22100 10525 22100 0 E2BEGb[2]
rlabel metal1 9476 21862 9476 21862 0 E2BEGb[3]
rlabel metal1 9752 21862 9752 21862 0 E2BEGb[4]
rlabel metal3 10709 22916 10709 22916 0 E2BEGb[5]
rlabel metal3 10433 23188 10433 23188 0 E2BEGb[6]
rlabel metal3 10709 23460 10709 23460 0 E2BEGb[7]
rlabel metal3 10433 28084 10433 28084 0 E6BEG[0]
rlabel metal1 9660 31926 9660 31926 0 E6BEG[10]
rlabel metal1 9430 31926 9430 31926 0 E6BEG[11]
rlabel metal3 10387 28356 10387 28356 0 E6BEG[1]
rlabel metal3 10893 28628 10893 28628 0 E6BEG[2]
rlabel metal3 10755 28900 10755 28900 0 E6BEG[3]
rlabel metal3 10571 29172 10571 29172 0 E6BEG[4]
rlabel metal3 10479 29444 10479 29444 0 E6BEG[5]
rlabel metal3 10387 29716 10387 29716 0 E6BEG[6]
rlabel metal3 10709 29988 10709 29988 0 E6BEG[7]
rlabel metal3 10571 30260 10571 30260 0 E6BEG[8]
rlabel metal3 10433 30532 10433 30532 0 E6BEG[9]
rlabel metal3 10433 23732 10433 23732 0 EE4BEG[0]
rlabel metal3 10985 26452 10985 26452 0 EE4BEG[10]
rlabel metal3 10249 26724 10249 26724 0 EE4BEG[11]
rlabel metal3 10709 26996 10709 26996 0 EE4BEG[12]
rlabel metal3 10433 27268 10433 27268 0 EE4BEG[13]
rlabel metal3 10801 27540 10801 27540 0 EE4BEG[14]
rlabel metal3 10709 27812 10709 27812 0 EE4BEG[15]
rlabel metal3 10709 24004 10709 24004 0 EE4BEG[1]
rlabel metal3 10433 24276 10433 24276 0 EE4BEG[2]
rlabel metal1 9752 24378 9752 24378 0 EE4BEG[3]
rlabel metal3 10709 24820 10709 24820 0 EE4BEG[4]
rlabel metal3 10433 25092 10433 25092 0 EE4BEG[5]
rlabel metal3 10387 25364 10387 25364 0 EE4BEG[6]
rlabel metal3 10709 25636 10709 25636 0 EE4BEG[7]
rlabel metal3 10433 25908 10433 25908 0 EE4BEG[8]
rlabel metal3 10755 26180 10755 26180 0 EE4BEG[9]
rlabel metal3 666 15572 666 15572 0 FrameData[0]
rlabel metal3 758 23732 758 23732 0 FrameData[10]
rlabel metal3 758 24548 758 24548 0 FrameData[11]
rlabel metal3 758 25364 758 25364 0 FrameData[12]
rlabel metal3 390 26180 390 26180 0 FrameData[13]
rlabel metal3 758 26996 758 26996 0 FrameData[14]
rlabel metal3 758 27812 758 27812 0 FrameData[15]
rlabel metal3 252 28628 252 28628 0 FrameData[16]
rlabel metal3 758 29444 758 29444 0 FrameData[17]
rlabel metal3 459 30260 459 30260 0 FrameData[18]
rlabel metal1 1196 31790 1196 31790 0 FrameData[19]
rlabel metal3 758 16388 758 16388 0 FrameData[1]
rlabel metal3 804 31892 804 31892 0 FrameData[20]
rlabel metal3 436 32708 436 32708 0 FrameData[21]
rlabel metal3 252 33524 252 33524 0 FrameData[22]
rlabel metal3 528 34340 528 34340 0 FrameData[23]
rlabel metal3 804 35156 804 35156 0 FrameData[24]
rlabel metal3 804 35972 804 35972 0 FrameData[25]
rlabel metal3 804 36788 804 36788 0 FrameData[26]
rlabel metal3 804 37604 804 37604 0 FrameData[27]
rlabel metal3 436 38420 436 38420 0 FrameData[28]
rlabel metal3 804 39236 804 39236 0 FrameData[29]
rlabel metal3 390 17204 390 17204 0 FrameData[2]
rlabel metal3 804 40052 804 40052 0 FrameData[30]
rlabel metal3 804 40868 804 40868 0 FrameData[31]
rlabel metal3 758 18020 758 18020 0 FrameData[3]
rlabel metal3 758 18836 758 18836 0 FrameData[4]
rlabel metal3 758 19652 758 19652 0 FrameData[5]
rlabel metal3 482 20468 482 20468 0 FrameData[6]
rlabel metal3 758 21284 758 21284 0 FrameData[7]
rlabel metal3 758 22100 758 22100 0 FrameData[8]
rlabel metal3 758 22916 758 22916 0 FrameData[9]
rlabel metal3 10433 31348 10433 31348 0 FrameData_O[0]
rlabel metal3 10801 34068 10801 34068 0 FrameData_O[10]
rlabel metal3 10709 34340 10709 34340 0 FrameData_O[11]
rlabel metal3 10387 34612 10387 34612 0 FrameData_O[12]
rlabel metal3 10571 34884 10571 34884 0 FrameData_O[13]
rlabel metal3 10433 35156 10433 35156 0 FrameData_O[14]
rlabel metal3 10847 35428 10847 35428 0 FrameData_O[15]
rlabel metal3 10893 35700 10893 35700 0 FrameData_O[16]
rlabel metal3 10755 35972 10755 35972 0 FrameData_O[17]
rlabel metal3 11077 36244 11077 36244 0 FrameData_O[18]
rlabel metal3 10663 36516 10663 36516 0 FrameData_O[19]
rlabel metal3 10410 31620 10410 31620 0 FrameData_O[1]
rlabel metal3 10847 36788 10847 36788 0 FrameData_O[20]
rlabel metal3 10617 37060 10617 37060 0 FrameData_O[21]
rlabel metal3 10571 37332 10571 37332 0 FrameData_O[22]
rlabel metal3 10709 37604 10709 37604 0 FrameData_O[23]
rlabel metal3 10755 37876 10755 37876 0 FrameData_O[24]
rlabel metal3 10801 38148 10801 38148 0 FrameData_O[25]
rlabel metal3 10663 38420 10663 38420 0 FrameData_O[26]
rlabel metal3 10985 38692 10985 38692 0 FrameData_O[27]
rlabel metal3 10709 38964 10709 38964 0 FrameData_O[28]
rlabel metal3 10433 39236 10433 39236 0 FrameData_O[29]
rlabel metal3 10801 31892 10801 31892 0 FrameData_O[2]
rlabel metal3 10893 39508 10893 39508 0 FrameData_O[30]
rlabel metal3 10801 39780 10801 39780 0 FrameData_O[31]
rlabel metal3 10709 32164 10709 32164 0 FrameData_O[3]
rlabel metal3 10709 32436 10709 32436 0 FrameData_O[4]
rlabel metal3 10433 32708 10433 32708 0 FrameData_O[5]
rlabel metal3 10939 32980 10939 32980 0 FrameData_O[6]
rlabel metal3 10663 33252 10663 33252 0 FrameData_O[7]
rlabel metal3 10893 33524 10893 33524 0 FrameData_O[8]
rlabel metal3 10571 33796 10571 33796 0 FrameData_O[9]
rlabel metal2 1426 2571 1426 2571 0 FrameStrobe[0]
rlabel metal2 6026 55 6026 55 0 FrameStrobe[10]
rlabel metal2 6486 599 6486 599 0 FrameStrobe[11]
rlabel metal1 6256 41650 6256 41650 0 FrameStrobe[12]
rlabel metal1 8832 41582 8832 41582 0 FrameStrobe[13]
rlabel metal3 10212 13260 10212 13260 0 FrameStrobe[14]
rlabel metal1 9706 40358 9706 40358 0 FrameStrobe[15]
rlabel metal1 10120 18734 10120 18734 0 FrameStrobe[16]
rlabel metal2 9246 599 9246 599 0 FrameStrobe[17]
rlabel metal2 9706 55 9706 55 0 FrameStrobe[18]
rlabel metal2 10166 667 10166 667 0 FrameStrobe[19]
rlabel metal2 1886 2112 1886 2112 0 FrameStrobe[1]
rlabel metal2 2346 1228 2346 1228 0 FrameStrobe[2]
rlabel metal2 2806 1296 2806 1296 0 FrameStrobe[3]
rlabel metal2 3266 1058 3266 1058 0 FrameStrobe[4]
rlabel metal2 3726 667 3726 667 0 FrameStrobe[5]
rlabel metal2 828 32572 828 32572 0 FrameStrobe[6]
rlabel metal2 4646 599 4646 599 0 FrameStrobe[7]
rlabel metal2 5106 667 5106 667 0 FrameStrobe[8]
rlabel metal2 5566 1330 5566 1330 0 FrameStrobe[9]
rlabel metal1 1564 42330 1564 42330 0 FrameStrobe_O[0]
rlabel metal2 6026 43644 6026 43644 0 FrameStrobe_O[10]
rlabel metal1 6624 42330 6624 42330 0 FrameStrobe_O[11]
rlabel metal1 7130 42330 7130 42330 0 FrameStrobe_O[12]
rlabel metal1 7544 42330 7544 42330 0 FrameStrobe_O[13]
rlabel metal2 8418 42908 8418 42908 0 FrameStrobe_O[14]
rlabel metal1 8694 42058 8694 42058 0 FrameStrobe_O[15]
rlabel metal1 9154 42330 9154 42330 0 FrameStrobe_O[16]
rlabel metal2 6762 42160 6762 42160 0 FrameStrobe_O[17]
rlabel metal1 7866 41480 7866 41480 0 FrameStrobe_O[18]
rlabel metal1 9752 41786 9752 41786 0 FrameStrobe_O[19]
rlabel metal1 2024 42330 2024 42330 0 FrameStrobe_O[1]
rlabel metal1 2484 42330 2484 42330 0 FrameStrobe_O[2]
rlabel metal1 2898 42330 2898 42330 0 FrameStrobe_O[3]
rlabel metal2 3450 42891 3450 42891 0 FrameStrobe_O[4]
rlabel metal1 3818 42330 3818 42330 0 FrameStrobe_O[5]
rlabel metal1 4278 42330 4278 42330 0 FrameStrobe_O[6]
rlabel metal1 4738 42330 4738 42330 0 FrameStrobe_O[7]
rlabel metal1 5198 42330 5198 42330 0 FrameStrobe_O[8]
rlabel metal1 5612 42330 5612 42330 0 FrameStrobe_O[9]
rlabel metal2 138 30124 138 30124 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 10074 33201 10074 33201 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal1 4416 30090 4416 30090 0 Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 3634 31076 3634 31076 0 Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal1 3266 21862 3266 21862 0 Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal1 2668 22406 2668 22406 0 Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 8418 36890 8418 36890 0 Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 7866 37468 7866 37468 0 Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal1 3726 21114 3726 21114 0 Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 8878 21454 8878 21454 0 Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal1 8050 33422 8050 33422 0 Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 8786 33694 8786 33694 0 Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal1 6762 8330 6762 8330 0 Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 6302 7786 6302 7786 0 Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal1 3082 12682 3082 12682 0 Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal1 9384 8942 9384 8942 0 Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal1 8464 8942 8464 8942 0 Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 8464 6766 8464 6766 0 Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 8878 7854 8878 7854 0 Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal1 9154 7174 9154 7174 0 Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 5658 12444 5658 12444 0 Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 6210 12342 6210 12342 0 Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal1 7130 12920 7130 12920 0 Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal1 6532 12818 6532 12818 0 Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal1 5198 10132 5198 10132 0 Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal1 3726 12410 3726 12410 0 Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal1 6486 10132 6486 10132 0 Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal1 5014 10574 5014 10574 0 Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 2806 16898 2806 16898 0 Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal1 4094 17034 4094 17034 0 Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal1 7498 20026 7498 20026 0 Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal1 7912 20570 7912 20570 0 Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 8326 31450 8326 31450 0 Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 8878 31790 8878 31790 0 Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 8418 30396 8418 30396 0 Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 7590 29954 7590 29954 0 Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 3082 33252 3082 33252 0 Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 3542 33626 3542 33626 0 Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 5382 38556 5382 38556 0 Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal1 4646 38454 4646 38454 0 Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 3266 26724 3266 26724 0 Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal1 4186 26792 4186 26792 0 Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal1 4508 34034 4508 34034 0 Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 4462 34510 4462 34510 0 Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 3726 36108 3726 36108 0 Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal1 3036 35598 3036 35598 0 Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 5658 6732 5658 6732 0 Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal1 7958 28730 7958 28730 0 Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal1 7682 28186 7682 28186 0 Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal1 7912 14926 7912 14926 0 Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal1 8786 14824 8786 14824 0 Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 8786 17476 8786 17476 0 Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal1 8050 17102 8050 17102 0 Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 5290 22270 5290 22270 0 Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel via2 5474 21675 5474 21675 0 Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal1 3588 27914 3588 27914 0 Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 2714 28458 2714 28458 0 Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal1 6302 6834 6302 6834 0 Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 3910 24106 3910 24106 0 Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 4462 23868 4462 23868 0 Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 4830 7514 4830 7514 0 Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel viali 5382 7306 5382 7306 0 Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal1 8970 16014 8970 16014 0 Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal1 8188 16014 8188 16014 0 Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 8786 18462 8786 18462 0 Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal1 7636 18258 7636 18258 0 Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal1 7222 33014 7222 33014 0 Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal1 7176 32538 7176 32538 0 Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal1 2668 23834 2668 23834 0 Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal1 3864 23290 3864 23290 0 Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 5566 34085 5566 34085 0 Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 4968 31858 4968 31858 0 Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 4094 19482 4094 19482 0 Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal1 3174 19278 3174 19278 0 Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 8878 35802 8878 35802 0 Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal1 8280 35258 8280 35258 0 Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 2898 11458 2898 11458 0 Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal1 4462 11662 4462 11662 0 Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 3542 14042 3542 14042 0 Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 5014 16218 5014 16218 0 Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal1 5658 15572 5658 15572 0 Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 8326 10098 8326 10098 0 Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal1 8372 10234 8372 10234 0 Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal1 8096 23834 8096 23834 0 Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal1 8280 24378 8280 24378 0 Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 6302 26860 6302 26860 0 Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal1 5704 26486 5704 26486 0 Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal1 2484 30906 2484 30906 0 Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 2990 32164 2990 32164 0 Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 4094 13974 4094 13974 0 Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal1 4094 37706 4094 37706 0 Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal1 3036 37774 3036 37774 0 Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 3082 15810 3082 15810 0 Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal1 3312 15130 3312 15130 0 Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal1 7820 19210 7820 19210 0 Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal1 8970 19278 8970 19278 0 Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal1 8372 25806 8372 25806 0 Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal1 9016 25466 9016 25466 0 Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal1 4370 5780 4370 5780 0 Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 6394 22950 6394 22950 0 Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 8878 22746 8878 22746 0 Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal1 9476 28186 9476 28186 0 Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal1 6670 24310 6670 24310 0 Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 5842 24650 5842 24650 0 Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 5198 29478 5198 29478 0 Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal1 5198 28730 5198 28730 0 Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal1 5106 18802 5106 18802 0 Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal1 3772 18122 3772 18122 0 Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal1 3680 5202 3680 5202 0 Inst_W_IO_switch_matrix.E1BEG0
rlabel metal2 6026 22780 6026 22780 0 Inst_W_IO_switch_matrix.E1BEG1
rlabel metal1 9660 22610 9660 22610 0 Inst_W_IO_switch_matrix.E1BEG2
rlabel metal1 7866 29716 7866 29716 0 Inst_W_IO_switch_matrix.E1BEG3
rlabel metal1 5842 24378 5842 24378 0 Inst_W_IO_switch_matrix.E2BEG0
rlabel metal2 6486 30022 6486 30022 0 Inst_W_IO_switch_matrix.E2BEG1
rlabel metal1 4094 18938 4094 18938 0 Inst_W_IO_switch_matrix.E2BEG2
rlabel metal2 8234 32572 8234 32572 0 Inst_W_IO_switch_matrix.E2BEG3
rlabel metal1 4646 14042 4646 14042 0 Inst_W_IO_switch_matrix.E2BEG4
rlabel metal2 4370 15674 4370 15674 0 Inst_W_IO_switch_matrix.E2BEG5
rlabel metal1 9016 19482 9016 19482 0 Inst_W_IO_switch_matrix.E2BEG6
rlabel metal2 8602 25466 8602 25466 0 Inst_W_IO_switch_matrix.E2BEG7
rlabel metal2 5198 24140 5198 24140 0 Inst_W_IO_switch_matrix.E2BEGb0
rlabel metal2 4370 32198 4370 32198 0 Inst_W_IO_switch_matrix.E2BEGb1
rlabel metal2 2898 19652 2898 19652 0 Inst_W_IO_switch_matrix.E2BEGb2
rlabel metal1 8464 32402 8464 32402 0 Inst_W_IO_switch_matrix.E2BEGb3
rlabel metal1 4968 11730 4968 11730 0 Inst_W_IO_switch_matrix.E2BEGb4
rlabel metal1 6026 15470 6026 15470 0 Inst_W_IO_switch_matrix.E2BEGb5
rlabel metal1 8924 10778 8924 10778 0 Inst_W_IO_switch_matrix.E2BEGb6
rlabel metal2 8602 24378 8602 24378 0 Inst_W_IO_switch_matrix.E2BEGb7
rlabel metal1 6532 21998 6532 21998 0 Inst_W_IO_switch_matrix.E6BEG0
rlabel metal2 2438 28288 2438 28288 0 Inst_W_IO_switch_matrix.E6BEG1
rlabel metal1 8786 21658 8786 21658 0 Inst_W_IO_switch_matrix.E6BEG10
rlabel metal1 8832 33626 8832 33626 0 Inst_W_IO_switch_matrix.E6BEG11
rlabel metal1 5290 23834 5290 23834 0 Inst_W_IO_switch_matrix.E6BEG2
rlabel metal1 5520 31314 5520 31314 0 Inst_W_IO_switch_matrix.E6BEG3
rlabel metal1 4692 12818 4692 12818 0 Inst_W_IO_switch_matrix.E6BEG4
rlabel metal1 4416 17170 4416 17170 0 Inst_W_IO_switch_matrix.E6BEG5
rlabel metal1 8556 20434 8556 20434 0 Inst_W_IO_switch_matrix.E6BEG6
rlabel metal1 9062 31450 9062 31450 0 Inst_W_IO_switch_matrix.E6BEG7
rlabel metal2 4094 21114 4094 21114 0 Inst_W_IO_switch_matrix.E6BEG8
rlabel metal1 7958 36890 7958 36890 0 Inst_W_IO_switch_matrix.E6BEG9
rlabel metal2 6946 26758 6946 26758 0 Inst_W_IO_switch_matrix.EE4BEG0
rlabel metal2 1794 32130 1794 32130 0 Inst_W_IO_switch_matrix.EE4BEG1
rlabel metal1 3266 27098 3266 27098 0 Inst_W_IO_switch_matrix.EE4BEG10
rlabel metal1 5704 33966 5704 33966 0 Inst_W_IO_switch_matrix.EE4BEG11
rlabel metal2 4370 36278 4370 36278 0 Inst_W_IO_switch_matrix.EE4BEG12
rlabel metal2 8602 28730 8602 28730 0 Inst_W_IO_switch_matrix.EE4BEG13
rlabel metal1 7636 15130 7636 15130 0 Inst_W_IO_switch_matrix.EE4BEG14
rlabel metal1 8878 17306 8878 17306 0 Inst_W_IO_switch_matrix.EE4BEG15
rlabel metal2 4370 38454 4370 38454 0 Inst_W_IO_switch_matrix.EE4BEG2
rlabel metal1 9430 30294 9430 30294 0 Inst_W_IO_switch_matrix.EE4BEG3
rlabel metal1 6762 6970 6762 6970 0 Inst_W_IO_switch_matrix.EE4BEG4
rlabel metal1 6762 7344 6762 7344 0 Inst_W_IO_switch_matrix.EE4BEG5
rlabel metal1 9292 14382 9292 14382 0 Inst_W_IO_switch_matrix.EE4BEG6
rlabel metal1 8740 17646 8740 17646 0 Inst_W_IO_switch_matrix.EE4BEG7
rlabel metal2 2438 33762 2438 33762 0 Inst_W_IO_switch_matrix.EE4BEG8
rlabel metal1 5888 38522 5888 38522 0 Inst_W_IO_switch_matrix.EE4BEG9
rlabel metal1 1196 10982 1196 10982 0 UserCLK
rlabel via2 1357 30260 1357 30260 0 UserCLK_regs
rlabel metal2 1426 42534 1426 42534 0 UserCLKo
rlabel metal3 10479 5236 10479 5236 0 W1END[0]
rlabel metal3 10433 5508 10433 5508 0 W1END[1]
rlabel metal3 10939 5780 10939 5780 0 W1END[2]
rlabel metal3 10479 6052 10479 6052 0 W1END[3]
rlabel metal3 10433 8500 10433 8500 0 W2END[0]
rlabel metal3 10525 8772 10525 8772 0 W2END[1]
rlabel metal3 10479 9044 10479 9044 0 W2END[2]
rlabel metal3 11077 9316 11077 9316 0 W2END[3]
rlabel metal3 10617 9588 10617 9588 0 W2END[4]
rlabel metal3 10433 9860 10433 9860 0 W2END[5]
rlabel metal3 10985 10132 10985 10132 0 W2END[6]
rlabel metal3 10479 10404 10479 10404 0 W2END[7]
rlabel metal3 10479 6324 10479 6324 0 W2MID[0]
rlabel metal3 10433 6596 10433 6596 0 W2MID[1]
rlabel metal3 10571 6868 10571 6868 0 W2MID[2]
rlabel metal3 10433 7140 10433 7140 0 W2MID[3]
rlabel metal3 10525 7412 10525 7412 0 W2MID[4]
rlabel metal3 10479 7684 10479 7684 0 W2MID[5]
rlabel metal3 10433 7956 10433 7956 0 W2MID[6]
rlabel metal3 10571 8228 10571 8228 0 W2MID[7]
rlabel metal3 9973 15028 9973 15028 0 W6END[0]
rlabel metal3 10479 17748 10479 17748 0 W6END[10]
rlabel metal3 10525 18020 10525 18020 0 W6END[11]
rlabel metal3 10847 15300 10847 15300 0 W6END[1]
rlabel metal3 10479 15572 10479 15572 0 W6END[2]
rlabel metal3 10433 15844 10433 15844 0 W6END[3]
rlabel metal3 10525 16116 10525 16116 0 W6END[4]
rlabel metal3 10479 16388 10479 16388 0 W6END[5]
rlabel metal3 10433 16660 10433 16660 0 W6END[6]
rlabel metal3 10433 16932 10433 16932 0 W6END[7]
rlabel metal3 10479 17204 10479 17204 0 W6END[8]
rlabel metal3 10433 17476 10433 17476 0 W6END[9]
rlabel metal3 10019 10676 10019 10676 0 WW4END[0]
rlabel metal3 11077 13396 11077 13396 0 WW4END[10]
rlabel metal3 10571 13668 10571 13668 0 WW4END[11]
rlabel metal3 10755 13940 10755 13940 0 WW4END[12]
rlabel metal3 10939 14212 10939 14212 0 WW4END[13]
rlabel metal3 10019 14484 10019 14484 0 WW4END[14]
rlabel metal3 10479 14756 10479 14756 0 WW4END[15]
rlabel metal3 10525 10948 10525 10948 0 WW4END[1]
rlabel metal3 10571 11220 10571 11220 0 WW4END[2]
rlabel metal3 10479 11492 10479 11492 0 WW4END[3]
rlabel metal3 10479 11764 10479 11764 0 WW4END[4]
rlabel metal3 10433 12036 10433 12036 0 WW4END[5]
rlabel metal3 10525 12308 10525 12308 0 WW4END[6]
rlabel metal3 10709 12580 10709 12580 0 WW4END[7]
rlabel metal3 10479 12852 10479 12852 0 WW4END[8]
rlabel metal3 10433 13124 10433 13124 0 WW4END[9]
rlabel metal2 6854 13124 6854 13124 0 _000_
rlabel metal1 7038 11866 7038 11866 0 _001_
rlabel metal1 8165 8942 8165 8942 0 _002_
rlabel metal2 9522 8602 9522 8602 0 _003_
rlabel via1 8717 6154 8717 6154 0 _004_
rlabel metal1 5658 10030 5658 10030 0 _005_
rlabel metal2 7314 12070 7314 12070 0 _006_
rlabel metal1 6992 12138 6992 12138 0 _007_
rlabel metal1 6808 12410 6808 12410 0 _008_
rlabel metal1 6624 12682 6624 12682 0 _009_
rlabel metal2 9338 13498 9338 13498 0 _010_
rlabel metal1 9338 12954 9338 12954 0 _011_
rlabel metal1 8832 13158 8832 13158 0 _012_
rlabel metal1 8924 8602 8924 8602 0 _013_
rlabel metal2 9246 8058 9246 8058 0 _014_
rlabel metal2 6946 8568 6946 8568 0 _015_
rlabel metal1 8970 7854 8970 7854 0 _016_
rlabel metal1 9062 10982 9062 10982 0 _017_
rlabel metal2 9246 11356 9246 11356 0 _018_
rlabel metal1 9384 7854 9384 7854 0 _019_
rlabel metal2 8510 7854 8510 7854 0 _020_
rlabel metal1 7866 6902 7866 6902 0 _021_
rlabel metal1 8096 6834 8096 6834 0 _022_
rlabel metal2 8602 6902 8602 6902 0 _023_
rlabel metal1 9016 6834 9016 6834 0 _024_
rlabel metal2 8786 7038 8786 7038 0 _025_
rlabel metal1 5566 9928 5566 9928 0 _026_
rlabel metal2 4738 9860 4738 9860 0 _027_
rlabel metal2 5014 9758 5014 9758 0 _028_
rlabel metal1 6348 9350 6348 9350 0 _029_
rlabel metal1 5428 9690 5428 9690 0 _030_
rlabel metal2 5474 9486 5474 9486 0 _031_
rlabel metal2 6394 37638 6394 37638 0 clknet_0_UserCLK
rlabel metal2 7498 35802 7498 35802 0 clknet_0_UserCLK_regs
rlabel metal1 6486 36754 6486 36754 0 clknet_1_0__leaf_UserCLK
rlabel metal2 4278 36516 4278 36516 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal1 6256 35054 6256 35054 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal1 1426 33354 1426 33354 0 net1
rlabel metal1 1150 29274 1150 29274 0 net10
rlabel metal1 2070 6324 2070 6324 0 net100
rlabel metal1 1702 9588 1702 9588 0 net101
rlabel metal2 1012 12206 1012 12206 0 net102
rlabel metal1 1702 11084 1702 11084 0 net103
rlabel metal1 920 12410 920 12410 0 net104
rlabel metal1 1702 7310 1702 7310 0 net105
rlabel metal2 4830 9146 4830 9146 0 net106
rlabel metal1 1564 6630 1564 6630 0 net107
rlabel metal1 1932 6426 1932 6426 0 net108
rlabel metal1 4738 5066 4738 5066 0 net109
rlabel metal2 5382 32436 5382 32436 0 net11
rlabel metal2 1104 17068 1104 17068 0 net110
rlabel metal2 3726 7055 3726 7055 0 net111
rlabel metal1 7866 18394 7866 18394 0 net112
rlabel via1 6877 21998 6877 21998 0 net113
rlabel metal2 9062 29665 9062 29665 0 net114
rlabel metal2 9798 25772 9798 25772 0 net115
rlabel metal3 9407 20468 9407 20468 0 net116
rlabel metal1 6164 19482 6164 19482 0 net117
rlabel metal1 10028 19822 10028 19822 0 net118
rlabel metal3 8878 19380 8878 19380 0 net119
rlabel metal1 2024 6766 2024 6766 0 net12
rlabel metal1 4324 15674 4324 15674 0 net120
rlabel metal2 8786 20468 8786 20468 0 net121
rlabel metal1 9798 20910 9798 20910 0 net122
rlabel metal2 8510 22746 8510 22746 0 net123
rlabel metal3 9085 21964 9085 21964 0 net124
rlabel metal2 4554 20434 4554 20434 0 net125
rlabel metal1 8970 21998 8970 21998 0 net126
rlabel metal2 9384 19482 9384 19482 0 net127
rlabel metal2 5842 21692 5842 21692 0 net128
rlabel metal2 8556 20876 8556 20876 0 net129
rlabel metal1 2392 11730 2392 11730 0 net13
rlabel metal1 8970 23698 8970 23698 0 net130
rlabel metal1 9384 29138 9384 29138 0 net131
rlabel metal1 8372 22202 8372 22202 0 net132
rlabel metal1 8924 31790 8924 31790 0 net133
rlabel metal2 3634 28968 3634 28968 0 net134
rlabel metal2 9384 29478 9384 29478 0 net135
rlabel metal1 9154 30192 9154 30192 0 net136
rlabel metal2 11178 18870 11178 18870 0 net137
rlabel metal3 5980 24820 5980 24820 0 net138
rlabel metal2 8602 23732 8602 23732 0 net139
rlabel metal1 1472 17850 1472 17850 0 net14
rlabel metal2 8786 31178 8786 31178 0 net140
rlabel metal1 7406 30634 7406 30634 0 net141
rlabel metal2 8464 30702 8464 30702 0 net142
rlabel metal1 9522 23732 9522 23732 0 net143
rlabel metal1 9522 27472 9522 27472 0 net144
rlabel metal1 9430 34034 9430 34034 0 net145
rlabel via3 7245 31756 7245 31756 0 net146
rlabel metal1 9154 28050 9154 28050 0 net147
rlabel via3 9453 27676 9453 27676 0 net148
rlabel metal1 8970 17850 8970 17850 0 net149
rlabel metal1 1426 32198 1426 32198 0 net15
rlabel metal1 3220 32198 3220 32198 0 net150
rlabel metal3 7222 32028 7222 32028 0 net151
rlabel metal1 9246 31110 9246 31110 0 net152
rlabel metal2 10856 17204 10856 17204 0 net153
rlabel metal3 5244 14892 5244 14892 0 net154
rlabel via2 9338 14603 9338 14603 0 net155
rlabel metal1 8786 17544 8786 17544 0 net156
rlabel metal1 3680 33830 3680 33830 0 net157
rlabel metal3 7889 35156 7889 35156 0 net158
rlabel metal1 4508 32538 4508 32538 0 net159
rlabel metal4 2576 21420 2576 21420 0 net16
rlabel metal1 2346 33048 2346 33048 0 net160
rlabel metal1 1380 34102 1380 34102 0 net161
rlabel metal1 9016 36142 9016 36142 0 net162
rlabel metal1 8510 35020 8510 35020 0 net163
rlabel metal1 1150 25466 1150 25466 0 net164
rlabel metal2 1978 26333 1978 26333 0 net165
rlabel metal1 6808 35802 6808 35802 0 net166
rlabel metal2 6578 35938 6578 35938 0 net167
rlabel metal2 4186 36992 4186 36992 0 net168
rlabel metal2 5934 36686 5934 36686 0 net169
rlabel metal1 1426 21318 1426 21318 0 net17
rlabel metal1 5014 30906 5014 30906 0 net170
rlabel metal2 1058 7191 1058 7191 0 net171
rlabel metal3 8096 15980 8096 15980 0 net172
rlabel metal4 4324 17340 4324 17340 0 net173
rlabel metal3 6325 16524 6325 16524 0 net174
rlabel metal3 8763 38692 8763 38692 0 net175
rlabel metal3 9131 39372 9131 39372 0 net176
rlabel via2 5934 18955 5934 18955 0 net177
rlabel via2 5106 21131 5106 21131 0 net178
rlabel metal2 460 33422 460 33422 0 net179
rlabel metal1 1472 32946 1472 32946 0 net18
rlabel metal3 1173 10948 1173 10948 0 net180
rlabel metal1 1610 8602 1610 8602 0 net181
rlabel metal1 2346 37128 2346 37128 0 net182
rlabel metal2 3910 39032 3910 39032 0 net183
rlabel metal1 1012 8398 1012 8398 0 net184
rlabel via3 2461 8228 2461 8228 0 net185
rlabel metal3 1633 7956 1633 7956 0 net186
rlabel via2 6302 17867 6302 17867 0 net187
rlabel metal1 6670 36074 6670 36074 0 net188
rlabel metal1 8326 34918 8326 34918 0 net189
rlabel metal1 7544 17646 7544 17646 0 net19
rlabel metal1 7544 32198 7544 32198 0 net190
rlabel metal1 1472 42194 1472 42194 0 net191
rlabel metal1 6486 41242 6486 41242 0 net192
rlabel metal2 6578 41990 6578 41990 0 net193
rlabel metal2 7498 41990 7498 41990 0 net194
rlabel metal1 8234 41786 8234 41786 0 net195
rlabel metal2 8602 41797 8602 41797 0 net196
rlabel metal1 9384 42126 9384 42126 0 net197
rlabel metal1 8924 42262 8924 42262 0 net198
rlabel metal1 7682 41650 7682 41650 0 net199
rlabel metal1 1472 6426 1472 6426 0 net2
rlabel metal1 6854 18258 6854 18258 0 net20
rlabel metal1 8142 41242 8142 41242 0 net200
rlabel metal1 9292 41582 9292 41582 0 net201
rlabel metal1 2208 42058 2208 42058 0 net202
rlabel metal1 2392 42194 2392 42194 0 net203
rlabel metal1 3588 42262 3588 42262 0 net204
rlabel metal1 3634 42092 3634 42092 0 net205
rlabel metal1 4094 42228 4094 42228 0 net206
rlabel metal1 4554 42126 4554 42126 0 net207
rlabel metal1 6302 41480 6302 41480 0 net208
rlabel metal2 5474 41956 5474 41956 0 net209
rlabel metal1 5796 18734 5796 18734 0 net21
rlabel metal1 5842 42160 5842 42160 0 net210
rlabel metal1 3542 41582 3542 41582 0 net211
rlabel metal4 2668 17952 2668 17952 0 net22
rlabel metal3 2024 21556 2024 21556 0 net23
rlabel metal1 1932 10030 1932 10030 0 net24
rlabel metal1 2254 8466 2254 8466 0 net25
rlabel metal1 2254 18700 2254 18700 0 net26
rlabel metal1 2346 37230 2346 37230 0 net27
rlabel metal1 2300 12206 2300 12206 0 net28
rlabel metal2 2346 7616 2346 7616 0 net29
rlabel metal1 2576 17714 2576 17714 0 net3
rlabel metal1 2346 7378 2346 7378 0 net30
rlabel metal1 6072 17646 6072 17646 0 net31
rlabel metal1 1610 20808 1610 20808 0 net32
rlabel via3 7107 21828 7107 21828 0 net33
rlabel metal1 6854 25908 6854 25908 0 net34
rlabel metal1 3128 2618 3128 2618 0 net35
rlabel metal4 11040 12420 11040 12420 0 net36
rlabel metal1 7682 21420 7682 21420 0 net37
rlabel metal3 3542 12716 3542 12716 0 net38
rlabel metal2 4186 6477 4186 6477 0 net39
rlabel metal1 1840 21930 1840 21930 0 net4
rlabel metal2 6762 17204 6762 17204 0 net40
rlabel metal1 5934 8398 5934 8398 0 net41
rlabel metal1 4738 16014 4738 16014 0 net42
rlabel metal1 4830 11186 4830 11186 0 net43
rlabel metal1 2622 5814 2622 5814 0 net44
rlabel metal1 4094 28526 4094 28526 0 net45
rlabel metal2 5014 27438 5014 27438 0 net46
rlabel metal1 7084 9486 7084 9486 0 net47
rlabel metal1 2530 33320 2530 33320 0 net48
rlabel metal1 1886 14518 1886 14518 0 net49
rlabel metal1 2254 23052 2254 23052 0 net5
rlabel metal1 1886 33524 1886 33524 0 net50
rlabel metal1 2300 8398 2300 8398 0 net51
rlabel metal1 1518 28730 1518 28730 0 net52
rlabel metal1 4278 22644 4278 22644 0 net53
rlabel metal1 6486 18258 6486 18258 0 net54
rlabel metal1 4646 14348 4646 14348 0 net55
rlabel metal1 2070 10540 2070 10540 0 net56
rlabel metal2 1426 20315 1426 20315 0 net57
rlabel metal2 2622 30430 2622 30430 0 net58
rlabel metal4 7176 20740 7176 20740 0 net59
rlabel metal1 1610 25160 1610 25160 0 net6
rlabel metal1 5106 7956 5106 7956 0 net60
rlabel metal3 6095 31756 6095 31756 0 net61
rlabel metal1 5842 12274 5842 12274 0 net62
rlabel metal3 7429 20332 7429 20332 0 net63
rlabel metal1 7314 13838 7314 13838 0 net64
rlabel metal1 7176 7514 7176 7514 0 net65
rlabel metal1 7728 7514 7728 7514 0 net66
rlabel metal3 7383 32300 7383 32300 0 net67
rlabel metal2 7590 18428 7590 18428 0 net68
rlabel metal1 7728 7786 7728 7786 0 net69
rlabel metal1 1334 26554 1334 26554 0 net7
rlabel metal3 6785 21284 6785 21284 0 net70
rlabel metal2 9798 19125 9798 19125 0 net71
rlabel metal3 6693 18292 6693 18292 0 net72
rlabel metal1 8050 18938 8050 18938 0 net73
rlabel via1 9982 14603 9982 14603 0 net74
rlabel via1 3805 26894 3805 26894 0 net75
rlabel metal1 3749 35598 3749 35598 0 net76
rlabel metal1 6670 16762 6670 16762 0 net77
rlabel via1 3345 21454 3345 21454 0 net78
rlabel metal1 9016 16218 9016 16218 0 net79
rlabel metal1 2300 19822 2300 19822 0 net8
rlabel metal2 9522 18241 9522 18241 0 net80
rlabel metal1 10097 16762 10097 16762 0 net81
rlabel metal2 7636 17850 7636 17850 0 net82
rlabel metal3 9545 19244 9545 19244 0 net83
rlabel metal1 4140 20978 4140 20978 0 net84
rlabel metal1 4117 13838 4117 13838 0 net85
rlabel metal1 9982 12682 9982 12682 0 net86
rlabel metal1 5290 12818 5290 12818 0 net87
rlabel metal3 5819 26588 5819 26588 0 net88
rlabel metal1 5635 24242 5635 24242 0 net89
rlabel metal2 1702 20434 1702 20434 0 net9
rlabel metal1 7544 19346 7544 19346 0 net90
rlabel metal1 2484 16082 2484 16082 0 net91
rlabel metal2 3082 11441 3082 11441 0 net92
rlabel metal3 6049 16116 6049 16116 0 net93
rlabel metal1 5796 18802 5796 18802 0 net94
rlabel metal3 4784 18020 4784 18020 0 net95
rlabel metal1 8878 12342 8878 12342 0 net96
rlabel via2 7774 13515 7774 13515 0 net97
rlabel metal2 8234 20553 8234 20553 0 net98
rlabel metal1 2254 5202 2254 5202 0 net99
<< properties >>
string FIXED_BBOX 0 0 11250 45000
<< end >>
