* NGSPICE file created from LUT4AB.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd1_1 abstract view
.subckt sg13g2_dlygate4sd1_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VSS VDD B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_inv_16 abstract view
.subckt sg13g2_inv_16 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dfrbp_1 abstract view
.subckt sg13g2_dfrbp_1 CLK RESET_B D Q_N Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_4 abstract view
.subckt sg13g2_buf_4 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_2 abstract view
.subckt sg13g2_mux2_2 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
X_3086_ E6END[5] net138 VPWR VGND sg13g2_buf_1
X_3155_ net1097 net196 VPWR VGND sg13g2_buf_1
XFILLER_39_288 VPWR VGND sg13g2_fill_2
XFILLER_39_255 VPWR VGND sg13g2_fill_2
XFILLER_39_233 VPWR VGND sg13g2_decap_4
X_2106_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q _0746_ _0747_ VPWR VGND sg13g2_nor2_1
X_2037_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0199_ _0683_ VPWR VGND sg13g2_mux4_1
X_2939_ net1171 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_420 VPWR VGND sg13g2_fill_1
Xrebuffer7 Inst_LUT4AB_switch_matrix.JS2BEG4 net380 VPWR VGND sg13g2_dlygate4sd1_1
X_1270_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q _1100_ _1101_ VPWR VGND sg13g2_nor2_1
XFILLER_32_431 VPWR VGND sg13g2_fill_2
X_1606_ _0269_ net987 net1004 VPWR VGND sg13g2_nand2b_1
X_2655_ net1159 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2724_ net1144 net1104 Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_317 VPWR VGND sg13g2_fill_2
X_3207_ NN4END[12] net263 VPWR VGND sg13g2_buf_1
X_1468_ _0134_ VPWR _0135_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q net936 sg13g2_o21ai_1
X_1537_ _0201_ _0149_ _0199_ VPWR VGND sg13g2_nand2_1
X_1399_ VGND VPWR _0057_ _0069_ _0061_ _0068_ sg13g2_a21oi_2
X_2586_ net1177 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q VPWR VGND sg13g2_dlhq_1
X_3138_ net1151 net180 VPWR VGND sg13g2_buf_1
XFILLER_27_258 VPWR VGND sg13g2_decap_8
XFILLER_27_236 VPWR VGND sg13g2_fill_1
XFILLER_27_225 VPWR VGND sg13g2_decap_8
X_3069_ Inst_LUT4AB_switch_matrix.E2BEG2 net119 VPWR VGND sg13g2_buf_1
XFILLER_50_272 VPWR VGND sg13g2_fill_1
XFILLER_37_62 VPWR VGND sg13g2_fill_1
X_2440_ net1175 net1060 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
X_1253_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q net46 net17 net74 net101 Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q
+ _1084_ VPWR VGND sg13g2_mux4_1
X_1322_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q net79 _1150_ _1149_ sg13g2_a21oi_1
X_2371_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q net37 net52 net1211 net963 Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ Inst_LUT4AB_switch_matrix.N4BEG0 VPWR VGND sg13g2_mux4_1
X_1184_ VPWR _1017_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q VGND sg13g2_inv_1
Xoutput253 net253 NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput242 net242 N4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput231 net231 N2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput220 net220 N2BEG[3] VPWR VGND sg13g2_buf_1
X_2569_ net1142 net1083 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
Xoutput264 net264 NN4BEG[9] VPWR VGND sg13g2_buf_1
X_2638_ net1122 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q VPWR VGND sg13g2_dlhq_1
Xoutput275 net275 S2BEG[6] VPWR VGND sg13g2_buf_1
Xoutput286 net286 S4BEG[10] VPWR VGND sg13g2_buf_1
X_2707_ net1199 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q VPWR VGND sg13g2_dlhq_1
Xoutput297 net297 S4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_11_456 VPWR VGND sg13g2_fill_2
XFILLER_23_31 VPWR VGND sg13g2_fill_2
XFILLER_23_42 VPWR VGND sg13g2_fill_1
XFILLER_38_309 VPWR VGND sg13g2_fill_1
XFILLER_2_198 VPWR VGND sg13g2_fill_1
XFILLER_2_176 VPWR VGND sg13g2_fill_1
XFILLER_0_46 VPWR VGND sg13g2_fill_1
X_1940_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q _0585_ net981 _0588_ _0587_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
+ _0590_ VPWR VGND sg13g2_mux4_1
X_1871_ _0523_ net105 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VPWR VGND sg13g2_nand2_1
X_2423_ Inst_LF_LUT4c_frame_config_dffesr.c_reset_value _0496_ _1005_ _1006_ VPWR
+ VGND sg13g2_mux2_1
X_2285_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q net953 net936 net931 net929 Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0909_ VPWR VGND sg13g2_mux4_1
XFILLER_37_342 VPWR VGND sg13g2_decap_4
XFILLER_37_331 VPWR VGND sg13g2_decap_8
X_1236_ _1068_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1067_ VPWR VGND sg13g2_nand2_2
X_1305_ VPWR _1134_ _1133_ VGND sg13g2_inv_1
X_2354_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q net950 _0237_ Inst_LUT4AB_switch_matrix.JS2BEG0
+ net376 Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q Inst_LUT4AB_switch_matrix.W1BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_20_231 VPWR VGND sg13g2_decap_4
XFILLER_3_452 VPWR VGND sg13g2_fill_2
X_2070_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q net974 net969 net939 net945 Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ _0713_ VPWR VGND sg13g2_mux4_1
X_2972_ net1168 net1051 Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1923_ _0574_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q net13 VPWR VGND sg13g2_nand2b_1
X_1854_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q _0506_ _0507_ VPWR VGND sg13g2_and2_1
X_1785_ net984 net1009 net40 net1216 net11 Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ _0441_ VPWR VGND sg13g2_mux4_1
X_2406_ _0993_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q net925 VPWR VGND sg13g2_nand2_1
X_1219_ VPWR _1052_ net935 VGND sg13g2_inv_1
X_2337_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q _0953_ _0954_ VPWR VGND sg13g2_nor2_1
X_2268_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q VPWR _0893_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ _0148_ sg13g2_o21ai_1
X_2199_ net1002 net1210 _0834_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_194 VPWR VGND sg13g2_decap_8
XFILLER_25_378 VPWR VGND sg13g2_decap_8
XFILLER_45_62 VPWR VGND sg13g2_fill_2
X_3240_ S4END[9] net296 VPWR VGND sg13g2_buf_1
X_1570_ net20 Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0233_ VPWR VGND sg13g2_nor2b_1
Xfanout1050 net1052 net1050 VPWR VGND sg13g2_buf_1
Xfanout1083 net1085 net1083 VPWR VGND sg13g2_buf_1
X_3171_ Inst_LUT4AB_switch_matrix.JN2BEG4 net221 VPWR VGND sg13g2_buf_2
Xfanout1072 net1073 net1072 VPWR VGND sg13g2_buf_1
X_2122_ _0758_ _0697_ _0752_ _0762_ VPWR VGND sg13g2_mux2_1
X_2053_ _0696_ _0697_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q Inst_LUT4AB_switch_matrix.M_AD
+ VPWR VGND sg13g2_mux2_1
Xfanout1061 net1062 net1061 VPWR VGND sg13g2_buf_1
Xfanout1094 net1095 net1094 VPWR VGND sg13g2_buf_1
XFILLER_20_4 VPWR VGND sg13g2_fill_2
X_2955_ net1129 net1052 Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_120 VPWR VGND sg13g2_decap_8
X_1837_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0487_ _0491_ VPWR VGND sg13g2_mux4_1
X_1906_ net48 net19 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q _0557_ VPWR VGND sg13g2_mux2_1
X_1768_ _0423_ VPWR _0424_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q _0420_ sg13g2_o21ai_1
X_2886_ net1135 net1033 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1699_ _0357_ VPWR _0358_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q net93 sg13g2_o21ai_1
XFILLER_25_120 VPWR VGND sg13g2_fill_1
XFILLER_40_189 VPWR VGND sg13g2_fill_2
XFILLER_40_167 VPWR VGND sg13g2_fill_1
XFILLER_48_223 VPWR VGND sg13g2_fill_2
X_2740_ net1196 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q VPWR VGND sg13g2_dlhq_1
X_1622_ VGND VPWR _0283_ _0284_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q Inst_LUT4AB_switch_matrix.E2BEG3
+ sg13g2_a21oi_2
X_2671_ net1119 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q VPWR VGND sg13g2_dlhq_1
X_3223_ Inst_LUT4AB_switch_matrix.JS2BEG4 net273 VPWR VGND sg13g2_buf_1
X_1553_ _0216_ VPWR _0217_ VGND net997 net941 sg13g2_o21ai_1
X_1484_ _0150_ net990 net966 VPWR VGND sg13g2_nand2b_1
XFILLER_54_237 VPWR VGND sg13g2_fill_2
X_3085_ E6END[4] net137 VPWR VGND sg13g2_buf_1
X_2036_ _0678_ _0681_ _0679_ _0682_ VPWR VGND sg13g2_nor3_2
X_2105_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q _0743_ _0746_ _0745_ sg13g2_a21oi_1
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_3154_ net1102 net195 VPWR VGND sg13g2_buf_1
X_2938_ net1177 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_329 VPWR VGND sg13g2_fill_2
XFILLER_22_167 VPWR VGND sg13g2_decap_8
X_2869_ net1192 net1036 Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q VPWR VGND sg13g2_dlhq_1
XFILLER_45_237 VPWR VGND sg13g2_fill_1
Xrebuffer8 _0640_ net381 VPWR VGND sg13g2_buf_2
XFILLER_42_63 VPWR VGND sg13g2_fill_1
X_2723_ net1148 net1107 Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_0 VPWR VGND sg13g2_fill_2
X_1605_ _0265_ _0267_ _0268_ VPWR VGND sg13g2_nor2_1
X_1536_ _0149_ _0199_ _0200_ VPWR VGND sg13g2_nor2_1
X_2585_ net1180 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2654_ net1162 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q VPWR VGND sg13g2_dlhq_1
X_3206_ NN4END[11] net262 VPWR VGND sg13g2_buf_1
X_1467_ _0134_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_switch_matrix.M_EF
+ VPWR VGND sg13g2_nand2b_1
X_3137_ net1154 net179 VPWR VGND sg13g2_buf_1
X_1398_ VGND VPWR _1160_ _0052_ _0067_ _0050_ _0068_ _0049_ sg13g2_a221oi_1
X_2019_ _0667_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_nand2_1
X_3068_ net382 net118 VPWR VGND sg13g2_buf_1
XFILLER_23_432 VPWR VGND sg13g2_fill_1
XFILLER_53_73 VPWR VGND sg13g2_fill_1
XFILLER_5_174 VPWR VGND sg13g2_fill_1
X_2370_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q net38 net53 net1213 net958 Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ Inst_LUT4AB_switch_matrix.N4BEG1 VPWR VGND sg13g2_mux4_1
X_1252_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q net16 net73 net100 Inst_LUT4AB_switch_matrix.E2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q _1083_ VPWR VGND sg13g2_mux4_1
X_1321_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q net67 _1149_ VPWR VGND sg13g2_nor2b_1
X_1183_ VPWR _1016_ net1217 VGND sg13g2_inv_1
X_2706_ net1202 net1104 Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_20_424 VPWR VGND sg13g2_fill_1
Xoutput210 net210 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_2568_ net1176 net1083 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
Xoutput254 Inst_LUT4AB_switch_matrix.NN4BEG2 NN4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput232 net232 N2BEGb[7] VPWR VGND sg13g2_buf_1
X_1519_ _0183_ VPWR _0184_ VGND net60 net988 sg13g2_o21ai_1
Xoutput243 net243 N4BEG[4] VPWR VGND sg13g2_buf_1
X_2637_ net1123 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q VPWR VGND sg13g2_dlhq_1
Xoutput221 net221 N2BEG[4] VPWR VGND sg13g2_buf_1
X_2499_ net1148 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
Xoutput265 net265 S1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput276 net276 S2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput298 net298 S4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput287 net287 S4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_55_376 VPWR VGND sg13g2_fill_1
X_1870_ _0522_ net78 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VPWR VGND sg13g2_nand2b_1
X_2422_ _1005_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q net925 VPWR VGND sg13g2_nand2_1
X_2353_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q net934 Inst_LUT4AB_switch_matrix.JS2BEG1
+ net980 _0623_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q Inst_LUT4AB_switch_matrix.W1BEG2
+ VPWR VGND sg13g2_mux4_1
X_2284_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q _1158_ _0196_ _0276_ _0556_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0908_ VPWR VGND sg13g2_mux4_1
X_1235_ net934 net928 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1067_ VPWR VGND sg13g2_mux2_1
X_1304_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q net57 net24 net1217 net1212 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ _1133_ VPWR VGND sg13g2_mux4_1
X_1999_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q VPWR _0647_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q
+ _0538_ sg13g2_o21ai_1
XFILLER_43_357 VPWR VGND sg13g2_fill_1
XFILLER_50_96 VPWR VGND sg13g2_fill_2
XFILLER_7_269 VPWR VGND sg13g2_fill_1
Xfanout1210 net1211 net1210 VPWR VGND sg13g2_buf_1
X_2971_ net1171 net1051 Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1922_ _0572_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q _0573_ VPWR VGND sg13g2_nor2b_1
X_1853_ _0505_ VPWR _0506_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0504_ sg13g2_o21ai_1
X_1784_ VGND VPWR _0439_ _0440_ _0433_ _1039_ sg13g2_a21oi_2
XFILLER_41_0 VPWR VGND sg13g2_fill_1
X_2336_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q net1010 net87 net1217 net973 Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
+ _0953_ VPWR VGND sg13g2_mux4_1
X_2405_ _0992_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q net927 VPWR VGND sg13g2_nand2b_1
X_1218_ net951 _1051_ VPWR VGND sg13g2_inv_16
X_2198_ VGND VPWR _1028_ net1002 _0833_ _0832_ sg13g2_a21oi_1
X_2267_ _0887_ _0892_ Inst_LUT4AB_switch_matrix.SS4BEG1 VPWR VGND sg13g2_nor2_1
Xhold20 Inst_LF_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net393 sg13g2_dlygate4sd3_1
XFILLER_0_423 VPWR VGND sg13g2_fill_1
XFILLER_45_52 VPWR VGND sg13g2_fill_1
XFILLER_45_41 VPWR VGND sg13g2_fill_1
XFILLER_43_154 VPWR VGND sg13g2_decap_4
XFILLER_43_143 VPWR VGND sg13g2_decap_4
XFILLER_31_316 VPWR VGND sg13g2_decap_8
XFILLER_16_357 VPWR VGND sg13g2_fill_1
Xfanout1040 net1041 net1040 VPWR VGND sg13g2_buf_1
X_3170_ Inst_LUT4AB_switch_matrix.JN2BEG3 net220 VPWR VGND sg13g2_buf_1
Xfanout1084 net1085 net1084 VPWR VGND sg13g2_buf_1
Xfanout1051 net1052 net1051 VPWR VGND sg13g2_buf_1
X_2121_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0760_ _0759_ _0761_ VPWR VGND
+ sg13g2_nor3_2
X_2052_ _0696_ net930 _0693_ _0697_ VPWR VGND sg13g2_mux2_1
Xfanout1073 net1074 net1073 VPWR VGND sg13g2_buf_1
Xfanout1095 FrameStrobe[12] net1095 VPWR VGND sg13g2_buf_1
XFILLER_13_4 VPWR VGND sg13g2_fill_1
Xfanout1062 FrameStrobe[18] net1062 VPWR VGND sg13g2_buf_1
X_1905_ _0554_ VPWR _0556_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q _0555_ sg13g2_o21ai_1
X_2954_ net1132 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q VPWR VGND sg13g2_dlhq_1
X_2885_ net1138 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_305 VPWR VGND sg13g2_decap_4
X_1836_ _0490_ _0486_ _0487_ VPWR VGND sg13g2_nand2_1
X_1698_ _0357_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q _1030_ VPWR VGND sg13g2_nand2_1
X_1767_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q _0422_ _0421_ _0423_ VPWR VGND sg13g2_nand3_1
X_2319_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q net1008 net61 net1215 net960 Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ _0938_ VPWR VGND sg13g2_mux4_1
XFILLER_15_22 VPWR VGND sg13g2_fill_2
Xinput110 WW4END[2] net110 VPWR VGND sg13g2_buf_1
XFILLER_48_268 VPWR VGND sg13g2_fill_2
XFILLER_44_452 VPWR VGND sg13g2_fill_2
XFILLER_31_168 VPWR VGND sg13g2_fill_1
XFILLER_31_124 VPWR VGND sg13g2_fill_1
X_1552_ _0216_ net997 net946 VPWR VGND sg13g2_nand2b_1
X_2670_ net1120 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1621_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q net81 _0283_ VPWR VGND sg13g2_nor2b_1
X_2104_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VPWR _0745_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ _0744_ sg13g2_o21ai_1
X_1483_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q _0147_ _0148_ _0130_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q
+ _0149_ VPWR VGND sg13g2_mux4_1
X_3153_ net1106 net194 VPWR VGND sg13g2_buf_1
X_3222_ Inst_LUT4AB_switch_matrix.JS2BEG3 net272 VPWR VGND sg13g2_buf_1
X_3084_ E6END[3] net136 VPWR VGND sg13g2_buf_1
X_2035_ _0680_ _0676_ _0681_ VPWR VGND sg13g2_nor2b_1
X_2937_ net1180 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2868_ net1195 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_179 VPWR VGND sg13g2_fill_1
X_2799_ net1119 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1819_ _0473_ _0470_ _0472_ _0469_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q VPWR
+ VGND sg13g2_a22oi_1
XFILLER_53_260 VPWR VGND sg13g2_fill_1
XFILLER_26_98 VPWR VGND sg13g2_fill_1
Xrebuffer9 Inst_LUT4AB_switch_matrix.E2BEG1 net382 VPWR VGND sg13g2_dlygate4sd1_1
X_2722_ net1151 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_319 VPWR VGND sg13g2_fill_1
X_2584_ net1185 net1085 Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1604_ _1042_ VPWR _0267_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0266_ sg13g2_o21ai_1
X_1535_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q _0197_ _0198_ _0170_ _0169_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q
+ _0199_ VPWR VGND sg13g2_mux4_1
X_2653_ net1166 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3205_ NN4END[10] net261 VPWR VGND sg13g2_buf_1
X_1466_ net959 net954 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q _0133_ VPWR VGND sg13g2_mux2_1
X_3136_ net1157 net178 VPWR VGND sg13g2_buf_1
X_1397_ _0067_ _0064_ _0066_ _0063_ _0062_ VPWR VGND sg13g2_a22oi_1
X_3067_ Inst_LUT4AB_switch_matrix.E2BEG0 net117 VPWR VGND sg13g2_buf_2
X_2018_ VGND VPWR _0659_ _0666_ _0665_ _0661_ sg13g2_a21oi_2
XFILLER_2_359 VPWR VGND sg13g2_fill_1
X_1320_ VGND VPWR _1147_ _1025_ _1145_ _1024_ _1148_ _1143_ sg13g2_a221oi_1
X_1251_ _1082_ _1019_ _1075_ Inst_LUT4AB_switch_matrix.E2BEG3 VPWR VGND sg13g2_a21o_2
X_1182_ VPWR _1015_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VGND sg13g2_inv_1
XFILLER_24_208 VPWR VGND sg13g2_fill_2
Xoutput200 net200 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_2636_ net1127 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q VPWR VGND sg13g2_dlhq_1
X_2705_ net1204 net1104 Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q VPWR VGND sg13g2_dlhq_1
Xoutput255 Inst_LUT4AB_switch_matrix.NN4BEG3 NN4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput244 net244 N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput211 net211 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_2567_ net1208 net1086 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
Xoutput222 Inst_LUT4AB_switch_matrix.JN2BEG5 N2BEG[5] VPWR VGND sg13g2_buf_1
X_1518_ _0183_ net988 net68 VPWR VGND sg13g2_nand2b_1
Xoutput233 net233 N4BEG[0] VPWR VGND sg13g2_buf_1
X_2498_ net1150 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
Xoutput266 net266 S1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput277 net277 S2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput299 net299 S4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput288 net288 S4BEG[12] VPWR VGND sg13g2_buf_1
X_1449_ net975 net970 net993 _0117_ VPWR VGND sg13g2_mux2_1
X_3119_ net1117 net191 VPWR VGND sg13g2_buf_1
XFILLER_7_418 VPWR VGND sg13g2_fill_2
XFILLER_11_458 VPWR VGND sg13g2_fill_1
XFILLER_2_167 VPWR VGND sg13g2_fill_2
X_2421_ _1004_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q net927 VPWR VGND sg13g2_nand2b_1
X_2283_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q
+ _0906_ _0902_ _0907_ _0905_ sg13g2_a221oi_1
X_1303_ _1131_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q _1132_ VPWR VGND sg13g2_nor2b_1
X_2352_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q A _1159_ Inst_LUT4AB_switch_matrix.JS2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q Inst_LUT4AB_switch_matrix.W1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_49_193 VPWR VGND sg13g2_fill_2
XFILLER_37_355 VPWR VGND sg13g2_fill_1
X_1234_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q net55 net65 net8 net92 Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q
+ _1066_ VPWR VGND sg13g2_mux4_1
XFILLER_52_369 VPWR VGND sg13g2_fill_1
X_1998_ _0556_ _0561_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q _0646_ VPWR VGND sg13g2_mux2_1
X_2619_ net1172 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_28_322 VPWR VGND sg13g2_fill_2
Xfanout1200 FrameData[12] net1200 VPWR VGND sg13g2_buf_1
Xfanout1211 E6END[1] net1211 VPWR VGND sg13g2_buf_1
XFILLER_3_454 VPWR VGND sg13g2_fill_1
XFILLER_19_300 VPWR VGND sg13g2_fill_1
X_2970_ net1177 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1921_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0570_ _0572_ _0571_ sg13g2_a21oi_1
X_1852_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0503_ _0505_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q
+ sg13g2_a21oi_1
X_1783_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VPWR _0439_ VGND _0438_ _0437_ sg13g2_o21ai_1
X_2335_ VPWR _0952_ _0951_ VGND sg13g2_inv_1
X_2266_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q _0888_ _0892_ _0891_
+ sg13g2_a21oi_1
X_2404_ net394 _0991_ _0990_ _0001_ VPWR VGND sg13g2_mux2_1
X_1217_ VPWR _1050_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q VGND sg13g2_inv_1
XFILLER_25_325 VPWR VGND sg13g2_fill_1
X_2197_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q VPWR _0832_ VGND net91 net1001 sg13g2_o21ai_1
XFILLER_0_457 VPWR VGND sg13g2_fill_2
Xhold21 Inst_LA_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net394 sg13g2_dlygate4sd3_1
XFILLER_45_64 VPWR VGND sg13g2_fill_1
XFILLER_43_188 VPWR VGND sg13g2_fill_2
X_2120_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0757_ _0760_ VPWR VGND sg13g2_nor2_1
Xfanout1074 net1076 net1074 VPWR VGND sg13g2_buf_1
Xfanout1052 FrameStrobe[2] net1052 VPWR VGND sg13g2_buf_1
Xfanout1063 net1064 net1063 VPWR VGND sg13g2_buf_1
Xfanout1041 FrameStrobe[4] net1041 VPWR VGND sg13g2_buf_1
XFILLER_20_6 VPWR VGND sg13g2_fill_1
Xfanout1030 net1031 net1030 VPWR VGND sg13g2_buf_1
X_2051_ net942 net948 _0695_ _0696_ VPWR VGND sg13g2_mux2_1
Xfanout1096 net1097 net1096 VPWR VGND sg13g2_buf_1
Xfanout1085 net1086 net1085 VPWR VGND sg13g2_buf_1
X_1904_ net18 net75 Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q _0555_ VPWR VGND sg13g2_mux2_1
X_1835_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0487_ _0489_ VPWR VGND sg13g2_mux4_1
X_2953_ net1141 net1049 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q VPWR VGND sg13g2_dlhq_1
X_2884_ net1146 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1697_ VGND VPWR _0356_ _0355_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q sg13g2_or2_1
X_1766_ _0422_ net106 Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VPWR VGND sg13g2_nand2b_1
XFILLER_57_214 VPWR VGND sg13g2_fill_2
X_2318_ _0933_ _0936_ _0937_ VPWR VGND sg13g2_nor2_1
X_2249_ VGND VPWR _0876_ _0877_ _0875_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q sg13g2_a21oi_2
XFILLER_31_66 VPWR VGND sg13g2_fill_2
Xinput111 WW4END[3] net111 VPWR VGND sg13g2_buf_1
XFILLER_0_221 VPWR VGND sg13g2_fill_1
Xinput100 W2MID[2] net100 VPWR VGND sg13g2_buf_1
XFILLER_56_41 VPWR VGND sg13g2_fill_2
X_1551_ _0211_ _0214_ _0215_ VPWR VGND sg13g2_nor2_1
X_1482_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q net46 net17 net74 net101 Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q
+ _0148_ VPWR VGND sg13g2_mux4_1
X_1620_ net57 net8 Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q _0282_ VPWR VGND sg13g2_mux2_1
X_3152_ net1015 net212 VPWR VGND sg13g2_buf_1
X_3083_ E6END[2] net133 VPWR VGND sg13g2_buf_1
X_2103_ net59 net61 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q _0744_ VPWR VGND sg13g2_mux2_1
X_3221_ Inst_LUT4AB_switch_matrix.JS2BEG2 net271 VPWR VGND sg13g2_buf_1
XFILLER_47_280 VPWR VGND sg13g2_fill_1
X_2034_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0199_ _0680_ VPWR VGND sg13g2_mux4_1
X_2867_ net1200 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2798_ net1122 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q VPWR VGND sg13g2_dlhq_1
X_2936_ net1183 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1818_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q _0471_ _0472_ VPWR VGND sg13g2_nor2_1
X_1749_ _0406_ net985 net929 VPWR VGND sg13g2_nand2b_1
XFILLER_42_21 VPWR VGND sg13g2_fill_1
XFILLER_51_209 VPWR VGND sg13g2_fill_2
XFILLER_36_228 VPWR VGND sg13g2_decap_8
X_2721_ net1153 net1107 Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2652_ net1168 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_2 VPWR VGND sg13g2_fill_1
X_3204_ NN4END[9] net260 VPWR VGND sg13g2_buf_1
X_1465_ _0132_ _0131_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR VGND sg13g2_nand2b_1
X_2583_ net1188 net1085 Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VPWR VGND sg13g2_dlhq_1
X_1603_ net1008 net41 net987 _0266_ VPWR VGND sg13g2_mux2_1
X_1534_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q net48 net19 net76 net103 Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q
+ _0198_ VPWR VGND sg13g2_mux4_1
X_2017_ _0655_ _0664_ _0665_ VPWR VGND sg13g2_nor2b_1
X_3135_ net1160 net177 VPWR VGND sg13g2_buf_1
X_1396_ _1085_ _0065_ _0066_ VPWR VGND sg13g2_and2_1
X_2919_ net1207 net1046 Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_41_242 VPWR VGND sg13g2_decap_8
XFILLER_37_87 VPWR VGND sg13g2_decap_8
X_3049__369 VPWR VGND net369 sg13g2_tiehi
XFILLER_41_275 VPWR VGND sg13g2_fill_1
XFILLER_41_253 VPWR VGND sg13g2_fill_1
X_1250_ VGND VPWR _1080_ _1081_ _1082_ _1077_ sg13g2_a21oi_1
X_1181_ VPWR _1014_ net1213 VGND sg13g2_inv_1
Xoutput201 net201 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput212 net212 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_2635_ net1129 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q VPWR VGND sg13g2_dlhq_1
Xoutput234 net234 N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput223 net223 N2BEG[6] VPWR VGND sg13g2_buf_1
X_2704_ net1114 net1104 Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VPWR VGND sg13g2_dlhq_1
Xoutput256 net256 NN4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput245 net245 N4BEG[6] VPWR VGND sg13g2_buf_1
X_2566_ net1137 net1081 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_55_301 VPWR VGND sg13g2_fill_2
X_1517_ _1035_ _0181_ _0182_ VPWR VGND sg13g2_nor2_1
X_2497_ net1154 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
Xoutput289 net289 S4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput267 Inst_LUT4AB_switch_matrix.S1BEG2 S1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput278 net278 S2BEGb[1] VPWR VGND sg13g2_buf_1
X_1448_ _0115_ VPWR _0116_ VGND net993 net945 sg13g2_o21ai_1
X_3118_ net1121 net190 VPWR VGND sg13g2_buf_1
XFILLER_55_367 VPWR VGND sg13g2_fill_2
X_1379_ _0049_ _0048_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VPWR VGND sg13g2_nand2_2
X_3049_ UserCLK net369 _0002_ _3049_/Q_N Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
XFILLER_23_12 VPWR VGND sg13g2_fill_2
X_2420_ net396 _1003_ _1001_ _0005_ VPWR VGND sg13g2_mux2_1
X_2282_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q net941 net946 net965 net958 Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0906_ VPWR VGND sg13g2_mux4_1
X_2351_ _0963_ _0965_ Inst_LUT4AB_switch_matrix.NN4BEG0 VPWR VGND sg13g2_nor2_1
X_1302_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q _1130_ _1131_ VPWR VGND sg13g2_nor2_1
X_1233_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q net24 net81 net97 Inst_LUT4AB_switch_matrix.E2BEG1
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q _1065_ VPWR VGND sg13g2_mux4_1
X_1997_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0642_ _0644_ _0645_ VPWR VGND sg13g2_or3_1
XFILLER_20_256 VPWR VGND sg13g2_fill_2
X_2549_ net1193 net1077 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
X_2618_ net1178 net1092 Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_28_345 VPWR VGND sg13g2_fill_2
XFILLER_18_45 VPWR VGND sg13g2_fill_1
XFILLER_55_164 VPWR VGND sg13g2_fill_2
XFILLER_43_337 VPWR VGND sg13g2_fill_2
XFILLER_50_98 VPWR VGND sg13g2_fill_1
XFILLER_3_400 VPWR VGND sg13g2_fill_1
XFILLER_59_30 VPWR VGND sg13g2_fill_1
Xfanout1201 net1203 net1201 VPWR VGND sg13g2_buf_1
Xfanout1212 net1213 net1212 VPWR VGND sg13g2_buf_1
X_1920_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR _0571_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ _0568_ sg13g2_o21ai_1
X_1851_ net976 net972 net996 _0504_ VPWR VGND sg13g2_mux2_1
X_1782_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VPWR _0438_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ _0435_ sg13g2_o21ai_1
X_2403_ Inst_LA_LUT4c_frame_config_dffesr.c_reset_value _0069_ _0989_ _0991_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_57_407 VPWR VGND sg13g2_fill_2
X_1216_ VPWR _1049_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VGND sg13g2_inv_1
X_2334_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q VPWR _0951_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
+ _0950_ sg13g2_o21ai_1
XFILLER_27_0 VPWR VGND sg13g2_fill_2
X_2265_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q VPWR _0891_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ _0890_ sg13g2_o21ai_1
X_2196_ _0830_ VPWR _0831_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0829_ sg13g2_o21ai_1
Xhold22 Inst_LB_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net395 sg13g2_dlygate4sd3_1
XFILLER_43_123 VPWR VGND sg13g2_fill_2
XFILLER_28_197 VPWR VGND sg13g2_fill_2
XFILLER_28_164 VPWR VGND sg13g2_decap_8
XFILLER_28_131 VPWR VGND sg13g2_fill_2
XFILLER_16_304 VPWR VGND sg13g2_decap_8
XFILLER_16_315 VPWR VGND sg13g2_fill_2
Xfanout1086 FrameStrobe[14] net1086 VPWR VGND sg13g2_buf_1
X_2050_ _0694_ VPWR _0695_ VGND _0693_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q
+ sg13g2_o21ai_1
Xfanout1075 net1076 net1075 VPWR VGND sg13g2_buf_1
Xfanout1020 FrameStrobe[8] net1020 VPWR VGND sg13g2_buf_1
Xfanout1097 FrameStrobe[12] net1097 VPWR VGND sg13g2_buf_1
Xfanout1053 net1054 net1053 VPWR VGND sg13g2_buf_1
Xfanout1031 FrameStrobe[6] net1031 VPWR VGND sg13g2_buf_1
Xfanout1064 net1065 net1064 VPWR VGND sg13g2_buf_1
Xfanout1042 net1043 net1042 VPWR VGND sg13g2_buf_1
X_2952_ net1174 net1048 Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VPWR VGND sg13g2_dlhq_1
XFILLER_19_175 VPWR VGND sg13g2_fill_2
X_1834_ _0486_ _0487_ _0488_ VPWR VGND sg13g2_nor2_1
X_1903_ Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ _0553_ _0554_ VPWR VGND sg13g2_a21o_1
XFILLER_30_362 VPWR VGND sg13g2_fill_2
X_1765_ _0421_ Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_nand2_2
X_2883_ net1149 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1696_ net1211 net66 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q _0355_ VPWR VGND sg13g2_mux2_1
X_2317_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q VPWR _0936_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
+ _0935_ sg13g2_o21ai_1
X_2248_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VPWR _0876_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ _0873_ sg13g2_o21ai_1
X_2179_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VPWR _0815_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ _0813_ sg13g2_o21ai_1
X_3297_ W6END[11] net349 VPWR VGND sg13g2_buf_1
Xinput101 W2MID[3] net101 VPWR VGND sg13g2_buf_1
XFILLER_44_454 VPWR VGND sg13g2_fill_1
XFILLER_12_395 VPWR VGND sg13g2_fill_2
X_1550_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VPWR _0214_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ _0213_ sg13g2_o21ai_1
X_1481_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q net45 net100 net16 Inst_LUT4AB_switch_matrix.E2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q _0147_ VPWR VGND sg13g2_mux4_1
X_3220_ Inst_LUT4AB_switch_matrix.JS2BEG1 net270 VPWR VGND sg13g2_buf_1
X_3151_ net1018 net211 VPWR VGND sg13g2_buf_1
XFILLER_39_237 VPWR VGND sg13g2_fill_1
X_2102_ _0742_ VPWR _0743_ VGND net83 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q sg13g2_o21ai_1
X_3082_ net21 net132 VPWR VGND sg13g2_buf_1
X_2033_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q _0452_ _0454_ _0430_ _0424_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q
+ _0679_ VPWR VGND sg13g2_mux4_1
X_2935_ net1186 net1046 Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2866_ net1203 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2797_ net1125 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1748_ VGND VPWR _0404_ _0405_ _1051_ net985 sg13g2_a21oi_2
X_1817_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q _0329_ _0471_ VPWR VGND sg13g2_nor2_1
X_1679_ _0336_ VPWR _0339_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q _0338_ sg13g2_o21ai_1
XFILLER_38_270 VPWR VGND sg13g2_fill_1
XFILLER_26_454 VPWR VGND sg13g2_fill_1
XFILLER_13_148 VPWR VGND sg13g2_fill_1
XFILLER_3_49 VPWR VGND sg13g2_fill_2
XFILLER_17_432 VPWR VGND sg13g2_fill_1
X_2582_ net1191 net1084 Inst_LH_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
X_1602_ VGND VPWR net12 net987 _0265_ _0264_ sg13g2_a21oi_1
X_2651_ net1171 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2720_ net1157 net1107 Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3203_ NN4END[8] net259 VPWR VGND sg13g2_buf_1
X_1464_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q net976 net972 net942 net947 Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0131_ VPWR VGND sg13g2_mux4_1
X_1533_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q net47 net18 net75 net380 Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q
+ _0197_ VPWR VGND sg13g2_mux4_1
X_1395_ _0065_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 net982 VPWR
+ VGND sg13g2_nand2b_1
X_2016_ _0645_ _0663_ net381 _0664_ VPWR VGND sg13g2_nand3_1
X_3134_ net1163 net176 VPWR VGND sg13g2_buf_1
XFILLER_35_240 VPWR VGND sg13g2_fill_1
XFILLER_27_207 VPWR VGND sg13g2_fill_1
X_2918_ net1135 net1038 Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q VPWR VGND sg13g2_dlhq_1
X_2849_ net1154 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_37_55 VPWR VGND sg13g2_decap_8
XFILLER_49_387 VPWR VGND sg13g2_fill_1
X_1180_ VPWR _1013_ net4 VGND sg13g2_inv_1
Xoutput257 net257 NN4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput235 net235 N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput202 net202 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_2565_ net1140 net1079 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_57_0 VPWR VGND sg13g2_fill_2
X_1516_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0179_ _0181_ _0180_ sg13g2_a21oi_1
Xoutput246 net246 N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput224 net224 N2BEG[7] VPWR VGND sg13g2_buf_1
X_2634_ net1132 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q VPWR VGND sg13g2_dlhq_1
Xoutput213 Inst_LUT4AB_switch_matrix.N1BEG0 N1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput268 Inst_LUT4AB_switch_matrix.S1BEG3 S1BEG[3] VPWR VGND sg13g2_buf_1
X_2703_ net1117 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q VPWR VGND sg13g2_dlhq_1
X_3117_ net1124 net189 VPWR VGND sg13g2_buf_1
X_2496_ net1158 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
Xoutput279 net279 S2BEGb[2] VPWR VGND sg13g2_buf_1
X_1378_ _0047_ VPWR _0048_ VGND _0044_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q sg13g2_o21ai_1
X_1447_ _0115_ net993 net964 VPWR VGND sg13g2_nand2b_1
X_3048_ UserCLK net370 _0001_ _3048_/Q_N Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
X_3048__370 VPWR VGND net370 sg13g2_tiehi
XFILLER_23_232 VPWR VGND sg13g2_fill_1
XFILLER_11_438 VPWR VGND sg13g2_fill_1
XFILLER_46_346 VPWR VGND sg13g2_fill_2
X_2281_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q _0904_ _0905_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q
+ sg13g2_a21oi_1
X_2350_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q _0964_ _0965_ VPWR VGND sg13g2_nor2_1
XFILLER_29_4 VPWR VGND sg13g2_fill_2
X_1301_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q net975 net944 net939 net962 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ _1130_ VPWR VGND sg13g2_mux4_1
X_1232_ VPWR _1064_ net383 VGND sg13g2_inv_1
X_1996_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q _0643_ _0644_ VPWR VGND sg13g2_nor2_1
XFILLER_20_202 VPWR VGND sg13g2_fill_1
XFILLER_20_224 VPWR VGND sg13g2_decap_8
X_2548_ net1196 net1079 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
X_2617_ net1181 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2479_ net1117 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_327 VPWR VGND sg13g2_fill_2
XFILLER_36_390 VPWR VGND sg13g2_fill_2
Xfanout1202 net1203 net1202 VPWR VGND sg13g2_buf_1
Xfanout1213 E6END[0] net1213 VPWR VGND sg13g2_buf_1
XFILLER_46_165 VPWR VGND sg13g2_fill_2
XFILLER_46_143 VPWR VGND sg13g2_fill_1
X_1850_ _0502_ VPWR _0503_ VGND net996 net942 sg13g2_o21ai_1
X_1781_ VGND VPWR _0436_ _0437_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_switch_matrix.M_AD
+ sg13g2_a21oi_2
X_2333_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q _0308_ _0950_ _0949_ sg13g2_a21oi_1
X_2402_ _0990_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q net927 VPWR VGND sg13g2_nand2b_1
X_1215_ VPWR _1048_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VGND sg13g2_inv_1
X_2264_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q _1157_ _0890_ _0889_
+ sg13g2_a21oi_1
X_2195_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0827_ _0830_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q
+ sg13g2_a21oi_1
XFILLER_52_179 VPWR VGND sg13g2_fill_2
XFILLER_37_187 VPWR VGND sg13g2_decap_8
X_1979_ net378 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0565_ _0628_ VPWR VGND sg13g2_mux4_1
X_3052__366 VPWR VGND net366 sg13g2_tiehi
Xhold23 Inst_LE_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net396 sg13g2_dlygate4sd3_1
XFILLER_45_99 VPWR VGND sg13g2_fill_1
XFILLER_28_143 VPWR VGND sg13g2_decap_4
Xfanout1076 FrameStrobe[16] net1076 VPWR VGND sg13g2_buf_1
Xfanout1098 net1099 net1098 VPWR VGND sg13g2_buf_1
Xfanout1032 net1033 net1032 VPWR VGND sg13g2_buf_1
Xfanout1087 net1092 net1087 VPWR VGND sg13g2_buf_1
Xfanout1021 net1022 net1021 VPWR VGND sg13g2_buf_1
Xfanout1010 net31 net1010 VPWR VGND sg13g2_buf_1
Xfanout1065 FrameStrobe[18] net1065 VPWR VGND sg13g2_buf_1
Xfanout1043 net1046 net1043 VPWR VGND sg13g2_buf_1
Xfanout1054 net1055 net1054 VPWR VGND sg13g2_buf_1
X_1902_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q VPWR _0553_ VGND _1026_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ sg13g2_o21ai_1
XFILLER_34_179 VPWR VGND sg13g2_fill_2
XFILLER_34_113 VPWR VGND sg13g2_fill_2
X_2951_ net1207 net1048 Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VPWR VGND sg13g2_dlhq_1
X_1833_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q _0307_ _0309_ _0290_ _0286_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
+ _0487_ VPWR VGND sg13g2_mux4_1
X_1764_ _0419_ VPWR _0420_ VGND _1012_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q sg13g2_o21ai_1
X_2882_ net1152 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_57_216 VPWR VGND sg13g2_fill_1
X_1695_ _0354_ _1031_ _0353_ VPWR VGND sg13g2_nand2_1
X_2316_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q _1084_ _0935_ _0934_
+ sg13g2_a21oi_1
X_3296_ W6END[10] net348 VPWR VGND sg13g2_buf_1
X_2247_ _0874_ VPWR _0875_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q _0556_ sg13g2_o21ai_1
X_2178_ net91 net107 net995 _0814_ VPWR VGND sg13g2_mux2_1
XFILLER_40_127 VPWR VGND sg13g2_fill_2
XFILLER_31_68 VPWR VGND sg13g2_fill_1
XFILLER_56_43 VPWR VGND sg13g2_fill_1
Xinput102 W2MID[4] net102 VPWR VGND sg13g2_buf_1
XFILLER_56_87 VPWR VGND sg13g2_fill_2
XFILLER_8_367 VPWR VGND sg13g2_fill_2
X_3150_ net1025 net210 VPWR VGND sg13g2_buf_1
X_1480_ Inst_LUT4AB_switch_matrix.E2BEG4 _0140_ _0146_ _0132_ _0138_ VPWR VGND sg13g2_a22oi_1
X_3081_ net20 net131 VPWR VGND sg13g2_buf_1
X_2032_ _0676_ _0677_ _0678_ VPWR VGND sg13g2_nor2_1
X_2101_ _0742_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q net108 VPWR VGND sg13g2_nand2b_1
X_2865_ net1206 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q VPWR VGND sg13g2_dlhq_1
X_2934_ net1189 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2796_ net1126 net30 Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1747_ net985 net955 _0404_ VPWR VGND sg13g2_nor2_2
XFILLER_7_70 VPWR VGND sg13g2_fill_1
X_1816_ _0470_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q _0334_ VPWR VGND sg13g2_nand2_1
X_1678_ _0337_ VPWR _0338_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q _0329_ sg13g2_o21ai_1
X_3279_ Inst_LUT4AB_switch_matrix.JW2BEG7 net329 VPWR VGND sg13g2_buf_1
XFILLER_45_219 VPWR VGND sg13g2_fill_1
XFILLER_26_411 VPWR VGND sg13g2_fill_1
XFILLER_26_57 VPWR VGND sg13g2_fill_2
XFILLER_26_35 VPWR VGND sg13g2_fill_1
XFILLER_9_109 VPWR VGND sg13g2_fill_1
XFILLER_32_458 VPWR VGND sg13g2_fill_1
X_2581_ net1194 net1083 Inst_LH_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_1601_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q VPWR _0264_ VGND _1013_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ sg13g2_o21ai_1
X_1532_ _0193_ VPWR _0196_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q _0195_ sg13g2_o21ai_1
X_2650_ net1177 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q VPWR VGND sg13g2_dlhq_1
X_3202_ NN4END[7] net258 VPWR VGND sg13g2_buf_1
X_3133_ net1166 net175 VPWR VGND sg13g2_buf_1
X_1394_ _0064_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 net982 VPWR
+ VGND sg13g2_nand2_1
X_1463_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q net37 net8 net65 net110 Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q
+ _0130_ VPWR VGND sg13g2_mux4_1
X_2015_ VPWR _0663_ _0662_ VGND sg13g2_inv_1
XFILLER_50_222 VPWR VGND sg13g2_fill_2
XFILLER_50_211 VPWR VGND sg13g2_fill_1
X_3064_ Inst_LUT4AB_switch_matrix.E1BEG1 net114 VPWR VGND sg13g2_buf_1
X_2848_ net1157 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2917_ net1138 net1038 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q VPWR VGND sg13g2_dlhq_1
X_2779_ net1173 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_2_307 VPWR VGND sg13g2_fill_2
XFILLER_14_436 VPWR VGND sg13g2_fill_2
XFILLER_1_362 VPWR VGND sg13g2_fill_1
X_2702_ net1121 net1107 Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q VPWR VGND sg13g2_dlhq_1
Xoutput203 net203 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_2564_ net1145 net1081 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_59_108 VPWR VGND sg13g2_fill_2
Xoutput247 net247 N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput258 net258 NN4BEG[3] VPWR VGND sg13g2_buf_1
X_1515_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VPWR _0180_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ _0177_ sg13g2_o21ai_1
Xoutput225 net225 N2BEGb[0] VPWR VGND sg13g2_buf_1
X_2633_ net1141 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VPWR VGND sg13g2_dlhq_1
Xoutput236 net236 N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput214 net214 N1BEG[1] VPWR VGND sg13g2_buf_1
X_2495_ net1161 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
Xoutput269 net269 S2BEG[0] VPWR VGND sg13g2_buf_1
X_3116_ net1127 net188 VPWR VGND sg13g2_buf_1
XFILLER_55_325 VPWR VGND sg13g2_fill_1
XFILLER_55_303 VPWR VGND sg13g2_fill_1
X_1377_ _0045_ _0046_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q _0047_ VPWR VGND sg13g2_nand3_1
X_1446_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0111_ _0114_ _0113_ sg13g2_a21oi_1
X_3047_ UserCLK net371 _0000_ _3047_/Q_N Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
XFILLER_23_200 VPWR VGND sg13g2_decap_4
XFILLER_14_233 VPWR VGND sg13g2_fill_1
XFILLER_14_255 VPWR VGND sg13g2_fill_1
X_2280_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q net971 _0904_ _0903_ sg13g2_a21oi_1
X_1300_ _1128_ VPWR _1129_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _1126_ sg13g2_o21ai_1
X_1231_ _1056_ VPWR Inst_LUT4AB_switch_matrix.E2BEG1 VGND _1058_ _1063_ sg13g2_o21ai_1
X_1995_ _0520_ _0525_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q _0643_ VPWR VGND sg13g2_mux2_1
X_2616_ net1184 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2547_ net1199 net1077 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
X_1429_ _0073_ VPWR _0098_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0081_ sg13g2_o21ai_1
X_2478_ net1121 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_55_166 VPWR VGND sg13g2_fill_1
XFILLER_55_111 VPWR VGND sg13g2_fill_2
XFILLER_28_347 VPWR VGND sg13g2_fill_1
XFILLER_28_303 VPWR VGND sg13g2_fill_2
XFILLER_11_247 VPWR VGND sg13g2_decap_4
Xfanout1214 net5 net1214 VPWR VGND sg13g2_buf_1
XFILLER_59_87 VPWR VGND sg13g2_fill_2
Xfanout1203 FrameData[11] net1203 VPWR VGND sg13g2_buf_1
XFILLER_19_325 VPWR VGND sg13g2_decap_4
X_1780_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q VPWR _0436_ VGND net984 net933 sg13g2_o21ai_1
XFILLER_57_409 VPWR VGND sg13g2_fill_1
X_2332_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q net943 _0949_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_295 VPWR VGND sg13g2_fill_2
X_2401_ _0989_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q net925 VPWR VGND sg13g2_nand2_1
X_1214_ VPWR _1047_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q VGND sg13g2_inv_1
X_2263_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q net932 _0889_ VPWR VGND sg13g2_nor2_1
X_2194_ VGND VPWR net52 net1001 _0829_ _0828_ sg13g2_a21oi_1
X_1978_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q _0617_ _0622_ _0626_ _0624_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q
+ _0627_ VPWR VGND sg13g2_mux4_1
Xhold24 Inst_LH_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net397 sg13g2_dlygate4sd3_1
XFILLER_28_122 VPWR VGND sg13g2_fill_1
XFILLER_43_158 VPWR VGND sg13g2_fill_2
XFILLER_43_125 VPWR VGND sg13g2_fill_1
XFILLER_43_114 VPWR VGND sg13g2_fill_2
XFILLER_31_309 VPWR VGND sg13g2_decap_8
Xfanout1022 net30 net1022 VPWR VGND sg13g2_buf_1
Xfanout1011 FrameStrobe[9] net1011 VPWR VGND sg13g2_buf_1
Xfanout1000 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q net1000 VPWR VGND sg13g2_buf_1
XFILLER_3_276 VPWR VGND sg13g2_fill_1
XFILLER_59_291 VPWR VGND sg13g2_fill_1
Xfanout1077 net1078 net1077 VPWR VGND sg13g2_buf_1
Xfanout1044 net1046 net1044 VPWR VGND sg13g2_buf_1
Xfanout1088 net1089 net1088 VPWR VGND sg13g2_buf_1
Xfanout1055 net1058 net1055 VPWR VGND sg13g2_buf_1
Xfanout1099 net1100 net1099 VPWR VGND sg13g2_buf_1
Xfanout1033 net1034 net1033 VPWR VGND sg13g2_buf_1
Xfanout1066 net1067 net1066 VPWR VGND sg13g2_buf_1
X_1901_ _0545_ _0552_ Inst_LUT4AB_switch_matrix.JS2BEG6 VPWR VGND sg13g2_nor2_2
X_1832_ _0486_ _0485_ VPWR VGND _0483_ sg13g2_nand2b_2
XFILLER_30_364 VPWR VGND sg13g2_fill_1
X_2950_ net1135 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q VPWR VGND sg13g2_dlhq_1
X_2881_ net1155 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_309 VPWR VGND sg13g2_fill_1
X_1694_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q net38 net54 net3 net9 Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ _0353_ VPWR VGND sg13g2_mux4_1
XFILLER_30_386 VPWR VGND sg13g2_fill_1
X_1763_ _0419_ net83 Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VPWR VGND sg13g2_nand2_1
X_2315_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q net954 _0934_ VPWR VGND sg13g2_nor2b_1
X_2246_ _0874_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q _0023_ VPWR VGND sg13g2_nand2_1
XFILLER_32_0 VPWR VGND sg13g2_fill_2
X_3295_ W6END[9] net347 VPWR VGND sg13g2_buf_1
XFILLER_38_453 VPWR VGND sg13g2_fill_2
X_2177_ VGND VPWR net64 net994 _0813_ _0812_ sg13g2_a21oi_1
XFILLER_33_191 VPWR VGND sg13g2_decap_8
Xinput103 W2MID[5] net103 VPWR VGND sg13g2_buf_1
X_3080_ net19 net130 VPWR VGND sg13g2_buf_1
X_2100_ _0741_ _0740_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VPWR VGND sg13g2_nand2b_1
XFILLER_54_209 VPWR VGND sg13g2_fill_2
X_2031_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0199_ _0677_ VPWR VGND sg13g2_mux4_1
X_2933_ net1192 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2795_ net1129 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2864_ net1116 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1815_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q _0315_ _0469_ _0468_ sg13g2_a21oi_1
X_1746_ _0403_ _0402_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR VGND sg13g2_nand2b_1
XFILLER_7_60 VPWR VGND sg13g2_fill_2
X_1677_ _0337_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q _0334_ VPWR VGND sg13g2_nand2_1
X_2229_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q _0308_ _0860_ _0859_
+ sg13g2_a21oi_1
X_3278_ Inst_LUT4AB_switch_matrix.JW2BEG6 net328 VPWR VGND sg13g2_buf_8
XFILLER_41_448 VPWR VGND sg13g2_fill_2
X_2580_ net1196 net1083 Inst_LH_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
X_1600_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q VPWR _0263_ VGND _0261_ _0262_ sg13g2_o21ai_1
X_1531_ _0194_ VPWR _0195_ VGND _1021_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q sg13g2_o21ai_1
XFILLER_4_360 VPWR VGND sg13g2_fill_2
X_1462_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q net53 net8 net97 Inst_LUT4AB_switch_matrix.E2BEG2
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q _0129_ VPWR VGND sg13g2_mux4_1
X_3201_ NN4END[6] net257 VPWR VGND sg13g2_buf_1
X_3132_ net1169 net174 VPWR VGND sg13g2_buf_1
X_1393_ VGND VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _1121_
+ _0063_ _1085_ sg13g2_a21oi_1
X_3063_ Inst_LUT4AB_switch_matrix.E1BEG0 net113 VPWR VGND sg13g2_buf_1
X_2014_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ net379 _0662_ VPWR VGND sg13g2_mux4_1
XFILLER_50_234 VPWR VGND sg13g2_fill_1
X_2778_ net1179 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q VPWR VGND sg13g2_dlhq_1
X_2847_ net1160 net1027 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2916_ net1146 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1729_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0384_ _0387_ _0386_ sg13g2_a21oi_1
XFILLER_41_223 VPWR VGND sg13g2_fill_2
XFILLER_26_297 VPWR VGND sg13g2_decap_8
XFILLER_17_253 VPWR VGND sg13g2_fill_2
X_2632_ net1176 net1097 Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2701_ net1124 net1105 Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q VPWR VGND sg13g2_dlhq_1
Xoutput204 net204 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput259 net259 NN4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput248 net248 N4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput226 net226 N2BEGb[1] VPWR VGND sg13g2_buf_1
X_2563_ net1148 net1081 Inst_LG_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
X_1514_ _0178_ VPWR _0179_ VGND net989 net936 sg13g2_o21ai_1
Xoutput237 net237 N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput215 Inst_LUT4AB_switch_matrix.N1BEG2 N1BEG[2] VPWR VGND sg13g2_buf_1
X_2494_ net1163 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
X_1445_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VPWR _0113_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ _0112_ sg13g2_o21ai_1
X_3115_ net1129 net187 VPWR VGND sg13g2_buf_1
X_1376_ _0046_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q net99 VPWR VGND sg13g2_nand2_1
X_3046_ net1137 net1110 Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_245 VPWR VGND sg13g2_decap_8
XFILLER_46_348 VPWR VGND sg13g2_fill_1
X_1230_ _1062_ _1060_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q _1063_ VPWR VGND sg13g2_a21o_1
X_1994_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q _0527_ _0642_ _0641_ sg13g2_a21oi_1
X_2615_ net1187 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2546_ net1202 net1079 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
X_1428_ _0091_ _0096_ _0097_ VPWR VGND sg13g2_and2_1
X_2477_ net1124 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_36_392 VPWR VGND sg13g2_fill_1
X_1359_ net67 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0030_ VPWR VGND sg13g2_nor2_1
X_3029_ net1192 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_35 VPWR VGND sg13g2_fill_2
XFILLER_50_24 VPWR VGND sg13g2_fill_1
Xfanout1204 FrameData[10] net1204 VPWR VGND sg13g2_buf_1
XFILLER_46_167 VPWR VGND sg13g2_fill_1
XFILLER_46_101 VPWR VGND sg13g2_fill_1
Xfanout1215 net4 net1215 VPWR VGND sg13g2_buf_1
XFILLER_19_348 VPWR VGND sg13g2_decap_4
X_2400_ _0975_ VPWR _0000_ VGND _0988_ _0987_ sg13g2_o21ai_1
X_1213_ VPWR _1046_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VGND sg13g2_inv_1
X_2331_ _0946_ _0947_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q _0948_ VPWR VGND sg13g2_nand3_1
X_2262_ _0197_ _0316_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q _0888_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_37_134 VPWR VGND sg13g2_decap_4
XFILLER_25_318 VPWR VGND sg13g2_decap_8
X_2193_ net1001 net36 _0828_ VPWR VGND sg13g2_nor2b_1
X_1977_ VPWR _0626_ _0625_ VGND sg13g2_inv_1
X_2529_ net1154 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_56_454 VPWR VGND sg13g2_fill_1
XFILLER_28_178 VPWR VGND sg13g2_fill_2
Xfanout1023 net1024 net1023 VPWR VGND sg13g2_buf_1
Xfanout1045 net1046 net1045 VPWR VGND sg13g2_buf_1
Xfanout1056 net1058 net1056 VPWR VGND sg13g2_buf_1
Xfanout1012 FrameStrobe[9] net1012 VPWR VGND sg13g2_buf_1
Xfanout1034 net29 net1034 VPWR VGND sg13g2_buf_1
Xfanout1001 net1002 net1001 VPWR VGND sg13g2_buf_1
XFILLER_47_432 VPWR VGND sg13g2_fill_1
Xfanout1078 net1079 net1078 VPWR VGND sg13g2_buf_1
Xfanout1089 net1091 net1089 VPWR VGND sg13g2_buf_1
Xfanout1067 net1068 net1067 VPWR VGND sg13g2_buf_1
X_1900_ VGND VPWR _0551_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q _0550_ _1044_ _0552_
+ _0546_ sg13g2_a221oi_1
X_1831_ _0484_ VPWR _0485_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q _0276_ sg13g2_o21ai_1
X_2880_ net1156 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1693_ _0351_ VPWR _0352_ VGND _1031_ _0350_ sg13g2_o21ai_1
X_1762_ Inst_LUT4AB_switch_matrix.JW2BEG2 _0417_ _0418_ _0403_ _0410_ VPWR VGND sg13g2_a22oi_1
X_2314_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q _0529_ _0933_ _0932_
+ sg13g2_a21oi_1
X_2245_ _0872_ VPWR _0873_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q net967 sg13g2_o21ai_1
XFILLER_25_0 VPWR VGND sg13g2_fill_2
X_3294_ W6END[8] net346 VPWR VGND sg13g2_buf_1
X_2176_ net995 net1210 _0812_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_129 VPWR VGND sg13g2_fill_1
XFILLER_15_49 VPWR VGND sg13g2_fill_2
XFILLER_21_310 VPWR VGND sg13g2_fill_1
Xinput104 W2MID[6] net104 VPWR VGND sg13g2_buf_1
XFILLER_8_369 VPWR VGND sg13g2_fill_1
X_2030_ _0676_ _0672_ _0675_ _0208_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_a22oi_1
X_2932_ net1197 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q VPWR VGND sg13g2_dlhq_1
X_2794_ net1132 net1024 Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_30_173 VPWR VGND sg13g2_decap_4
X_2863_ net1119 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1745_ net985 net975 net968 net944 net961 Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0402_ VPWR VGND sg13g2_mux4_1
X_1814_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q _0316_ _0468_ VPWR VGND sg13g2_nor2_1
XFILLER_7_391 VPWR VGND sg13g2_fill_1
X_1676_ _0335_ VPWR _0336_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q _0316_ sg13g2_o21ai_1
XFILLER_38_251 VPWR VGND sg13g2_decap_8
X_2228_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q net939 _0859_ VPWR VGND sg13g2_nor2b_1
X_2159_ net994 net955 _0795_ VPWR VGND sg13g2_nor2b_1
X_3277_ net377 net327 VPWR VGND sg13g2_buf_1
XFILLER_13_107 VPWR VGND sg13g2_fill_2
XFILLER_3_19 VPWR VGND sg13g2_fill_2
XFILLER_32_91 VPWR VGND sg13g2_decap_4
XFILLER_8_111 VPWR VGND sg13g2_fill_2
X_3200_ NN4END[5] net256 VPWR VGND sg13g2_buf_1
X_1530_ _0194_ net18 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q VPWR VGND sg13g2_nand2_1
X_1392_ _0062_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _1121_ VPWR
+ VGND sg13g2_nand2b_1
X_1461_ VGND VPWR _0122_ _0128_ Inst_LUT4AB_switch_matrix.E2BEG2 _0120_ sg13g2_a21oi_1
X_2013_ _0645_ net381 _0660_ _0661_ VPWR VGND sg13g2_a21o_1
X_3131_ net1172 net173 VPWR VGND sg13g2_buf_1
X_2915_ net1149 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1728_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR _0386_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0385_ sg13g2_o21ai_1
X_2777_ net1182 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2846_ net1163 net1030 Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_2_309 VPWR VGND sg13g2_fill_1
XFILLER_58_324 VPWR VGND sg13g2_fill_1
X_1659_ _0319_ VPWR _0320_ VGND _0317_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q sg13g2_o21ai_1
XFILLER_58_379 VPWR VGND sg13g2_fill_2
XFILLER_5_114 VPWR VGND sg13g2_fill_1
XFILLER_32_268 VPWR VGND sg13g2_fill_1
Xoutput205 net205 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_2562_ net1151 net1079 Inst_LG_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
Xoutput216 Inst_LUT4AB_switch_matrix.N1BEG3 N1BEG[3] VPWR VGND sg13g2_buf_1
X_2631_ net1208 net1097 Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2700_ net1126 net1105 Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q VPWR VGND sg13g2_dlhq_1
Xoutput249 net249 NN4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput238 net238 N4BEG[14] VPWR VGND sg13g2_buf_1
X_1513_ _0178_ net989 net928 VPWR VGND sg13g2_nand2b_1
Xoutput227 net227 N2BEGb[2] VPWR VGND sg13g2_buf_1
X_2493_ net1166 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
X_1375_ _0045_ net72 Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q VPWR VGND sg13g2_nand2b_1
X_1444_ net957 net952 net993 _0112_ VPWR VGND sg13g2_mux2_1
X_3114_ net1133 net186 VPWR VGND sg13g2_buf_1
X_3045_ net1139 net1110 Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q VPWR VGND sg13g2_dlhq_1
X_2829_ net1124 net1030 Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q VPWR VGND sg13g2_dlhq_1
XFILLER_58_121 VPWR VGND sg13g2_fill_2
X_1993_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q VPWR _0641_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q
+ _0528_ sg13g2_o21ai_1
XFILLER_20_249 VPWR VGND sg13g2_fill_2
XFILLER_55_0 VPWR VGND sg13g2_fill_2
X_2545_ net1205 net1077 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
X_2614_ net1190 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1358_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0028_ _0029_ VPWR VGND sg13g2_nor2b_1
X_1427_ _0073_ _0092_ _0093_ _0095_ _0096_ VPWR VGND sg13g2_or4_1
XFILLER_18_38 VPWR VGND sg13g2_fill_2
X_2476_ net1128 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
X_3028_ net1195 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q VPWR VGND sg13g2_dlhq_1
X_1289_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q net58 net108 net82 Inst_LUT4AB_switch_matrix.JN2BEG1
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q _1118_ VPWR VGND sg13g2_mux4_1
Xfanout1216 net3 net1216 VPWR VGND sg13g2_buf_1
Xfanout1205 FrameData[10] net1205 VPWR VGND sg13g2_buf_1
XFILLER_46_113 VPWR VGND sg13g2_fill_2
XFILLER_6_297 VPWR VGND sg13g2_fill_1
X_2330_ _0947_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q _0130_ VPWR VGND sg13g2_nand2b_1
X_1212_ VPWR _1045_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VGND sg13g2_inv_1
X_2192_ net1214 net7 net1002 _0827_ VPWR VGND sg13g2_mux2_1
X_2261_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q _0886_ _0887_ VPWR VGND sg13g2_nor2_1
XFILLER_18_360 VPWR VGND sg13g2_fill_1
X_1976_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q net36 net64 net25 net91 Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q
+ _0625_ VPWR VGND sg13g2_mux4_1
X_2528_ net1158 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_43_116 VPWR VGND sg13g2_fill_1
X_2459_ net1172 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_24_330 VPWR VGND sg13g2_decap_4
Xfanout1079 FrameStrobe[15] net1079 VPWR VGND sg13g2_buf_1
Xfanout1057 net1058 net1057 VPWR VGND sg13g2_buf_1
Xfanout1024 net1025 net1024 VPWR VGND sg13g2_buf_1
Xfanout1035 net1036 net1035 VPWR VGND sg13g2_buf_1
Xfanout1013 net1014 net1013 VPWR VGND sg13g2_buf_1
Xfanout1046 FrameStrobe[3] net1046 VPWR VGND sg13g2_buf_1
Xfanout1068 FrameStrobe[17] net1068 VPWR VGND sg13g2_buf_1
Xfanout1002 Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q net1002 VPWR VGND sg13g2_buf_1
XFILLER_34_149 VPWR VGND sg13g2_fill_1
XFILLER_34_127 VPWR VGND sg13g2_fill_1
XFILLER_42_160 VPWR VGND sg13g2_fill_1
X_1830_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q _0277_ _0484_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q
+ sg13g2_a21oi_1
X_1761_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q _0415_ _0418_ VPWR VGND sg13g2_nor2_1
X_1692_ _0351_ _1031_ _0349_ VPWR VGND sg13g2_nand2b_1
X_2313_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q VPWR _0932_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ _0148_ sg13g2_o21ai_1
X_2244_ _0872_ _0276_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q VPWR VGND sg13g2_nand2_2
X_3293_ W6END[7] net345 VPWR VGND sg13g2_buf_1
X_2175_ _0810_ VPWR _0811_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0809_ sg13g2_o21ai_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
XFILLER_33_171 VPWR VGND sg13g2_fill_2
XFILLER_25_138 VPWR VGND sg13g2_fill_2
XFILLER_25_116 VPWR VGND sg13g2_decap_4
XFILLER_21_300 VPWR VGND sg13g2_fill_2
X_1959_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0607_ _0609_ _0608_ sg13g2_a21oi_1
Xinput105 W2MID[7] net105 VPWR VGND sg13g2_buf_1
XFILLER_8_304 VPWR VGND sg13g2_fill_1
XFILLER_8_326 VPWR VGND sg13g2_fill_2
XFILLER_12_377 VPWR VGND sg13g2_fill_1
X_2931_ net1198 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2793_ net1141 net1024 Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1813_ _0467_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ C VPWR VGND sg13g2_mux2_1
X_2862_ net1120 net1033 Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1744_ VGND VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 net926
+ _0401_ _0400_ sg13g2_a21oi_1
X_3276_ Inst_LUT4AB_switch_matrix.JW2BEG4 net326 VPWR VGND sg13g2_buf_1
X_1675_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q _0315_ _0335_ _1043_ sg13g2_a21oi_1
X_2089_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VPWR _0731_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ _0730_ sg13g2_o21ai_1
X_2227_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q _0171_ _0858_ _0857_
+ sg13g2_a21oi_1
X_2158_ _0794_ VPWR Inst_LUT4AB_switch_matrix.JS2BEG0 VGND _0785_ _0786_ sg13g2_o21ai_1
XFILLER_44_255 VPWR VGND sg13g2_fill_1
XFILLER_8_189 VPWR VGND sg13g2_fill_1
XFILLER_12_163 VPWR VGND sg13g2_fill_2
X_3130_ net1178 net171 VPWR VGND sg13g2_buf_1
XFILLER_4_384 VPWR VGND sg13g2_fill_1
XFILLER_4_362 VPWR VGND sg13g2_fill_1
X_1391_ _0061_ _0060_ _1160_ VPWR VGND sg13g2_nand2b_1
X_1460_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q _0127_ _0128_ VPWR VGND sg13g2_nor2_1
X_2012_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0649_ _0660_ VPWR VGND sg13g2_mux4_1
X_2845_ net1167 net1030 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2914_ net1152 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q VPWR VGND sg13g2_dlhq_1
X_1727_ net60 net68 net999 _0385_ VPWR VGND sg13g2_mux2_1
X_2776_ net1184 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1658_ _0319_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0318_ VPWR VGND sg13g2_nand2b_1
X_3259_ SS4END[12] net315 VPWR VGND sg13g2_buf_1
X_1589_ _0250_ _0251_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q _0252_ VPWR VGND sg13g2_nand3_1
XFILLER_53_36 VPWR VGND sg13g2_fill_1
XFILLER_26_277 VPWR VGND sg13g2_fill_2
XFILLER_17_255 VPWR VGND sg13g2_fill_1
XFILLER_17_277 VPWR VGND sg13g2_fill_1
Xoutput206 net206 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput228 net228 N2BEGb[3] VPWR VGND sg13g2_buf_1
X_1512_ net958 net954 net988 _0177_ VPWR VGND sg13g2_mux2_1
Xoutput239 Inst_LUT4AB_switch_matrix.N4BEG3 N4BEG[15] VPWR VGND sg13g2_buf_1
X_2561_ net1154 net1081 Inst_LG_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
Xoutput217 net217 N2BEG[0] VPWR VGND sg13g2_buf_1
X_2630_ net1137 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q VPWR VGND sg13g2_dlhq_1
X_2492_ net1169 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
X_3113_ net1141 net183 VPWR VGND sg13g2_buf_1
X_1374_ net44 net15 Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q _0044_ VPWR VGND sg13g2_mux2_1
X_1443_ _0110_ VPWR _0111_ VGND net993 net935 sg13g2_o21ai_1
XFILLER_48_380 VPWR VGND sg13g2_fill_2
X_3044_ net1144 net1110 Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_225 VPWR VGND sg13g2_decap_8
X_2828_ net1126 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_23_269 VPWR VGND sg13g2_decap_8
X_2759_ net1208 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_457 VPWR VGND sg13g2_fill_2
X_1992_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux VPWR _0640_ VGND _0638_ _0591_ sg13g2_o21ai_1
X_2544_ net1115 net1080 Inst_LF_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
X_2475_ net1131 net1067 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
X_2613_ net1193 net1092 Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q VPWR VGND sg13g2_dlhq_1
X_1357_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q net1008 net10 net39 net1212 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ _0028_ VPWR VGND sg13g2_mux4_1
X_1288_ Inst_LUT4AB_switch_matrix.JN2BEG1 _1110_ _1117_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
+ _1108_ VPWR VGND sg13g2_a22oi_1
X_1426_ _0094_ VPWR _0095_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0083_ sg13g2_o21ai_1
X_3027_ net1198 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q VPWR VGND sg13g2_dlhq_1
Xfanout1206 FrameData[10] net1206 VPWR VGND sg13g2_buf_1
Xfanout1217 net2 net1217 VPWR VGND sg13g2_buf_1
XFILLER_24_82 VPWR VGND sg13g2_fill_1
XFILLER_6_254 VPWR VGND sg13g2_fill_2
X_1211_ VPWR _1044_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VGND sg13g2_inv_1
X_2260_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q net1007 net1214 net1003 net975
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q _0886_ VPWR VGND sg13g2_mux4_1
X_2191_ _0825_ VPWR _0826_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0818_ sg13g2_o21ai_1
X_1975_ VPWR _0624_ _0623_ VGND sg13g2_inv_1
X_2527_ net1160 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
X_1409_ _0075_ _0074_ _0078_ VPWR VGND sg13g2_nor2b_1
X_2458_ net1178 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_36_180 VPWR VGND sg13g2_decap_4
X_2389_ _0390_ _0237_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0978_ VPWR VGND sg13g2_mux2_1
XFILLER_3_235 VPWR VGND sg13g2_fill_2
Xfanout1003 net89 net1003 VPWR VGND sg13g2_buf_1
XFILLER_47_401 VPWR VGND sg13g2_fill_1
Xfanout1058 FrameStrobe[1] net1058 VPWR VGND sg13g2_buf_1
Xfanout1014 net1015 net1014 VPWR VGND sg13g2_buf_1
Xfanout1025 net30 net1025 VPWR VGND sg13g2_buf_1
Xfanout1036 net29 net1036 VPWR VGND sg13g2_buf_1
Xfanout1069 net1070 net1069 VPWR VGND sg13g2_buf_1
Xfanout1047 net1049 net1047 VPWR VGND sg13g2_buf_1
XFILLER_19_60 VPWR VGND sg13g2_fill_2
XFILLER_15_320 VPWR VGND sg13g2_fill_2
X_1691_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q net960 net954 net936 net928 Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ _0350_ VPWR VGND sg13g2_mux4_1
X_1760_ _0417_ _0416_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR VGND sg13g2_nand2b_1
X_2312_ _0931_ _0930_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q Inst_LUT4AB_switch_matrix.EE4BEG1
+ VPWR VGND sg13g2_mux2_1
X_3292_ W6END[6] net344 VPWR VGND sg13g2_buf_1
XFILLER_38_434 VPWR VGND sg13g2_fill_2
X_2243_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q _0870_ _0871_ VPWR VGND sg13g2_nor2_1
X_2174_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0807_ _0810_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
+ sg13g2_a21oi_1
XFILLER_33_150 VPWR VGND sg13g2_fill_1
X_1958_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR _0608_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ _0605_ sg13g2_o21ai_1
X_1889_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q VPWR _0541_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ net933 sg13g2_o21ai_1
XFILLER_29_401 VPWR VGND sg13g2_fill_2
Xinput106 W6END[0] net106 VPWR VGND sg13g2_buf_1
XFILLER_56_297 VPWR VGND sg13g2_fill_2
XFILLER_24_172 VPWR VGND sg13g2_fill_2
XFILLER_21_83 VPWR VGND sg13g2_fill_1
XFILLER_50_418 VPWR VGND sg13g2_fill_2
XFILLER_50_407 VPWR VGND sg13g2_fill_2
X_2930_ net1201 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2861_ net1123 net1033 Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q VPWR VGND sg13g2_dlhq_1
XFILLER_30_186 VPWR VGND sg13g2_fill_1
X_1674_ _0333_ VPWR _0334_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q _0330_ sg13g2_o21ai_1
XFILLER_7_96 VPWR VGND sg13g2_fill_2
X_2792_ net1174 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VPWR VGND sg13g2_dlhq_1
XFILLER_7_371 VPWR VGND sg13g2_fill_2
X_1743_ _0203_ _0399_ _0400_ VPWR VGND _0202_ sg13g2_nand3b_1
X_1812_ _0466_ _0457_ _0463_ _0467_ VPWR VGND sg13g2_a21o_1
X_2226_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q VPWR _0857_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ net980 sg13g2_o21ai_1
X_3275_ Inst_LUT4AB_switch_matrix.JW2BEG3 net325 VPWR VGND sg13g2_buf_1
X_2088_ net59 net63 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q _0730_ VPWR VGND sg13g2_mux2_1
XFILLER_13_109 VPWR VGND sg13g2_fill_1
X_2157_ _0793_ VPWR _0794_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0787_ sg13g2_o21ai_1
XFILLER_42_38 VPWR VGND sg13g2_fill_2
XFILLER_44_278 VPWR VGND sg13g2_fill_1
XFILLER_8_113 VPWR VGND sg13g2_fill_1
X_1390_ _0059_ _0058_ _1085_ _0060_ VPWR VGND sg13g2_mux2_1
X_2011_ _0659_ _0654_ _0655_ _0658_ VPWR VGND sg13g2_and3_1
X_2844_ net1169 net1028 Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2913_ net1155 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1726_ _0383_ VPWR _0384_ VGND net1006 net999 sg13g2_o21ai_1
X_1588_ _0251_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q net95 VPWR VGND sg13g2_nand2_1
X_1657_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q net966 net953 net937 net928 Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0318_ VPWR VGND sg13g2_mux4_1
X_2775_ net1187 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q VPWR VGND sg13g2_dlhq_1
X_3258_ SS4END[11] net314 VPWR VGND sg13g2_buf_1
X_3189_ N4END[10] net245 VPWR VGND sg13g2_buf_1
X_2209_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q net939 net944 net963 net956 Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0843_ VPWR VGND sg13g2_mux4_1
XFILLER_1_333 VPWR VGND sg13g2_fill_1
XFILLER_27_82 VPWR VGND sg13g2_fill_2
Xoutput207 net207 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_1511_ _0175_ VPWR _0176_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0174_ sg13g2_o21ai_1
Xoutput218 net218 N2BEG[1] VPWR VGND sg13g2_buf_8
X_2560_ net1157 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
Xoutput229 net229 N2BEGb[4] VPWR VGND sg13g2_buf_1
X_2491_ net1172 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
X_1442_ _0110_ net993 net931 VPWR VGND sg13g2_nand2b_1
X_3112_ net1176 net172 VPWR VGND sg13g2_buf_1
X_1373_ _0039_ _0042_ _0043_ VPWR VGND sg13g2_nor2_1
X_3043_ net1147 net1112 Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q VPWR VGND sg13g2_dlhq_1
X_2758_ net1137 net1015 Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q VPWR VGND sg13g2_dlhq_1
X_2827_ net1131 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2689_ net1155 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1709_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q VPWR _0367_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
+ _0366_ sg13g2_o21ai_1
XFILLER_14_226 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_1
Xfanout990 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q net990 VPWR VGND sg13g2_buf_1
X_1991_ VGND VPWR _0639_ net387 _0591_ sg13g2_or2_1
X_2612_ net1195 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q VPWR VGND sg13g2_dlhq_1
X_2543_ net1118 net1078 Inst_LF_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_1425_ VGND VPWR _0094_ _0076_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sg13g2_or2_1
X_2474_ net1134 net1067 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
X_3026_ net1203 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_362 VPWR VGND sg13g2_fill_2
X_1356_ _0026_ VPWR _0027_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0024_ sg13g2_o21ai_1
X_1287_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q _1116_ _1117_ VPWR VGND sg13g2_nor2_1
XFILLER_34_39 VPWR VGND sg13g2_fill_1
XFILLER_59_69 VPWR VGND sg13g2_fill_1
Xfanout1207 net1209 net1207 VPWR VGND sg13g2_buf_1
XFILLER_19_318 VPWR VGND sg13g2_decap_8
XFILLER_19_329 VPWR VGND sg13g2_fill_2
X_1210_ VPWR _1043_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q VGND sg13g2_inv_1
X_2190_ _0824_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q _0825_ VPWR VGND sg13g2_nor2b_1
X_1974_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q net55 net90 net1213 Inst_LUT4AB_switch_matrix.JW2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q _0623_ VPWR VGND sg13g2_mux4_1
Xhold17 Inst_LG_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net390 sg13g2_dlygate4sd3_1
X_2526_ net1163 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_28_104 VPWR VGND sg13g2_fill_2
X_2457_ net1181 net1060 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
X_1408_ _0073_ VPWR _0077_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0076_ sg13g2_o21ai_1
X_2388_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _1104_ _0977_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ sg13g2_a21oi_1
XFILLER_56_435 VPWR VGND sg13g2_fill_1
XFILLER_36_192 VPWR VGND sg13g2_fill_2
X_1339_ _0011_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0009_ VPWR VGND sg13g2_nand2b_1
X_3009_ net1153 net1055 Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q VPWR VGND sg13g2_dlhq_1
Xfanout1004 net1005 net1004 VPWR VGND sg13g2_buf_1
Xfanout1015 FrameStrobe[9] net1015 VPWR VGND sg13g2_buf_1
Xfanout1026 net1028 net1026 VPWR VGND sg13g2_buf_1
Xfanout1048 net1049 net1048 VPWR VGND sg13g2_buf_1
Xfanout1037 FrameStrobe[4] net1037 VPWR VGND sg13g2_buf_1
Xfanout1059 net28 net1059 VPWR VGND sg13g2_buf_1
XFILLER_15_354 VPWR VGND sg13g2_fill_1
X_1690_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q net978 net973 net948 net967 Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ _0349_ VPWR VGND sg13g2_mux4_1
X_2311_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q net1007 net1214 net62 net978 Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ _0931_ VPWR VGND sg13g2_mux4_1
X_2242_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q net1009 net1216 net88 D Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ _0870_ VPWR VGND sg13g2_mux4_1
X_3291_ W6END[5] net343 VPWR VGND sg13g2_buf_1
X_2173_ VGND VPWR net36 net994 _0809_ _0808_ sg13g2_a21oi_1
XFILLER_18_181 VPWR VGND sg13g2_fill_1
X_1957_ _0606_ VPWR _0607_ VGND net70 net983 sg13g2_o21ai_1
XFILLER_21_335 VPWR VGND sg13g2_decap_4
XFILLER_21_379 VPWR VGND sg13g2_fill_2
X_1888_ net965 net958 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q _0540_ VPWR VGND sg13g2_mux2_1
X_2509_ net1125 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_56_59 VPWR VGND sg13g2_fill_2
Xinput107 W6END[1] net107 VPWR VGND sg13g2_buf_1
XFILLER_56_287 VPWR VGND sg13g2_fill_2
XFILLER_24_195 VPWR VGND sg13g2_fill_2
XFILLER_8_328 VPWR VGND sg13g2_fill_1
XFILLER_30_132 VPWR VGND sg13g2_fill_2
XFILLER_7_20 VPWR VGND sg13g2_fill_1
X_2791_ net1207 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2860_ net1126 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_15_162 VPWR VGND sg13g2_fill_1
X_1811_ _0464_ _0465_ _0203_ _0466_ VPWR VGND sg13g2_mux2_1
X_1673_ _0331_ _0332_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q _0333_ VPWR VGND sg13g2_nand3_1
X_1742_ _0399_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 net926 VPWR
+ VGND sg13g2_nand2b_1
X_2225_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q _0851_ _0852_ _0854_ _0856_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q
+ Inst_LUT4AB_switch_matrix.WW4BEG3 VPWR VGND sg13g2_mux4_1
X_3274_ Inst_LUT4AB_switch_matrix.JW2BEG2 net324 VPWR VGND sg13g2_buf_1
X_2087_ _0728_ VPWR _0729_ VGND net87 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q sg13g2_o21ai_1
X_2156_ VGND VPWR _0789_ _0792_ _0793_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q sg13g2_a21oi_1
X_2989_ net1123 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_165 VPWR VGND sg13g2_fill_2
X_2010_ _0645_ _0657_ net381 _0658_ VPWR VGND sg13g2_nand3_1
X_2912_ net1156 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1725_ _0383_ net999 net89 VPWR VGND sg13g2_nand2b_1
X_2774_ net1190 net1020 Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2843_ net1171 net1028 Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1587_ _0250_ net84 Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q VPWR VGND sg13g2_nand2b_1
X_1656_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q net977 net972 net942 net947 Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0317_ VPWR VGND sg13g2_mux4_1
X_3257_ SS4END[10] net313 VPWR VGND sg13g2_buf_1
X_3188_ N4END[9] net244 VPWR VGND sg13g2_buf_1
X_2208_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q net1215 net1004 net974 net969 Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0842_ VPWR VGND sg13g2_mux4_1
X_2139_ _0773_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q _0776_ _0777_ VPWR VGND sg13g2_a21o_1
XFILLER_41_249 VPWR VGND sg13g2_decap_4
XFILLER_26_279 VPWR VGND sg13g2_fill_1
XFILLER_22_452 VPWR VGND sg13g2_fill_2
XFILLER_40_293 VPWR VGND sg13g2_decap_8
XFILLER_40_260 VPWR VGND sg13g2_decap_8
XFILLER_9_456 VPWR VGND sg13g2_fill_2
XFILLER_13_430 VPWR VGND sg13g2_fill_1
XFILLER_13_452 VPWR VGND sg13g2_fill_2
Xoutput219 net219 N2BEG[2] VPWR VGND sg13g2_buf_8
Xoutput208 net208 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
X_1510_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q _0175_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ _0173_ sg13g2_a21oi_2
X_2490_ net1178 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_4_172 VPWR VGND sg13g2_fill_2
X_1441_ _0109_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ B VPWR VGND sg13g2_mux2_1
X_3111_ net1208 net161 VPWR VGND sg13g2_buf_1
X_1372_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q _0040_ _0041_ _0042_ VPWR VGND sg13g2_nor3_1
X_3042_ net1150 net1112 Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2757_ net1140 net1015 Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_282 VPWR VGND sg13g2_fill_2
X_1708_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q net58 net69 net12 net96 Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q
+ _0366_ VPWR VGND sg13g2_mux4_1
X_2688_ net1158 net1100 Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2826_ net1134 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q VPWR VGND sg13g2_dlhq_1
X_1639_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0299_ _0301_ _0300_ sg13g2_a21oi_1
X_3309_ WW4END[13] net365 VPWR VGND sg13g2_buf_1
Xfanout980 _0586_ net980 VPWR VGND sg13g2_buf_1
Xfanout991 Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q net991 VPWR VGND sg13g2_buf_1
X_1990_ VGND VPWR net378 _0488_ net374 net386 _0638_ _0490_ sg13g2_a221oi_1
XFILLER_13_260 VPWR VGND sg13g2_decap_4
X_2542_ net1121 net1081 Inst_LF_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
X_2611_ net1198 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1424_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0081_ _0093_ VPWR
+ VGND sg13g2_nor2_1
X_1355_ _0026_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0025_ VPWR VGND sg13g2_nand2b_1
X_2473_ net1143 net1067 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
X_3025_ net1204 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1286_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q _1114_ _1116_ _1115_ sg13g2_a21oi_1
X_2809_ net1180 net1025 Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_1_8 VPWR VGND sg13g2_fill_2
Xfanout1208 net1209 net1208 VPWR VGND sg13g2_buf_1
XFILLER_42_311 VPWR VGND sg13g2_fill_2
XFILLER_10_274 VPWR VGND sg13g2_fill_2
XFILLER_52_119 VPWR VGND sg13g2_fill_1
XFILLER_37_138 VPWR VGND sg13g2_fill_1
XFILLER_33_377 VPWR VGND sg13g2_fill_2
X_1973_ _0621_ VPWR _0622_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q _0618_ sg13g2_o21ai_1
XFILLER_53_0 VPWR VGND sg13g2_fill_2
X_2525_ net1166 net1073 Inst_LE_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
Xhold18 Inst_LD_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net391 sg13g2_dlygate4sd3_1
X_1338_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q net974 net944 net938 net962 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ _0010_ VPWR VGND sg13g2_mux4_1
X_2456_ net1184 net1060 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
X_1407_ _0076_ _0075_ _0074_ VPWR VGND sg13g2_nand2b_1
X_2387_ _0976_ net385 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VPWR VGND sg13g2_nand2b_1
XFILLER_45_39 VPWR VGND sg13g2_fill_2
X_1269_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q _1095_ _1096_ _1099_ _1097_ _1015_
+ _1100_ VPWR VGND sg13g2_mux4_1
X_3008_ net1156 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q VPWR VGND sg13g2_dlhq_1
Xfanout1016 net1020 net1016 VPWR VGND sg13g2_buf_1
Xfanout1005 W1END[2] net1005 VPWR VGND sg13g2_buf_1
XFILLER_3_237 VPWR VGND sg13g2_fill_1
Xfanout1027 net1028 net1027 VPWR VGND sg13g2_buf_1
Xfanout1038 FrameStrobe[4] net1038 VPWR VGND sg13g2_buf_1
XFILLER_47_458 VPWR VGND sg13g2_fill_1
Xfanout1049 FrameStrobe[2] net1049 VPWR VGND sg13g2_buf_1
XFILLER_34_108 VPWR VGND sg13g2_fill_1
XFILLER_19_62 VPWR VGND sg13g2_fill_1
XFILLER_19_73 VPWR VGND sg13g2_fill_1
XFILLER_19_95 VPWR VGND sg13g2_fill_1
XFILLER_27_193 VPWR VGND sg13g2_decap_8
X_2241_ _0868_ _0869_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q Inst_LUT4AB_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux2_1
X_2310_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q net937 _1157_ _0197_ _0239_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ _0930_ VPWR VGND sg13g2_mux4_1
X_3290_ W6END[4] net342 VPWR VGND sg13g2_buf_1
XFILLER_2_270 VPWR VGND sg13g2_fill_2
X_2172_ net994 net1007 _0808_ VPWR VGND sg13g2_nor2b_1
XFILLER_53_417 VPWR VGND sg13g2_fill_1
X_1956_ _0606_ net983 net1003 VPWR VGND sg13g2_nand2b_1
X_1887_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q net976 net971 net941 net946 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ _0539_ VPWR VGND sg13g2_mux4_1
X_2508_ net1127 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
Xinput108 WW4END[0] net108 VPWR VGND sg13g2_buf_1
XFILLER_56_299 VPWR VGND sg13g2_fill_1
XFILLER_56_222 VPWR VGND sg13g2_fill_2
XFILLER_56_200 VPWR VGND sg13g2_fill_1
XFILLER_44_406 VPWR VGND sg13g2_fill_2
XFILLER_29_458 VPWR VGND sg13g2_fill_1
XFILLER_29_447 VPWR VGND sg13g2_fill_1
XFILLER_29_403 VPWR VGND sg13g2_fill_1
X_2439_ net1209 net1060 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_24_130 VPWR VGND sg13g2_decap_4
XFILLER_21_41 VPWR VGND sg13g2_fill_2
XFILLER_50_409 VPWR VGND sg13g2_fill_1
XFILLER_35_417 VPWR VGND sg13g2_fill_2
XFILLER_30_199 VPWR VGND sg13g2_decap_4
XFILLER_7_54 VPWR VGND sg13g2_fill_2
X_1810_ _0202_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0395_ _0465_ VPWR VGND sg13g2_mux4_1
X_1741_ _0396_ _0397_ _0206_ _0398_ VPWR VGND sg13g2_nand3_1
X_2790_ net1136 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1672_ _0332_ net99 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VPWR VGND sg13g2_nand2_1
XFILLER_7_373 VPWR VGND sg13g2_fill_1
XFILLER_38_244 VPWR VGND sg13g2_decap_8
X_2224_ _0855_ VPWR _0856_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0556_
+ sg13g2_o21ai_1
XFILLER_26_19 VPWR VGND sg13g2_fill_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
X_2155_ _0791_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0792_ VPWR VGND sg13g2_nor2b_1
X_3273_ Inst_LUT4AB_switch_matrix.JW2BEG1 net323 VPWR VGND sg13g2_buf_1
XFILLER_53_258 VPWR VGND sg13g2_fill_2
X_2086_ _0728_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q net1004 VPWR VGND sg13g2_nand2b_1
X_1939_ VPWR _0589_ _0588_ VGND sg13g2_inv_1
X_2988_ net1126 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q VPWR VGND sg13g2_dlhq_1
Xinput90 W2END[0] net90 VPWR VGND sg13g2_buf_1
XFILLER_21_188 VPWR VGND sg13g2_decap_4
XFILLER_29_255 VPWR VGND sg13g2_fill_2
XFILLER_29_222 VPWR VGND sg13g2_fill_2
XFILLER_32_95 VPWR VGND sg13g2_fill_1
X_2911_ net1161 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2773_ net1194 net1018 Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q VPWR VGND sg13g2_dlhq_1
X_1724_ _0381_ VPWR _0382_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0380_ sg13g2_o21ai_1
X_2842_ net1178 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q VPWR VGND sg13g2_dlhq_1
X_3256_ SS4END[9] net312 VPWR VGND sg13g2_buf_1
X_1586_ net40 net11 Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q _0249_ VPWR VGND sg13g2_mux2_1
X_1655_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q net57 net7 net64 net91 Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q
+ _0316_ VPWR VGND sg13g2_mux4_1
X_3187_ N4END[8] net243 VPWR VGND sg13g2_buf_1
X_2207_ VGND VPWR _0840_ _0841_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0838_ sg13g2_a21oi_2
XFILLER_26_214 VPWR VGND sg13g2_fill_2
X_2138_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VPWR _0776_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ _0775_ sg13g2_o21ai_1
X_2069_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q net963 net951 net956 net930 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ _0712_ VPWR VGND sg13g2_mux4_1
XFILLER_32_217 VPWR VGND sg13g2_fill_1
XFILLER_9_424 VPWR VGND sg13g2_fill_1
Xoutput209 net209 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_1371_ net43 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q _0041_ VPWR VGND sg13g2_nor2_1
X_1440_ VGND VPWR _0108_ _0109_ _0085_ _0097_ sg13g2_a21oi_2
X_3041_ net1153 net1112 Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VPWR VGND sg13g2_dlhq_1
X_2825_ net1143 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q VPWR VGND sg13g2_dlhq_1
X_2756_ net1145 net1015 Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1638_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VPWR _0300_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0297_ sg13g2_o21ai_1
X_2687_ net1161 net1100 Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q VPWR VGND sg13g2_dlhq_1
X_1707_ VGND VPWR _0365_ _0364_ _0362_ sg13g2_or2_1
X_3239_ S4END[8] net295 VPWR VGND sg13g2_buf_1
X_1569_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0230_ _0232_ _0231_ sg13g2_a21oi_1
X_3308_ WW4END[12] net364 VPWR VGND sg13g2_buf_1
XFILLER_54_375 VPWR VGND sg13g2_fill_2
Xfanout992 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q net992 VPWR VGND sg13g2_buf_1
XFILLER_49_158 VPWR VGND sg13g2_fill_2
Xfanout981 _0586_ net981 VPWR VGND sg13g2_buf_1
Xfanout970 B net970 VPWR VGND sg13g2_buf_8
X_2610_ net1201 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2541_ net1125 net1078 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_2472_ net1175 net1067 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
X_1354_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q net955 net950 net934 net930 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ _0025_ VPWR VGND sg13g2_mux4_1
X_1285_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VPWR _1115_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ _1112_ sg13g2_o21ai_1
X_1423_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0078_ _0092_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_36_364 VPWR VGND sg13g2_fill_1
X_3024_ net1114 net1110 Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2808_ net1184 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2739_ net1199 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q VPWR VGND sg13g2_dlhq_1
Xfanout1209 FrameData[0] net1209 VPWR VGND sg13g2_buf_1
XFILLER_39_191 VPWR VGND sg13g2_fill_2
XFILLER_27_331 VPWR VGND sg13g2_fill_2
XFILLER_33_345 VPWR VGND sg13g2_fill_2
X_1972_ _0619_ _0620_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q _0621_ VPWR VGND sg13g2_nand3_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_2524_ net1169 net1073 Inst_LE_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_2455_ net1187 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
X_2386_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q net397 _0975_ VPWR VGND _0973_ sg13g2_nand3b_1
X_1337_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q net955 net950 net934 net928 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ _0009_ VPWR VGND sg13g2_mux4_1
X_1268_ VGND VPWR _1012_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1099_ _1098_ sg13g2_a21oi_1
X_1406_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q _1157_ _1159_ _1141_ _1140_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
+ _0075_ VPWR VGND sg13g2_mux4_1
Xhold19 Inst_LC_LUT4c_frame_config_dffesr.LUT_flop VPWR VGND net392 sg13g2_dlygate4sd3_1
XFILLER_51_164 VPWR VGND sg13g2_fill_2
XFILLER_24_334 VPWR VGND sg13g2_fill_1
X_1199_ VPWR _1032_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VGND sg13g2_inv_1
X_3007_ net1159 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_21 VPWR VGND sg13g2_fill_2
Xfanout1017 net1018 net1017 VPWR VGND sg13g2_buf_1
Xfanout1039 net1040 net1039 VPWR VGND sg13g2_buf_1
Xfanout1006 net88 net1006 VPWR VGND sg13g2_buf_1
Xfanout1028 FrameStrobe[6] net1028 VPWR VGND sg13g2_buf_1
XFILLER_10_87 VPWR VGND sg13g2_fill_2
XFILLER_15_312 VPWR VGND sg13g2_decap_4
XFILLER_19_106 VPWR VGND sg13g2_fill_2
XFILLER_42_131 VPWR VGND sg13g2_fill_1
X_2240_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q net953 _1084_ _0148_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ _0869_ VPWR VGND sg13g2_mux4_1
X_2171_ net52 net23 net995 _0807_ VPWR VGND sg13g2_mux2_1
X_1955_ net60 net62 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q _0605_ VPWR VGND sg13g2_mux2_1
X_1886_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q net56 net68 net11 net95 Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q
+ _0538_ VPWR VGND sg13g2_mux4_1
X_2507_ net1129 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
X_2438_ net1136 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
Xinput109 WW4END[1] net109 VPWR VGND sg13g2_buf_1
XFILLER_0_219 VPWR VGND sg13g2_fill_2
XFILLER_56_278 VPWR VGND sg13g2_fill_1
X_2369_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q net35 net54 net107 net951 Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ Inst_LUT4AB_switch_matrix.N4BEG2 VPWR VGND sg13g2_mux4_1
XFILLER_24_197 VPWR VGND sg13g2_fill_1
XFILLER_47_289 VPWR VGND sg13g2_fill_1
X_1671_ _0331_ net72 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VPWR VGND sg13g2_nand2b_1
XFILLER_7_352 VPWR VGND sg13g2_fill_2
X_1740_ _0397_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 net926 VPWR
+ VGND sg13g2_nand2b_1
X_3272_ Inst_LUT4AB_switch_matrix.JW2BEG0 net322 VPWR VGND sg13g2_buf_1
X_2085_ _0726_ VPWR _0727_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0724_ sg13g2_o21ai_1
X_2223_ _0855_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _1141_ VPWR VGND sg13g2_nand2_1
X_2154_ VGND VPWR _1028_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _0791_ _0790_ sg13g2_a21oi_1
XFILLER_42_19 VPWR VGND sg13g2_fill_2
XFILLER_34_440 VPWR VGND sg13g2_fill_2
X_2987_ net1131 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR VGND sg13g2_dlhq_1
Xinput80 S4END[1] net80 VPWR VGND sg13g2_buf_1
X_1938_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q net38 net83 net9 net93 Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q
+ _0588_ VPWR VGND sg13g2_mux4_1
X_1869_ net50 net21 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q _0521_ VPWR VGND sg13g2_mux2_1
Xinput91 W2END[1] net91 VPWR VGND sg13g2_buf_1
XFILLER_44_237 VPWR VGND sg13g2_fill_1
XFILLER_16_64 VPWR VGND sg13g2_fill_1
XFILLER_16_86 VPWR VGND sg13g2_fill_2
XFILLER_32_30 VPWR VGND sg13g2_decap_8
X_2910_ net1162 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q VPWR VGND sg13g2_dlhq_1
X_2841_ net1181 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VPWR VGND sg13g2_dlhq_1
X_1723_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0379_ _0381_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q
+ sg13g2_a21oi_1
X_2772_ net1197 net1018 Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_7_182 VPWR VGND sg13g2_fill_1
X_1654_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q _1040_ _1030_ _1022_ _0037_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q
+ _0315_ VPWR VGND sg13g2_mux4_1
X_3255_ SS4END[8] net311 VPWR VGND sg13g2_buf_1
X_2206_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q VPWR _0840_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
+ _0839_ sg13g2_o21ai_1
X_1585_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q net52 net84 net94 Inst_LUT4AB_switch_matrix.JS2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q _0248_ VPWR VGND sg13g2_mux4_1
X_3186_ N4END[7] net242 VPWR VGND sg13g2_buf_1
X_2068_ VGND VPWR _1046_ _0711_ Inst_LUT4AB_switch_matrix.JS2BEG7 _0704_ sg13g2_a21oi_1
XFILLER_26_237 VPWR VGND sg13g2_fill_2
X_2137_ VGND VPWR net80 net986 _0775_ _0774_ sg13g2_a21oi_1
XFILLER_22_454 VPWR VGND sg13g2_fill_1
XFILLER_13_410 VPWR VGND sg13g2_fill_2
XFILLER_9_458 VPWR VGND sg13g2_fill_1
XFILLER_4_78 VPWR VGND sg13g2_fill_2
X_1370_ net14 Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q _0040_ VPWR VGND sg13g2_nor2b_1
X_3040_ net1156 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_284 VPWR VGND sg13g2_fill_1
X_2824_ net1175 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q VPWR VGND sg13g2_dlhq_1
XFILLER_16_281 VPWR VGND sg13g2_decap_8
X_1637_ _0298_ VPWR _0299_ VGND net69 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q sg13g2_o21ai_1
X_2686_ net1162 net1100 Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1706_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q Inst_LUT4AB_switch_matrix.JN2BEG2
+ _0364_ _0363_ sg13g2_a21oi_1
X_2755_ net1147 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q VPWR VGND sg13g2_dlhq_1
X_3238_ S4END[7] net294 VPWR VGND sg13g2_buf_1
X_1568_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q VPWR _0231_ VGND net104 Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q
+ sg13g2_o21ai_1
X_1499_ net66 net82 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q _0165_ VPWR VGND sg13g2_mux2_1
X_3169_ Inst_LUT4AB_switch_matrix.JN2BEG2 net219 VPWR VGND sg13g2_buf_8
X_3307_ WW4END[11] net363 VPWR VGND sg13g2_buf_1
XFILLER_13_98 VPWR VGND sg13g2_fill_1
Xfanout960 F net960 VPWR VGND sg13g2_buf_1
Xfanout971 net972 net971 VPWR VGND sg13g2_buf_1
XFILLER_38_62 VPWR VGND sg13g2_decap_4
Xfanout982 _1121_ net982 VPWR VGND sg13g2_buf_8
Xfanout993 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q net993 VPWR VGND sg13g2_buf_1
X_2540_ net1127 net1077 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_2471_ net1209 net1067 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
X_1422_ VGND VPWR Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0089_ _0091_ _0090_ sg13g2_a21oi_1
X_1353_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q net974 net968 net938 net961 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ _0024_ VPWR VGND sg13g2_mux4_1
X_3023_ net1117 net1110 Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1284_ _1113_ VPWR _1114_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q net92 sg13g2_o21ai_1
XFILLER_51_302 VPWR VGND sg13g2_fill_2
X_2738_ net1202 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2807_ net1187 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_28 VPWR VGND sg13g2_fill_2
X_2669_ net1123 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1971_ _0620_ net99 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VPWR VGND sg13g2_nand2_1
X_2385_ _0974_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0973_ VPWR VGND sg13g2_nand2b_1
X_2523_ net1172 net1073 Inst_LE_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
X_2454_ net1190 net1061 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
X_1405_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q _1083_ _1084_ _1066_ _1065_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q
+ _0074_ VPWR VGND sg13g2_mux4_1
X_1198_ VPWR _1031_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VGND sg13g2_inv_1
XFILLER_28_118 VPWR VGND sg13g2_decap_4
X_1267_ net39 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1098_ VPWR VGND sg13g2_nor2_1
Xinput1 Ci net1 VPWR VGND sg13g2_buf_2
X_1336_ _1160_ _1162_ _0008_ VPWR VGND sg13g2_nor2_1
X_3006_ net1162 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_173 VPWR VGND sg13g2_decap_8
Xfanout1007 net34 net1007 VPWR VGND sg13g2_buf_1
Xfanout1018 net1020 net1018 VPWR VGND sg13g2_buf_1
Xfanout1029 net1030 net1029 VPWR VGND sg13g2_buf_1
Xoutput360 net360 WW4BEG[4] VPWR VGND sg13g2_buf_1
X_2170_ _0800_ _0805_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q _0806_ VPWR VGND sg13g2_nand3_1
X_1954_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q _0603_ _0604_ VPWR VGND sg13g2_and2_1
XFILLER_33_198 VPWR VGND sg13g2_decap_8
X_1885_ _0536_ VPWR _0537_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q _0533_ sg13g2_o21ai_1
X_2506_ net1133 net1074 Inst_LD_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
X_2437_ net1139 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
X_2368_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q net36 net106 net51 net935 Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ Inst_LUT4AB_switch_matrix.N4BEG3 VPWR VGND sg13g2_mux4_1
X_2299_ _0920_ VPWR _0921_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q net967
+ sg13g2_o21ai_1
X_1319_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1146_ _1147_ _1024_ sg13g2_a21oi_1
Xoutput190 net190 FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_46_51 VPWR VGND sg13g2_fill_1
X_1670_ net44 net15 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q _0330_ VPWR VGND sg13g2_mux2_1
X_2222_ VGND VPWR _0853_ _0854_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0276_
+ sg13g2_a21oi_2
XFILLER_38_268 VPWR VGND sg13g2_fill_2
X_2084_ _0726_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0725_ VPWR VGND sg13g2_nand2b_1
XFILLER_16_2 VPWR VGND sg13g2_fill_1
X_2153_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q VPWR _0790_ VGND net91 net991 sg13g2_o21ai_1
X_1937_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q net53 net92 net85 Inst_LUT4AB_switch_matrix.E2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q _0587_ VPWR VGND sg13g2_mux4_1
X_2986_ net1134 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q VPWR VGND sg13g2_dlhq_1
Xinput81 S4END[2] net81 VPWR VGND sg13g2_buf_1
Xinput70 S2END[7] net70 VPWR VGND sg13g2_buf_1
X_1868_ _0518_ VPWR _0520_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q _0519_ sg13g2_o21ai_1
Xinput92 W2END[2] net92 VPWR VGND sg13g2_buf_1
X_1799_ VPWR _0454_ _0453_ VGND sg13g2_inv_1
XFILLER_44_205 VPWR VGND sg13g2_fill_1
XFILLER_29_268 VPWR VGND sg13g2_fill_2
XFILLER_4_312 VPWR VGND sg13g2_fill_1
XFILLER_35_238 VPWR VGND sg13g2_fill_2
XFILLER_35_216 VPWR VGND sg13g2_fill_1
X_2771_ net1199 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2840_ net1184 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1722_ net32 net40 net999 _0380_ VPWR VGND sg13g2_mux2_1
X_1653_ _0313_ _0247_ _0314_ VPWR VGND sg13g2_nor2b_1
X_1584_ _0247_ _0246_ _0240_ VPWR VGND sg13g2_nand2_2
X_3185_ N4END[6] net241 VPWR VGND sg13g2_buf_1
X_3254_ SS4END[7] net310 VPWR VGND sg13g2_buf_1
Xfanout1190 net1191 net1190 VPWR VGND sg13g2_buf_1
X_2205_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q net953 net935 net931 net929 Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0839_ VPWR VGND sg13g2_mux4_1
XFILLER_53_19 VPWR VGND sg13g2_fill_2
XFILLER_26_249 VPWR VGND sg13g2_decap_8
X_2067_ VGND VPWR _1045_ _0705_ _0711_ _0710_ sg13g2_a21oi_1
X_2136_ net986 net64 _0774_ VPWR VGND sg13g2_nor2b_1
X_2969_ net1180 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_1_315 VPWR VGND sg13g2_fill_1
XFILLER_27_64 VPWR VGND sg13g2_fill_1
XFILLER_25_282 VPWR VGND sg13g2_fill_2
XFILLER_4_120 VPWR VGND sg13g2_fill_1
XFILLER_48_352 VPWR VGND sg13g2_fill_2
XFILLER_48_330 VPWR VGND sg13g2_fill_1
XFILLER_48_396 VPWR VGND sg13g2_fill_2
XFILLER_16_260 VPWR VGND sg13g2_decap_8
X_2823_ net1207 net1027 Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2754_ net1150 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q VPWR VGND sg13g2_dlhq_1
X_1705_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q VPWR _0363_ VGND _1023_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q
+ sg13g2_o21ai_1
X_1567_ Inst_LUT4AB_switch_matrix.JN2BEG5 _0230_ VPWR VGND sg13g2_inv_2
X_1636_ _0298_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q net1005 VPWR VGND sg13g2_nand2b_1
X_2685_ net1165 net1099 Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q VPWR VGND sg13g2_dlhq_1
X_3306_ WW4END[10] net362 VPWR VGND sg13g2_buf_1
X_3237_ S4END[6] net293 VPWR VGND sg13g2_buf_1
X_2119_ _0758_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0759_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_352 VPWR VGND sg13g2_fill_2
X_1498_ _0163_ VPWR _0164_ VGND net93 Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q sg13g2_o21ai_1
X_3168_ Inst_LUT4AB_switch_matrix.JN2BEG1 net218 VPWR VGND sg13g2_buf_8
XFILLER_54_377 VPWR VGND sg13g2_fill_1
X_3099_ EE4END[8] net155 VPWR VGND sg13g2_buf_1
XFILLER_14_219 VPWR VGND sg13g2_decap_8
Xfanout972 net973 net972 VPWR VGND sg13g2_buf_1
Xfanout983 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q net983 VPWR VGND sg13g2_buf_1
Xfanout950 net952 net950 VPWR VGND sg13g2_buf_1
Xfanout961 net963 net961 VPWR VGND sg13g2_buf_1
Xfanout994 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q net994 VPWR VGND sg13g2_buf_1
X_3054__372 VPWR VGND net372 sg13g2_tiehi
X_1421_ Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0086_ _0090_ VPWR VGND sg13g2_nor2b_1
X_2470_ net1136 net1064 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_48_193 VPWR VGND sg13g2_fill_2
XFILLER_36_311 VPWR VGND sg13g2_fill_1
X_1352_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q net35 net63 net6 net111 Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q
+ _0023_ VPWR VGND sg13g2_mux4_1
X_3022_ net1120 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1283_ _1113_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q net106 VPWR VGND sg13g2_nand2b_1
X_2806_ net1189 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2737_ net1204 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q VPWR VGND sg13g2_dlhq_1
X_2668_ net1128 net1102 Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1619_ VPWR _0281_ _0280_ VGND sg13g2_inv_1
X_2599_ net1207 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_355 VPWR VGND sg13g2_fill_2
XFILLER_27_333 VPWR VGND sg13g2_fill_1
XFILLER_40_20 VPWR VGND sg13g2_fill_2
XFILLER_2_454 VPWR VGND sg13g2_fill_1
XFILLER_6_248 VPWR VGND sg13g2_fill_1
XFILLER_49_51 VPWR VGND sg13g2_fill_1
XFILLER_45_185 VPWR VGND sg13g2_decap_4
XFILLER_45_163 VPWR VGND sg13g2_decap_4
X_1970_ _0619_ net72 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VPWR VGND sg13g2_nand2b_1
X_2522_ net1179 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_1335_ _1085_ _1161_ _1162_ VPWR VGND sg13g2_nor2_1
X_1404_ _0071_ VPWR _0073_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q _0072_
+ sg13g2_o21ai_1
X_2453_ net1193 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
X_2384_ _0971_ VPWR _0973_ VGND _0972_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q sg13g2_o21ai_1
X_3005_ net1165 net1055 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q VPWR VGND sg13g2_dlhq_1
X_1266_ net1215 net10 net1000 _1097_ VPWR VGND sg13g2_mux2_1
X_1197_ VPWR _1030_ net109 VGND sg13g2_inv_1
Xinput2 E1END[0] net2 VPWR VGND sg13g2_buf_1
XFILLER_51_166 VPWR VGND sg13g2_fill_1
XFILLER_51_144 VPWR VGND sg13g2_fill_2
XFILLER_10_67 VPWR VGND sg13g2_fill_2
Xoutput361 net361 WW4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput350 net350 WW4BEG[0] VPWR VGND sg13g2_buf_1
Xfanout1008 net33 net1008 VPWR VGND sg13g2_buf_1
Xfanout1019 net1020 net1019 VPWR VGND sg13g2_buf_1
XFILLER_19_43 VPWR VGND sg13g2_fill_2
XFILLER_35_20 VPWR VGND sg13g2_fill_2
X_1953_ _0602_ VPWR _0603_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0601_ sg13g2_o21ai_1
X_1884_ _0534_ _0535_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q _0536_ VPWR VGND sg13g2_nand3_1
XFILLER_21_306 VPWR VGND sg13g2_decap_4
XFILLER_21_328 VPWR VGND sg13g2_decap_4
XFILLER_21_339 VPWR VGND sg13g2_fill_2
XFILLER_51_0 VPWR VGND sg13g2_fill_2
X_2505_ net1142 net1074 Inst_LD_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_2298_ _0920_ _0276_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q VPWR VGND sg13g2_nand2_2
X_2436_ net1144 net28 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
X_1318_ net934 net931 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q _1146_ VPWR VGND sg13g2_mux2_1
X_2367_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q net945 Inst_LUT4AB_switch_matrix.JN2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q Inst_LUT4AB_switch_matrix.E1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1249_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1078_ _1081_ _1018_ sg13g2_a21oi_1
XFILLER_20_383 VPWR VGND sg13g2_fill_2
Xoutput180 net180 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput191 net191 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_21_88 VPWR VGND sg13g2_fill_1
XFILLER_7_398 VPWR VGND sg13g2_fill_2
X_2221_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q net966 _0853_ VPWR VGND sg13g2_nor2_1
X_3270_ Inst_LUT4AB_switch_matrix.W1BEG2 net320 VPWR VGND sg13g2_buf_1
X_2152_ _0788_ VPWR _0789_ VGND net64 net991 sg13g2_o21ai_1
XFILLER_38_258 VPWR VGND sg13g2_fill_2
X_2083_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q net966 net953 net959 net929 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ _0725_ VPWR VGND sg13g2_mux4_1
X_1867_ net49 net20 Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q _0519_ VPWR VGND sg13g2_mux2_1
X_1936_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q net46 net17 net74 net101 Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q
+ _0586_ VPWR VGND sg13g2_mux4_1
X_2985_ net1143 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q VPWR VGND sg13g2_dlhq_1
Xinput82 S4END[3] net82 VPWR VGND sg13g2_buf_1
Xinput71 S2MID[0] net71 VPWR VGND sg13g2_buf_1
Xinput60 S1END[1] net60 VPWR VGND sg13g2_buf_1
X_1798_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q net44 net15 net72 net99 Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q
+ _0453_ VPWR VGND sg13g2_mux4_1
Xinput93 W2END[3] net93 VPWR VGND sg13g2_buf_1
XFILLER_44_217 VPWR VGND sg13g2_fill_2
X_2419_ Inst_LE_LUT4c_frame_config_dffesr.c_reset_value net389 _1002_ _1003_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_52_294 VPWR VGND sg13g2_fill_2
XFILLER_37_280 VPWR VGND sg13g2_fill_1
XFILLER_4_302 VPWR VGND sg13g2_fill_2
X_2770_ net1203 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q VPWR VGND sg13g2_dlhq_1
X_1721_ _0378_ VPWR _0379_ VGND net999 net1216 sg13g2_o21ai_1
X_1652_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0310_ _0313_ VPWR VGND sg13g2_mux4_1
X_1583_ _0245_ VPWR _0246_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q _0242_ sg13g2_o21ai_1
X_3184_ N4END[5] net240 VPWR VGND sg13g2_buf_1
X_3253_ SS4END[6] net309 VPWR VGND sg13g2_buf_1
Xfanout1180 net1182 net1180 VPWR VGND sg13g2_buf_1
Xfanout1191 FrameData[15] net1191 VPWR VGND sg13g2_buf_1
X_2204_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q _1158_ _0196_ _0276_ _0556_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0838_ VPWR VGND sg13g2_mux4_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
X_2135_ net91 net107 net986 _0773_ VPWR VGND sg13g2_mux2_1
XFILLER_34_261 VPWR VGND sg13g2_fill_2
X_2066_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q _0707_ _0710_ _0709_ sg13g2_a21oi_1
XFILLER_22_434 VPWR VGND sg13g2_fill_1
X_1919_ _0569_ VPWR _0570_ VGND net992 net936 sg13g2_o21ai_1
X_2899_ net1198 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2968_ net1183 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_253 VPWR VGND sg13g2_decap_8
X_2753_ net1154 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_297 VPWR VGND sg13g2_decap_4
X_2822_ net1136 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q VPWR VGND sg13g2_dlhq_1
X_2684_ net1168 net1099 Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1704_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q _0361_ _0362_ VPWR VGND sg13g2_nor2_1
X_1566_ _0229_ VPWR _0230_ VGND _0221_ _0215_ sg13g2_o21ai_1
X_1635_ net59 net61 Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q _0297_ VPWR VGND sg13g2_mux2_1
X_1497_ _0163_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q net107 VPWR VGND sg13g2_nand2b_1
X_3305_ WW4END[9] net361 VPWR VGND sg13g2_buf_1
X_3236_ S4END[5] net292 VPWR VGND sg13g2_buf_1
X_2049_ _0694_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0669_ VPWR VGND sg13g2_nand2_1
X_2118_ _0757_ net929 _0753_ _0758_ VPWR VGND sg13g2_mux2_1
X_3098_ EE4END[7] net154 VPWR VGND sg13g2_buf_1
X_3167_ Inst_LUT4AB_switch_matrix.JN2BEG0 net217 VPWR VGND sg13g2_buf_2
Xfanout984 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q net984 VPWR VGND sg13g2_buf_1
Xfanout995 Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q net995 VPWR VGND sg13g2_buf_1
Xfanout962 net962 net963 VPWR VGND sg13g2_buf_16
Xfanout973 B net973 VPWR VGND sg13g2_buf_1
Xfanout951 net951 net952 VPWR VGND sg13g2_buf_16
Xfanout940 C net940 VPWR VGND sg13g2_buf_1
XFILLER_13_253 VPWR VGND sg13g2_decap_8
X_1420_ _0089_ _0088_ _0087_ VPWR VGND sg13g2_nand2_2
X_1351_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q _1012_ _1014_ _1022_ _0021_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q
+ _0022_ VPWR VGND sg13g2_mux4_1
XFILLER_51_304 VPWR VGND sg13g2_fill_1
X_3021_ net1123 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1282_ _1111_ VPWR _1112_ VGND _1014_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q sg13g2_o21ai_1
X_2805_ net1192 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q VPWR VGND sg13g2_dlhq_1
X_1618_ _0255_ _0279_ _0280_ VPWR VGND sg13g2_nor2b_1
X_2736_ net1115 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2667_ net1130 net1102 Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q VPWR VGND sg13g2_dlhq_1
X_1549_ VGND VPWR net997 _1051_ _0213_ _0212_ sg13g2_a21oi_1
X_3219_ Inst_LUT4AB_switch_matrix.JS2BEG0 net269 VPWR VGND sg13g2_buf_1
X_2598_ net1135 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_76 VPWR VGND sg13g2_decap_8
XFILLER_2_422 VPWR VGND sg13g2_fill_1
XFILLER_2_400 VPWR VGND sg13g2_fill_1
XFILLER_41_381 VPWR VGND sg13g2_fill_1
X_2521_ net1182 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_1265_ net94 net106 net1000 _1096_ VPWR VGND sg13g2_mux2_1
X_1334_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ net982 _1161_ VPWR VGND sg13g2_mux2_1
X_1403_ _0043_ _0048_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q _0072_ VPWR VGND
+ sg13g2_mux2_1
X_2452_ net1196 net1061 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
X_2383_ _0972_ _0969_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q _0967_ _0966_ VPWR
+ VGND sg13g2_a22oi_1
X_3004_ net1168 net1057 Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_131 VPWR VGND sg13g2_decap_8
X_1196_ VPWR _1029_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VGND sg13g2_inv_1
Xinput3 E1END[1] net3 VPWR VGND sg13g2_buf_1
Xfanout1009 net32 net1009 VPWR VGND sg13g2_buf_1
X_2719_ net1161 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q VPWR VGND sg13g2_dlhq_1
Xoutput362 net362 WW4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_10_46 VPWR VGND sg13g2_fill_1
Xoutput351 net351 WW4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput340 Inst_LUT4AB_switch_matrix.W6BEG1 W6BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_59_289 VPWR VGND sg13g2_fill_2
XFILLER_51_75 VPWR VGND sg13g2_fill_2
XFILLER_33_123 VPWR VGND sg13g2_decap_4
X_1952_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0600_ _0602_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q
+ sg13g2_a21oi_1
X_1883_ _0535_ net111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q VPWR VGND sg13g2_nand2b_1
XFILLER_44_0 VPWR VGND sg13g2_fill_2
X_2504_ net1176 net1074 Inst_LD_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
X_2435_ net1147 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
X_2297_ _0918_ VPWR _0919_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q _0556_
+ sg13g2_o21ai_1
X_1248_ _1080_ _1017_ _1079_ VPWR VGND sg13g2_nand2_1
X_1317_ _1145_ _1144_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q VPWR VGND sg13g2_nand2b_1
X_2366_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q net964 _0237_ Inst_LUT4AB_switch_matrix.JN2BEG0
+ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q Inst_LUT4AB_switch_matrix.E1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1179_ VPWR _1012_ net51 VGND sg13g2_inv_1
Xoutput192 net192 FrameData_O[9] VPWR VGND sg13g2_buf_1
Xoutput170 net170 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput181 net181 FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_55_281 VPWR VGND sg13g2_fill_2
XFILLER_47_226 VPWR VGND sg13g2_decap_4
XFILLER_15_123 VPWR VGND sg13g2_fill_1
X_2082_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q net977 net972 net942 net947 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ _0724_ VPWR VGND sg13g2_mux4_1
X_2220_ net1006 net945 Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0852_ VPWR VGND
+ sg13g2_mux2_1
X_2151_ VGND VPWR _1036_ net991 _0788_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q sg13g2_a21oi_1
X_2984_ net1174 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q VPWR VGND sg13g2_dlhq_1
Xinput72 S2MID[1] net72 VPWR VGND sg13g2_buf_2
Xinput61 S1END[2] net61 VPWR VGND sg13g2_buf_1
X_1935_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q net45 net100 net73 Inst_LUT4AB_switch_matrix.E2BEG6
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q _0585_ VPWR VGND sg13g2_mux4_1
X_1866_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q VPWR _0518_ VGND _0517_ _0516_ sg13g2_o21ai_1
Xinput50 N2MID[7] net50 VPWR VGND sg13g2_buf_1
X_1797_ _0450_ VPWR _0452_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q _0451_ sg13g2_o21ai_1
Xinput83 SS4END[0] net83 VPWR VGND sg13g2_buf_1
X_2418_ _1002_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q net925 VPWR VGND sg13g2_nand2_1
Xinput94 W2END[4] net94 VPWR VGND sg13g2_buf_1
X_2349_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q net1008 net1005 net1215 net960 Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ _0964_ VPWR VGND sg13g2_mux4_1
XFILLER_52_251 VPWR VGND sg13g2_fill_1
XFILLER_32_66 VPWR VGND sg13g2_decap_4
X_1720_ _0378_ net999 net11 VPWR VGND sg13g2_nand2b_1
X_1651_ _0281_ _0310_ _0312_ VPWR VGND sg13g2_nor2_1
X_3252_ SS4END[5] net308 VPWR VGND sg13g2_buf_1
X_1582_ VGND VPWR Inst_LE_LUT4c_frame_config_dffesr.c_I0mux _0245_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q
+ _0244_ sg13g2_a21oi_2
Xfanout1181 net1182 net1181 VPWR VGND sg13g2_buf_1
X_3183_ N4END[4] net233 VPWR VGND sg13g2_buf_1
Xfanout1170 FrameData[21] net1170 VPWR VGND sg13g2_buf_1
Xfanout1192 net1194 net1192 VPWR VGND sg13g2_buf_1
X_2065_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VPWR _0709_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0708_ sg13g2_o21ai_1
X_2134_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q net1007 net7 net36 net1210 net986
+ _0772_ VPWR VGND sg13g2_mux4_1
X_2203_ _0826_ VPWR Inst_LUT4AB_switch_matrix.JN2BEG0 VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q
+ _0837_ sg13g2_o21ai_1
X_2967_ net1186 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_284 VPWR VGND sg13g2_fill_1
X_2898_ net1201 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q VPWR VGND sg13g2_dlhq_1
X_1918_ _0569_ net992 net931 VPWR VGND sg13g2_nand2b_1
X_1849_ _0502_ net996 net947 VPWR VGND sg13g2_nand2b_1
XFILLER_43_21 VPWR VGND sg13g2_fill_2
XFILLER_48_398 VPWR VGND sg13g2_fill_1
XFILLER_48_354 VPWR VGND sg13g2_fill_1
XFILLER_0_361 VPWR VGND sg13g2_fill_2
X_2821_ net1139 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_232 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_fill_1
XFILLER_16_295 VPWR VGND sg13g2_fill_1
X_2752_ net1157 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1634_ _0296_ _0295_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VPWR VGND sg13g2_nand2b_1
X_2683_ net1171 net1099 Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1703_ net9 net86 Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q _0361_ VPWR VGND sg13g2_mux2_1
X_3235_ S4END[4] net285 VPWR VGND sg13g2_buf_1
X_1565_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q _0223_ _0228_ _0229_ VPWR VGND sg13g2_or3_1
X_1496_ net990 net58 net1216 net9 net1211 Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ _0162_ VPWR VGND sg13g2_mux4_1
X_3304_ WW4END[8] net360 VPWR VGND sg13g2_buf_1
X_3097_ EE4END[6] net153 VPWR VGND sg13g2_buf_1
X_2117_ VGND VPWR _0756_ _0757_ _0755_ net932 sg13g2_a21oi_2
X_2048_ _0693_ _0692_ _0690_ VPWR VGND sg13g2_nand2_2
XFILLER_10_416 VPWR VGND sg13g2_fill_2
XFILLER_57_140 VPWR VGND sg13g2_fill_1
Xfanout930 net930 Inst_LUT4AB_switch_matrix.M_AB VPWR VGND sg13g2_buf_4
Xfanout996 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q net996 VPWR VGND sg13g2_buf_1
Xfanout952 G net952 VPWR VGND sg13g2_buf_8
Xfanout941 net942 net941 VPWR VGND sg13g2_buf_1
XFILLER_38_98 VPWR VGND sg13g2_decap_8
Xfanout985 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q net985 VPWR VGND sg13g2_buf_1
Xfanout974 net974 net975 VPWR VGND sg13g2_buf_16
Xfanout963 net963 net964 VPWR VGND sg13g2_buf_16
XFILLER_9_269 VPWR VGND sg13g2_fill_2
X_1281_ _1111_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q net65 VPWR VGND sg13g2_nand2_1
X_1350_ VPWR Inst_LUT4AB_switch_matrix.JW2BEG1 _0021_ VGND sg13g2_inv_1
XFILLER_51_327 VPWR VGND sg13g2_fill_2
XFILLER_36_324 VPWR VGND sg13g2_decap_4
X_3020_ net1126 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q VPWR VGND sg13g2_dlhq_1
X_2804_ net1195 net1024 Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q VPWR VGND sg13g2_dlhq_1
X_1617_ _0278_ VPWR _0279_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q _0276_ sg13g2_o21ai_1
X_2666_ net1133 net1102 Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q VPWR VGND sg13g2_dlhq_1
X_2735_ net1117 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q VPWR VGND sg13g2_dlhq_1
X_2597_ net1138 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q VPWR VGND sg13g2_dlhq_1
X_1479_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q _0145_ _0146_ VPWR VGND sg13g2_nor2_1
X_1548_ net997 net965 _0212_ VPWR VGND sg13g2_nor2_1
XFILLER_39_184 VPWR VGND sg13g2_decap_8
X_3149_ net1030 net209 VPWR VGND sg13g2_buf_1
XFILLER_27_357 VPWR VGND sg13g2_fill_1
XFILLER_24_23 VPWR VGND sg13g2_fill_2
XFILLER_10_268 VPWR VGND sg13g2_fill_2
XFILLER_1_27 VPWR VGND sg13g2_fill_1
XFILLER_1_49 VPWR VGND sg13g2_fill_1
XFILLER_33_338 VPWR VGND sg13g2_decap_8
X_2520_ net1185 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_1402_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q _0022_ _0070_ _0071_ VPWR VGND
+ sg13g2_a21o_1
X_2451_ net1199 net1061 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
X_3003_ net1171 net1057 Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_110 VPWR VGND sg13g2_decap_4
X_1264_ net1212 net67 net1000 _1095_ VPWR VGND sg13g2_mux2_1
Xinput4 E1END[2] net4 VPWR VGND sg13g2_buf_1
X_2382_ _0971_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0970_ VPWR VGND sg13g2_nand2_1
X_1333_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q _1157_ _1159_ _1141_ _1140_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
+ _1160_ VPWR VGND sg13g2_mux4_1
XFILLER_51_146 VPWR VGND sg13g2_fill_1
XFILLER_36_143 VPWR VGND sg13g2_decap_4
X_1195_ VPWR _1028_ net107 VGND sg13g2_inv_1
XFILLER_24_305 VPWR VGND sg13g2_decap_4
X_2718_ net1163 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q VPWR VGND sg13g2_dlhq_1
Xoutput352 net352 WW4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput363 net363 WW4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput330 net330 W2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_10_69 VPWR VGND sg13g2_fill_1
Xoutput341 net341 W6BEG[1] VPWR VGND sg13g2_buf_1
X_2649_ net1180 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_35_22 VPWR VGND sg13g2_fill_1
XFILLER_51_21 VPWR VGND sg13g2_fill_1
XFILLER_23_360 VPWR VGND sg13g2_decap_4
XFILLER_4_0 VPWR VGND sg13g2_fill_2
XFILLER_2_220 VPWR VGND sg13g2_fill_1
XFILLER_38_408 VPWR VGND sg13g2_fill_1
X_1951_ net976 net971 net983 _0601_ VPWR VGND sg13g2_mux2_1
X_1882_ _0534_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q net380 VPWR VGND sg13g2_nand2_1
X_2503_ net1208 net1074 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_2434_ net1150 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
X_2365_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q net957 Inst_LUT4AB_switch_matrix.JN2BEG1
+ net980 _0623_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q Inst_LUT4AB_switch_matrix.E1BEG2
+ VPWR VGND sg13g2_mux4_1
X_2296_ _0918_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q _1119_ VPWR VGND sg13g2_nand2_1
X_1247_ net1212 net67 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1079_ VPWR VGND sg13g2_mux2_1
X_1316_ net955 net950 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q _1144_ VPWR VGND sg13g2_mux2_1
XFILLER_20_385 VPWR VGND sg13g2_fill_1
Xoutput193 net193 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput182 net182 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput171 net171 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput160 net160 EE4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_28_452 VPWR VGND sg13g2_fill_2
XFILLER_15_113 VPWR VGND sg13g2_fill_2
XFILLER_11_330 VPWR VGND sg13g2_fill_2
XFILLER_7_389 VPWR VGND sg13g2_fill_2
XFILLER_19_452 VPWR VGND sg13g2_fill_2
X_2150_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q net56 net7 net1214 net1210 Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ _0787_ VPWR VGND sg13g2_mux4_1
X_2081_ Inst_LUT4AB_switch_matrix.JW2BEG7 _0717_ _0723_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
+ _0715_ VPWR VGND sg13g2_a22oi_1
X_1934_ Inst_LUT4AB_switch_matrix.E2BEG6 _0578_ _0584_ _0573_ _0567_ VPWR VGND sg13g2_a22oi_1
X_2983_ net1207 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VPWR VGND sg13g2_dlhq_1
Xinput84 SS4END[1] net84 VPWR VGND sg13g2_buf_1
Xinput73 S2MID[2] net73 VPWR VGND sg13g2_buf_1
Xinput62 S1END[3] net62 VPWR VGND sg13g2_buf_1
X_1865_ net77 Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q _0517_ VPWR VGND sg13g2_nor2_1
Xinput95 W2END[5] net95 VPWR VGND sg13g2_buf_1
Xinput40 N2END[5] net40 VPWR VGND sg13g2_buf_1
Xinput51 N4END[0] net51 VPWR VGND sg13g2_buf_1
X_1796_ net43 net71 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q _0451_ VPWR VGND sg13g2_mux2_1
X_2348_ _0959_ _0962_ _0963_ VPWR VGND sg13g2_nor2_1
X_2417_ _1001_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q net927 VPWR VGND sg13g2_nand2b_1
X_2279_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q net978 _0903_ VPWR VGND sg13g2_nor2b_1
XFILLER_44_219 VPWR VGND sg13g2_fill_1
XFILLER_52_296 VPWR VGND sg13g2_fill_1
XFILLER_32_23 VPWR VGND sg13g2_decap_8
XFILLER_43_285 VPWR VGND sg13g2_decap_4
XFILLER_31_458 VPWR VGND sg13g2_fill_1
X_1650_ _0311_ _0281_ _0310_ VPWR VGND sg13g2_nand2_1
X_1581_ VGND VPWR _0243_ _0244_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q _0238_ sg13g2_a21oi_2
XFILLER_11_182 VPWR VGND sg13g2_fill_2
XFILLER_11_193 VPWR VGND sg13g2_fill_1
X_3251_ SS4END[4] net301 VPWR VGND sg13g2_buf_1
X_3182_ net50 net232 VPWR VGND sg13g2_buf_1
X_2202_ _0831_ VPWR _0837_ VGND _0833_ _0836_ sg13g2_o21ai_1
Xfanout1182 FrameData[18] net1182 VPWR VGND sg13g2_buf_1
Xfanout1171 net1173 net1171 VPWR VGND sg13g2_buf_1
Xfanout1193 net1194 net1193 VPWR VGND sg13g2_buf_1
Xfanout1160 net1161 net1160 VPWR VGND sg13g2_buf_1
X_2064_ net59 net63 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q _0708_ VPWR VGND sg13g2_mux2_1
XFILLER_26_208 VPWR VGND sg13g2_fill_1
X_2133_ _0770_ VPWR _0771_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0763_ sg13g2_o21ai_1
X_2897_ net1206 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1917_ net966 net960 net992 _0568_ VPWR VGND sg13g2_mux2_1
X_2966_ net1189 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1848_ VGND VPWR _0501_ _0498_ _0500_ sg13g2_or2_1
X_1779_ VGND VPWR net984 _1051_ _0435_ _0434_ sg13g2_a21oi_1
XFILLER_57_377 VPWR VGND sg13g2_fill_1
X_2751_ net1160 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2820_ net1144 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_16_274 VPWR VGND sg13g2_decap_8
X_1702_ Inst_LUT4AB_switch_matrix.JN2BEG2 _0354_ _0360_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
+ _0352_ VPWR VGND sg13g2_a22oi_1
X_1633_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q net1008 net41 net1215 net12 Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0295_ VPWR VGND sg13g2_mux4_1
X_2682_ net1177 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1564_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0225_ _0228_ _0227_ sg13g2_a21oi_1
X_1495_ _1038_ _0154_ _0161_ VPWR VGND sg13g2_nor2_1
X_3234_ net78 net284 VPWR VGND sg13g2_buf_1
X_3303_ WW4END[7] net359 VPWR VGND sg13g2_buf_1
X_3096_ EE4END[5] net152 VPWR VGND sg13g2_buf_1
X_2116_ net954 _0755_ _0756_ VPWR VGND sg13g2_nor2_2
X_2047_ _0691_ VPWR _0692_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q _0275_ sg13g2_o21ai_1
X_2949_ net1138 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q VPWR VGND sg13g2_dlhq_1
Xfanout942 net942 net943 VPWR VGND sg13g2_buf_16
Xfanout931 Inst_LUT4AB_switch_matrix.M_AD net931 VPWR VGND sg13g2_buf_1
Xfanout997 net998 net997 VPWR VGND sg13g2_buf_1
XFILLER_38_66 VPWR VGND sg13g2_fill_1
Xfanout953 net954 net953 VPWR VGND sg13g2_buf_1
Xfanout964 E net964 VPWR VGND sg13g2_buf_8
Xfanout986 Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q net986 VPWR VGND sg13g2_buf_1
Xfanout975 net975 A VPWR VGND sg13g2_buf_16
X_3047__371 VPWR VGND net371 sg13g2_tiehi
X_1280_ _1110_ _1109_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VPWR VGND sg13g2_nand2b_1
X_2803_ net1200 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2734_ net1121 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1547_ VGND VPWR net997 Inst_LUT4AB_switch_matrix.M_AD _0211_ _0210_ sg13g2_a21oi_1
X_1616_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q _0277_ _0278_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q
+ sg13g2_a21oi_1
X_2596_ net1146 net1085 Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q VPWR VGND sg13g2_dlhq_1
X_2665_ net1143 net1102 Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1478_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0142_ _0145_ _0144_ sg13g2_a21oi_1
XFILLER_39_130 VPWR VGND sg13g2_fill_1
X_3148_ net1036 net208 VPWR VGND sg13g2_buf_1
XFILLER_27_325 VPWR VGND sg13g2_fill_1
X_3079_ net18 net129 VPWR VGND sg13g2_buf_1
XFILLER_49_43 VPWR VGND sg13g2_fill_1
XFILLER_18_358 VPWR VGND sg13g2_fill_2
XFILLER_41_361 VPWR VGND sg13g2_fill_1
XFILLER_5_284 VPWR VGND sg13g2_fill_2
X_1401_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q VPWR _0070_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q
+ _0023_ sg13g2_o21ai_1
X_2450_ net1202 net1061 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
X_2381_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q Inst_LUT4AB_switch_matrix.JN2BEG2
+ Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_switch_matrix.E2BEG2 net384 Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q
+ _0970_ VPWR VGND sg13g2_mux4_1
X_3002_ net1177 net1057 Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1332_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q net48 net19 net76 net103 Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q
+ _1159_ VPWR VGND sg13g2_mux4_1
X_1263_ VGND VPWR _1093_ _1094_ _1086_ _1015_ sg13g2_a21oi_2
X_1194_ VPWR _1027_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VGND sg13g2_inv_1
Xinput5 E1END[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_51_136 VPWR VGND sg13g2_fill_2
XFILLER_51_103 VPWR VGND sg13g2_fill_2
X_2717_ net1166 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2579_ net1200 net1084 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
Xoutput331 net331 W2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput320 net320 W1BEG[2] VPWR VGND sg13g2_buf_1
X_2648_ net1183 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q VPWR VGND sg13g2_dlhq_1
Xoutput353 net353 WW4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput364 net364 WW4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput342 net342 W6BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_42_136 VPWR VGND sg13g2_fill_2
XFILLER_51_77 VPWR VGND sg13g2_fill_1
X_3051__367 VPWR VGND net367 sg13g2_tiehi
XFILLER_2_276 VPWR VGND sg13g2_fill_2
XFILLER_18_133 VPWR VGND sg13g2_fill_2
X_1950_ _0599_ VPWR _0600_ VGND net983 net941 sg13g2_o21ai_1
X_1881_ net1211 net80 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q _0533_ VPWR VGND sg13g2_mux2_1
X_2502_ net1136 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_2433_ net1153 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 VPWR
+ VGND sg13g2_dlhq_1
X_1315_ VPWR _1143_ _1142_ VGND sg13g2_inv_1
X_2364_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q net952 _1159_ Inst_LUT4AB_switch_matrix.JN2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q Inst_LUT4AB_switch_matrix.E1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_52_434 VPWR VGND sg13g2_fill_2
XFILLER_37_431 VPWR VGND sg13g2_fill_1
X_2295_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q _0916_ _0917_ VPWR VGND sg13g2_nor2_1
X_1246_ net94 net106 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1078_ VPWR VGND sg13g2_mux2_1
XFILLER_24_125 VPWR VGND sg13g2_fill_2
XFILLER_20_364 VPWR VGND sg13g2_fill_2
Xoutput150 Inst_LUT4AB_switch_matrix.EE4BEG2 EE4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput161 net161 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput183 net183 FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput194 net194 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput172 net172 FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_55_283 VPWR VGND sg13g2_fill_1
XFILLER_46_99 VPWR VGND sg13g2_fill_2
XFILLER_30_128 VPWR VGND sg13g2_decap_4
XFILLER_30_117 VPWR VGND sg13g2_decap_8
X_2080_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q _0722_ _0723_ VPWR VGND sg13g2_nor2_1
X_1933_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q _0583_ _0584_ VPWR VGND sg13g2_nor2_1
X_2982_ net1135 net1048 Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q VPWR VGND sg13g2_dlhq_1
Xinput85 SS4END[2] net85 VPWR VGND sg13g2_buf_1
Xinput63 S2END[0] net63 VPWR VGND sg13g2_buf_1
Xinput74 S2MID[3] net74 VPWR VGND sg13g2_buf_1
X_1864_ Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q
+ _0516_ VPWR VGND sg13g2_nor2b_1
Xinput52 N4END[1] net52 VPWR VGND sg13g2_buf_1
Xinput30 FrameStrobe[7] net30 VPWR VGND sg13g2_buf_1
Xinput41 N2END[6] net41 VPWR VGND sg13g2_buf_1
X_1795_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q VPWR _0450_ VGND _0449_ _0448_ sg13g2_o21ai_1
Xinput96 W2END[6] net96 VPWR VGND sg13g2_buf_1
X_2347_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q VPWR _0962_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
+ _0961_ sg13g2_o21ai_1
X_2278_ _0901_ VPWR _0902_ VGND _1013_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q sg13g2_o21ai_1
X_2416_ net391 _1000_ _0998_ _0004_ VPWR VGND sg13g2_mux2_1
XFILLER_29_228 VPWR VGND sg13g2_fill_2
X_1229_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _1061_ _1062_ _1020_ sg13g2_a21oi_1
XFILLER_16_47 VPWR VGND sg13g2_fill_2
XFILLER_57_10 VPWR VGND sg13g2_fill_2
XFILLER_57_87 VPWR VGND sg13g2_fill_2
XFILLER_31_448 VPWR VGND sg13g2_fill_1
X_1580_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q _0239_ _0243_ VPWR VGND sg13g2_nor2b_1
Xfanout1172 net1173 net1172 VPWR VGND sg13g2_buf_1
X_3181_ net49 net231 VPWR VGND sg13g2_buf_1
Xfanout1183 net1185 net1183 VPWR VGND sg13g2_buf_1
Xfanout1161 FrameData[24] net1161 VPWR VGND sg13g2_buf_1
Xfanout1150 net1151 net1150 VPWR VGND sg13g2_buf_1
X_3250_ Inst_LUT4AB_switch_matrix.S4BEG3 net291 VPWR VGND sg13g2_buf_1
X_2132_ _0769_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q _0770_ VPWR VGND sg13g2_nor2b_1
X_2201_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VPWR _0836_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ _0835_ sg13g2_o21ai_1
XFILLER_21_4 VPWR VGND sg13g2_fill_2
Xfanout1194 FrameData[14] net1194 VPWR VGND sg13g2_buf_1
XFILLER_34_253 VPWR VGND sg13g2_fill_2
X_2063_ _0706_ VPWR _0707_ VGND net87 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q sg13g2_o21ai_1
X_1916_ _0567_ _0566_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR VGND sg13g2_nand2b_1
X_1847_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR _0500_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ _0499_ sg13g2_o21ai_1
X_2965_ net1192 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2896_ net1116 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1778_ net984 net958 _0434_ VPWR VGND sg13g2_nor2_1
XFILLER_43_23 VPWR VGND sg13g2_fill_1
XFILLER_40_267 VPWR VGND sg13g2_fill_1
XFILLER_40_223 VPWR VGND sg13g2_fill_1
X_1701_ VGND VPWR _0356_ _0359_ _0360_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q sg13g2_a21oi_1
X_2750_ net1163 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q VPWR VGND sg13g2_dlhq_1
X_2681_ net1180 net1099 Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_256 VPWR VGND sg13g2_fill_1
X_1632_ _0293_ VPWR _0294_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0291_ sg13g2_o21ai_1
X_1563_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VPWR _0227_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ _0226_ sg13g2_o21ai_1
X_1494_ _0159_ VPWR _0160_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0156_ sg13g2_o21ai_1
X_3302_ WW4END[6] net358 VPWR VGND sg13g2_buf_1
X_3233_ net77 net283 VPWR VGND sg13g2_buf_1
X_2115_ _0754_ VPWR _0755_ VGND _0753_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q
+ sg13g2_o21ai_1
X_3095_ EE4END[4] net145 VPWR VGND sg13g2_buf_1
X_3164_ Inst_LUT4AB_switch_matrix.N1BEG1 net214 VPWR VGND sg13g2_buf_1
XFILLER_12_0 VPWR VGND sg13g2_fill_2
X_2046_ VGND VPWR _1047_ _0691_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q Inst_LUT4AB_switch_matrix.JW2BEG5
+ sg13g2_a21oi_2
X_2879_ net1159 net1033 Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_10_418 VPWR VGND sg13g2_fill_1
X_2948_ net1146 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VPWR VGND sg13g2_dlhq_1
Xfanout965 net966 net965 VPWR VGND sg13g2_buf_1
Xfanout954 G net954 VPWR VGND sg13g2_buf_1
Xfanout976 net977 net976 VPWR VGND sg13g2_buf_1
Xfanout932 _1052_ net932 VPWR VGND sg13g2_buf_1
Xfanout943 C net943 VPWR VGND sg13g2_buf_8
XFILLER_54_44 VPWR VGND sg13g2_fill_2
Xfanout987 Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q net987 VPWR VGND sg13g2_buf_1
Xfanout998 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q net998 VPWR VGND sg13g2_buf_1
XFILLER_13_201 VPWR VGND sg13g2_fill_1
XFILLER_48_186 VPWR VGND sg13g2_decap_8
XFILLER_51_329 VPWR VGND sg13g2_fill_1
X_2802_ net1201 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2733_ net1124 net1012 Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2664_ net1175 net1102 Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q VPWR VGND sg13g2_dlhq_1
X_1477_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR _0144_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0143_ sg13g2_o21ai_1
X_1546_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q VPWR _0210_ VGND net998 net933 sg13g2_o21ai_1
X_1615_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q net48 net19 net76 net103 Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q
+ _0277_ VPWR VGND sg13g2_mux4_1
X_2595_ net1149 net1085 Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_167 VPWR VGND sg13g2_fill_1
X_3078_ net17 net128 VPWR VGND sg13g2_buf_1
X_3216_ Inst_LUT4AB_switch_matrix.S1BEG1 net266 VPWR VGND sg13g2_buf_1
X_3147_ net1041 net207 VPWR VGND sg13g2_buf_1
X_2029_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux _0674_ _0675_ VPWR VGND sg13g2_nor2b_1
XFILLER_45_167 VPWR VGND sg13g2_fill_1
X_1331_ VPWR _1158_ _1157_ VGND sg13g2_inv_1
X_2380_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0334_ _0969_ _0968_ sg13g2_a21oi_1
X_1400_ _0069_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ A VPWR VGND sg13g2_mux2_2
X_3001_ net1182 net1057 Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q VPWR VGND sg13g2_dlhq_1
X_1193_ VPWR _1026_ net102 VGND sg13g2_inv_1
Xinput6 E2END[0] net6 VPWR VGND sg13g2_buf_1
X_1262_ _1093_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q _1092_ VPWR VGND sg13g2_nand2b_1
Xoutput310 net310 SS4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput321 Inst_LUT4AB_switch_matrix.W1BEG3 W1BEG[3] VPWR VGND sg13g2_buf_1
Xoutput332 net332 W2BEGb[2] VPWR VGND sg13g2_buf_1
X_2647_ net1186 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q VPWR VGND sg13g2_dlhq_1
Xoutput343 net343 W6BEG[3] VPWR VGND sg13g2_buf_1
X_2716_ net1169 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2578_ net1202 net1084 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_1529_ net380 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q _0192_ _0193_ VPWR VGND sg13g2_a21o_1
Xoutput354 net354 WW4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput365 net365 WW4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_55_421 VPWR VGND sg13g2_fill_2
X_1880_ _0530_ _0531_ Inst_LG_LUT4c_frame_config_dffesr.c_I0mux _0532_ VPWR VGND sg13g2_mux2_1
XFILLER_33_148 VPWR VGND sg13g2_fill_2
X_2501_ net1140 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_2294_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q net1009 net1216 net60 net948 Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ _0916_ VPWR VGND sg13g2_mux4_1
X_2432_ net1157 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
X_2363_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q net962 Inst_LUT4AB_switch_matrix.E2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q Inst_LUT4AB_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1314_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q net974 net968 net938 net961 Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ _1142_ VPWR VGND sg13g2_mux4_1
XFILLER_52_457 VPWR VGND sg13g2_fill_2
X_1245_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q _1076_ _1077_ VPWR VGND sg13g2_nor2_1
Xoutput195 net195 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput184 net184 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput162 net162 FrameData_O[10] VPWR VGND sg13g2_buf_1
Xoutput151 Inst_LUT4AB_switch_matrix.EE4BEG3 EE4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput173 net173 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput140 net140 E6BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_21_48 VPWR VGND sg13g2_fill_1
XFILLER_28_454 VPWR VGND sg13g2_fill_1
XFILLER_11_332 VPWR VGND sg13g2_fill_1
XFILLER_19_454 VPWR VGND sg13g2_fill_1
X_1932_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0580_ _0583_ _0582_ sg13g2_a21oi_1
X_1863_ Inst_LUT4AB_switch_matrix.JN2BEG6 _0509_ _0515_ _0507_ _0501_ VPWR VGND sg13g2_a22oi_1
X_2981_ net1138 net1048 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q VPWR VGND sg13g2_dlhq_1
Xinput31 N1END[0] net31 VPWR VGND sg13g2_buf_1
Xinput20 E2MID[6] net20 VPWR VGND sg13g2_buf_1
Xinput64 S2END[1] net64 VPWR VGND sg13g2_buf_1
Xinput75 S2MID[4] net75 VPWR VGND sg13g2_buf_1
Xinput86 SS4END[3] net86 VPWR VGND sg13g2_buf_1
XFILLER_42_0 VPWR VGND sg13g2_fill_2
X_2415_ Inst_LD_LUT4c_frame_config_dffesr.c_reset_value _0688_ _0999_ _1000_ VPWR
+ VGND sg13g2_mux2_1
Xinput53 N4END[2] net53 VPWR VGND sg13g2_buf_1
Xinput97 W2END[7] net97 VPWR VGND sg13g2_buf_1
Xinput42 N2END[7] net42 VPWR VGND sg13g2_buf_1
X_1794_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q net98 _0449_ VPWR VGND sg13g2_nor2_1
X_2346_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q _1084_ _0961_ _0960_ sg13g2_a21oi_1
X_2277_ VGND VPWR net1004 Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q _0901_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ sg13g2_a21oi_1
XFILLER_29_218 VPWR VGND sg13g2_decap_4
X_1228_ net92 net111 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q _1061_ VPWR VGND sg13g2_mux2_1
XFILLER_20_162 VPWR VGND sg13g2_fill_1
XFILLER_16_402 VPWR VGND sg13g2_fill_1
XFILLER_11_184 VPWR VGND sg13g2_fill_1
Xfanout1140 FrameData[30] net1140 VPWR VGND sg13g2_buf_1
Xfanout1184 net1185 net1184 VPWR VGND sg13g2_buf_1
Xfanout1173 FrameData[20] net1173 VPWR VGND sg13g2_buf_1
Xfanout1195 net1197 net1195 VPWR VGND sg13g2_buf_1
X_3180_ net48 net230 VPWR VGND sg13g2_buf_1
Xfanout1162 net1164 net1162 VPWR VGND sg13g2_buf_1
Xfanout1151 FrameData[27] net1151 VPWR VGND sg13g2_buf_1
X_2062_ _0706_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q net1004 VPWR VGND sg13g2_nand2b_1
X_2131_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q _0767_ _0769_ _0768_ sg13g2_a21oi_1
X_2200_ VGND VPWR net84 net1002 _0835_ _0834_ sg13g2_a21oi_1
X_2964_ net1195 net1050 Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_34_243 VPWR VGND sg13g2_fill_2
X_1915_ net992 net978 net973 net943 D Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0566_
+ VPWR VGND sg13g2_mux4_1
X_1846_ net965 net959 net996 _0499_ VPWR VGND sg13g2_mux2_1
X_1777_ net984 net976 net971 net941 net946 Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ _0433_ VPWR VGND sg13g2_mux4_1
X_2895_ net1119 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VPWR VGND sg13g2_dlhq_1
X_2329_ VGND VPWR _0946_ net980 Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q sg13g2_or2_1
X_1700_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0358_ _0359_ _1031_ sg13g2_a21oi_1
X_1631_ _0293_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0292_ VPWR VGND sg13g2_nand2b_1
X_2680_ net1183 net1099 Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1562_ net61 net69 net997 _0226_ VPWR VGND sg13g2_mux2_1
X_1493_ VGND VPWR _1037_ _0159_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0158_ sg13g2_a21oi_2
X_3232_ net76 net282 VPWR VGND sg13g2_buf_1
X_3301_ WW4END[5] net357 VPWR VGND sg13g2_buf_1
XFILLER_54_327 VPWR VGND sg13g2_fill_1
XFILLER_54_305 VPWR VGND sg13g2_fill_1
X_2114_ _0754_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0670_ VPWR VGND sg13g2_nand2_1
X_2045_ _0689_ VPWR _0690_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q _0230_ sg13g2_o21ai_1
X_2947_ net1149 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1829_ VGND VPWR _0482_ _0483_ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q sg13g2_a21oi_2
X_2878_ net1162 net1036 Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q VPWR VGND sg13g2_dlhq_1
Xfanout999 Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q net999 VPWR VGND sg13g2_buf_1
Xfanout966 net967 net966 VPWR VGND sg13g2_buf_1
Xfanout933 _1052_ net933 VPWR VGND sg13g2_buf_1
Xfanout977 net979 net977 VPWR VGND sg13g2_buf_1
Xfanout988 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q net988 VPWR VGND sg13g2_buf_1
Xfanout955 net955 net956 VPWR VGND sg13g2_buf_16
Xfanout944 net945 net944 VPWR VGND sg13g2_buf_2
XFILLER_53_382 VPWR VGND sg13g2_fill_1
XFILLER_13_268 VPWR VGND sg13g2_fill_1
X_2801_ net1206 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1614_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q _1021_ _1026_ _1034_ _0275_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q
+ _0276_ VPWR VGND sg13g2_mux4_1
X_2732_ net1128 net1012 Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q VPWR VGND sg13g2_dlhq_1
X_2594_ net1152 net1086 Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2663_ net1209 net1102 Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q VPWR VGND sg13g2_dlhq_1
X_1476_ net60 net62 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q _0143_ VPWR VGND sg13g2_mux2_1
X_1545_ _0201_ VPWR _0209_ VGND _0208_ _0200_ sg13g2_o21ai_1
X_3215_ Inst_LUT4AB_switch_matrix.S1BEG0 net265 VPWR VGND sg13g2_buf_1
X_3146_ net1044 net206 VPWR VGND sg13g2_buf_1
X_3077_ net16 net127 VPWR VGND sg13g2_buf_1
XFILLER_39_154 VPWR VGND sg13g2_decap_4
X_2028_ _0673_ VPWR _0674_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q _0389_ sg13g2_o21ai_1
XFILLER_14_92 VPWR VGND sg13g2_fill_2
XFILLER_30_80 VPWR VGND sg13g2_fill_2
XFILLER_5_286 VPWR VGND sg13g2_fill_1
X_1261_ VGND VPWR _1091_ _1092_ _1090_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q sg13g2_a21oi_2
X_1330_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q net47 net18 net102 Inst_LUT4AB_switch_matrix.JS2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q _1157_ VPWR VGND sg13g2_mux4_1
XFILLER_51_105 VPWR VGND sg13g2_fill_1
X_3000_ net1183 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q VPWR VGND sg13g2_dlhq_1
Xinput7 E2END[1] net7 VPWR VGND sg13g2_buf_1
X_1192_ VPWR _1025_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VGND sg13g2_inv_1
XFILLER_51_138 VPWR VGND sg13g2_fill_1
X_2577_ net1205 net1083 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
Xoutput300 net300 S4BEG[9] VPWR VGND sg13g2_buf_1
X_2646_ net1189 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q VPWR VGND sg13g2_dlhq_1
Xoutput311 net311 SS4BEG[4] VPWR VGND sg13g2_buf_1
X_2715_ net1172 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q VPWR VGND sg13g2_dlhq_1
Xoutput333 net333 W2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput355 net355 WW4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput344 net344 W6BEG[4] VPWR VGND sg13g2_buf_1
Xoutput322 net322 W2BEG[0] VPWR VGND sg13g2_buf_1
X_1528_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q VPWR _0192_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ _1034_ sg13g2_o21ai_1
XFILLER_19_37 VPWR VGND sg13g2_fill_1
X_1459_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0124_ _0127_ _0126_ sg13g2_a21oi_1
X_3129_ net1181 net170 VPWR VGND sg13g2_buf_1
XFILLER_27_146 VPWR VGND sg13g2_decap_4
XFILLER_18_135 VPWR VGND sg13g2_fill_1
X_2500_ net1144 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2431_ net1160 net1059 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_271 VPWR VGND sg13g2_fill_2
X_2293_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q _0912_ _0913_ _0914_ _0915_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
+ Inst_LUT4AB_switch_matrix.E6BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_2_84 VPWR VGND sg13g2_fill_1
X_1244_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q net1008 net39 net51 net10 Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q
+ _1076_ VPWR VGND sg13g2_mux4_1
X_2362_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q net957 _0237_ Inst_LUT4AB_switch_matrix.E2BEG0
+ net376 Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q Inst_LUT4AB_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1313_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q net39 net67 net22 net94 Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q
+ _1141_ VPWR VGND sg13g2_mux4_1
Xoutput196 net196 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput141 net141 E6BEG[6] VPWR VGND sg13g2_buf_1
Xoutput185 net185 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput174 net174 FrameData_O[21] VPWR VGND sg13g2_buf_1
Xoutput163 net163 FrameData_O[11] VPWR VGND sg13g2_buf_1
Xoutput130 net130 E2BEGb[5] VPWR VGND sg13g2_buf_1
X_2629_ net1140 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q VPWR VGND sg13g2_dlhq_1
Xoutput152 net152 EE4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_28_433 VPWR VGND sg13g2_fill_2
XFILLER_2_0 VPWR VGND sg13g2_fill_2
X_2980_ net1146 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1931_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR _0582_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ _0581_ sg13g2_o21ai_1
X_1862_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q _0514_ _0515_ VPWR VGND sg13g2_nor2_1
Xinput10 E2END[4] net10 VPWR VGND sg13g2_buf_1
Xinput21 E2MID[7] net21 VPWR VGND sg13g2_buf_1
Xinput54 N4END[3] net54 VPWR VGND sg13g2_buf_1
Xinput43 N2MID[0] net43 VPWR VGND sg13g2_buf_1
X_1793_ Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
+ _0448_ VPWR VGND sg13g2_nor2b_1
Xinput32 N1END[1] net32 VPWR VGND sg13g2_buf_1
Xinput65 S2END[2] net65 VPWR VGND sg13g2_buf_1
Xinput76 S2MID[5] net76 VPWR VGND sg13g2_buf_1
X_2414_ _0999_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q net925 VPWR VGND sg13g2_nand2_1
XFILLER_35_0 VPWR VGND sg13g2_fill_2
Xinput98 W2MID[0] net98 VPWR VGND sg13g2_buf_1
Xinput87 W1END[0] net87 VPWR VGND sg13g2_buf_1
X_2345_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q net954 _0960_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_263 VPWR VGND sg13g2_decap_4
X_2276_ _0898_ _0900_ Inst_LUT4AB_switch_matrix.SS4BEG0 VPWR VGND sg13g2_nor2_2
X_1227_ _1060_ _1059_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q VPWR VGND sg13g2_nand2b_1
XFILLER_32_37 VPWR VGND sg13g2_decap_4
XFILLER_57_67 VPWR VGND sg13g2_fill_2
XFILLER_57_12 VPWR VGND sg13g2_fill_1
XFILLER_28_241 VPWR VGND sg13g2_fill_1
Xfanout1196 net1197 net1196 VPWR VGND sg13g2_buf_1
Xfanout1185 FrameData[17] net1185 VPWR VGND sg13g2_buf_1
Xfanout1163 net1164 net1163 VPWR VGND sg13g2_buf_1
Xfanout1130 FrameData[4] net1130 VPWR VGND sg13g2_buf_1
Xfanout1141 FrameData[2] net1141 VPWR VGND sg13g2_buf_1
Xfanout1152 FrameData[27] net1152 VPWR VGND sg13g2_buf_1
X_2061_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q net1010 net35 net1217 net6 Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0705_ VPWR VGND sg13g2_mux4_1
X_2130_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VPWR _0768_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ _0765_ sg13g2_o21ai_1
XFILLER_21_6 VPWR VGND sg13g2_fill_1
Xfanout1174 net1176 net1174 VPWR VGND sg13g2_buf_1
X_2963_ net1200 net1051 Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1914_ _0564_ VPWR _0565_ VGND _0562_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q sg13g2_o21ai_1
X_1845_ VGND VPWR _0497_ _0498_ Inst_LUT4AB_switch_matrix.M_AH net996 sg13g2_a21oi_2
X_2894_ net1120 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1776_ VGND VPWR _0431_ _0432_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q _0425_
+ sg13g2_a21oi_2
X_2328_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q _0940_ _0941_ _0943_ _0945_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q
+ Inst_LUT4AB_switch_matrix.NN4BEG3 VPWR VGND sg13g2_mux4_1
X_2259_ _0883_ _0885_ Inst_LUT4AB_switch_matrix.SS4BEG2 VPWR VGND sg13g2_nor2_1
XFILLER_4_19 VPWR VGND sg13g2_fill_1
XFILLER_0_332 VPWR VGND sg13g2_fill_2
XFILLER_16_288 VPWR VGND sg13g2_decap_8
X_1630_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q net967 net953 net937 net930 Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0292_ VPWR VGND sg13g2_mux4_1
X_3231_ net75 net281 VPWR VGND sg13g2_buf_1
X_1561_ _0224_ VPWR _0225_ VGND net997 net87 sg13g2_o21ai_1
X_1492_ _0157_ VPWR _0158_ VGND net990 net937 sg13g2_o21ai_1
X_3162_ net1059 net203 VPWR VGND sg13g2_buf_1
X_3300_ WW4END[4] net350 VPWR VGND sg13g2_buf_1
X_3093_ Inst_LUT4AB_switch_matrix.E6BEG0 net134 VPWR VGND sg13g2_buf_1
X_2113_ _0752_ _0693_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0753_ VPWR VGND
+ sg13g2_mux2_1
X_2044_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q Inst_LUT4AB_switch_matrix.E2BEG5
+ _0689_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q sg13g2_a21oi_1
X_2877_ net1165 net1036 Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2946_ net1152 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_247 VPWR VGND sg13g2_fill_2
X_1828_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q VPWR _0482_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q
+ _0253_ sg13g2_o21ai_1
X_1759_ net985 net1009 net38 net25 net1210 Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0416_ VPWR VGND sg13g2_mux4_1
Xfanout989 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q net989 VPWR VGND sg13g2_buf_1
Xfanout978 net979 net978 VPWR VGND sg13g2_buf_1
Xfanout967 E net967 VPWR VGND sg13g2_buf_1
Xfanout956 net956 net957 VPWR VGND sg13g2_buf_16
Xfanout934 net934 net935 VPWR VGND sg13g2_buf_16
Xfanout945 D net945 VPWR VGND sg13g2_buf_1
XFILLER_53_350 VPWR VGND sg13g2_fill_2
XFILLER_13_247 VPWR VGND sg13g2_fill_2
XFILLER_48_133 VPWR VGND sg13g2_fill_2
XFILLER_36_328 VPWR VGND sg13g2_fill_2
XFILLER_44_90 VPWR VGND sg13g2_fill_2
X_2731_ net1130 net1012 Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2800_ net1114 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1613_ VPWR Inst_LUT4AB_switch_matrix.JS2BEG5 _0275_ VGND sg13g2_inv_1
X_2593_ net1155 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1544_ VGND VPWR _0206_ _0208_ _0204_ _0207_ sg13g2_a21oi_2
X_2662_ net1135 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3145_ net1052 net205 VPWR VGND sg13g2_buf_1
X_1475_ _0141_ VPWR _0142_ VGND net68 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q sg13g2_o21ai_1
XFILLER_39_122 VPWR VGND sg13g2_fill_1
XFILLER_39_100 VPWR VGND sg13g2_fill_1
X_2027_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q _0391_ _0673_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q
+ sg13g2_a21oi_1
X_3076_ net15 net126 VPWR VGND sg13g2_buf_1
X_2929_ net1206 net1045 Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_37 VPWR VGND sg13g2_fill_2
XFILLER_49_79 VPWR VGND sg13g2_fill_2
XFILLER_53_191 VPWR VGND sg13g2_fill_2
XFILLER_53_180 VPWR VGND sg13g2_fill_1
Xinput8 E2END[2] net8 VPWR VGND sg13g2_buf_1
X_1260_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VPWR _1091_ VGND _1088_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ sg13g2_o21ai_1
X_1191_ VPWR _1024_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VGND sg13g2_inv_1
XFILLER_24_309 VPWR VGND sg13g2_fill_1
X_2714_ net1178 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q VPWR VGND sg13g2_dlhq_1
X_2576_ net1114 net1084 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_1527_ Inst_LUT4AB_switch_matrix.JS2BEG4 _0191_ _1035_ _0176_ _0182_ VPWR VGND sg13g2_a22oi_1
X_2645_ net1192 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q VPWR VGND sg13g2_dlhq_1
Xoutput334 net334 W2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput312 net312 SS4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput301 net301 SS4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput356 Inst_LUT4AB_switch_matrix.WW4BEG3 WW4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput323 net323 W2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput345 net345 W6BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_59_239 VPWR VGND sg13g2_fill_2
X_3128_ net1185 net169 VPWR VGND sg13g2_buf_1
X_1389_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ net982 _0059_ VPWR VGND sg13g2_mux2_1
X_1458_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VPWR _0126_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ _0125_ sg13g2_o21ai_1
XFILLER_35_37 VPWR VGND sg13g2_fill_2
XFILLER_23_353 VPWR VGND sg13g2_fill_2
XFILLER_23_364 VPWR VGND sg13g2_fill_1
XFILLER_51_47 VPWR VGND sg13g2_fill_2
XFILLER_18_103 VPWR VGND sg13g2_fill_1
XFILLER_14_397 VPWR VGND sg13g2_fill_1
X_2430_ _1008_ VPWR _0007_ VGND _1010_ _1011_ sg13g2_o21ai_1
X_2361_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q net952 net382 net980 _0623_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q
+ Inst_LUT4AB_switch_matrix.S1BEG2 VPWR VGND sg13g2_mux4_1
X_2292_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q _1084_ _0148_ _0308_ net981 Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0915_ VPWR VGND sg13g2_mux4_1
XFILLER_37_412 VPWR VGND sg13g2_fill_2
X_1243_ VGND VPWR _1074_ _1019_ _1072_ _1070_ _1075_ _1068_ sg13g2_a221oi_1
X_1312_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q net52 net1210 net107 Inst_LUT4AB_switch_matrix.JS2BEG1
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q _1140_ VPWR VGND sg13g2_mux4_1
XFILLER_52_415 VPWR VGND sg13g2_fill_2
XFILLER_20_301 VPWR VGND sg13g2_decap_8
XFILLER_20_334 VPWR VGND sg13g2_decap_4
Xoutput197 net197 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput186 net186 FrameData_O[3] VPWR VGND sg13g2_buf_1
Xoutput164 net164 FrameData_O[12] VPWR VGND sg13g2_buf_1
X_2559_ net1160 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
Xoutput142 net142 E6BEG[7] VPWR VGND sg13g2_buf_1
Xoutput153 net153 EE4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput175 net175 FrameData_O[22] VPWR VGND sg13g2_buf_1
X_2628_ net1145 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q VPWR VGND sg13g2_dlhq_1
Xoutput131 net131 E2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput120 net120 E2BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_23_150 VPWR VGND sg13g2_fill_2
X_1930_ net60 net62 net992 _0581_ VPWR VGND sg13g2_mux2_1
Xinput77 S2MID[6] net77 VPWR VGND sg13g2_buf_1
Xinput66 S2END[3] net66 VPWR VGND sg13g2_buf_1
X_1861_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0511_ _0514_ _0513_ sg13g2_a21oi_1
X_1792_ _0447_ _0440_ Inst_LUT4AB_switch_matrix.JW2BEG4 VPWR VGND sg13g2_nor2_2
Xinput22 EE4END[0] net22 VPWR VGND sg13g2_buf_1
Xinput11 E2END[5] net11 VPWR VGND sg13g2_buf_1
Xinput44 N2MID[1] net44 VPWR VGND sg13g2_buf_8
Xinput55 NN4END[0] net55 VPWR VGND sg13g2_buf_1
Xinput33 N1END[2] net33 VPWR VGND sg13g2_buf_1
Xinput88 W1END[1] net88 VPWR VGND sg13g2_buf_1
X_2344_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q _0589_ _0959_ _0958_ sg13g2_a21oi_1
X_2413_ _0998_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q net927 VPWR VGND sg13g2_nand2b_1
Xinput99 W2MID[1] net99 VPWR VGND sg13g2_buf_1
XFILLER_37_220 VPWR VGND sg13g2_fill_1
XFILLER_25_415 VPWR VGND sg13g2_fill_2
X_2275_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q _0899_ _0900_ VPWR VGND sg13g2_nor2_2
X_1226_ net1212 net65 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q _1059_ VPWR VGND sg13g2_mux2_1
XFILLER_43_289 VPWR VGND sg13g2_fill_1
XFILLER_43_223 VPWR VGND sg13g2_fill_2
XFILLER_28_275 VPWR VGND sg13g2_decap_4
Xfanout1120 net1122 net1120 VPWR VGND sg13g2_buf_1
Xfanout1131 FrameData[4] net1131 VPWR VGND sg13g2_buf_1
Xfanout1164 FrameData[23] net1164 VPWR VGND sg13g2_buf_1
Xfanout1197 FrameData[13] net1197 VPWR VGND sg13g2_buf_1
Xfanout1186 net1188 net1186 VPWR VGND sg13g2_buf_1
Xfanout1142 FrameData[2] net1142 VPWR VGND sg13g2_buf_1
X_2060_ VGND VPWR _1045_ _0702_ _0704_ _0703_ sg13g2_a21oi_1
Xfanout1153 FrameData[26] net1153 VPWR VGND sg13g2_buf_1
XFILLER_19_253 VPWR VGND sg13g2_fill_1
XFILLER_19_286 VPWR VGND sg13g2_decap_4
Xfanout1175 net1176 net1175 VPWR VGND sg13g2_buf_1
X_2962_ net1201 net1051 Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q VPWR VGND sg13g2_dlhq_1
X_1913_ _0537_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q _0563_ _0564_ VPWR VGND sg13g2_a21o_1
X_2893_ net1123 net1037 Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1844_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q VPWR _0497_ VGND net996 net933 sg13g2_o21ai_1
X_1775_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q VPWR _0431_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q
+ _0430_ sg13g2_o21ai_1
X_2327_ _0944_ VPWR _0945_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0556_
+ sg13g2_o21ai_1
X_2258_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q _0884_ _0885_ VPWR VGND sg13g2_nor2_1
X_1209_ VPWR _1042_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VGND sg13g2_inv_1
X_2189_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0822_ _0824_ _0823_ sg13g2_a21oi_1
XFILLER_16_267 VPWR VGND sg13g2_decap_8
X_1560_ _0224_ net997 net1004 VPWR VGND sg13g2_nand2b_1
XFILLER_39_304 VPWR VGND sg13g2_decap_4
X_1491_ _0157_ net990 Inst_LUT4AB_switch_matrix.M_AB VPWR VGND sg13g2_nand2b_1
X_2112_ _0751_ VPWR _0752_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q _0748_ sg13g2_o21ai_1
X_3230_ net74 net280 VPWR VGND sg13g2_buf_1
X_3161_ net1065 net202 VPWR VGND sg13g2_buf_1
X_3092_ E6END[11] net144 VPWR VGND sg13g2_buf_1
X_2043_ _0688_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ D VPWR VGND sg13g2_mux2_2
X_2876_ net1170 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1827_ _0481_ _0480_ _0476_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux _0479_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_30_292 VPWR VGND sg13g2_decap_4
X_2945_ net1155 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1689_ _0348_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ E VPWR VGND sg13g2_mux2_1
X_1758_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q _0413_ _0415_ _0414_ sg13g2_a21oi_1
Xfanout935 H net935 VPWR VGND sg13g2_buf_8
Xfanout957 net957 F VPWR VGND sg13g2_buf_16
Xfanout946 net946 net947 VPWR VGND sg13g2_buf_16
Xfanout979 A net979 VPWR VGND sg13g2_buf_1
Xfanout968 net970 net968 VPWR VGND sg13g2_buf_1
XFILLER_53_340 VPWR VGND sg13g2_fill_2
X_2730_ net1134 net1012 Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q VPWR VGND sg13g2_dlhq_1
X_2661_ net1139 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q VPWR VGND sg13g2_dlhq_1
X_1474_ _0141_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q net1006 VPWR VGND sg13g2_nand2b_1
X_1612_ _0274_ VPWR _0275_ VGND _0263_ _0257_ sg13g2_o21ai_1
XFILLER_8_296 VPWR VGND sg13g2_fill_2
X_1543_ _0083_ _0089_ _0080_ _0207_ VPWR VGND sg13g2_a21o_1
X_2592_ net1156 net1086 Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q VPWR VGND sg13g2_dlhq_1
X_3144_ net1058 net204 VPWR VGND sg13g2_buf_1
X_3075_ net14 net125 VPWR VGND sg13g2_buf_1
XFILLER_54_159 VPWR VGND sg13g2_fill_2
XFILLER_54_148 VPWR VGND sg13g2_fill_1
X_2026_ _0365_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q _0671_ _0672_ VPWR VGND sg13g2_a21o_1
X_2859_ net1131 net29 Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2928_ net1116 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_30_82 VPWR VGND sg13g2_fill_1
Xinput9 E2END[3] net9 VPWR VGND sg13g2_buf_1
X_1190_ VPWR _1023_ net110 VGND sg13g2_inv_1
X_2644_ net1195 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q VPWR VGND sg13g2_dlhq_1
X_2713_ net1181 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2575_ net1118 net1084 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
XFILLER_58_0 VPWR VGND sg13g2_fill_2
X_1526_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0190_ _0188_ _0184_ _0186_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q
+ _0191_ VPWR VGND sg13g2_mux4_1
Xoutput313 net313 SS4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput357 net357 WW4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput302 net302 SS4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput335 net335 W2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput346 net346 W6BEG[6] VPWR VGND sg13g2_buf_1
Xoutput324 net324 W2BEG[2] VPWR VGND sg13g2_buf_1
X_1457_ net1210 net66 net993 _0125_ VPWR VGND sg13g2_mux2_1
X_3127_ net1188 net168 VPWR VGND sg13g2_buf_1
X_1388_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _1121_ _0058_ VPWR VGND sg13g2_mux2_1
X_2009_ VPWR _0657_ _0656_ VGND sg13g2_inv_1
XFILLER_23_310 VPWR VGND sg13g2_fill_1
XFILLER_2_247 VPWR VGND sg13g2_fill_2
XFILLER_2_225 VPWR VGND sg13g2_fill_1
XFILLER_58_284 VPWR VGND sg13g2_fill_2
X_2291_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q net953 net936 net930 net928 Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0914_ VPWR VGND sg13g2_mux4_1
X_1311_ _1132_ _1129_ _1139_ Inst_LUT4AB_switch_matrix.JS2BEG1 VPWR VGND sg13g2_a21o_1
X_2360_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q net934 _1159_ Inst_LUT4AB_switch_matrix.E2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q Inst_LUT4AB_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_49_273 VPWR VGND sg13g2_fill_1
XFILLER_37_457 VPWR VGND sg13g2_fill_2
X_1242_ VGND VPWR _1017_ _1073_ _1074_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q sg13g2_a21oi_1
XFILLER_2_20 VPWR VGND sg13g2_fill_2
Xoutput143 net143 E6BEG[8] VPWR VGND sg13g2_buf_1
X_2627_ net1148 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q VPWR VGND sg13g2_dlhq_1
Xoutput132 net132 E2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput121 net121 E2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput198 net198 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput165 net165 FrameData_O[13] VPWR VGND sg13g2_buf_1
X_1509_ net976 net971 net989 _0174_ VPWR VGND sg13g2_mux2_1
X_2558_ net1163 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
Xoutput187 net187 FrameData_O[4] VPWR VGND sg13g2_buf_1
Xoutput176 net176 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput154 net154 EE4BEG[3] VPWR VGND sg13g2_buf_1
X_2489_ net1181 net1069 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_11_302 VPWR VGND sg13g2_fill_2
XFILLER_11_379 VPWR VGND sg13g2_fill_2
XFILLER_2_2 VPWR VGND sg13g2_fill_1
XFILLER_46_221 VPWR VGND sg13g2_decap_8
X_1860_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR _0513_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ _0512_ sg13g2_o21ai_1
XFILLER_14_173 VPWR VGND sg13g2_fill_2
Xinput67 S2END[4] net67 VPWR VGND sg13g2_buf_1
Xinput78 S2MID[7] net78 VPWR VGND sg13g2_buf_1
X_1791_ VGND VPWR _0446_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q _0445_ _1039_ _0447_
+ _0441_ sg13g2_a221oi_1
Xinput23 EE4END[1] net23 VPWR VGND sg13g2_buf_1
Xinput12 E2END[6] net12 VPWR VGND sg13g2_buf_1
Xinput45 N2MID[2] net45 VPWR VGND sg13g2_buf_1
Xinput56 NN4END[1] net56 VPWR VGND sg13g2_buf_1
Xinput34 N1END[3] net34 VPWR VGND sg13g2_buf_1
Xinput89 W1END[3] net89 VPWR VGND sg13g2_buf_1
X_2343_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q VPWR _0958_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ _0148_ sg13g2_o21ai_1
XFILLER_35_2 VPWR VGND sg13g2_fill_1
X_2412_ net392 _0997_ _0995_ _0003_ VPWR VGND sg13g2_mux2_1
X_2274_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q net1008 net1005 net1215 net957
+ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _0899_ VPWR VGND sg13g2_mux4_1
XFILLER_37_276 VPWR VGND sg13g2_decap_4
X_1225_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _1057_ _1058_ VPWR VGND sg13g2_nor2_1
X_1989_ _0637_ VPWR G VGND _0636_ Inst_LG_LUT4c_frame_config_dffesr.c_out_mux sg13g2_o21ai_1
XFILLER_40_419 VPWR VGND sg13g2_fill_2
XFILLER_57_69 VPWR VGND sg13g2_fill_1
Xfanout1121 net1122 net1121 VPWR VGND sg13g2_buf_1
Xfanout1165 net1167 net1165 VPWR VGND sg13g2_buf_1
Xfanout1132 FrameData[3] net1132 VPWR VGND sg13g2_buf_1
Xfanout1154 net1155 net1154 VPWR VGND sg13g2_buf_1
Xfanout1143 FrameData[2] net1143 VPWR VGND sg13g2_buf_1
Xfanout1110 net1112 net1110 VPWR VGND sg13g2_buf_1
Xfanout1198 net1200 net1198 VPWR VGND sg13g2_buf_1
Xfanout1187 net1188 net1187 VPWR VGND sg13g2_buf_1
Xfanout1176 net26 net1176 VPWR VGND sg13g2_buf_1
X_2961_ net1206 net1051 Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1843_ _0496_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ F VPWR VGND sg13g2_mux2_2
X_2892_ net1127 net1041 Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1912_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q VPWR _0563_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q
+ _0538_ sg13g2_o21ai_1
XFILLER_8_63 VPWR VGND sg13g2_fill_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_1774_ _0429_ VPWR _0430_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q _0426_ sg13g2_o21ai_1
XFILLER_57_338 VPWR VGND sg13g2_fill_1
X_2326_ _0944_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _1066_ VPWR VGND sg13g2_nand2_1
X_1208_ VPWR _1041_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VGND sg13g2_inv_1
X_2257_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q net31 net87 net1217 net970 Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ _0884_ VPWR VGND sg13g2_mux4_1
XFILLER_33_290 VPWR VGND sg13g2_fill_2
X_2188_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VPWR _0823_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ _0820_ sg13g2_o21ai_1
XFILLER_0_334 VPWR VGND sg13g2_fill_1
XFILLER_56_371 VPWR VGND sg13g2_fill_1
XFILLER_33_93 VPWR VGND sg13g2_decap_4
X_1490_ VGND VPWR net990 _1051_ _0156_ _0155_ sg13g2_a21oi_1
XFILLER_8_456 VPWR VGND sg13g2_fill_2
X_3091_ E6END[10] net143 VPWR VGND sg13g2_buf_1
X_2042_ _0687_ _0684_ _0682_ _0688_ VPWR VGND sg13g2_a21o_1
X_2111_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q _0750_ _0749_ _0751_ VPWR VGND sg13g2_nand3_1
X_3160_ FrameStrobe[17] net201 VPWR VGND sg13g2_buf_1
X_2875_ net1173 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1826_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q _0478_ _0480_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux
+ sg13g2_a21oi_1
X_2944_ net1156 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q VPWR VGND sg13g2_dlhq_1
Xfanout925 _0985_ net925 VPWR VGND sg13g2_buf_2
Xfanout947 net947 net948 VPWR VGND sg13g2_buf_16
Xfanout936 net937 net936 VPWR VGND sg13g2_buf_1
Xfanout958 net959 net958 VPWR VGND sg13g2_buf_2
X_1688_ _0348_ _0347_ _0342_ VPWR VGND sg13g2_nand2b_1
X_1757_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR _0414_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0411_ sg13g2_o21ai_1
X_2309_ Inst_LUT4AB_switch_matrix.EE4BEG2 _0927_ _0929_ _0925_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ VPWR VGND sg13g2_a22oi_1
X_3289_ W6END[3] net341 VPWR VGND sg13g2_buf_1
Xfanout969 net969 net970 VPWR VGND sg13g2_buf_16
XFILLER_48_135 VPWR VGND sg13g2_fill_1
XFILLER_0_175 VPWR VGND sg13g2_fill_1
XFILLER_0_197 VPWR VGND sg13g2_fill_1
XFILLER_44_374 VPWR VGND sg13g2_fill_1
X_1611_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q _0268_ _0273_ _0274_ VPWR VGND sg13g2_or3_1
X_2660_ net1146 net1095 Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q VPWR VGND sg13g2_dlhq_1
X_1473_ _0140_ _0139_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR VGND sg13g2_nand2b_1
X_3212_ Inst_LUT4AB_switch_matrix.NN4BEG1 net253 VPWR VGND sg13g2_buf_1
X_2591_ net1159 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q VPWR VGND sg13g2_dlhq_1
X_1542_ VPWR _0206_ _0205_ VGND sg13g2_inv_1
X_2025_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q VPWR _0671_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
+ _0366_ sg13g2_o21ai_1
X_3143_ FrameStrobe[0] net193 VPWR VGND sg13g2_buf_1
X_2927_ net1119 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VPWR VGND sg13g2_dlhq_1
XFILLER_40_39 VPWR VGND sg13g2_fill_1
X_2858_ net1132 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q VPWR VGND sg13g2_dlhq_1
X_1809_ _0202_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ net926 _0464_ VPWR VGND sg13g2_mux4_1
X_2789_ net1138 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_53_193 VPWR VGND sg13g2_fill_1
XFILLER_41_300 VPWR VGND sg13g2_decap_4
XFILLER_26_385 VPWR VGND sg13g2_decap_4
XFILLER_41_355 VPWR VGND sg13g2_fill_1
XFILLER_30_61 VPWR VGND sg13g2_fill_2
XFILLER_5_256 VPWR VGND sg13g2_fill_2
X_2574_ net1122 net1084 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
Xoutput303 net303 SS4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput314 net314 SS4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput325 net325 W2BEG[3] VPWR VGND sg13g2_buf_1
X_2643_ net1198 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q VPWR VGND sg13g2_dlhq_1
X_2712_ net1184 net1107 Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1525_ _0189_ VPWR _0190_ VGND net1009 net988 sg13g2_o21ai_1
X_1387_ VGND VPWR _1160_ _0053_ _0056_ _1124_ _0057_ _0008_ sg13g2_a221oi_1
Xoutput336 net336 W2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput347 net347 W6BEG[7] VPWR VGND sg13g2_buf_1
Xoutput358 net358 WW4BEG[2] VPWR VGND sg13g2_buf_1
X_1456_ _0123_ VPWR _0124_ VGND net93 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q sg13g2_o21ai_1
X_2008_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0649_ _0656_ VPWR VGND sg13g2_mux4_1
XFILLER_55_403 VPWR VGND sg13g2_fill_1
XFILLER_35_39 VPWR VGND sg13g2_fill_1
X_3126_ net1190 net167 VPWR VGND sg13g2_buf_1
XFILLER_23_355 VPWR VGND sg13g2_fill_1
XFILLER_41_174 VPWR VGND sg13g2_decap_4
X_2290_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q net943 net948 net965 net960 Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0913_ VPWR VGND sg13g2_mux4_1
X_1241_ net974 net968 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1073_ VPWR VGND sg13g2_mux2_1
X_1310_ VGND VPWR _1138_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q _1136_ _1027_ _1139_
+ _1134_ sg13g2_a221oi_1
XFILLER_32_163 VPWR VGND sg13g2_fill_1
Xoutput144 net144 E6BEG[9] VPWR VGND sg13g2_buf_1
Xoutput133 net133 E6BEG[0] VPWR VGND sg13g2_buf_1
X_2557_ net1166 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
Xoutput166 net166 FrameData_O[14] VPWR VGND sg13g2_buf_1
Xoutput177 net177 FrameData_O[24] VPWR VGND sg13g2_buf_1
X_2626_ net1152 net1089 Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q VPWR VGND sg13g2_dlhq_1
Xoutput155 net155 EE4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput122 Inst_LUT4AB_switch_matrix.E2BEG5 E2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput199 net199 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_1508_ _0172_ VPWR _0173_ VGND net989 net941 sg13g2_o21ai_1
Xoutput188 net188 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_46_49 VPWR VGND sg13g2_fill_2
X_2488_ net1184 net1070 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
X_1439_ _0091_ _0102_ _0107_ _0108_ VPWR VGND sg13g2_nor3_1
XFILLER_55_244 VPWR VGND sg13g2_fill_2
XFILLER_46_200 VPWR VGND sg13g2_fill_2
XFILLER_36_82 VPWR VGND sg13g2_fill_2
XFILLER_36_60 VPWR VGND sg13g2_fill_1
X_1790_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q _0443_ _0446_ _1039_ sg13g2_a21oi_1
Xinput13 E2END[7] net13 VPWR VGND sg13g2_buf_1
XFILLER_14_196 VPWR VGND sg13g2_fill_2
Xinput79 S4END[0] net79 VPWR VGND sg13g2_buf_1
Xinput68 S2END[5] net68 VPWR VGND sg13g2_buf_1
Xinput24 EE4END[2] net24 VPWR VGND sg13g2_buf_1
X_2411_ Inst_LC_LUT4c_frame_config_dffesr.c_reset_value _0467_ _0996_ _0997_ VPWR
+ VGND sg13g2_mux2_1
Xinput57 NN4END[2] net57 VPWR VGND sg13g2_buf_1
Xinput46 N2MID[3] net46 VPWR VGND sg13g2_buf_1
Xinput35 N2END[0] net35 VPWR VGND sg13g2_buf_1
X_2342_ _0957_ VPWR Inst_LUT4AB_switch_matrix.NN4BEG1 VGND _1050_ _0955_ sg13g2_o21ai_1
X_2273_ _0894_ _0897_ _0898_ VPWR VGND sg13g2_nor2_1
X_1224_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q net31 net37 net53 net8 Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ _1057_ VPWR VGND sg13g2_mux4_1
X_1988_ _0637_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_122 VPWR VGND sg13g2_fill_2
X_2609_ net1205 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_51 VPWR VGND sg13g2_fill_1
Xfanout1199 net1200 net1199 VPWR VGND sg13g2_buf_1
Xfanout1122 FrameData[7] net1122 VPWR VGND sg13g2_buf_1
Xfanout1177 net1179 net1177 VPWR VGND sg13g2_buf_1
Xfanout1166 net1167 net1166 VPWR VGND sg13g2_buf_1
Xfanout1188 FrameData[16] net1188 VPWR VGND sg13g2_buf_1
Xfanout1133 FrameData[3] net1133 VPWR VGND sg13g2_buf_1
Xfanout1144 FrameData[29] net1144 VPWR VGND sg13g2_buf_1
XFILLER_0_0 VPWR VGND sg13g2_fill_2
Xfanout1155 FrameData[26] net1155 VPWR VGND sg13g2_buf_1
Xfanout1100 net1101 net1100 VPWR VGND sg13g2_buf_1
Xfanout1111 net1112 net1111 VPWR VGND sg13g2_buf_1
X_2960_ net1116 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1911_ _0556_ _0561_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q _0562_ VPWR VGND sg13g2_mux2_1
X_2891_ net1129 net1041 Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VPWR VGND sg13g2_dlhq_1
X_1842_ _0492_ _0495_ _0473_ _0496_ VPWR VGND sg13g2_mux2_1
X_1773_ _0427_ _0428_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q _0429_ VPWR VGND sg13g2_nand3_1
X_2325_ VGND VPWR _0942_ _0943_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0276_
+ sg13g2_a21oi_2
X_1207_ VPWR _1040_ net25 VGND sg13g2_inv_1
X_2256_ _0879_ _0882_ _0883_ VPWR VGND sg13g2_nor2_1
X_2187_ _0821_ VPWR _0822_ VGND net1001 net932 sg13g2_o21ai_1
XFILLER_21_431 VPWR VGND sg13g2_fill_2
XFILLER_4_118 VPWR VGND sg13g2_fill_2
XFILLER_8_424 VPWR VGND sg13g2_fill_2
XFILLER_8_435 VPWR VGND sg13g2_fill_2
XFILLER_3_140 VPWR VGND sg13g2_fill_2
X_3090_ E6END[9] net142 VPWR VGND sg13g2_buf_1
X_2041_ _0679_ _0686_ _0687_ VPWR VGND sg13g2_and2_1
X_2110_ _0750_ Inst_LUT4AB_switch_matrix.JS2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_2943_ net1159 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VPWR VGND sg13g2_dlhq_1
X_2874_ net1177 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1825_ _0209_ _0311_ _0312_ _0479_ VPWR VGND sg13g2_a21o_1
X_1756_ _0412_ VPWR _0413_ VGND net93 net985 sg13g2_o21ai_1
Xfanout937 H net937 VPWR VGND sg13g2_buf_1
Xfanout948 net948 D VPWR VGND sg13g2_buf_16
Xfanout959 net960 net959 VPWR VGND sg13g2_buf_2
X_1687_ _0344_ _0346_ _0339_ _0347_ VPWR VGND sg13g2_nand3_1
X_2308_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q _0928_ _0929_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ sg13g2_a21oi_1
Xfanout926 _0395_ net926 VPWR VGND sg13g2_buf_1
XFILLER_57_158 VPWR VGND sg13g2_fill_2
XFILLER_53_342 VPWR VGND sg13g2_fill_1
X_2239_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q net33 net61 net1004 net959 Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ _0868_ VPWR VGND sg13g2_mux4_1
X_3288_ W6END[2] net338 VPWR VGND sg13g2_buf_1
XFILLER_21_272 VPWR VGND sg13g2_fill_2
XFILLER_36_309 VPWR VGND sg13g2_fill_2
X_1610_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0270_ _0273_ _0272_ sg13g2_a21oi_1
XFILLER_8_298 VPWR VGND sg13g2_fill_1
X_2590_ net1162 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1472_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q net32 net40 net1216 net11 Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0139_ VPWR VGND sg13g2_mux4_1
X_3211_ Inst_LUT4AB_switch_matrix.NN4BEG0 net252 VPWR VGND sg13g2_buf_1
X_1541_ _0205_ _0202_ _0203_ VPWR VGND sg13g2_nand2_1
X_3142_ net1137 net185 VPWR VGND sg13g2_buf_1
XFILLER_54_128 VPWR VGND sg13g2_fill_2
X_3073_ Inst_LUT4AB_switch_matrix.E2BEG6 net123 VPWR VGND sg13g2_buf_2
X_2024_ net965 net958 _0670_ Inst_LUT4AB_switch_matrix.M_EF VPWR VGND sg13g2_mux2_2
X_2857_ net1141 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q VPWR VGND sg13g2_dlhq_1
X_2926_ net1120 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1808_ _0401_ _0462_ _0460_ _0463_ VPWR VGND _0457_ sg13g2_nor4_2
X_1739_ _0396_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 net926 VPWR
+ VGND sg13g2_nand2_1
X_2788_ net1144 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_49_49 VPWR VGND sg13g2_fill_2
XFILLER_41_367 VPWR VGND sg13g2_fill_2
X_2711_ net1187 net1105 Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_58_2 VPWR VGND sg13g2_fill_1
X_2573_ net1124 net1083 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
X_1524_ _0189_ net988 net40 VPWR VGND sg13g2_nand2b_1
Xoutput337 net337 W2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput315 net315 SS4BEG[8] VPWR VGND sg13g2_buf_1
X_2642_ net1201 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q VPWR VGND sg13g2_dlhq_1
Xoutput304 Inst_LUT4AB_switch_matrix.SS4BEG0 SS4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput348 net348 W6BEG[8] VPWR VGND sg13g2_buf_1
Xoutput359 net359 WW4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput326 net326 W2BEG[4] VPWR VGND sg13g2_buf_1
X_1386_ _0055_ _0054_ _1085_ _0056_ VPWR VGND sg13g2_mux2_1
X_3125_ net1193 net166 VPWR VGND sg13g2_buf_1
X_1455_ _0123_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q net107 VPWR VGND sg13g2_nand2b_1
X_2007_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q _0617_ _0622_ _0626_ _0624_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q
+ _0655_ VPWR VGND sg13g2_mux4_1
X_2909_ net1165 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_41_120 VPWR VGND sg13g2_fill_2
XFILLER_26_172 VPWR VGND sg13g2_fill_2
X_1240_ _1072_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1071_ VPWR VGND sg13g2_nand2_1
XFILLER_37_437 VPWR VGND sg13g2_fill_2
XFILLER_32_153 VPWR VGND sg13g2_fill_1
Xoutput189 net189 FrameData_O[6] VPWR VGND sg13g2_buf_1
Xoutput112 net112 Co VPWR VGND sg13g2_buf_1
X_1507_ _0172_ net989 net946 VPWR VGND sg13g2_nand2b_1
Xoutput134 net134 E6BEG[10] VPWR VGND sg13g2_buf_1
X_2556_ net1169 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
Xoutput167 net167 FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput178 net178 FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput156 net156 EE4BEG[5] VPWR VGND sg13g2_buf_1
X_2625_ net1155 net1089 Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q VPWR VGND sg13g2_dlhq_1
Xoutput145 net145 EE4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput123 net123 E2BEG[6] VPWR VGND sg13g2_buf_1
X_2487_ net1187 net1068 Inst_LC_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
X_3108_ Inst_LUT4AB_switch_matrix.EE4BEG1 net149 VPWR VGND sg13g2_buf_1
XFILLER_28_426 VPWR VGND sg13g2_fill_2
X_1369_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q _0037_ _0039_ _0038_ sg13g2_a21oi_1
X_1438_ _0073_ _0103_ _0104_ _0106_ _0107_ VPWR VGND sg13g2_nor4_1
XFILLER_43_429 VPWR VGND sg13g2_fill_1
XFILLER_11_304 VPWR VGND sg13g2_fill_1
X_3039_ net1159 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_46_245 VPWR VGND sg13g2_fill_2
XFILLER_36_50 VPWR VGND sg13g2_decap_4
XFILLER_52_82 VPWR VGND sg13g2_fill_1
Xinput25 EE4END[3] net25 VPWR VGND sg13g2_buf_1
Xinput14 E2MID[0] net14 VPWR VGND sg13g2_buf_1
Xinput36 N2END[1] net36 VPWR VGND sg13g2_buf_1
Xinput69 S2END[6] net69 VPWR VGND sg13g2_buf_1
X_2341_ _0957_ _1050_ _0956_ VPWR VGND sg13g2_nand2_1
Xinput58 NN4END[3] net58 VPWR VGND sg13g2_buf_1
Xinput47 N2MID[4] net47 VPWR VGND sg13g2_buf_1
X_2410_ _0996_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q net925 VPWR VGND sg13g2_nand2_1
XFILLER_37_201 VPWR VGND sg13g2_decap_4
X_2272_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q VPWR _0897_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ _0896_ sg13g2_o21ai_1
X_1223_ _1056_ _1055_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VPWR VGND sg13g2_nand2_2
XFILLER_37_267 VPWR VGND sg13g2_fill_1
X_1987_ VGND VPWR _0630_ _0636_ _0635_ _0632_ sg13g2_a21oi_2
X_2539_ net1129 net1077 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_2608_ net1116 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q VPWR VGND sg13g2_dlhq_1
XFILLER_43_259 VPWR VGND sg13g2_fill_2
XFILLER_59_381 VPWR VGND sg13g2_fill_1
Xfanout1178 net1179 net1178 VPWR VGND sg13g2_buf_1
Xfanout1123 net1125 net1123 VPWR VGND sg13g2_buf_1
Xfanout1189 net1191 net1189 VPWR VGND sg13g2_buf_1
Xfanout1167 FrameData[22] net1167 VPWR VGND sg13g2_buf_1
Xfanout1134 FrameData[3] net1134 VPWR VGND sg13g2_buf_1
Xfanout1156 net1158 net1156 VPWR VGND sg13g2_buf_1
Xfanout1145 FrameData[29] net1145 VPWR VGND sg13g2_buf_1
Xfanout1101 net1102 net1101 VPWR VGND sg13g2_buf_1
Xfanout1112 FrameStrobe[0] net1112 VPWR VGND sg13g2_buf_1
X_2890_ net1132 net1041 Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q VPWR VGND sg13g2_dlhq_1
X_1910_ _0560_ VPWR _0561_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q _0557_ sg13g2_o21ai_1
XFILLER_34_215 VPWR VGND sg13g2_fill_1
X_1841_ _0493_ _0494_ _0486_ _0495_ VPWR VGND sg13g2_mux2_1
X_1772_ _0428_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q net90 VPWR VGND sg13g2_nand2_1
XFILLER_6_160 VPWR VGND sg13g2_fill_1
X_2324_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q net967 _0942_ VPWR VGND sg13g2_nor2_1
XFILLER_40_2 VPWR VGND sg13g2_fill_1
XFILLER_26_0 VPWR VGND sg13g2_fill_2
X_1206_ VPWR _1039_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VGND sg13g2_inv_1
XFILLER_27_19 VPWR VGND sg13g2_fill_1
X_2255_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q VPWR _0882_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
+ _0881_ sg13g2_o21ai_1
X_2186_ _0821_ net1001 net930 VPWR VGND sg13g2_nand2_1
XFILLER_8_458 VPWR VGND sg13g2_fill_1
X_2040_ _0686_ _0676_ _0685_ VPWR VGND sg13g2_nand2b_1
X_2873_ net1180 net1035 Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2942_ net1162 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_22_207 VPWR VGND sg13g2_fill_2
X_1686_ _0346_ _0247_ _0345_ VPWR VGND sg13g2_nand2b_1
X_1824_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q _0238_ _0478_ _0477_ sg13g2_a21oi_1
X_1755_ _0412_ _1028_ net985 VPWR VGND sg13g2_nand2_1
Xfanout927 _0973_ net927 VPWR VGND sg13g2_buf_8
X_2238_ _0867_ VPWR Inst_LUT4AB_switch_matrix.WW4BEG1 VGND _1048_ _0865_ sg13g2_o21ai_1
X_3287_ net105 net337 VPWR VGND sg13g2_buf_1
X_2307_ net59 net973 Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0928_ VPWR VGND sg13g2_mux2_1
Xfanout938 net939 net938 VPWR VGND sg13g2_buf_2
X_2169_ _0804_ VPWR _0805_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0803_ sg13g2_o21ai_1
XFILLER_0_155 VPWR VGND sg13g2_fill_2
X_1540_ VGND VPWR _0204_ _0203_ _0202_ sg13g2_or2_1
XFILLER_8_266 VPWR VGND sg13g2_fill_1
X_3141_ net1140 net184 VPWR VGND sg13g2_buf_1
X_1471_ _0137_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q _0138_ VPWR VGND sg13g2_nor2b_1
X_3210_ NN4END[15] net251 VPWR VGND sg13g2_buf_1
XFILLER_39_126 VPWR VGND sg13g2_decap_4
X_2023_ _0668_ _0669_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0670_ VPWR VGND
+ sg13g2_mux2_1
X_2856_ net26 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q VPWR VGND sg13g2_dlhq_1
X_1807_ _0398_ VPWR _0462_ VGND _0204_ _0461_ sg13g2_o21ai_1
X_2925_ net1123 net1042 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1738_ _0394_ _0207_ Inst_LC_LUT4c_frame_config_dffesr.c_I0mux _0395_ VPWR VGND sg13g2_mux2_1
X_2787_ net1147 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1669_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q net14 net71 net98 net377 Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q
+ _0329_ VPWR VGND sg13g2_mux4_1
XFILLER_5_258 VPWR VGND sg13g2_fill_1
XFILLER_49_457 VPWR VGND sg13g2_fill_2
XFILLER_32_324 VPWR VGND sg13g2_decap_4
X_2710_ net1190 net1105 Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2572_ net1127 net1084 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
X_1523_ _0187_ VPWR _0188_ VGND net1216 net988 sg13g2_o21ai_1
Xoutput305 net305 SS4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput316 net316 SS4BEG[9] VPWR VGND sg13g2_buf_1
X_2641_ net1206 net1093 Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q VPWR VGND sg13g2_dlhq_1
Xoutput327 net327 W2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput338 net338 W6BEG[0] VPWR VGND sg13g2_buf_1
X_1454_ _0122_ _1032_ _0121_ VPWR VGND sg13g2_nand2_1
Xoutput349 net349 W6BEG[9] VPWR VGND sg13g2_buf_1
X_3124_ net1196 net165 VPWR VGND sg13g2_buf_1
X_1385_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ net982 _0055_ VPWR VGND sg13g2_mux2_1
X_2006_ _0645_ net388 _0653_ _0654_ VPWR VGND sg13g2_a21o_1
X_2908_ net1168 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2839_ net1187 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_26_195 VPWR VGND sg13g2_decap_4
XFILLER_49_221 VPWR VGND sg13g2_fill_1
XFILLER_32_110 VPWR VGND sg13g2_fill_2
XFILLER_17_140 VPWR VGND sg13g2_fill_1
X_2624_ net1158 net1089 Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q VPWR VGND sg13g2_dlhq_1
XFILLER_20_338 VPWR VGND sg13g2_fill_1
XFILLER_56_0 VPWR VGND sg13g2_fill_2
X_2555_ net1172 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
Xoutput135 Inst_LUT4AB_switch_matrix.E6BEG1 E6BEG[11] VPWR VGND sg13g2_buf_1
Xoutput157 net157 EE4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput146 net146 EE4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput179 net179 FrameData_O[26] VPWR VGND sg13g2_buf_1
Xoutput168 net168 FrameData_O[16] VPWR VGND sg13g2_buf_1
Xoutput124 Inst_LUT4AB_switch_matrix.E2BEG7 E2BEG[7] VPWR VGND sg13g2_buf_1
X_1506_ VPWR _0171_ _0170_ VGND sg13g2_inv_1
X_2486_ net1190 net1068 Inst_LC_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_1437_ _0105_ VPWR _0106_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0083_ sg13g2_o21ai_1
Xoutput113 net113 E1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_55_246 VPWR VGND sg13g2_fill_1
X_3107_ Inst_LUT4AB_switch_matrix.EE4BEG0 net148 VPWR VGND sg13g2_buf_1
X_3038_ net1164 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1299_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _1127_ _1128_ _1027_ sg13g2_a21oi_1
X_1368_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VPWR _0038_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ net71 sg13g2_o21ai_1
XFILLER_23_143 VPWR VGND sg13g2_decap_8
XFILLER_36_84 VPWR VGND sg13g2_fill_1
Xinput59 S1END[0] net59 VPWR VGND sg13g2_buf_1
Xinput26 FrameData[1] net26 VPWR VGND sg13g2_buf_1
Xinput48 N2MID[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_6_320 VPWR VGND sg13g2_fill_1
XFILLER_6_342 VPWR VGND sg13g2_fill_1
Xinput37 N2END[2] net37 VPWR VGND sg13g2_buf_1
Xinput15 net15 E2MID[1] VPWR VGND sg13g2_buf_16
X_2340_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q net1007 net1214 net1003 net978 Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ _0956_ VPWR VGND sg13g2_mux4_1
X_2271_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _1084_ _0896_ _0895_
+ sg13g2_a21oi_1
X_1222_ _1053_ _1054_ _1020_ _1055_ VPWR VGND sg13g2_mux2_1
XFILLER_52_249 VPWR VGND sg13g2_fill_2
X_1986_ _0627_ _0634_ _0635_ VPWR VGND sg13g2_nor2_1
X_2607_ net1118 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VPWR VGND sg13g2_dlhq_1
X_2538_ net1133 net1077 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2469_ net1139 net1064 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_28_279 VPWR VGND sg13g2_fill_1
XFILLER_28_268 VPWR VGND sg13g2_decap_8
Xfanout1113 FrameStrobe[0] net1113 VPWR VGND sg13g2_buf_1
XFILLER_0_2 VPWR VGND sg13g2_fill_1
Xfanout1102 net27 net1102 VPWR VGND sg13g2_buf_1
Xfanout1179 FrameData[19] net1179 VPWR VGND sg13g2_buf_1
Xfanout1124 net1125 net1124 VPWR VGND sg13g2_buf_1
Xfanout1168 net1170 net1168 VPWR VGND sg13g2_buf_1
Xfanout1157 net1158 net1157 VPWR VGND sg13g2_buf_1
Xfanout1146 FrameData[29] net1146 VPWR VGND sg13g2_buf_1
Xfanout1135 net1136 net1135 VPWR VGND sg13g2_buf_1
XFILLER_19_235 VPWR VGND sg13g2_fill_1
XFILLER_19_279 VPWR VGND sg13g2_decap_8
X_1840_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0487_ _0494_ VPWR VGND sg13g2_mux4_1
X_1771_ _0427_ net63 Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q VPWR VGND sg13g2_nand2b_1
X_2323_ net1006 net948 Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0941_ VPWR VGND
+ sg13g2_mux2_1
X_2254_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q _0308_ _0881_ _0880_ sg13g2_a21oi_1
X_1205_ VPWR _1038_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VGND sg13g2_inv_1
XFILLER_25_238 VPWR VGND sg13g2_fill_2
XFILLER_19_0 VPWR VGND sg13g2_fill_2
X_2185_ VGND VPWR net1001 net951 _0820_ _0819_ sg13g2_a21oi_1
X_1969_ net44 net15 Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q _0618_ VPWR VGND sg13g2_mux2_1
XFILLER_8_426 VPWR VGND sg13g2_fill_1
XFILLER_8_437 VPWR VGND sg13g2_fill_1
XFILLER_3_153 VPWR VGND sg13g2_fill_2
XFILLER_3_142 VPWR VGND sg13g2_fill_1
X_1823_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q _0239_ _0477_ VPWR VGND sg13g2_nor2b_1
X_2941_ net1165 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2872_ net1183 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q VPWR VGND sg13g2_dlhq_1
X_1685_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0310_ _0345_ VPWR VGND sg13g2_mux4_1
X_1754_ net82 net86 Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q _0411_ VPWR VGND sg13g2_mux2_1
X_3286_ net104 net336 VPWR VGND sg13g2_buf_1
Xfanout928 Inst_LUT4AB_switch_matrix.M_AH net928 VPWR VGND sg13g2_buf_1
X_2237_ _0867_ _1048_ _0866_ VPWR VGND sg13g2_nand2_1
X_2306_ _0926_ VPWR _0927_ VGND net1010 Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ sg13g2_o21ai_1
Xfanout939 net940 net939 VPWR VGND sg13g2_buf_2
X_2099_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q net1010 net35 net1217 net6 Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ _0740_ VPWR VGND sg13g2_mux4_1
X_2168_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0801_ _0804_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
+ sg13g2_a21oi_1
XFILLER_21_274 VPWR VGND sg13g2_fill_1
XFILLER_29_385 VPWR VGND sg13g2_fill_1
XFILLER_44_388 VPWR VGND sg13g2_fill_1
X_1470_ VGND VPWR _0136_ _0137_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0135_ sg13g2_a21oi_2
X_3140_ net1145 net182 VPWR VGND sg13g2_buf_1
X_3071_ Inst_LUT4AB_switch_matrix.E2BEG4 net121 VPWR VGND sg13g2_buf_2
X_2022_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_switch_matrix.JW2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q _0669_ VPWR VGND sg13g2_mux4_1
XFILLER_35_399 VPWR VGND sg13g2_fill_1
XFILLER_35_300 VPWR VGND sg13g2_decap_8
X_2855_ net1208 net1034 Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2786_ net1150 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2924_ net1126 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1806_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ net926 _0461_ VPWR VGND sg13g2_mux2_1
X_1599_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VPWR _0262_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0259_ sg13g2_o21ai_1
X_1668_ Inst_LUT4AB_switch_matrix.JW2BEG5 _0322_ _0328_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
+ _0320_ VPWR VGND sg13g2_a22oi_1
X_1737_ _0394_ _0393_ _0368_ VPWR VGND sg13g2_nand2b_1
XFILLER_53_130 VPWR VGND sg13g2_fill_2
XFILLER_26_355 VPWR VGND sg13g2_fill_2
X_3269_ Inst_LUT4AB_switch_matrix.W1BEG1 net319 VPWR VGND sg13g2_buf_1
XFILLER_41_369 VPWR VGND sg13g2_fill_1
XFILLER_5_215 VPWR VGND sg13g2_fill_1
XFILLER_32_314 VPWR VGND sg13g2_fill_1
XFILLER_29_193 VPWR VGND sg13g2_decap_4
XFILLER_17_322 VPWR VGND sg13g2_decap_8
XFILLER_17_333 VPWR VGND sg13g2_fill_1
X_2640_ net1116 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q VPWR VGND sg13g2_dlhq_1
Xoutput317 net317 UserCLKo VPWR VGND sg13g2_buf_1
X_2571_ net1130 net1083 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
X_1522_ _0187_ net988 net11 VPWR VGND sg13g2_nand2b_1
Xoutput306 net306 SS4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput328 net328 W2BEG[6] VPWR VGND sg13g2_buf_1
X_1453_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q net1009 net54 net38 net9 net993 _0121_
+ VPWR VGND sg13g2_mux4_1
Xoutput339 Inst_LUT4AB_switch_matrix.W6BEG0 W6BEG[10] VPWR VGND sg13g2_buf_1
X_2005_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ net379 _0653_ VPWR VGND sg13g2_mux4_1
X_3123_ net1199 net164 VPWR VGND sg13g2_buf_1
X_3054_ UserCLK net372 _0007_ _3054_/Q_N Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
X_1384_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ net982 _0054_ VPWR VGND sg13g2_mux2_1
X_2907_ net1171 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_19 VPWR VGND sg13g2_fill_2
XFILLER_50_188 VPWR VGND sg13g2_fill_2
X_2769_ net1204 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q VPWR VGND sg13g2_dlhq_1
X_2838_ net1190 net1030 Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_41_111 VPWR VGND sg13g2_fill_1
XFILLER_41_199 VPWR VGND sg13g2_fill_2
XFILLER_25_75 VPWR VGND sg13g2_fill_1
XFILLER_37_439 VPWR VGND sg13g2_fill_1
XFILLER_32_133 VPWR VGND sg13g2_fill_2
X_2554_ net1179 net1081 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
X_2623_ net1160 net1089 Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q VPWR VGND sg13g2_dlhq_1
Xoutput125 net125 E2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput114 net114 E1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_49_0 VPWR VGND sg13g2_fill_2
Xoutput169 net169 FrameData_O[17] VPWR VGND sg13g2_buf_1
Xoutput147 net147 EE4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput136 net136 E6BEG[1] VPWR VGND sg13g2_buf_1
Xoutput158 net158 EE4BEG[7] VPWR VGND sg13g2_buf_1
X_1505_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q net39 net10 net85 net94 Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q
+ _0170_ VPWR VGND sg13g2_mux4_1
X_1367_ VPWR Inst_LUT4AB_switch_matrix.JW2BEG3 _0037_ VGND sg13g2_inv_1
X_1436_ _0105_ _0078_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_nand2b_1
X_2485_ net1193 net1068 Inst_LC_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
X_3106_ EE4END[15] net147 VPWR VGND sg13g2_buf_1
XFILLER_46_19 VPWR VGND sg13g2_fill_2
X_3037_ net1167 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_28_428 VPWR VGND sg13g2_fill_1
X_1298_ net935 net929 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _1127_ VPWR VGND sg13g2_mux2_1
XFILLER_23_177 VPWR VGND sg13g2_fill_2
XFILLER_46_247 VPWR VGND sg13g2_fill_1
Xinput38 N2END[3] net38 VPWR VGND sg13g2_buf_1
Xinput49 N2MID[6] net49 VPWR VGND sg13g2_buf_1
Xinput27 FrameStrobe[11] net27 VPWR VGND sg13g2_buf_1
Xinput16 E2MID[2] net16 VPWR VGND sg13g2_buf_1
X_2270_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q net952 _0895_ VPWR VGND sg13g2_nor2b_1
X_1221_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q net975 net945 net940 net962 Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ _1054_ VPWR VGND sg13g2_mux4_1
X_1985_ _0532_ _0633_ _0634_ VPWR VGND sg13g2_nor2_1
X_2606_ net1120 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q VPWR VGND sg13g2_dlhq_1
X_2537_ net1142 net1077 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2399_ _0974_ VPWR _0988_ VGND Inst_LH_LUT4c_frame_config_dffesr.c_reset_value _0986_
+ sg13g2_o21ai_1
X_1419_ _1085_ VPWR _0088_ VGND net1 _1160_ sg13g2_o21ai_1
X_2468_ net1144 net1065 Inst_LB_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
XFILLER_22_87 VPWR VGND sg13g2_fill_1
Xfanout1125 FrameData[6] net1125 VPWR VGND sg13g2_buf_1
Xfanout1114 FrameData[9] net1114 VPWR VGND sg13g2_buf_1
Xfanout1147 net1148 net1147 VPWR VGND sg13g2_buf_1
XFILLER_3_335 VPWR VGND sg13g2_fill_2
Xfanout1103 net1104 net1103 VPWR VGND sg13g2_buf_1
Xfanout1136 net1137 net1136 VPWR VGND sg13g2_buf_1
Xfanout1169 net1170 net1169 VPWR VGND sg13g2_buf_1
Xfanout1158 FrameData[25] net1158 VPWR VGND sg13g2_buf_1
XFILLER_42_283 VPWR VGND sg13g2_fill_2
X_1770_ net35 net23 Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q _0426_ VPWR VGND sg13g2_mux2_1
X_2322_ net1009 net1216 Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0940_ VPWR VGND
+ sg13g2_mux2_1
X_1204_ VPWR _1037_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VGND sg13g2_inv_1
X_2184_ net1001 net956 _0819_ VPWR VGND sg13g2_nor2b_1
X_2253_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q net940 _0880_ VPWR VGND sg13g2_nor2b_1
X_1899_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q _0548_ _0551_ _1044_ sg13g2_a21oi_1
X_1968_ _0615_ VPWR _0617_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q _0616_ sg13g2_o21ai_1
XFILLER_33_97 VPWR VGND sg13g2_fill_1
X_2940_ net1168 net1044 Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1822_ VGND VPWR _0476_ _0475_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q sg13g2_or2_1
XFILLER_30_231 VPWR VGND sg13g2_fill_1
X_1753_ _0409_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q _0410_ VPWR VGND sg13g2_nor2b_1
X_2871_ net1186 net1032 Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q VPWR VGND sg13g2_dlhq_1
Xfanout929 Inst_LUT4AB_switch_matrix.M_EF net929 VPWR VGND sg13g2_buf_2
X_1684_ VGND VPWR _0344_ _0343_ _0247_ sg13g2_or2_1
X_2236_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q net1007 net62 net1003 net977 Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ _0866_ VPWR VGND sg13g2_mux4_1
X_3285_ net103 net335 VPWR VGND sg13g2_buf_1
X_2305_ VGND VPWR _1016_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0926_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ sg13g2_a21oi_1
X_2167_ VGND VPWR net994 net938 _0803_ _0802_ sg13g2_a21oi_1
X_2098_ _0738_ VPWR _0739_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0736_ sg13g2_o21ai_1
XFILLER_0_157 VPWR VGND sg13g2_fill_1
XFILLER_29_331 VPWR VGND sg13g2_fill_2
XFILLER_4_452 VPWR VGND sg13g2_fill_2
X_2021_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q Inst_LUT4AB_switch_matrix.JN2BEG6
+ Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_switch_matrix.JW2BEG6
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q _0668_ VPWR VGND sg13g2_mux4_1
X_3070_ Inst_LUT4AB_switch_matrix.E2BEG3 net120 VPWR VGND sg13g2_buf_1
XFILLER_35_367 VPWR VGND sg13g2_fill_2
X_2923_ net1131 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2785_ net1153 net1020 Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q VPWR VGND sg13g2_dlhq_1
X_1736_ _0392_ VPWR _0393_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q _0389_
+ sg13g2_o21ai_1
X_2854_ net1136 net1031 Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1805_ VGND VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 net926
+ _0460_ _0459_ sg13g2_a21oi_1
X_3053__373 VPWR VGND net373 sg13g2_tiehi
XFILLER_49_19 VPWR VGND sg13g2_fill_1
X_1598_ _0260_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0261_ VPWR VGND sg13g2_nor2b_1
X_1667_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q _0327_ _0328_ VPWR VGND sg13g2_nor2_1
X_3199_ NN4END[4] net249 VPWR VGND sg13g2_buf_1
XFILLER_41_304 VPWR VGND sg13g2_fill_2
X_2219_ net1009 net60 Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0851_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_26_378 VPWR VGND sg13g2_decap_8
X_3268_ Inst_LUT4AB_switch_matrix.W1BEG0 net318 VPWR VGND sg13g2_buf_1
XFILLER_5_249 VPWR VGND sg13g2_fill_2
XFILLER_39_96 VPWR VGND sg13g2_decap_4
X_2570_ net1132 net1083 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
Xoutput307 Inst_LUT4AB_switch_matrix.SS4BEG3 SS4BEG[15] VPWR VGND sg13g2_buf_1
X_3122_ net1202 net163 VPWR VGND sg13g2_buf_1
X_1521_ _0185_ VPWR _0186_ VGND net1006 net989 sg13g2_o21ai_1
X_1383_ VGND VPWR _0049_ _0050_ _0053_ _0052_ sg13g2_a21oi_1
Xoutput329 net329 W2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput318 net318 W1BEG[0] VPWR VGND sg13g2_buf_1
X_1452_ _1033_ _0114_ _0119_ _0120_ VPWR VGND sg13g2_nor3_1
X_2004_ _0649_ _0650_ _0652_ VPWR VGND sg13g2_nor2_2
X_3053_ UserCLK net373 _0006_ _3053_/Q_N Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
X_2906_ net1177 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1719_ _0376_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q _0377_ VPWR VGND sg13g2_nor2b_1
X_2768_ net1115 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q VPWR VGND sg13g2_dlhq_1
X_2837_ net1193 net1030 Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2699_ net1131 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_46_407 VPWR VGND sg13g2_fill_2
XFILLER_41_167 VPWR VGND sg13g2_decap_8
XFILLER_41_53 VPWR VGND sg13g2_fill_1
XFILLER_1_252 VPWR VGND sg13g2_fill_2
X_2553_ net1182 net1080 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
Xoutput148 net148 EE4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput137 net137 E6BEG[2] VPWR VGND sg13g2_buf_1
X_2622_ net1164 net1089 Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q VPWR VGND sg13g2_dlhq_1
Xoutput159 net159 EE4BEG[8] VPWR VGND sg13g2_buf_1
X_1504_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q net56 net23 net80 Inst_LUT4AB_switch_matrix.JS2BEG2
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q _0169_ VPWR VGND sg13g2_mux4_1
Xoutput115 Inst_LUT4AB_switch_matrix.E1BEG2 E1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput126 net126 E2BEGb[1] VPWR VGND sg13g2_buf_1
X_3105_ EE4END[14] net146 VPWR VGND sg13g2_buf_1
X_1366_ _0027_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q _0036_ _0037_ VPWR VGND sg13g2_a21o_2
X_1435_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0081_ _0104_ VPWR
+ VGND sg13g2_nor2_1
X_2484_ net1196 net1067 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_237 VPWR VGND sg13g2_fill_2
XFILLER_51_432 VPWR VGND sg13g2_fill_2
X_3036_ net1170 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1297_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q net951 _1126_ _1125_ sg13g2_a21oi_1
XFILLER_11_67 VPWR VGND sg13g2_fill_2
XFILLER_36_31 VPWR VGND sg13g2_fill_2
XFILLER_52_41 VPWR VGND sg13g2_fill_2
Xinput39 N2END[4] net39 VPWR VGND sg13g2_buf_1
XFILLER_6_377 VPWR VGND sg13g2_fill_1
Xinput28 FrameStrobe[19] net28 VPWR VGND sg13g2_buf_1
Xinput17 E2MID[3] net17 VPWR VGND sg13g2_buf_1
X_1220_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q net957 net950 net935 net930 Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q
+ _1053_ VPWR VGND sg13g2_mux4_1
X_1984_ net378 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ net374 _0633_ VPWR VGND sg13g2_mux4_1
X_2605_ net1125 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2536_ net26 net1078 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 VPWR
+ VGND sg13g2_dlhq_1
X_2467_ net1147 net1065 Inst_LB_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_2398_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q _0659_ _0985_ _0665_ _0987_
+ _0661_ sg13g2_a221oi_1
X_1418_ _0087_ net1 _1160_ VPWR VGND sg13g2_nand2_1
X_1349_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q _0012_ _0020_ _0021_ VPWR VGND sg13g2_a21o_2
XFILLER_36_281 VPWR VGND sg13g2_decap_8
X_3019_ net1131 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q VPWR VGND sg13g2_dlhq_1
Xfanout1137 FrameData[31] net1137 VPWR VGND sg13g2_buf_1
Xfanout1115 FrameData[9] net1115 VPWR VGND sg13g2_buf_1
Xfanout1159 net1161 net1159 VPWR VGND sg13g2_buf_1
Xfanout1148 net1149 net1148 VPWR VGND sg13g2_buf_1
Xfanout1126 net1128 net1126 VPWR VGND sg13g2_buf_1
Xfanout1104 net1105 net1104 VPWR VGND sg13g2_buf_1
XFILLER_30_435 VPWR VGND sg13g2_fill_2
XFILLER_8_68 VPWR VGND sg13g2_fill_1
X_2321_ _0937_ _0939_ Inst_LUT4AB_switch_matrix.EE4BEG0 VPWR VGND sg13g2_nor2_1
XFILLER_33_4 VPWR VGND sg13g2_fill_2
X_1203_ VPWR _1036_ net80 VGND sg13g2_inv_1
XFILLER_19_2 VPWR VGND sg13g2_fill_1
X_2183_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q net968 net944 net938 net961 net1001
+ _0818_ VPWR VGND sg13g2_mux4_1
X_2252_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q _0430_ _0879_ _0878_ sg13g2_a21oi_1
XFILLER_33_284 VPWR VGND sg13g2_fill_2
XFILLER_18_270 VPWR VGND sg13g2_fill_2
XFILLER_21_424 VPWR VGND sg13g2_fill_2
X_1898_ VGND VPWR _0550_ _0549_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q sg13g2_or2_1
X_1967_ net43 net14 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q _0616_ VPWR VGND sg13g2_mux2_1
XFILLER_21_457 VPWR VGND sg13g2_fill_2
X_2519_ net1188 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_44 VPWR VGND sg13g2_fill_1
XFILLER_17_66 VPWR VGND sg13g2_fill_1
X_2870_ net1189 net1036 Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1683_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0310_ _0343_ VPWR VGND sg13g2_mux4_1
X_1821_ _0474_ VPWR _0475_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q _0236_ sg13g2_o21ai_1
X_1752_ VGND VPWR _0408_ _0409_ _0407_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q sg13g2_a21oi_2
X_3284_ net102 net334 VPWR VGND sg13g2_buf_1
X_2304_ VPWR _0925_ _0924_ VGND sg13g2_inv_1
XFILLER_24_0 VPWR VGND sg13g2_fill_2
X_2235_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q net932 _1158_ _0196_ _0253_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ _0865_ VPWR VGND sg13g2_mux4_1
X_2097_ _0738_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0737_ VPWR VGND sg13g2_nand2b_1
X_2166_ net994 net968 _0802_ VPWR VGND sg13g2_nor2b_1
X_2999_ net1186 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VPWR VGND sg13g2_dlhq_1
XFILLER_44_368 VPWR VGND sg13g2_fill_2
XFILLER_29_365 VPWR VGND sg13g2_fill_2
X_2020_ _0667_ VPWR H VGND _0666_ Inst_LH_LUT4c_frame_config_dffesr.c_out_mux sg13g2_o21ai_1
XFILLER_47_162 VPWR VGND sg13g2_fill_2
XFILLER_39_118 VPWR VGND sg13g2_decap_4
X_2922_ net1134 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q VPWR VGND sg13g2_dlhq_1
X_2853_ net1139 net1031 Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q VPWR VGND sg13g2_dlhq_1
X_1666_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0324_ _0327_ _0326_ sg13g2_a21oi_1
X_2784_ net1158 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1735_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q _0391_ _0392_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q
+ sg13g2_a21oi_1
X_1804_ _0458_ _0202_ _0459_ VPWR VGND _0203_ sg13g2_nand3b_1
X_3267_ UserCLK net317 VPWR VGND sg13g2_buf_1
X_1597_ net936 Inst_LUT4AB_switch_matrix.M_EF net987 _0260_ VPWR VGND sg13g2_mux2_1
XFILLER_38_140 VPWR VGND sg13g2_fill_1
X_2218_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q _0847_ _0848_ _0849_ _0850_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
+ Inst_LUT4AB_switch_matrix.W6BEG0 VPWR VGND sg13g2_mux4_1
X_2149_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VPWR _0786_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q
+ _0779_ sg13g2_o21ai_1
XFILLER_29_173 VPWR VGND sg13g2_fill_2
XFILLER_44_143 VPWR VGND sg13g2_fill_1
X_1520_ _0185_ net988 net89 VPWR VGND sg13g2_nand2b_1
Xoutput308 net308 SS4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput319 net319 W1BEG[1] VPWR VGND sg13g2_buf_1
X_3121_ net1204 net162 VPWR VGND sg13g2_buf_1
X_1382_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q _0022_ _0052_ _0051_ sg13g2_a21oi_1
X_1451_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0116_ _0119_ _0118_ sg13g2_a21oi_1
X_2003_ _0651_ _0649_ _0650_ VPWR VGND sg13g2_nand2_1
X_3052_ UserCLK net366 _0005_ _3052_/Q_N Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
XFILLER_35_121 VPWR VGND sg13g2_fill_1
X_2905_ net1180 net1041 Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_168 VPWR VGND sg13g2_fill_2
X_2836_ net1196 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q VPWR VGND sg13g2_dlhq_1
X_2767_ net1117 net1018 Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1718_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0374_ _0376_ _0375_ sg13g2_a21oi_1
X_1649_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q _0307_ _0309_ _0290_ _0286_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
+ _0310_ VPWR VGND sg13g2_mux4_1
X_2698_ net1134 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_32_135 VPWR VGND sg13g2_fill_1
XFILLER_9_331 VPWR VGND sg13g2_fill_1
XFILLER_9_364 VPWR VGND sg13g2_fill_2
XFILLER_20_308 VPWR VGND sg13g2_fill_1
Xoutput138 net138 E6BEG[3] VPWR VGND sg13g2_buf_1
X_2552_ net1185 net1079 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
Xoutput149 net149 EE4BEG[13] VPWR VGND sg13g2_buf_1
X_2621_ net1166 net1088 Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VPWR VGND sg13g2_dlhq_1
X_1503_ Inst_LUT4AB_switch_matrix.JS2BEG2 _0168_ _1038_ _0160_ _0161_ VPWR VGND sg13g2_a22oi_1
Xoutput127 net127 E2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput116 Inst_LUT4AB_switch_matrix.E1BEG3 E1BEG[3] VPWR VGND sg13g2_buf_1
X_2483_ net1199 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_3104_ EE4END[13] net160 VPWR VGND sg13g2_buf_1
X_3035_ net1173 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1434_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0076_ _0103_ VPWR
+ VGND sg13g2_nor2_1
X_1365_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q _0029_ _0035_ _0036_ VPWR VGND sg13g2_nor3_1
X_1296_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q net956 _1125_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_190 VPWR VGND sg13g2_fill_2
X_2819_ net1147 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_54 VPWR VGND sg13g2_fill_1
XFILLER_36_43 VPWR VGND sg13g2_decap_8
XFILLER_14_135 VPWR VGND sg13g2_fill_1
Xinput18 E2MID[4] net18 VPWR VGND sg13g2_buf_1
Xinput29 FrameStrobe[5] net29 VPWR VGND sg13g2_buf_1
XFILLER_18_430 VPWR VGND sg13g2_fill_1
X_1983_ _0632_ _0532_ _0631_ VPWR VGND sg13g2_nand2b_1
X_2604_ net1127 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_0 VPWR VGND sg13g2_fill_2
X_2535_ net1209 net1078 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
X_2466_ net1150 net1065 Inst_LB_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
X_1417_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q _1102_ _1103_ _1119_ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q
+ _0086_ VPWR VGND sg13g2_mux4_1
X_2397_ _0986_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q _0985_ VPWR VGND sg13g2_nand2_1
X_3018_ net1134 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q VPWR VGND sg13g2_dlhq_1
X_1348_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q _0014_ _0019_ _0020_ VPWR VGND sg13g2_nor3_1
X_1279_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q net37 net2 net53 net8 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ _1109_ VPWR VGND sg13g2_mux4_1
XFILLER_3_337 VPWR VGND sg13g2_fill_1
Xfanout1116 FrameData[9] net1116 VPWR VGND sg13g2_buf_1
Xfanout1127 net1128 net1127 VPWR VGND sg13g2_buf_1
Xfanout1149 FrameData[28] net1149 VPWR VGND sg13g2_buf_1
Xfanout1138 net1139 net1138 VPWR VGND sg13g2_buf_1
Xfanout1105 net1108 net1105 VPWR VGND sg13g2_buf_1
X_2320_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q _0938_ _0939_ VPWR VGND sg13g2_nor2_1
X_2251_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q VPWR _0878_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ net980 sg13g2_o21ai_1
X_1202_ VPWR _1035_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VGND sg13g2_inv_1
X_2182_ _0806_ VPWR Inst_LUT4AB_switch_matrix.E2BEG0 VGND _0816_ _0817_ sg13g2_o21ai_1
X_1966_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VPWR _0615_ VGND _0614_ _0613_ sg13g2_o21ai_1
X_1897_ net62 net70 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q _0549_ VPWR VGND sg13g2_mux2_1
X_2518_ net1191 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2449_ net1204 net1062 Inst_LA_LUT4c_frame_config_dffesr.c_reset_value VPWR VGND
+ sg13g2_dlhq_1
XFILLER_56_333 VPWR VGND sg13g2_fill_2
XFILLER_47_399 VPWR VGND sg13g2_fill_2
X_1820_ _0474_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q _0237_ VPWR VGND sg13g2_nand2_1
X_1682_ _0341_ _0339_ _0314_ _0342_ VPWR VGND sg13g2_nor3_2
X_1751_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR _0408_ VGND _0405_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ sg13g2_o21ai_1
X_2303_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q net943 _0308_ net980 _0366_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ _0924_ VPWR VGND sg13g2_mux4_1
X_2234_ _0862_ _0864_ Inst_LUT4AB_switch_matrix.WW4BEG2 VPWR VGND sg13g2_nor2_1
X_3283_ net101 net333 VPWR VGND sg13g2_buf_1
XFILLER_53_303 VPWR VGND sg13g2_fill_2
X_2096_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q net966 net954 net960 net928 Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ _0737_ VPWR VGND sg13g2_mux4_1
X_2165_ net944 net961 net994 _0801_ VPWR VGND sg13g2_mux2_1
X_1949_ _0599_ net983 net946 VPWR VGND sg13g2_nand2b_1
X_2998_ net1189 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_200 VPWR VGND sg13g2_decap_4
XFILLER_21_222 VPWR VGND sg13g2_decap_8
XFILLER_28_22 VPWR VGND sg13g2_fill_2
XFILLER_4_454 VPWR VGND sg13g2_fill_1
XFILLER_47_185 VPWR VGND sg13g2_fill_1
X_2783_ net1161 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q VPWR VGND sg13g2_dlhq_1
X_1803_ _0458_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 net926 VPWR
+ VGND sg13g2_nand2b_1
X_2852_ net1146 net1031 Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q VPWR VGND sg13g2_dlhq_1
X_2921_ net1143 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1596_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q _1051_ _0259_ _0258_ sg13g2_a21oi_1
X_1665_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VPWR _0326_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0325_ sg13g2_o21ai_1
X_1734_ VPWR _0391_ _0390_ VGND sg13g2_inv_1
X_2217_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q _1084_ _0148_ _0308_ net981 Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0850_ VPWR VGND sg13g2_mux4_1
X_3197_ Inst_LUT4AB_switch_matrix.N4BEG2 net238 VPWR VGND sg13g2_buf_1
XFILLER_26_325 VPWR VGND sg13g2_fill_1
X_2079_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q _0720_ _0722_ _0721_ sg13g2_a21oi_1
X_2148_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q _0781_ _0785_ _0784_ sg13g2_a21oi_1
XFILLER_49_417 VPWR VGND sg13g2_fill_2
XFILLER_39_21 VPWR VGND sg13g2_fill_2
XFILLER_55_31 VPWR VGND sg13g2_fill_2
XFILLER_40_350 VPWR VGND sg13g2_fill_2
XFILLER_32_328 VPWR VGND sg13g2_fill_2
Xoutput309 net309 SS4BEG[2] VPWR VGND sg13g2_buf_1
X_1450_ _1032_ VPWR _0118_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0117_ sg13g2_o21ai_1
X_3120_ net1114 net192 VPWR VGND sg13g2_buf_1
X_3051_ UserCLK net367 _0004_ _3051_/Q_N Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
X_1381_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q VPWR _0051_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q
+ _0023_ sg13g2_o21ai_1
X_2002_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q _0585_ net981 _0588_ _0587_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
+ _0650_ VPWR VGND sg13g2_mux4_1
X_2766_ net1121 net1018 Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q VPWR VGND sg13g2_dlhq_1
X_2904_ net1183 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_372 VPWR VGND sg13g2_decap_8
X_2835_ net1198 net1026 Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1717_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR _0375_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0372_ sg13g2_o21ai_1
X_1648_ VPWR _0309_ _0308_ VGND sg13g2_inv_1
X_1579_ _0241_ VPWR _0242_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q _0236_ sg13g2_o21ai_1
X_2697_ net1143 net1104 Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_26_144 VPWR VGND sg13g2_fill_2
XFILLER_26_122 VPWR VGND sg13g2_decap_4
X_3249_ Inst_LUT4AB_switch_matrix.S4BEG2 net290 VPWR VGND sg13g2_buf_1
XFILLER_41_22 VPWR VGND sg13g2_fill_1
XFILLER_25_89 VPWR VGND sg13g2_fill_1
XFILLER_49_247 VPWR VGND sg13g2_fill_2
XFILLER_1_232 VPWR VGND sg13g2_fill_2
XFILLER_32_147 VPWR VGND sg13g2_fill_1
X_2620_ net1169 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2551_ net1187 net1077 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
Xoutput139 net139 E6BEG[4] VPWR VGND sg13g2_buf_1
X_1502_ VGND VPWR _1037_ _0162_ _0168_ _0167_ sg13g2_a21oi_1
Xoutput128 net128 E2BEGb[3] VPWR VGND sg13g2_buf_1
X_1433_ _0098_ _0099_ _0101_ _0102_ VPWR VGND sg13g2_nor3_1
Xoutput117 net117 E2BEG[0] VPWR VGND sg13g2_buf_1
X_2482_ net1202 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_239 VPWR VGND sg13g2_fill_1
X_3103_ EE4END[12] net159 VPWR VGND sg13g2_buf_1
X_3034_ net1179 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q VPWR VGND sg13g2_dlhq_1
X_1295_ _1122_ _1123_ _1085_ _1124_ VPWR VGND sg13g2_nand3_1
X_1364_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q _0033_ _0035_ _0034_ sg13g2_a21oi_1
XFILLER_51_456 VPWR VGND sg13g2_fill_2
XFILLER_51_434 VPWR VGND sg13g2_fill_1
XFILLER_23_125 VPWR VGND sg13g2_fill_1
X_2749_ net1167 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q VPWR VGND sg13g2_dlhq_1
X_2818_ net1150 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_33 VPWR VGND sg13g2_fill_1
XFILLER_52_43 VPWR VGND sg13g2_fill_1
XFILLER_10_331 VPWR VGND sg13g2_fill_1
XFILLER_10_364 VPWR VGND sg13g2_fill_1
Xinput19 E2MID[5] net19 VPWR VGND sg13g2_buf_1
XFILLER_28_8 VPWR VGND sg13g2_fill_2
X_1982_ net378 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ net374 _0631_ VPWR VGND sg13g2_mux4_1
XFILLER_45_283 VPWR VGND sg13g2_fill_1
X_2534_ net1137 net1076 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
X_2603_ net1129 net1091 Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q VPWR VGND sg13g2_dlhq_1
XFILLER_47_0 VPWR VGND sg13g2_fill_1
X_1347_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q _0017_ _0019_ _0018_ sg13g2_a21oi_1
X_2465_ net1153 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_1416_ _0084_ _0079_ _0082_ _0077_ _0085_ VPWR VGND sg13g2_or4_1
X_2396_ VGND VPWR _0979_ _0985_ _0984_ _0983_ sg13g2_a21oi_2
X_3017_ net1143 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1278_ _1107_ VPWR _1108_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _1106_ sg13g2_o21ai_1
XFILLER_11_128 VPWR VGND sg13g2_fill_1
Xfanout1117 FrameData[8] net1117 VPWR VGND sg13g2_buf_1
Xfanout1139 net1140 net1139 VPWR VGND sg13g2_buf_1
Xfanout1128 FrameData[5] net1128 VPWR VGND sg13g2_buf_1
Xfanout1106 net1107 net1106 VPWR VGND sg13g2_buf_1
XFILLER_42_297 VPWR VGND sg13g2_fill_2
XFILLER_30_437 VPWR VGND sg13g2_fill_1
XFILLER_27_272 VPWR VGND sg13g2_decap_8
X_1201_ VPWR _1034_ net75 VGND sg13g2_inv_1
X_2250_ _0871_ _0877_ Inst_LUT4AB_switch_matrix.SS4BEG3 VPWR VGND sg13g2_nor2_2
XFILLER_33_6 VPWR VGND sg13g2_fill_1
X_2181_ _0817_ _0811_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VPWR VGND sg13g2_nand2b_1
X_1965_ net98 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q _0614_ VPWR VGND sg13g2_nor2_1
XFILLER_21_426 VPWR VGND sg13g2_fill_1
X_1896_ _0547_ VPWR _0548_ VGND net1006 Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ sg13g2_o21ai_1
X_2517_ net1194 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_2448_ net1114 net1062 Inst_LA_LUT4c_frame_config_dffesr.c_I0mux VPWR VGND sg13g2_dlhq_1
X_2379_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0453_ _0968_ VPWR VGND sg13g2_nor2_1
XFILLER_58_64 VPWR VGND sg13g2_fill_1
XFILLER_59_150 VPWR VGND sg13g2_fill_1
X_1750_ _0406_ VPWR _0407_ VGND net985 net934 sg13g2_o21ai_1
X_1681_ _0247_ _0340_ _0341_ VPWR VGND sg13g2_nor2_1
X_3282_ net100 net332 VPWR VGND sg13g2_buf_1
X_2302_ _0917_ _0923_ Inst_LUT4AB_switch_matrix.EE4BEG3 VPWR VGND sg13g2_nor2_2
X_2233_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q _0863_ _0864_ VPWR VGND sg13g2_nor2_1
X_2164_ _0798_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0799_ _0800_ VPWR VGND sg13g2_a21o_1
X_2095_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q net978 net973 net943 net948 Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ _0736_ VPWR VGND sg13g2_mux4_1
X_1948_ VGND VPWR _0598_ _0595_ _0597_ sg13g2_or2_1
X_1879_ VGND VPWR net386 _0490_ _0531_ _0488_ sg13g2_a21oi_1
X_2997_ net1192 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q VPWR VGND sg13g2_dlhq_1
XFILLER_56_120 VPWR VGND sg13g2_fill_2
XFILLER_29_367 VPWR VGND sg13g2_fill_1
XFILLER_12_245 VPWR VGND sg13g2_decap_4
XFILLER_50_307 VPWR VGND sg13g2_fill_2
XFILLER_43_370 VPWR VGND sg13g2_fill_2
X_2920_ net1174 net1043 Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2782_ net1164 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1733_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q net50 net21 net78 net105 Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q
+ _0390_ VPWR VGND sg13g2_mux4_1
X_1802_ _0432_ _0456_ _0457_ VPWR VGND sg13g2_nor2b_2
X_2851_ net1149 net1031 Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q VPWR VGND sg13g2_dlhq_1
X_1595_ net987 net965 _0258_ VPWR VGND sg13g2_nor2_1
X_1664_ net59 net61 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q _0325_ VPWR VGND sg13g2_mux2_1
XFILLER_53_101 VPWR VGND sg13g2_fill_2
XFILLER_38_197 VPWR VGND sg13g2_fill_2
X_2216_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q net953 net937 Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0849_
+ VPWR VGND sg13g2_mux4_1
X_3196_ Inst_LUT4AB_switch_matrix.N4BEG1 net237 VPWR VGND sg13g2_buf_1
XFILLER_26_304 VPWR VGND sg13g2_decap_4
X_3265_ Inst_LUT4AB_switch_matrix.SS4BEG2 net306 VPWR VGND sg13g2_buf_1
X_2147_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VPWR _0784_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ _0783_ sg13g2_o21ai_1
XFILLER_53_178 VPWR VGND sg13g2_fill_2
X_2078_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VPWR _0721_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ _0718_ sg13g2_o21ai_1
XFILLER_32_307 VPWR VGND sg13g2_decap_8
XFILLER_29_175 VPWR VGND sg13g2_fill_1
XFILLER_17_304 VPWR VGND sg13g2_fill_1
X_1380_ VGND VPWR _1029_ _0043_ _0050_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q
+ sg13g2_a21oi_1
X_2001_ _0648_ VPWR _0649_ VGND _0646_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q sg13g2_o21ai_1
X_3050_ UserCLK net368 _0003_ _3050_/Q_N Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
+ VPWR VGND sg13g2_dfrbp_1
X_2903_ net1186 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VPWR VGND sg13g2_dlhq_1
X_1716_ _0373_ VPWR _0374_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q net936 sg13g2_o21ai_1
X_2834_ net1202 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q VPWR VGND sg13g2_dlhq_1
X_2696_ net1174 net1108 Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2765_ net1124 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q VPWR VGND sg13g2_dlhq_1
X_1578_ _0241_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q _0237_ VPWR VGND sg13g2_nand2_1
X_1647_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q net46 net17 net74 net101 Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q
+ _0308_ VPWR VGND sg13g2_mux4_1
X_3179_ net47 net229 VPWR VGND sg13g2_buf_1
X_3248_ Inst_LUT4AB_switch_matrix.S4BEG1 net289 VPWR VGND sg13g2_buf_1
XFILLER_25_57 VPWR VGND sg13g2_fill_2
XFILLER_2_39 VPWR VGND sg13g2_fill_2
XFILLER_32_159 VPWR VGND sg13g2_decap_4
X_2550_ net1191 net1079 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_13_373 VPWR VGND sg13g2_fill_1
X_1501_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0164_ _0167_ _0166_ sg13g2_a21oi_1
Xoutput129 net129 E2BEGb[4] VPWR VGND sg13g2_buf_1
X_1363_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VPWR _0034_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ _0031_ sg13g2_o21ai_1
X_1432_ _0100_ VPWR _0101_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0076_ sg13g2_o21ai_1
Xoutput118 net118 E2BEG[1] VPWR VGND sg13g2_buf_1
X_2481_ net1204 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_3102_ EE4END[11] net158 VPWR VGND sg13g2_buf_1
XFILLER_55_207 VPWR VGND sg13g2_fill_1
X_3033_ net1181 net1113 Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q VPWR VGND sg13g2_dlhq_1
X_1294_ _1123_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 net982 VPWR
+ VGND sg13g2_nand2_1
X_3050__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_31_192 VPWR VGND sg13g2_fill_1
X_2748_ net1170 net1015 Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2679_ net1186 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2817_ net1153 net1022 Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_54_273 VPWR VGND sg13g2_fill_2
XFILLER_54_251 VPWR VGND sg13g2_fill_1
XFILLER_39_281 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_fill_2
XFILLER_37_218 VPWR VGND sg13g2_fill_2
X_1981_ VGND VPWR _0629_ _0630_ _0593_ _0532_ sg13g2_a21oi_2
XFILLER_9_152 VPWR VGND sg13g2_fill_1
X_2533_ net1140 net1076 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
X_2602_ net1132 net1091 Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_5_380 VPWR VGND sg13g2_fill_2
X_1415_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0083_ _0084_ VPWR
+ VGND sg13g2_nor2_1
X_1346_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VPWR _0018_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ _0015_ sg13g2_o21ai_1
X_2464_ net1157 net1064 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_2395_ _0981_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q _0984_ VPWR VGND sg13g2_nor2b_1
X_3016_ net1174 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q VPWR VGND sg13g2_dlhq_1
X_1277_ _1107_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _1105_ VPWR VGND sg13g2_nand2b_1
XFILLER_51_276 VPWR VGND sg13g2_fill_2
Xfanout1129 FrameData[4] net1129 VPWR VGND sg13g2_buf_1
Xfanout1118 FrameData[8] net1118 VPWR VGND sg13g2_buf_1
Xfanout1107 net1108 net1107 VPWR VGND sg13g2_buf_1
XFILLER_42_276 VPWR VGND sg13g2_decap_8
X_2180_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0814_ _0816_ _0815_ sg13g2_a21oi_1
X_1200_ VPWR _1033_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VGND sg13g2_inv_1
X_1895_ _0547_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q net1003 VPWR VGND sg13g2_nand2b_1
X_1964_ Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ _0613_ VPWR VGND sg13g2_nor2b_1
X_2516_ net1197 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 VPWR
+ VGND sg13g2_dlhq_1
X_2447_ net1117 net1062 Inst_LA_LUT4c_frame_config_dffesr.c_out_mux VPWR VGND sg13g2_dlhq_1
XFILLER_56_335 VPWR VGND sg13g2_fill_1
X_1329_ _1156_ _1153_ _1148_ Inst_LUT4AB_switch_matrix.JS2BEG3 VPWR VGND sg13g2_a21o_2
X_2378_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0048_ _0967_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a21oi_1
XFILLER_59_140 VPWR VGND sg13g2_fill_2
XFILLER_47_302 VPWR VGND sg13g2_fill_2
Xoutput290 net290 S4BEG[14] VPWR VGND sg13g2_buf_1
X_1680_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0310_ _0340_ VPWR VGND sg13g2_mux4_1
X_2301_ VGND VPWR _0922_ _0923_ _0919_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q sg13g2_a21oi_2
XFILLER_53_305 VPWR VGND sg13g2_fill_1
X_2232_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q net1010 net87 net59 net969 Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ _0863_ VPWR VGND sg13g2_mux4_1
X_3281_ net99 net331 VPWR VGND sg13g2_buf_1
X_2163_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VPWR _0799_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ _0796_ sg13g2_o21ai_1
X_2094_ Inst_LUT4AB_switch_matrix.JN2BEG7 _0734_ _0735_ _0727_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_a22oi_1
X_1947_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR _0597_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ _0596_ sg13g2_o21ai_1
X_1878_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q _0520_ _0525_ _0529_ _0527_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q
+ _0530_ VPWR VGND sg13g2_mux4_1
X_2996_ net1195 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_56_198 VPWR VGND sg13g2_fill_2
XFILLER_20_290 VPWR VGND sg13g2_fill_1
X_2850_ net1151 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2781_ net1165 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q VPWR VGND sg13g2_dlhq_1
X_1732_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q net20 net104 net77 Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q _0389_ VPWR VGND sg13g2_mux4_1
X_1663_ _0323_ VPWR _0324_ VGND net69 Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q sg13g2_o21ai_1
X_1801_ _0455_ VPWR _0456_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q _0452_
+ sg13g2_o21ai_1
X_1594_ _1042_ _0256_ _0257_ VPWR VGND sg13g2_and2_1
X_3264_ Inst_LUT4AB_switch_matrix.SS4BEG1 net305 VPWR VGND sg13g2_buf_1
X_2215_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q net942 net947 net966 net959 Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0848_ VPWR VGND sg13g2_mux4_1
X_2077_ _0719_ VPWR _0720_ VGND net63 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q sg13g2_o21ai_1
X_3195_ Inst_LUT4AB_switch_matrix.N4BEG0 net236 VPWR VGND sg13g2_buf_1
X_2146_ VGND VPWR net991 net951 _0783_ _0782_ sg13g2_a21oi_1
X_2979_ net1149 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_39_23 VPWR VGND sg13g2_fill_1
XFILLER_29_154 VPWR VGND sg13g2_fill_2
XFILLER_55_33 VPWR VGND sg13g2_fill_1
XFILLER_32_319 VPWR VGND sg13g2_fill_1
XFILLER_25_371 VPWR VGND sg13g2_decap_8
X_2000_ _0537_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q _0647_ _0648_ VPWR VGND sg13g2_a21o_1
XFILLER_50_149 VPWR VGND sg13g2_fill_2
XFILLER_43_190 VPWR VGND sg13g2_fill_1
X_2902_ net1189 net1040 Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q VPWR VGND sg13g2_dlhq_1
X_2833_ net1204 net1029 Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1715_ _0373_ net999 net930 VPWR VGND sg13g2_nand2b_1
X_1646_ _0306_ VPWR _0307_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q _0303_ sg13g2_o21ai_1
X_2695_ net1208 net1108 Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_60 VPWR VGND sg13g2_fill_2
XFILLER_6_82 VPWR VGND sg13g2_fill_1
X_2764_ net1126 net1016 Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q VPWR VGND sg13g2_dlhq_1
X_1577_ _0240_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux _0209_ VPWR VGND sg13g2_nand2_1
XFILLER_39_452 VPWR VGND sg13g2_fill_2
X_3247_ Inst_LUT4AB_switch_matrix.S4BEG0 net288 VPWR VGND sg13g2_buf_1
XFILLER_26_146 VPWR VGND sg13g2_fill_1
XFILLER_25_69 VPWR VGND sg13g2_fill_1
X_3178_ net46 net228 VPWR VGND sg13g2_buf_1
X_2129_ _0766_ VPWR _0767_ VGND net986 net932 sg13g2_o21ai_1
Xrebuffer10 Inst_LUT4AB_switch_matrix.E2BEG1 net383 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_1_234 VPWR VGND sg13g2_fill_1
XFILLER_49_249 VPWR VGND sg13g2_fill_1
XFILLER_40_160 VPWR VGND sg13g2_decap_8
X_1500_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VPWR _0166_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ _0165_ sg13g2_o21ai_1
Xoutput119 net119 E2BEG[2] VPWR VGND sg13g2_buf_1
X_2480_ net1114 net1066 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_3101_ EE4END[10] net157 VPWR VGND sg13g2_buf_1
X_1293_ _1122_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 net982 VPWR
+ VGND sg13g2_nand2b_1
X_1362_ _0032_ VPWR _0033_ VGND net94 Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q sg13g2_o21ai_1
X_1431_ _0100_ _0078_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 VPWR
+ VGND sg13g2_nand2b_1
X_3032_ net1183 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_458 VPWR VGND sg13g2_fill_1
X_2816_ net1156 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2747_ net1172 net1015 Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1629_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q net979 net973 net943 net948 Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0291_ VPWR VGND sg13g2_mux4_1
X_2678_ net1191 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_11_38 VPWR VGND sg13g2_fill_1
XFILLER_10_388 VPWR VGND sg13g2_fill_2
X_1980_ _0627_ VPWR _0629_ VGND _0628_ _0532_ sg13g2_o21ai_1
Xrebuffer1 _0565_ net374 VPWR VGND sg13g2_dlygate4sd1_1
X_2532_ net1145 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
X_2601_ net1141 net1090 Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q VPWR VGND sg13g2_dlhq_1
X_2463_ net1160 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_3015_ net1207 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q VPWR VGND sg13g2_dlhq_1
X_1345_ _0016_ VPWR _0017_ VGND net92 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q sg13g2_o21ai_1
X_1276_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q net975 D net940 net963 Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ _1106_ VPWR VGND sg13g2_mux4_1
X_1414_ VGND VPWR _0083_ _0075_ _0074_ sg13g2_or2_1
X_2394_ _0982_ VPWR _0983_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q Inst_LUT4AB_switch_matrix.JN2BEG1
+ sg13g2_o21ai_1
Xfanout1119 FrameData[8] net1119 VPWR VGND sg13g2_buf_1
Xfanout1108 FrameStrobe[10] net1108 VPWR VGND sg13g2_buf_1
XFILLER_47_56 VPWR VGND sg13g2_fill_2
XFILLER_42_244 VPWR VGND sg13g2_decap_8
XFILLER_6_189 VPWR VGND sg13g2_fill_1
XFILLER_18_263 VPWR VGND sg13g2_decap_8
X_1894_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q net34 net42 net5 net13 Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ _0546_ VPWR VGND sg13g2_mux4_1
X_1963_ Inst_LUT4AB_switch_matrix.JW2BEG6 _0611_ _0612_ _0604_ _0598_ VPWR VGND sg13g2_a22oi_1
XFILLER_52_0 VPWR VGND sg13g2_fill_2
X_2515_ net1199 net1072 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 VPWR
+ VGND sg13g2_dlhq_1
X_2446_ net1121 net1060 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_1328_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q _1155_ _1156_ VPWR VGND sg13g2_nor2_1
X_1259_ _1089_ VPWR _1090_ VGND net1000 net934 sg13g2_o21ai_1
X_2377_ _0966_ _0617_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VPWR VGND sg13g2_nand2b_1
XFILLER_12_439 VPWR VGND sg13g2_fill_2
XFILLER_24_277 VPWR VGND sg13g2_decap_8
XFILLER_59_196 VPWR VGND sg13g2_fill_2
Xoutput280 net280 S2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput291 net291 S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_30_258 VPWR VGND sg13g2_fill_1
XFILLER_7_454 VPWR VGND sg13g2_fill_1
X_2300_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VPWR _0922_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ _0921_ sg13g2_o21ai_1
X_2231_ _0858_ _0861_ _0862_ VPWR VGND sg13g2_nor2_1
X_3280_ net98 net330 VPWR VGND sg13g2_buf_1
X_2093_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q _0732_ _0735_ VPWR VGND sg13g2_nor2_1
X_2162_ _0797_ VPWR _0798_ VGND net995 net932 sg13g2_o21ai_1
X_2995_ net1198 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1946_ net965 net958 net983 _0596_ VPWR VGND sg13g2_mux2_1
X_1877_ VPWR _0529_ _0528_ VGND sg13g2_inv_1
X_2429_ _1007_ VPWR _1011_ VGND Inst_LG_LUT4c_frame_config_dffesr.c_reset_value _1009_
+ sg13g2_o21ai_1
XFILLER_28_47 VPWR VGND sg13g2_fill_2
XFILLER_29_358 VPWR VGND sg13g2_decap_8
XFILLER_43_372 VPWR VGND sg13g2_fill_1
X_1800_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q _0453_ _0455_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q
+ sg13g2_a21oi_1
X_1731_ Inst_LUT4AB_switch_matrix.JN2BEG4 _0382_ _0388_ _0370_ _0377_ VPWR VGND sg13g2_a22oi_1
X_2780_ net1170 net1019 Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1662_ _0323_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q net1004 VPWR VGND sg13g2_nand2b_1
X_3194_ N4END[15] net235 VPWR VGND sg13g2_buf_1
X_1593_ net987 net977 net971 net941 net946 Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0256_ VPWR VGND sg13g2_mux4_1
X_2214_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q net1214 net1003 net977 net972 Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0847_ VPWR VGND sg13g2_mux4_1
XFILLER_38_199 VPWR VGND sg13g2_fill_1
XFILLER_34_350 VPWR VGND sg13g2_fill_2
X_2076_ _0719_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q net87 VPWR VGND sg13g2_nand2b_1
XFILLER_15_0 VPWR VGND sg13g2_fill_1
X_2145_ net991 net956 _0782_ VPWR VGND sg13g2_nor2b_1
X_1929_ _0579_ VPWR _0580_ VGND net70 net992 sg13g2_o21ai_1
X_2978_ net1152 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_35_114 VPWR VGND sg13g2_decap_8
X_2763_ net1130 net1018 Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q VPWR VGND sg13g2_dlhq_1
X_2901_ net1192 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2832_ net1114 net1027 Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1576_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q net42 net70 net24 net97 Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q
+ _0239_ VPWR VGND sg13g2_mux4_1
X_1714_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q _1051_ _0372_ _0371_ sg13g2_a21oi_1
X_1645_ _0304_ _0305_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q _0306_ VPWR VGND sg13g2_nand3_1
X_2694_ net1135 net1100 Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q VPWR VGND sg13g2_dlhq_1
X_3246_ S4END[15] net287 VPWR VGND sg13g2_buf_1
XFILLER_54_412 VPWR VGND sg13g2_fill_1
X_3177_ net45 net227 VPWR VGND sg13g2_buf_1
Xrebuffer11 Inst_LUT4AB_switch_matrix.JW2BEG2 net384 VPWR VGND sg13g2_dlygate4sd1_1
X_2059_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VPWR _0703_ VGND _0699_ _0701_ sg13g2_o21ai_1
X_2128_ _0766_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q net931 VPWR VGND sg13g2_nand2_1
XFILLER_32_106 VPWR VGND sg13g2_decap_4
XFILLER_15_70 VPWR VGND sg13g2_fill_1
X_1430_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0083_ _0099_ VPWR
+ VGND sg13g2_nor2_1
X_3100_ EE4END[9] net156 VPWR VGND sg13g2_buf_1
X_1361_ _0032_ _1023_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q VPWR VGND sg13g2_nand2_1
X_1292_ _1120_ net1 Inst_LA_LUT4c_frame_config_dffesr.c_I0mux _1121_ VPWR VGND sg13g2_mux2_2
X_3031_ net1186 net1109 Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q VPWR VGND sg13g2_dlhq_1
X_2746_ net1178 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_161 VPWR VGND sg13g2_decap_8
X_2815_ net1159 net1021 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q VPWR VGND sg13g2_dlhq_1
X_1628_ VGND VPWR _1041_ _0289_ _0290_ _0288_ sg13g2_a21oi_1
X_1559_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0222_ _0223_ VPWR VGND sg13g2_nor2b_1
X_2677_ net1194 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VPWR VGND sg13g2_dlhq_1
X_3229_ net73 net279 VPWR VGND sg13g2_buf_1
XFILLER_54_275 VPWR VGND sg13g2_fill_1
XFILLER_7_2 VPWR VGND sg13g2_fill_1
XFILLER_18_412 VPWR VGND sg13g2_fill_2
XFILLER_18_445 VPWR VGND sg13g2_fill_2
XFILLER_18_456 VPWR VGND sg13g2_fill_2
X_2600_ net1174 net1087 Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q VPWR VGND sg13g2_dlhq_1
Xrebuffer2 _0248_ net375 VPWR VGND sg13g2_dlygate4sd1_1
X_2531_ net1148 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_382 VPWR VGND sg13g2_fill_1
XFILLER_5_360 VPWR VGND sg13g2_fill_2
X_1413_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0081_ _0082_ VPWR
+ VGND sg13g2_nor2_1
X_2462_ net1163 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2393_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _1064_ _0982_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ sg13g2_a21oi_1
XFILLER_3_51 VPWR VGND sg13g2_fill_1
X_1344_ _0016_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q net106 VPWR VGND sg13g2_nand2b_1
X_1275_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q net957 net951 net935 net931 Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ _1105_ VPWR VGND sg13g2_mux4_1
X_3014_ net1135 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q VPWR VGND sg13g2_dlhq_1
X_2729_ net1142 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q VPWR VGND sg13g2_dlhq_1
Xfanout1109 net1112 net1109 VPWR VGND sg13g2_buf_1
XFILLER_27_286 VPWR VGND sg13g2_fill_1
XFILLER_30_407 VPWR VGND sg13g2_decap_8
X_1962_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q _0609_ _0612_ VPWR VGND sg13g2_nor2_1
XFILLER_33_212 VPWR VGND sg13g2_fill_2
X_1893_ VGND VPWR _1044_ _0539_ _0545_ _0544_ sg13g2_a21oi_1
X_2376_ _0651_ VPWR net112 VGND _0652_ _0639_ sg13g2_o21ai_1
X_2514_ net1203 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_45_0 VPWR VGND sg13g2_fill_2
X_2445_ net1124 net1060 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_1258_ _1089_ net1000 net929 VPWR VGND sg13g2_nand2b_1
X_1327_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _1154_ _1155_ VPWR VGND sg13g2_nor2_1
X_1189_ VPWR _1022_ net79 VGND sg13g2_inv_1
XFILLER_17_38 VPWR VGND sg13g2_fill_1
Xoutput270 net270 S2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_47_304 VPWR VGND sg13g2_fill_1
Xoutput281 net281 S2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput292 net292 S4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_15_223 VPWR VGND sg13g2_fill_1
XFILLER_7_400 VPWR VGND sg13g2_fill_1
X_2230_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q VPWR _0861_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
+ _0860_ sg13g2_o21ai_1
XFILLER_38_337 VPWR VGND sg13g2_fill_2
X_2092_ _0734_ _0733_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VPWR VGND sg13g2_nand2b_1
X_2161_ _0797_ net995 net929 VPWR VGND sg13g2_nand2_1
X_1945_ VGND VPWR _0594_ _0595_ Inst_LUT4AB_switch_matrix.M_EF net983 sg13g2_a21oi_2
X_2994_ net1201 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_204 VPWR VGND sg13g2_fill_1
X_1876_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q net42 net13 net70 net108 Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q
+ _0528_ VPWR VGND sg13g2_mux4_1
X_2428_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q _0630_ net925 _0632_ _1010_
+ _0635_ sg13g2_a221oi_1
X_2359_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q net1210 net80 net65 net975 Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ Inst_LUT4AB_switch_matrix.S4BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_44_47 VPWR VGND sg13g2_fill_2
XFILLER_12_215 VPWR VGND sg13g2_fill_2
XFILLER_4_403 VPWR VGND sg13g2_fill_1
XFILLER_35_307 VPWR VGND sg13g2_fill_1
XFILLER_43_395 VPWR VGND sg13g2_fill_2
XFILLER_43_351 VPWR VGND sg13g2_fill_2
X_1730_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q _0387_ _0388_ VPWR VGND sg13g2_nor2_1
X_1592_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q _0248_ _0255_ _0254_ sg13g2_a21oi_1
X_1661_ _0322_ _0321_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VPWR VGND sg13g2_nand2b_1
X_3262_ SS4END[15] net303 VPWR VGND sg13g2_buf_1
X_3193_ N4END[14] net234 VPWR VGND sg13g2_buf_1
XFILLER_38_112 VPWR VGND sg13g2_fill_2
X_2213_ Inst_LUT4AB_switch_matrix.W6BEG1 _0846_ _0841_ VPWR VGND sg13g2_nand2b_1
X_2144_ _0780_ VPWR _0781_ VGND net991 net932 sg13g2_o21ai_1
XFILLER_53_137 VPWR VGND sg13g2_fill_2
X_2075_ net59 net61 Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q _0718_ VPWR VGND sg13g2_mux2_1
X_1928_ _0579_ net992 net1003 VPWR VGND sg13g2_nand2b_1
X_1859_ net62 net70 net996 _0512_ VPWR VGND sg13g2_mux2_1
X_2977_ net1155 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_17_329 VPWR VGND sg13g2_decap_4
X_2900_ net1197 net1039 Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q VPWR VGND sg13g2_dlhq_1
X_1713_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q net958 _0371_ VPWR VGND sg13g2_nor2_1
X_2762_ net1132 net1018 Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q VPWR VGND sg13g2_dlhq_1
XFILLER_43_181 VPWR VGND sg13g2_fill_2
XFILLER_31_365 VPWR VGND sg13g2_fill_2
X_2831_ net1117 net1027 Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q VPWR VGND sg13g2_dlhq_1
X_1644_ _0305_ net73 Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VPWR VGND sg13g2_nand2b_1
X_1575_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q net54 net93 net9 Inst_LUT4AB_switch_matrix.JN2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q _0238_ VPWR VGND sg13g2_mux4_1
X_3314_ Inst_LUT4AB_switch_matrix.WW4BEG2 net355 VPWR VGND sg13g2_buf_1
X_2693_ net1138 net1099 Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_62 VPWR VGND sg13g2_fill_1
X_3245_ S4END[14] net286 VPWR VGND sg13g2_buf_1
Xrebuffer12 _0520_ net385 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_39_454 VPWR VGND sg13g2_fill_1
XFILLER_26_137 VPWR VGND sg13g2_decap_8
XFILLER_26_126 VPWR VGND sg13g2_fill_1
X_3176_ net44 net226 VPWR VGND sg13g2_buf_1
X_2127_ VGND VPWR net986 net950 _0765_ _0764_ sg13g2_a21oi_1
X_2058_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q net974 net969 net939 net945 Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0702_ VPWR VGND sg13g2_mux4_1
XFILLER_22_365 VPWR VGND sg13g2_fill_1
XFILLER_57_262 VPWR VGND sg13g2_fill_2
XFILLER_45_402 VPWR VGND sg13g2_fill_2
XFILLER_25_181 VPWR VGND sg13g2_fill_1
X_1360_ VGND VPWR _1022_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0031_ _0030_ sg13g2_a21oi_1
X_1291_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q _1102_ _1103_ _1119_ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q
+ _1120_ VPWR VGND sg13g2_mux4_1
X_3030_ net1189 net1111 Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q VPWR VGND sg13g2_dlhq_1
XFILLER_36_457 VPWR VGND sg13g2_fill_2
X_2814_ net1164 net1023 Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_31_173 VPWR VGND sg13g2_fill_2
X_2745_ net1181 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q VPWR VGND sg13g2_dlhq_1
X_2676_ net1195 net27 Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q VPWR VGND sg13g2_dlhq_1
X_1627_ net38 net9 Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q _0289_ VPWR VGND sg13g2_mux2_1
X_1558_ net998 net33 net41 net4 net12 Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0222_
+ VPWR VGND sg13g2_mux4_1
X_1489_ net990 net959 _0155_ VPWR VGND sg13g2_nor2_1
X_3159_ net1075 net200 VPWR VGND sg13g2_buf_1
X_3228_ net72 net278 VPWR VGND sg13g2_buf_1
XFILLER_33_438 VPWR VGND sg13g2_fill_1
X_2530_ net1151 net1075 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
Xrebuffer3 _0248_ net376 VPWR VGND sg13g2_dlygate4sd1_1
X_1343_ net65 net81 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q _0015_ VPWR VGND sg13g2_mux2_1
X_1412_ _0081_ _0074_ _0075_ VPWR VGND sg13g2_nand2_1
X_2461_ net1166 net1064 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2392_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0021_ _0981_ _0980_ sg13g2_a21oi_1
XFILLER_36_221 VPWR VGND sg13g2_decap_8
X_3013_ net1138 net1054 Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q VPWR VGND sg13g2_dlhq_1
X_1274_ VPWR _1104_ _1103_ VGND sg13g2_inv_1
X_2728_ net1176 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VPWR VGND sg13g2_dlhq_1
X_2659_ net1147 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_59_379 VPWR VGND sg13g2_fill_2
XFILLER_59_357 VPWR VGND sg13g2_fill_1
XFILLER_47_58 VPWR VGND sg13g2_fill_1
XFILLER_42_202 VPWR VGND sg13g2_decap_4
XFILLER_27_265 VPWR VGND sg13g2_decap_8
XFILLER_6_158 VPWR VGND sg13g2_fill_2
XFILLER_10_143 VPWR VGND sg13g2_fill_1
XFILLER_5_0 VPWR VGND sg13g2_fill_1
XFILLER_37_80 VPWR VGND sg13g2_decap_8
X_1961_ _0611_ _0610_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR VGND sg13g2_nand2b_1
X_1892_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VPWR _0544_ VGND _0542_ _0543_ sg13g2_o21ai_1
XFILLER_33_257 VPWR VGND sg13g2_fill_2
XFILLER_52_2 VPWR VGND sg13g2_fill_1
X_2513_ net1205 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_38_0 VPWR VGND sg13g2_fill_2
X_2444_ net1128 net1060 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_1326_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q net39 net1215 net10 net1212 Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ _1154_ VPWR VGND sg13g2_mux4_1
X_2375_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q net939 Inst_LUT4AB_switch_matrix.JW2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q Inst_LUT4AB_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1188_ VPWR _1021_ net47 VGND sg13g2_inv_1
X_1257_ VGND VPWR _1087_ _1088_ _1051_ net1000 sg13g2_a21oi_2
XFILLER_59_110 VPWR VGND sg13g2_fill_1
Xoutput260 net260 NN4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput271 net271 S2BEG[2] VPWR VGND sg13g2_buf_1
Xoutput293 net293 S4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput282 net282 S2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_59_198 VPWR VGND sg13g2_fill_1
XFILLER_47_327 VPWR VGND sg13g2_fill_1
XFILLER_30_249 VPWR VGND sg13g2_decap_4
X_2160_ VGND VPWR net994 net950 _0796_ _0795_ sg13g2_a21oi_1
X_2091_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q net1010 net35 net1217 net22 Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ _0733_ VPWR VGND sg13g2_mux4_1
X_1944_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q VPWR _0594_ VGND net983 net933 sg13g2_o21ai_1
X_1875_ VPWR _0527_ _0526_ VGND sg13g2_inv_1
X_2993_ net1206 net1056 Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q VPWR VGND sg13g2_dlhq_1
X_2427_ _1009_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q net925 VPWR VGND sg13g2_nand2_1
X_2289_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q net1214 net1003 net978 net973 Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0912_ VPWR VGND sg13g2_mux4_1
X_1309_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _1137_ _1138_ _1027_ sg13g2_a21oi_1
X_2358_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q net1212 net81 net66 net970 Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ Inst_LUT4AB_switch_matrix.S4BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_12_238 VPWR VGND sg13g2_decap_8
XFILLER_12_249 VPWR VGND sg13g2_fill_1
X_1591_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q VPWR _0254_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q
+ _0253_ sg13g2_o21ai_1
X_1660_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q net1008 net41 net1215 net12 Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0321_ VPWR VGND sg13g2_mux4_1
XFILLER_7_242 VPWR VGND sg13g2_fill_1
X_3192_ N4END[13] net248 VPWR VGND sg13g2_buf_1
X_3261_ SS4END[14] net302 VPWR VGND sg13g2_buf_1
XFILLER_38_179 VPWR VGND sg13g2_fill_1
X_2212_ _0845_ VPWR _0846_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0842_ sg13g2_o21ai_1
X_2143_ _0780_ net991 net928 VPWR VGND sg13g2_nand2_1
X_2074_ _0717_ _0716_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VPWR VGND sg13g2_nand2b_1
X_1927_ _0577_ VPWR _0578_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0576_ sg13g2_o21ai_1
X_1858_ _0510_ VPWR _0511_ VGND net996 net1006 sg13g2_o21ai_1
X_2976_ net1156 net1049 Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VPWR VGND sg13g2_dlhq_1
X_1789_ VGND VPWR _0445_ _0444_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q sg13g2_or2_1
XFILLER_40_300 VPWR VGND sg13g2_fill_2
XFILLER_25_385 VPWR VGND sg13g2_fill_2
XFILLER_45_80 VPWR VGND sg13g2_fill_1
X_2830_ net1121 net1030 Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q VPWR VGND sg13g2_dlhq_1
X_1712_ _0370_ _0369_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR VGND sg13g2_nand2b_1
X_2761_ net1141 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q VPWR VGND sg13g2_dlhq_1
X_1643_ _0304_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q Inst_LUT4AB_switch_matrix.E2BEG5
+ VPWR VGND sg13g2_nand2_1
X_2692_ net1146 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q VPWR VGND sg13g2_dlhq_1
X_3244_ S4END[13] net300 VPWR VGND sg13g2_buf_1
X_3313_ Inst_LUT4AB_switch_matrix.WW4BEG1 net354 VPWR VGND sg13g2_buf_1
X_1574_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q net50 net21 net78 net105 Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q
+ _0237_ VPWR VGND sg13g2_mux4_1
XFILLER_54_458 VPWR VGND sg13g2_fill_1
Xrebuffer13 _0479_ net386 VPWR VGND sg13g2_buf_2
Xfanout1090 net1091 net1090 VPWR VGND sg13g2_buf_1
X_3175_ net43 net225 VPWR VGND sg13g2_buf_1
X_2126_ net986 net955 _0764_ VPWR VGND sg13g2_nor2b_1
X_2057_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VPWR _0701_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0700_ sg13g2_o21ai_1
XFILLER_25_39 VPWR VGND sg13g2_fill_1
X_2959_ net1119 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VPWR VGND sg13g2_dlhq_1
XFILLER_45_458 VPWR VGND sg13g2_fill_1
XFILLER_17_138 VPWR VGND sg13g2_fill_2
X_1290_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q net41 net86 net12 net96 Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q
+ _1119_ VPWR VGND sg13g2_mux4_1
X_2813_ net1167 net1024 Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q VPWR VGND sg13g2_dlhq_1
X_1626_ VGND VPWR _1030_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q _0288_ _0287_ sg13g2_a21oi_1
X_2744_ net1184 net1011 Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q VPWR VGND sg13g2_dlhq_1
X_2675_ net1198 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q VPWR VGND sg13g2_dlhq_1
X_1557_ _0221_ _0220_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q VPWR VGND sg13g2_nand2_2
X_1488_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0151_ _0154_ _0153_ sg13g2_a21oi_1
X_3227_ net71 net277 VPWR VGND sg13g2_buf_1
X_3158_ net1081 net199 VPWR VGND sg13g2_buf_1
XFILLER_54_211 VPWR VGND sg13g2_fill_1
XFILLER_54_200 VPWR VGND sg13g2_fill_1
XFILLER_39_274 VPWR VGND sg13g2_decap_8
X_2109_ _0749_ Inst_LUT4AB_switch_matrix.JW2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_nand2_2
X_3089_ E6END[8] net141 VPWR VGND sg13g2_buf_1
XFILLER_27_425 VPWR VGND sg13g2_fill_1
XFILLER_22_174 VPWR VGND sg13g2_fill_1
XFILLER_18_458 VPWR VGND sg13g2_fill_1
XFILLER_41_450 VPWR VGND sg13g2_fill_1
Xrebuffer4 Inst_LUT4AB_switch_matrix.JW2BEG5 net377 VPWR VGND sg13g2_dlygate4sd1_1
XFILLER_5_362 VPWR VGND sg13g2_fill_1
X_2460_ net1169 net1063 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_1273_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q net50 net21 net78 net105 Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q
+ _1103_ VPWR VGND sg13g2_mux4_1
X_1342_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0013_ _0014_ VPWR VGND sg13g2_nor2b_1
X_1411_ _0074_ _0075_ _0080_ VPWR VGND sg13g2_and2_1
X_2391_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q VPWR _0980_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ Inst_LUT4AB_switch_matrix.JS2BEG1 sg13g2_o21ai_1
X_3012_ net1144 net1055 Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_51_258 VPWR VGND sg13g2_fill_2
XFILLER_22_29 VPWR VGND sg13g2_fill_1
X_1609_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VPWR _0272_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0271_ sg13g2_o21ai_1
X_2727_ net1208 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q VPWR VGND sg13g2_dlhq_1
X_2658_ net1150 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2589_ net1165 net1082 Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_27_200 VPWR VGND sg13g2_decap_8
XFILLER_2_398 VPWR VGND sg13g2_fill_2
XFILLER_33_236 VPWR VGND sg13g2_fill_2
XFILLER_33_214 VPWR VGND sg13g2_fill_1
X_1960_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q net1007 net42 net1214 net13 Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ _0610_ VPWR VGND sg13g2_mux4_1
X_1891_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VPWR _0543_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ _0540_ sg13g2_o21ai_1
X_2512_ net1115 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 VPWR
+ VGND sg13g2_dlhq_1
X_2443_ net1131 net1060 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2374_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q net947 _0237_ Inst_LUT4AB_switch_matrix.JW2BEG0
+ net375 Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q Inst_LUT4AB_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1325_ _1152_ VPWR _1153_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1150_ sg13g2_o21ai_1
X_1256_ net1000 net955 _1087_ VPWR VGND sg13g2_nor2_1
X_1187_ VPWR _1020_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VGND sg13g2_inv_1
Xoutput261 net261 NN4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput250 net250 NN4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_58_36 VPWR VGND sg13g2_fill_2
Xoutput272 net272 S2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput283 net283 S2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput294 net294 S4BEG[3] VPWR VGND sg13g2_buf_1
X_2090_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q _0729_ _0732_ _0731_ sg13g2_a21oi_1
X_2992_ net1116 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1874_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q net54 net22 net82 Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q _0526_ VPWR VGND sg13g2_mux4_1
X_1943_ VPWR _0593_ _0592_ VGND sg13g2_inv_1
X_2426_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q net390 _1008_ VPWR VGND net927 sg13g2_nand3b_1
XFILLER_50_0 VPWR VGND sg13g2_fill_2
X_2288_ _0907_ _0911_ Inst_LUT4AB_switch_matrix.E6BEG1 VPWR VGND sg13g2_nor2_2
X_1239_ net939 net961 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1071_ VPWR VGND sg13g2_mux2_1
X_1308_ net92 net106 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _1137_ VPWR VGND sg13g2_mux2_1
X_2357_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q net63 net107 net82 net940 Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ Inst_LUT4AB_switch_matrix.S4BEG2 VPWR VGND sg13g2_mux4_1
XFILLER_44_49 VPWR VGND sg13g2_fill_1
XFILLER_18_61 VPWR VGND sg13g2_fill_2
XFILLER_43_397 VPWR VGND sg13g2_fill_1
X_3260_ SS4END[13] net316 VPWR VGND sg13g2_buf_1
X_1590_ _0252_ VPWR _0253_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q _0249_ sg13g2_o21ai_1
XFILLER_7_287 VPWR VGND sg13g2_fill_2
X_3191_ N4END[12] net247 VPWR VGND sg13g2_buf_1
X_2211_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0844_ _0845_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ sg13g2_a21oi_1
X_2142_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q net969 net944 net938 net964 net991
+ _0779_ VPWR VGND sg13g2_mux4_1
X_2073_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q net1010 net55 net1217 net6 Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ _0716_ VPWR VGND sg13g2_mux4_1
XFILLER_34_386 VPWR VGND sg13g2_fill_2
X_2975_ net1159 net1049 Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_14_19 VPWR VGND sg13g2_fill_1
X_1926_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0575_ _0577_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q
+ sg13g2_a21oi_1
X_1857_ _0510_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q net89 VPWR VGND sg13g2_nand2b_1
X_1788_ net60 net62 net984 _0444_ VPWR VGND sg13g2_mux2_1
X_2409_ _0995_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q net927 VPWR VGND sg13g2_nand2b_1
XFILLER_44_139 VPWR VGND sg13g2_decap_4
XFILLER_25_364 VPWR VGND sg13g2_decap_8
XFILLER_35_139 VPWR VGND sg13g2_fill_1
XFILLER_31_367 VPWR VGND sg13g2_fill_1
XFILLER_31_323 VPWR VGND sg13g2_decap_4
X_2760_ net1176 net1017 Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q VPWR VGND sg13g2_dlhq_1
X_1711_ net999 net976 net971 net941 net946 Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0369_ VPWR VGND sg13g2_mux4_1
X_1642_ net45 net16 Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q _0303_ VPWR VGND sg13g2_mux2_1
X_2691_ net1149 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_20 VPWR VGND sg13g2_fill_1
X_3243_ S4END[12] net299 VPWR VGND sg13g2_buf_1
X_1573_ _0232_ _0235_ _0236_ VPWR VGND sg13g2_nor2_1
X_3312_ Inst_LUT4AB_switch_matrix.WW4BEG0 net353 VPWR VGND sg13g2_buf_1
XFILLER_39_401 VPWR VGND sg13g2_fill_1
Xfanout1080 net1081 net1080 VPWR VGND sg13g2_buf_1
Xrebuffer14 _0638_ net387 VPWR VGND sg13g2_dlygate4sd1_1
X_3174_ Inst_LUT4AB_switch_matrix.JN2BEG7 net224 VPWR VGND sg13g2_buf_1
X_2125_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q net968 net944 net938 net961 net986
+ _0763_ VPWR VGND sg13g2_mux4_1
X_2056_ net963 net956 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q _0700_ VPWR VGND sg13g2_mux2_1
Xfanout1091 net1092 net1091 VPWR VGND sg13g2_buf_1
X_1909_ _0558_ _0559_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q _0560_ VPWR VGND sg13g2_nand3_1
X_2958_ net1120 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q VPWR VGND sg13g2_dlhq_1
X_2889_ net1141 net1041 Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q VPWR VGND sg13g2_dlhq_1
XFILLER_45_404 VPWR VGND sg13g2_fill_1
XFILLER_40_120 VPWR VGND sg13g2_decap_8
XFILLER_0_260 VPWR VGND sg13g2_fill_1
X_2812_ net1168 net1025 Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q VPWR VGND sg13g2_dlhq_1
X_2743_ net1188 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q VPWR VGND sg13g2_dlhq_1
X_1625_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VPWR _0287_ VGND net66 Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
+ sg13g2_o21ai_1
X_1556_ _0219_ VPWR _0220_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0218_ sg13g2_o21ai_1
X_2674_ net1201 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q VPWR VGND sg13g2_dlhq_1
X_3157_ net1084 net198 VPWR VGND sg13g2_buf_1
X_1487_ _1037_ VPWR _0153_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0152_ sg13g2_o21ai_1
X_3226_ Inst_LUT4AB_switch_matrix.JS2BEG7 net276 VPWR VGND sg13g2_buf_1
XFILLER_42_429 VPWR VGND sg13g2_fill_1
XFILLER_42_418 VPWR VGND sg13g2_fill_1
X_2039_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0199_ _0685_ VPWR VGND sg13g2_mux4_1
X_2108_ Inst_LUT4AB_switch_matrix.JN2BEG7 Inst_LUT4AB_switch_matrix.E2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ _0748_ VPWR VGND sg13g2_mux2_1
X_3088_ E6END[7] net140 VPWR VGND sg13g2_buf_1
Xrebuffer5 _0590_ net378 VPWR VGND sg13g2_buf_2
X_1410_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0078_ _0079_ VPWR
+ VGND sg13g2_nor2b_1
X_1272_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q net49 net77 net104 Inst_LUT4AB_switch_matrix.JN2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q _1102_ VPWR VGND sg13g2_mux4_1
X_1341_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q net1010 net8 net37 net1212 Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ _0013_ VPWR VGND sg13g2_mux4_1
X_3011_ net1147 net1055 Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q VPWR VGND sg13g2_dlhq_1
X_2390_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ _0978_ _0976_ _0979_ _0977_ sg13g2_a221oi_1
X_2726_ net1136 net1106 Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q VPWR VGND sg13g2_dlhq_1
X_1608_ net61 net69 net987 _0271_ VPWR VGND sg13g2_mux2_1
X_2588_ net1168 net1085 Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q VPWR VGND sg13g2_dlhq_1
X_1539_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q _0197_ _0198_ _0170_ _0169_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
+ _0203_ VPWR VGND sg13g2_mux4_1
X_2657_ net1153 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VPWR VGND sg13g2_dlhq_1
X_3209_ NN4END[14] net250 VPWR VGND sg13g2_buf_1
XFILLER_58_381 VPWR VGND sg13g2_fill_1
X_1890_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_switch_matrix.M_AB
+ _0542_ _0541_ sg13g2_a21oi_1
X_2511_ net1118 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 VPWR
+ VGND sg13g2_dlhq_1
XFILLER_38_2 VPWR VGND sg13g2_fill_1
X_2442_ net1134 net1061 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2373_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q net963 Inst_LUT4AB_switch_matrix.JW2BEG1
+ net980 _0623_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q Inst_LUT4AB_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
X_1255_ net1000 net974 net968 net938 net961 Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ _1086_ VPWR VGND sg13g2_mux4_1
X_1186_ VPWR _1019_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VGND sg13g2_inv_1
X_1324_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1151_ _1152_ _1024_ sg13g2_a21oi_1
X_2709_ net1193 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q VPWR VGND sg13g2_dlhq_1
Xoutput251 net251 NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput262 net262 NN4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput240 net240 N4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput295 net295 S4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput273 net273 S2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput284 net284 S2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_30_229 VPWR VGND sg13g2_fill_2
XFILLER_2_174 VPWR VGND sg13g2_fill_2
XFILLER_38_307 VPWR VGND sg13g2_fill_2
XFILLER_0_44 VPWR VGND sg13g2_fill_2
X_1942_ net378 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ net374 _0592_ VPWR VGND sg13g2_mux4_1
X_2991_ net1119 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VPWR VGND sg13g2_dlhq_1
XFILLER_21_229 VPWR VGND sg13g2_fill_1
X_1873_ _0524_ VPWR _0525_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q _0521_ sg13g2_o21ai_1
XFILLER_56_104 VPWR VGND sg13g2_fill_1
X_2425_ _1007_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q net927 VPWR VGND sg13g2_nand2b_1
XFILLER_43_0 VPWR VGND sg13g2_fill_2
X_2356_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q net64 net79 net106 net945 Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ Inst_LUT4AB_switch_matrix.S4BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_56_159 VPWR VGND sg13g2_fill_2
XFILLER_56_126 VPWR VGND sg13g2_fill_2
XFILLER_52_321 VPWR VGND sg13g2_fill_2
X_2287_ VGND VPWR _0910_ _0911_ _0909_ _1049_ sg13g2_a21oi_2
X_1238_ VGND VPWR _1017_ _1069_ _1070_ _1018_ sg13g2_a21oi_1
X_1307_ _1136_ _1135_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q VPWR VGND sg13g2_nand2b_1
XFILLER_11_251 VPWR VGND sg13g2_fill_2
X_3190_ N4END[11] net246 VPWR VGND sg13g2_buf_1
X_2210_ VPWR _0844_ _0843_ VGND sg13g2_inv_1
X_2141_ _0771_ VPWR Inst_LUT4AB_switch_matrix.JW2BEG0 VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
+ _0778_ sg13g2_o21ai_1
X_2072_ _0714_ VPWR _0715_ VGND _0713_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q sg13g2_o21ai_1
X_1925_ net1007 net42 Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q _0576_ VPWR VGND sg13g2_mux2_1
X_2974_ net1162 net1049 Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q VPWR VGND sg13g2_dlhq_1
X_1856_ _0509_ _0508_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR VGND sg13g2_nand2b_1
X_1787_ _0442_ VPWR _0443_ VGND net68 net984 sg13g2_o21ai_1
X_2339_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q net932 _1158_ _0196_ _0290_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ _0955_ VPWR VGND sg13g2_mux4_1
X_2408_ net395 _0994_ _0992_ _0002_ VPWR VGND sg13g2_mux2_1
XFILLER_20_41 VPWR VGND sg13g2_fill_2
XFILLER_31_379 VPWR VGND sg13g2_decap_8
X_1572_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q _0233_ _0234_ _0235_ VPWR VGND sg13g2_nor3_1
X_1641_ Inst_LUT4AB_switch_matrix.E2BEG5 _0296_ _0302_ _0294_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_a22oi_1
X_2690_ net1152 net1098 Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q VPWR VGND sg13g2_dlhq_1
X_1710_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q _0365_ _0368_ _0367_
+ sg13g2_a21oi_1
X_3311_ WW4END[15] net352 VPWR VGND sg13g2_buf_1
Xfanout1081 FrameStrobe[15] net1081 VPWR VGND sg13g2_buf_1
X_3242_ S4END[11] net298 VPWR VGND sg13g2_buf_1
X_3173_ Inst_LUT4AB_switch_matrix.JN2BEG6 net223 VPWR VGND sg13g2_buf_1
X_2124_ net979 net972 _0669_ Inst_LUT4AB_switch_matrix.M_AB VPWR VGND sg13g2_mux2_2
Xfanout1070 FrameStrobe[17] net1070 VPWR VGND sg13g2_buf_1
Xfanout1092 FrameStrobe[13] net1092 VPWR VGND sg13g2_buf_1
Xrebuffer15 _0640_ net388 VPWR VGND sg13g2_buf_2
X_2055_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q net931 _0699_ _0698_ sg13g2_a21oi_1
XFILLER_25_19 VPWR VGND sg13g2_fill_1
X_1839_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0487_ _0493_ VPWR VGND sg13g2_mux4_1
X_1908_ _0559_ net103 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VPWR VGND sg13g2_nand2_1
X_2957_ net1123 net1047 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q VPWR VGND sg13g2_dlhq_1
X_2888_ net1174 net1038 Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q VPWR VGND sg13g2_dlhq_1
XFILLER_0_294 VPWR VGND sg13g2_fill_1
XFILLER_16_162 VPWR VGND sg13g2_fill_1
X_2811_ net1173 net1025 Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q VPWR VGND sg13g2_dlhq_1
X_2742_ net1190 net1014 Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q VPWR VGND sg13g2_dlhq_1
X_1555_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0219_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ _0217_ sg13g2_a21oi_2
X_2673_ net1206 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q VPWR VGND sg13g2_dlhq_1
X_1624_ _0285_ VPWR _0286_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q _0282_ sg13g2_o21ai_1
X_3156_ net1090 net197 VPWR VGND sg13g2_buf_1
X_3225_ Inst_LUT4AB_switch_matrix.JS2BEG6 net275 VPWR VGND sg13g2_buf_1
X_3087_ E6END[6] net139 VPWR VGND sg13g2_buf_1
X_1486_ net978 net972 net990 _0152_ VPWR VGND sg13g2_mux2_1
X_2107_ Inst_LUT4AB_switch_matrix.E2BEG7 _0741_ _0747_ _0739_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_a22oi_1
X_2038_ VGND VPWR _0684_ _0683_ _0676_ sg13g2_or2_1
XFILLER_22_143 VPWR VGND sg13g2_decap_8
Xrebuffer6 _0649_ net379 VPWR VGND sg13g2_buf_2
X_1340_ _0011_ VPWR _0012_ VGND _0010_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q sg13g2_o21ai_1
X_1271_ _1101_ _1094_ Inst_LUT4AB_switch_matrix.JN2BEG3 VPWR VGND sg13g2_nor2_2
X_3010_ net1152 net1055 Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q VPWR VGND sg13g2_dlhq_1
X_2656_ net1157 net1094 Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q VPWR VGND sg13g2_dlhq_1
X_2725_ net1139 net1104 Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q VPWR VGND sg13g2_dlhq_1
X_1469_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR _0136_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0133_ sg13g2_o21ai_1
X_1607_ _0269_ VPWR _0270_ VGND net87 net987 sg13g2_o21ai_1
X_2587_ net1171 net1085 Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q VPWR VGND sg13g2_dlhq_1
X_1538_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q _0147_ _0148_ _0130_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q
+ _0202_ VPWR VGND sg13g2_mux4_1
X_3208_ NN4END[13] net264 VPWR VGND sg13g2_buf_1
X_3139_ net1148 net181 VPWR VGND sg13g2_buf_1
XFILLER_27_279 VPWR VGND sg13g2_decap_8
XFILLER_23_430 VPWR VGND sg13g2_fill_2
XFILLER_53_71 VPWR VGND sg13g2_fill_2
XFILLER_37_94 VPWR VGND sg13g2_fill_2
XFILLER_33_205 VPWR VGND sg13g2_decap_8
X_2510_ net1122 net1071 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_dlhq_1
X_2441_ net1143 net1061 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_1323_ net94 net110 Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q _1151_ VPWR VGND sg13g2_mux2_1
X_2372_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q net957 _1159_ net384 _1118_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q
+ Inst_LUT4AB_switch_matrix.N1BEG3 VPWR VGND sg13g2_mux4_1
X_1185_ VPWR _1018_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VGND sg13g2_inv_1
X_1254_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q _1083_ _1084_ _1066_ _1065_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q
+ _1085_ VPWR VGND sg13g2_mux4_1
XFILLER_24_227 VPWR VGND sg13g2_fill_2
Xoutput252 net252 NN4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput241 net241 N4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput230 net230 N2BEGb[5] VPWR VGND sg13g2_buf_1
X_2639_ net1119 net1096 Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VPWR VGND sg13g2_dlhq_1
X_2708_ net1196 net1103 Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VPWR VGND sg13g2_dlhq_1
XFILLER_58_38 VPWR VGND sg13g2_fill_1
Xoutput263 net263 NN4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput274 Inst_LUT4AB_switch_matrix.JS2BEG5 S2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput285 net285 S4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput296 net296 S4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_55_352 VPWR VGND sg13g2_fill_1
XFILLER_3_0 VPWR VGND sg13g2_fill_2
XFILLER_48_82 VPWR VGND sg13g2_fill_2
X_1941_ _0590_ _0565_ _0591_ VPWR VGND sg13g2_nor2_2
X_1872_ _0522_ _0523_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q _0524_ VPWR VGND sg13g2_nand3_1
X_2990_ net1120 net1053 Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q VPWR VGND sg13g2_dlhq_1
XFILLER_50_2 VPWR VGND sg13g2_fill_1
X_2424_ net393 _1006_ _1004_ _0006_ VPWR VGND sg13g2_mux2_1
X_2286_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q VPWR _0910_ VGND _1049_ _0908_ sg13g2_o21ai_1
XFILLER_36_0 VPWR VGND sg13g2_fill_2
X_2355_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q net955 Inst_LUT4AB_switch_matrix.JS2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q Inst_LUT4AB_switch_matrix.W1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1306_ net81 net85 Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _1135_ VPWR VGND sg13g2_mux2_1
X_1237_ net956 net950 Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1069_ VPWR VGND sg13g2_mux2_1
XFILLER_52_388 VPWR VGND sg13g2_fill_2
XFILLER_20_285 VPWR VGND sg13g2_fill_1
XFILLER_20_296 VPWR VGND sg13g2_fill_1
XFILLER_43_322 VPWR VGND sg13g2_fill_1
XFILLER_38_105 VPWR VGND sg13g2_decap_8
X_2140_ _0777_ VPWR _0778_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0772_ sg13g2_o21ai_1
XFILLER_46_193 VPWR VGND sg13g2_decap_8
XFILLER_19_352 VPWR VGND sg13g2_fill_1
X_2071_ _0714_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0712_ VPWR VGND sg13g2_nand2b_1
X_1924_ _0574_ VPWR _0575_ VGND net5 net992 sg13g2_o21ai_1
X_1855_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q net34 net42 net5 net13 Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ _0508_ VPWR VGND sg13g2_mux4_1
X_2973_ net1165 net1049 Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q VPWR VGND sg13g2_dlhq_1
X_1786_ _0442_ net984 net1006 VPWR VGND sg13g2_nand2b_1
XFILLER_39_29 VPWR VGND sg13g2_fill_2
X_2338_ VGND VPWR _0954_ Inst_LUT4AB_switch_matrix.NN4BEG2 _0948_ _0952_ sg13g2_a21oi_2
XFILLER_29_105 VPWR VGND sg13g2_fill_2
X_2269_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _0626_ _0894_ _0893_
+ sg13g2_a21oi_1
X_2407_ Inst_LB_LUT4c_frame_config_dffesr.c_reset_value _0109_ _0993_ _0994_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_40_314 VPWR VGND sg13g2_fill_1
XFILLER_29_40 VPWR VGND sg13g2_fill_1
XFILLER_0_421 VPWR VGND sg13g2_fill_2
XFILLER_45_50 VPWR VGND sg13g2_fill_2
XFILLER_28_171 VPWR VGND sg13g2_decap_8
XFILLER_16_311 VPWR VGND sg13g2_decap_4
XFILLER_16_355 VPWR VGND sg13g2_fill_2
X_1571_ net49 Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0234_ VPWR VGND sg13g2_nor2_1
X_1640_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q _0301_ _0302_ VPWR VGND sg13g2_nor2_1
X_3310_ WW4END[14] net351 VPWR VGND sg13g2_buf_1
X_3241_ S4END[10] net297 VPWR VGND sg13g2_buf_1
X_2123_ _0762_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0761_ Inst_LUT4AB_switch_matrix.M_AH
+ VPWR VGND sg13g2_a21o_1
Xfanout1071 net1073 net1071 VPWR VGND sg13g2_buf_1
Xrebuffer16 _0348_ net389 VPWR VGND sg13g2_dlygate4sd1_1
Xfanout1060 net1062 net1060 VPWR VGND sg13g2_buf_1
Xfanout1093 net1094 net1093 VPWR VGND sg13g2_buf_1
Xfanout1082 net1086 net1082 VPWR VGND sg13g2_buf_1
X_2054_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q VPWR _0698_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ _1051_ sg13g2_o21ai_1
X_1838_ _0489_ _0491_ _0486_ _0492_ VPWR VGND sg13g2_mux2_1
X_1907_ _0558_ net76 Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VPWR VGND sg13g2_nand2b_1
X_2956_ net1127 net1049 Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VPWR VGND sg13g2_dlhq_1
X_2887_ net1207 net1038 Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VPWR VGND sg13g2_dlhq_1
X_1769_ _0425_ _0424_ VPWR VGND sg13g2_inv_2
XFILLER_9_307 VPWR VGND sg13g2_fill_1
XFILLER_9_329 VPWR VGND sg13g2_fill_2
XFILLER_0_251 VPWR VGND sg13g2_fill_1
XFILLER_31_122 VPWR VGND sg13g2_fill_2
X_2810_ net1178 net1025 Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q VPWR VGND sg13g2_dlhq_1
X_2741_ net1193 net1013 Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q VPWR VGND sg13g2_dlhq_1
X_2672_ net1116 net1101 Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q VPWR VGND sg13g2_dlhq_1
X_1554_ net976 net971 net998 _0218_ VPWR VGND sg13g2_mux2_1
X_1485_ _0150_ VPWR _0151_ VGND net990 net947 sg13g2_o21ai_1
X_1623_ _0285_ _0284_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q VPWR VGND sg13g2_nand2_2
.ends

