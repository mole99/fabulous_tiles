* NGSPICE file created from S_CPU_IRQ.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

.subckt S_CPU_IRQ CONFIGURED_top Co FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] IRQ_top0 IRQ_top1
+ IRQ_top2 IRQ_top3 N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13]
+ N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7]
+ N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14]
+ NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7]
+ NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0] S2END[1] S2END[2]
+ S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3]
+ S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11] S4END[12] S4END[13]
+ S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5] S4END[6] S4END[7]
+ S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13] SS4END[14]
+ SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6] SS4END[7]
+ SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_9_148 VPWR VGND sg13g2_fill_2
XFILLER_5_387 VPWR VGND sg13g2_decap_8
XFILLER_5_343 VPWR VGND sg13g2_decap_4
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_2_324 VPWR VGND sg13g2_decap_8
XFILLER_5_140 VPWR VGND sg13g2_decap_8
X_062_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q VPWR _024_ VGND Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q
+ net42 sg13g2_o21ai_1
X_131_ FrameStrobe[10] net81 VPWR VGND sg13g2_buf_1
XFILLER_9_33 VPWR VGND sg13g2_decap_8
XFILLER_0_79 VPWR VGND sg13g2_decap_8
XFILLER_0_68 VPWR VGND sg13g2_decap_8
XFILLER_2_187 VPWR VGND sg13g2_decap_8
X_114_ net9 net65 VPWR VGND sg13g2_buf_1
X_045_ _001_ _008_ net100 VPWR VGND sg13g2_nor2_1
XFILLER_3_430 VPWR VGND sg13g2_decap_8
XFILLER_0_422 VPWR VGND sg13g2_decap_8
XANTENNA_5 VPWR VGND net63 sg13g2_antennanp
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XFILLER_1_219 VPWR VGND sg13g2_fill_1
Xoutput64 net66 FrameData_O[26] VPWR VGND sg13g2_buf_1
Xoutput86 net88 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput97 net99 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
XFILLER_8_374 VPWR VGND sg13g2_fill_1
Xoutput53 net55 FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_0_296 VPWR VGND sg13g2_decap_8
Xoutput75 net77 FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_5_366 VPWR VGND sg13g2_decap_8
XFILLER_5_322 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_decap_8
XFILLER_2_303 VPWR VGND sg13g2_decap_8
XFILLER_5_196 VPWR VGND sg13g2_decap_8
X_130_ FrameStrobe[9] net99 VPWR VGND sg13g2_buf_1
XFILLER_9_89 VPWR VGND sg13g2_fill_2
X_061_ net46 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q _023_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_25 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_6_450 VPWR VGND sg13g2_fill_1
XFILLER_4_409 VPWR VGND sg13g2_decap_8
XFILLER_7_236 VPWR VGND sg13g2_decap_8
X_113_ net8 net64 VPWR VGND sg13g2_buf_1
X_044_ net1 VPWR _008_ VGND _004_ _007_ sg13g2_o21ai_1
XFILLER_0_401 VPWR VGND sg13g2_decap_8
XANTENNA_6 VPWR VGND net64 sg13g2_antennanp
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_3_261 VPWR VGND sg13g2_decap_8
XFILLER_3_294 VPWR VGND sg13g2_decap_8
Xoutput65 net67 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput87 net89 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput54 net56 FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_0_275 VPWR VGND sg13g2_decap_8
Xoutput98 net100 IRQ_top0 VPWR VGND sg13g2_buf_1
Xoutput76 net78 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_8_397 VPWR VGND sg13g2_decap_4
XFILLER_5_301 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_2_359 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_8
XFILLER_1_381 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_fill_1
X_060_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q _020_ _021_ _022_ VPWR VGND sg13g2_nor3_1
XFILLER_7_429 VPWR VGND sg13g2_fill_2
XFILLER_7_407 VPWR VGND sg13g2_decap_4
XFILLER_2_145 VPWR VGND sg13g2_fill_1
XFILLER_9_68 VPWR VGND sg13g2_decap_8
X_189_ net43 net143 VPWR VGND sg13g2_buf_1
X_043_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q VPWR _007_ VGND _005_ _006_ sg13g2_o21ai_1
X_112_ net7 net63 VPWR VGND sg13g2_buf_1
XFILLER_6_292 VPWR VGND sg13g2_fill_2
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_4_229 VPWR VGND sg13g2_fill_1
XANTENNA_7 VPWR VGND FrameData[10] sg13g2_antennanp
XFILLER_6_14 VPWR VGND sg13g2_decap_8
Xoutput66 net68 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput88 net90 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput55 net57 FrameData_O[18] VPWR VGND sg13g2_buf_1
XFILLER_0_254 VPWR VGND sg13g2_decap_8
Xoutput99 net101 IRQ_top1 VPWR VGND sg13g2_buf_1
Xoutput77 net79 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_8_332 VPWR VGND sg13g2_decap_8
XFILLER_10_309 VPWR VGND sg13g2_decap_4
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_2_338 VPWR VGND sg13g2_decap_8
XFILLER_5_154 VPWR VGND sg13g2_decap_8
XFILLER_1_360 VPWR VGND sg13g2_decap_8
XFILLER_4_91 VPWR VGND sg13g2_decap_8
XFILLER_9_47 VPWR VGND sg13g2_decap_8
X_188_ net44 net142 VPWR VGND sg13g2_buf_1
XFILLER_9_290 VPWR VGND sg13g2_fill_1
X_042_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q VPWR _006_ VGND Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q
+ net40 sg13g2_o21ai_1
XFILLER_3_444 VPWR VGND sg13g2_decap_8
X_111_ net4 net62 VPWR VGND sg13g2_buf_1
XFILLER_1_81 VPWR VGND sg13g2_fill_1
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XANTENNA_8 VPWR VGND FrameData[11] sg13g2_antennanp
XFILLER_0_436 VPWR VGND sg13g2_fill_2
Xoutput67 net69 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput89 net91 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput78 net80 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput56 net58 FrameData_O[19] VPWR VGND sg13g2_buf_1
XFILLER_0_233 VPWR VGND sg13g2_decap_8
XFILLER_8_311 VPWR VGND sg13g2_fill_2
XFILLER_7_80 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_fill_1
XFILLER_5_336 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_8_185 VPWR VGND sg13g2_decap_8
XFILLER_5_133 VPWR VGND sg13g2_decap_8
XFILLER_2_317 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_9_26 VPWR VGND sg13g2_decap_8
X_187_ net45 net141 VPWR VGND sg13g2_buf_1
XFILLER_7_217 VPWR VGND sg13g2_fill_1
XFILLER_7_206 VPWR VGND sg13g2_decap_8
X_110_ net3 net61 VPWR VGND sg13g2_buf_1
X_041_ net44 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q _005_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_415 VPWR VGND sg13g2_decap_8
XFILLER_10_80 VPWR VGND sg13g2_decap_4
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_3_275 VPWR VGND sg13g2_fill_1
XANTENNA_9 VPWR VGND FrameData[18] sg13g2_antennanp
XFILLER_0_212 VPWR VGND sg13g2_decap_8
Xoutput46 net48 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput57 net59 FrameData_O[1] VPWR VGND sg13g2_buf_1
Xoutput79 net81 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
XFILLER_8_367 VPWR VGND sg13g2_decap_8
XFILLER_0_289 VPWR VGND sg13g2_decap_8
Xoutput68 net70 FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_5_359 VPWR VGND sg13g2_decap_8
XFILLER_5_315 VPWR VGND sg13g2_decap_8
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_8_131 VPWR VGND sg13g2_fill_1
XFILLER_4_381 VPWR VGND sg13g2_decap_8
XFILLER_5_189 VPWR VGND sg13g2_decap_8
XFILLER_5_112 VPWR VGND sg13g2_decap_8
X_186_ net46 net155 VPWR VGND sg13g2_buf_1
XFILLER_9_16 VPWR VGND sg13g2_fill_2
XFILLER_6_432 VPWR VGND sg13g2_decap_8
XFILLER_9_281 VPWR VGND sg13g2_decap_8
XFILLER_7_229 VPWR VGND sg13g2_decap_8
X_040_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q _002_ _003_ _004_ VPWR VGND sg13g2_nor3_1
XFILLER_10_280 VPWR VGND sg13g2_fill_1
X_169_ net39 net138 VPWR VGND sg13g2_buf_1
XFILLER_6_284 VPWR VGND sg13g2_fill_2
XFILLER_0_438 VPWR VGND sg13g2_fill_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_3_254 VPWR VGND sg13g2_decap_8
XFILLER_3_287 VPWR VGND sg13g2_decap_8
Xoutput69 net71 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput58 net60 FrameData_O[20] VPWR VGND sg13g2_buf_1
XFILLER_8_346 VPWR VGND sg13g2_fill_2
XFILLER_0_268 VPWR VGND sg13g2_decap_8
Xoutput47 net49 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_5_168 VPWR VGND sg13g2_decap_8
XFILLER_1_374 VPWR VGND sg13g2_decap_8
XFILLER_10_451 VPWR VGND sg13g2_fill_1
X_185_ net47 net154 VPWR VGND sg13g2_buf_1
XFILLER_2_138 VPWR VGND sg13g2_fill_2
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
X_099_ FrameData[10] net49 VPWR VGND sg13g2_buf_1
X_168_ S4END[8] net137 VPWR VGND sg13g2_buf_1
XFILLER_6_252 VPWR VGND sg13g2_decap_8
XFILLER_3_211 VPWR VGND sg13g2_decap_8
Xoutput59 net61 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_8_325 VPWR VGND sg13g2_decap_8
XFILLER_0_247 VPWR VGND sg13g2_decap_8
Xoutput48 net50 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_7_94 VPWR VGND sg13g2_decap_8
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_1_353 VPWR VGND sg13g2_decap_8
XFILLER_4_84 VPWR VGND sg13g2_decap_8
XFILLER_2_106 VPWR VGND sg13g2_fill_2
X_184_ SS4END[8] net153 VPWR VGND sg13g2_buf_1
XFILLER_6_412 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
X_167_ S4END[9] net136 VPWR VGND sg13g2_buf_1
X_098_ FrameData[9] net79 VPWR VGND sg13g2_buf_1
XFILLER_6_286 VPWR VGND sg13g2_fill_1
XFILLER_6_231 VPWR VGND sg13g2_decap_8
XFILLER_3_437 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_0_429 VPWR VGND sg13g2_decap_8
Xoutput49 net51 FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_0_226 VPWR VGND sg13g2_decap_8
XFILLER_7_73 VPWR VGND sg13g2_decap_8
XFILLER_5_329 VPWR VGND sg13g2_decap_8
XFILLER_4_395 VPWR VGND sg13g2_decap_8
XFILLER_5_126 VPWR VGND sg13g2_decap_8
XFILLER_1_332 VPWR VGND sg13g2_decap_8
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_4_181 VPWR VGND sg13g2_decap_8
X_183_ SS4END[9] net152 VPWR VGND sg13g2_buf_1
XFILLER_9_295 VPWR VGND sg13g2_fill_1
XFILLER_6_210 VPWR VGND sg13g2_decap_8
XFILLER_3_405 VPWR VGND sg13g2_fill_2
X_166_ S4END[10] net135 VPWR VGND sg13g2_buf_1
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_097_ FrameData[8] net78 VPWR VGND sg13g2_buf_1
XFILLER_10_73 VPWR VGND sg13g2_decap_8
XFILLER_0_408 VPWR VGND sg13g2_decap_8
XFILLER_3_268 VPWR VGND sg13g2_decap_8
XFILLER_10_84 VPWR VGND sg13g2_fill_1
X_149_ net31 net112 VPWR VGND sg13g2_buf_1
XFILLER_0_205 VPWR VGND sg13g2_decap_8
XFILLER_7_393 VPWR VGND sg13g2_fill_1
XFILLER_7_382 VPWR VGND sg13g2_fill_2
XFILLER_7_52 VPWR VGND sg13g2_decap_8
XFILLER_5_308 VPWR VGND sg13g2_decap_8
XFILLER_4_341 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_decap_8
XFILLER_5_105 VPWR VGND sg13g2_decap_8
XFILLER_1_311 VPWR VGND sg13g2_decap_8
XFILLER_1_388 VPWR VGND sg13g2_decap_4
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_4_160 VPWR VGND sg13g2_decap_8
X_182_ SS4END[10] net151 VPWR VGND sg13g2_buf_1
XFILLER_6_425 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_9_274 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_10_273 VPWR VGND sg13g2_decap_8
X_165_ S4END[11] net134 VPWR VGND sg13g2_buf_1
XFILLER_6_277 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
X_096_ FrameData[7] net77 VPWR VGND sg13g2_buf_1
XFILLER_10_52 VPWR VGND sg13g2_decap_8
X_148_ S2MID[4] net111 VPWR VGND sg13g2_buf_1
XFILLER_3_247 VPWR VGND sg13g2_decap_8
X_079_ net7 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q VPWR VGND sg13g2_dlhq_1
XFILLER_8_339 VPWR VGND sg13g2_decap_8
XFILLER_7_361 VPWR VGND sg13g2_decap_8
XFILLER_7_31 VPWR VGND sg13g2_decap_8
XFILLER_4_320 VPWR VGND sg13g2_decap_8
XFILLER_1_367 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_4_98 VPWR VGND sg13g2_decap_8
X_181_ SS4END[11] net150 VPWR VGND sg13g2_buf_1
XFILLER_1_142 VPWR VGND sg13g2_fill_1
XFILLER_1_175 VPWR VGND sg13g2_decap_8
X_164_ S4END[12] net133 VPWR VGND sg13g2_buf_1
XFILLER_6_245 VPWR VGND sg13g2_decap_8
XFILLER_1_99 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_4
X_095_ FrameData[6] net76 VPWR VGND sg13g2_buf_1
XFILLER_10_31 VPWR VGND sg13g2_decap_8
XFILLER_3_204 VPWR VGND sg13g2_decap_8
X_147_ S2MID[5] net110 VPWR VGND sg13g2_buf_1
X_078_ net4 net6 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q VPWR VGND sg13g2_dlhq_1
XFILLER_8_307 VPWR VGND sg13g2_decap_4
XFILLER_7_87 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_fill_2
XFILLER_7_192 VPWR VGND sg13g2_decap_8
XFILLER_1_346 VPWR VGND sg13g2_decap_8
XFILLER_4_77 VPWR VGND sg13g2_decap_8
XFILLER_4_195 VPWR VGND sg13g2_decap_8
X_180_ SS4END[12] net149 VPWR VGND sg13g2_buf_1
XFILLER_6_405 VPWR VGND sg13g2_decap_8
XFILLER_9_221 VPWR VGND sg13g2_decap_4
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XS_CPU_IRQ_155 VPWR VGND Co sg13g2_tielo
XFILLER_3_419 VPWR VGND sg13g2_decap_8
X_163_ S4END[13] net132 VPWR VGND sg13g2_buf_1
XFILLER_6_224 VPWR VGND sg13g2_decap_8
X_094_ FrameData[5] net75 VPWR VGND sg13g2_buf_1
XFILLER_1_56 VPWR VGND sg13g2_decap_8
X_146_ S2MID[6] net109 VPWR VGND sg13g2_buf_1
X_077_ net3 net6 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q VPWR VGND sg13g2_dlhq_1
XFILLER_2_282 VPWR VGND sg13g2_decap_8
XFILLER_0_219 VPWR VGND sg13g2_decap_8
XFILLER_7_352 VPWR VGND sg13g2_decap_4
XFILLER_7_66 VPWR VGND sg13g2_decap_8
X_129_ FrameStrobe[8] net98 VPWR VGND sg13g2_buf_1
XFILLER_4_388 VPWR VGND sg13g2_decap_8
XFILLER_7_160 VPWR VGND sg13g2_fill_1
XFILLER_5_119 VPWR VGND sg13g2_decap_8
XFILLER_1_325 VPWR VGND sg13g2_decap_8
XFILLER_0_380 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_4_174 VPWR VGND sg13g2_decap_8
XFILLER_9_244 VPWR VGND sg13g2_decap_8
XFILLER_6_439 VPWR VGND sg13g2_fill_2
XFILLER_9_288 VPWR VGND sg13g2_fill_2
XFILLER_5_450 VPWR VGND sg13g2_fill_1
X_162_ S4END[14] net131 VPWR VGND sg13g2_buf_1
XFILLER_6_203 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
X_093_ FrameData[4] net74 VPWR VGND sg13g2_buf_1
XFILLER_5_280 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_10_66 VPWR VGND sg13g2_decap_8
Xinput1 CONFIGURED_top net1 VPWR VGND sg13g2_buf_1
X_145_ S2MID[7] net108 VPWR VGND sg13g2_buf_1
X_076_ net2 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q VPWR VGND sg13g2_dlhq_1
XANTENNA_50 VPWR VGND FrameData[10] sg13g2_antennanp
X_059_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q net34 _021_ VPWR VGND sg13g2_nor2_1
XFILLER_7_375 VPWR VGND sg13g2_decap_8
XFILLER_7_331 VPWR VGND sg13g2_decap_8
XFILLER_7_45 VPWR VGND sg13g2_decap_8
X_128_ FrameStrobe[7] net97 VPWR VGND sg13g2_buf_1
XFILLER_4_334 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_1_304 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_4_153 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_1_123 VPWR VGND sg13g2_decap_4
XFILLER_9_267 VPWR VGND sg13g2_decap_8
XFILLER_9_212 VPWR VGND sg13g2_fill_1
X_161_ S4END[15] net124 VPWR VGND sg13g2_buf_1
XFILLER_6_259 VPWR VGND sg13g2_fill_1
XFILLER_1_14 VPWR VGND sg13g2_decap_8
X_092_ FrameData[3] net73 VPWR VGND sg13g2_buf_1
XFILLER_10_45 VPWR VGND sg13g2_decap_8
Xinput2 FrameData[20] net2 VPWR VGND sg13g2_buf_1
XFILLER_3_218 VPWR VGND sg13g2_fill_1
X_075_ _028_ _035_ net103 VPWR VGND sg13g2_nor2_1
X_144_ net16 net107 VPWR VGND sg13g2_buf_1
XFILLER_2_251 VPWR VGND sg13g2_fill_2
XANTENNA_40 VPWR VGND FrameData[10] sg13g2_antennanp
XANTENNA_51 VPWR VGND FrameData[11] sg13g2_antennanp
X_058_ net38 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q _020_ VPWR VGND sg13g2_nor2b_1
X_127_ FrameStrobe[6] net96 VPWR VGND sg13g2_buf_1
XFILLER_4_313 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_132 VPWR VGND sg13g2_decap_8
XFILLER_10_404 VPWR VGND sg13g2_decap_4
XFILLER_6_419 VPWR VGND sg13g2_fill_2
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_6_238 VPWR VGND sg13g2_decap_8
X_160_ net20 net123 VPWR VGND sg13g2_buf_1
X_091_ FrameData[2] net70 VPWR VGND sg13g2_buf_1
Xinput3 FrameData[21] net3 VPWR VGND sg13g2_buf_1
XFILLER_10_24 VPWR VGND sg13g2_decap_8
X_074_ net1 VPWR _035_ VGND _031_ _034_ sg13g2_o21ai_1
X_143_ net17 net106 VPWR VGND sg13g2_buf_1
XFILLER_2_296 VPWR VGND sg13g2_decap_8
XANTENNA_30 VPWR VGND FrameData[10] sg13g2_antennanp
XANTENNA_41 VPWR VGND FrameData[11] sg13g2_antennanp
XANTENNA_52 VPWR VGND FrameData[8] sg13g2_antennanp
X_057_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q _018_ _019_ VPWR VGND sg13g2_nor2_1
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_126_ FrameStrobe[5] net95 VPWR VGND sg13g2_buf_1
XFILLER_7_185 VPWR VGND sg13g2_decap_8
X_109_ net2 net60 VPWR VGND sg13g2_buf_1
XFILLER_3_380 VPWR VGND sg13g2_decap_8
XFILLER_3_391 VPWR VGND sg13g2_decap_8
XFILLER_1_339 VPWR VGND sg13g2_decap_8
XFILLER_0_394 VPWR VGND sg13g2_decap_8
XFILLER_4_188 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_5_91 VPWR VGND sg13g2_decap_8
XFILLER_0_191 VPWR VGND sg13g2_decap_8
XFILLER_6_217 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
X_090_ FrameData[1] net59 VPWR VGND sg13g2_buf_1
XFILLER_2_445 VPWR VGND sg13g2_decap_4
Xinput4 FrameData[22] net4 VPWR VGND sg13g2_buf_1
XFILLER_5_294 VPWR VGND sg13g2_decap_8
X_142_ net18 net105 VPWR VGND sg13g2_buf_1
X_073_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q VPWR _034_ VGND _032_ _033_ sg13g2_o21ai_1
XFILLER_2_253 VPWR VGND sg13g2_fill_1
XFILLER_2_275 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XANTENNA_53 VPWR VGND net63 sg13g2_antennanp
XANTENNA_20 VPWR VGND FrameData[11] sg13g2_antennanp
XANTENNA_31 VPWR VGND FrameData[11] sg13g2_antennanp
XANTENNA_42 VPWR VGND FrameData[8] sg13g2_antennanp
XFILLER_2_70 VPWR VGND sg13g2_decap_8
X_056_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q net18 net30 net22 net26 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q
+ _018_ VPWR VGND sg13g2_mux4_1
XFILLER_7_356 VPWR VGND sg13g2_fill_1
XFILLER_7_345 VPWR VGND sg13g2_decap_8
XFILLER_7_59 VPWR VGND sg13g2_decap_8
X_125_ FrameStrobe[4] net94 VPWR VGND sg13g2_buf_1
Xinput40 SS4END[2] net42 VPWR VGND sg13g2_buf_1
XFILLER_8_109 VPWR VGND sg13g2_fill_1
X_108_ FrameData[19] net58 VPWR VGND sg13g2_buf_1
X_039_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q net32 _003_ VPWR VGND sg13g2_nor2_1
XFILLER_1_318 VPWR VGND sg13g2_decap_8
XFILLER_0_373 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_4_112 VPWR VGND sg13g2_decap_8
XFILLER_4_167 VPWR VGND sg13g2_decap_8
XFILLER_9_237 VPWR VGND sg13g2_decap_8
XFILLER_1_137 VPWR VGND sg13g2_fill_1
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_0_170 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
Xinput5 FrameData[23] net7 VPWR VGND sg13g2_buf_1
XFILLER_5_273 VPWR VGND sg13g2_decap_8
XFILLER_10_59 VPWR VGND sg13g2_decap_8
X_072_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q VPWR _033_ VGND Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q
+ net43 sg13g2_o21ai_1
X_141_ net19 net104 VPWR VGND sg13g2_buf_1
XANTENNA_54 VPWR VGND net64 sg13g2_antennanp
XANTENNA_43 VPWR VGND net63 sg13g2_antennanp
XANTENNA_32 VPWR VGND FrameData[8] sg13g2_antennanp
XFILLER_2_82 VPWR VGND sg13g2_fill_2
XANTENNA_10 VPWR VGND FrameData[8] sg13g2_antennanp
XANTENNA_21 VPWR VGND FrameData[18] sg13g2_antennanp
Xoutput150 net152 NN4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_7_368 VPWR VGND sg13g2_decap_8
XFILLER_7_324 VPWR VGND sg13g2_decap_8
XFILLER_7_38 VPWR VGND sg13g2_decap_8
X_124_ FrameStrobe[3] net93 VPWR VGND sg13g2_buf_1
X_055_ _010_ _017_ net101 VPWR VGND sg13g2_nor2_1
Xinput41 SS4END[3] net43 VPWR VGND sg13g2_buf_1
Xinput30 S4END[0] net32 VPWR VGND sg13g2_buf_1
XFILLER_4_327 VPWR VGND sg13g2_decap_8
XFILLER_7_143 VPWR VGND sg13g2_fill_1
XFILLER_7_132 VPWR VGND sg13g2_decap_8
X_107_ FrameData[18] net57 VPWR VGND sg13g2_buf_1
X_038_ net36 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q _002_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_92 VPWR VGND sg13g2_decap_8
XFILLER_0_352 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_146 VPWR VGND sg13g2_decap_8
XFILLER_3_190 VPWR VGND sg13g2_decap_8
XFILLER_8_8 VPWR VGND sg13g2_decap_8
XFILLER_1_127 VPWR VGND sg13g2_fill_1
XFILLER_5_422 VPWR VGND sg13g2_decap_8
XFILLER_5_252 VPWR VGND sg13g2_decap_8
XFILLER_10_38 VPWR VGND sg13g2_decap_8
Xinput6 FrameData[24] net8 VPWR VGND sg13g2_buf_1
X_071_ net47 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q _032_ VPWR VGND sg13g2_nor2b_1
X_140_ FrameStrobe[19] net90 VPWR VGND sg13g2_buf_1
XANTENNA_11 VPWR VGND net63 sg13g2_antennanp
XANTENNA_33 VPWR VGND net63 sg13g2_antennanp
Xoutput140 net142 NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput151 net153 NN4BEG[7] VPWR VGND sg13g2_buf_1
XANTENNA_44 VPWR VGND net64 sg13g2_antennanp
XANTENNA_22 VPWR VGND FrameData[8] sg13g2_antennanp
Xinput31 S4END[1] net33 VPWR VGND sg13g2_buf_1
Xinput20 S2END[2] net22 VPWR VGND sg13g2_buf_1
X_123_ FrameStrobe[2] net92 VPWR VGND sg13g2_buf_1
X_054_ net1 VPWR _017_ VGND _013_ _016_ sg13g2_o21ai_1
Xinput42 SS4END[4] net44 VPWR VGND sg13g2_buf_1
XFILLER_6_391 VPWR VGND sg13g2_decap_8
XFILLER_4_306 VPWR VGND sg13g2_decap_8
XFILLER_7_199 VPWR VGND sg13g2_decap_8
XFILLER_7_166 VPWR VGND sg13g2_decap_4
X_106_ FrameData[17] net56 VPWR VGND sg13g2_buf_1
X_037_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit22.Q _000_ _001_ VPWR VGND sg13g2_nor2_1
XFILLER_8_71 VPWR VGND sg13g2_decap_8
XFILLER_0_331 VPWR VGND sg13g2_decap_8
XFILLER_4_125 VPWR VGND sg13g2_decap_8
XFILLER_1_117 VPWR VGND sg13g2_fill_2
XFILLER_1_106 VPWR VGND sg13g2_decap_8
XFILLER_5_401 VPWR VGND sg13g2_decap_8
XFILLER_8_283 VPWR VGND sg13g2_fill_2
XFILLER_5_231 VPWR VGND sg13g2_decap_8
XFILLER_2_415 VPWR VGND sg13g2_fill_2
Xinput7 FrameData[25] net9 VPWR VGND sg13g2_buf_1
X_070_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q _029_ _030_ _031_ VPWR VGND sg13g2_nor3_1
XFILLER_2_201 VPWR VGND sg13g2_decap_8
XFILLER_2_289 VPWR VGND sg13g2_decap_8
XFILLER_2_84 VPWR VGND sg13g2_fill_1
XANTENNA_12 VPWR VGND net64 sg13g2_antennanp
XANTENNA_23 VPWR VGND net63 sg13g2_antennanp
XANTENNA_45 VPWR VGND FrameData[10] sg13g2_antennanp
Xoutput141 net143 NN4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput152 net154 NN4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput130 net132 N4BEG[2] VPWR VGND sg13g2_buf_1
XANTENNA_34 VPWR VGND net64 sg13g2_antennanp
XFILLER_2_0 VPWR VGND sg13g2_decap_8
X_053_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q VPWR _016_ VGND _014_ _015_ sg13g2_o21ai_1
X_122_ FrameStrobe[1] net91 VPWR VGND sg13g2_buf_1
Xinput43 SS4END[5] net45 VPWR VGND sg13g2_buf_1
Xinput32 S4END[2] net34 VPWR VGND sg13g2_buf_1
Xinput21 S2END[3] net23 VPWR VGND sg13g2_buf_1
Xinput10 FrameData[28] net12 VPWR VGND sg13g2_buf_1
XFILLER_6_370 VPWR VGND sg13g2_fill_2
XFILLER_7_101 VPWR VGND sg13g2_decap_8
X_105_ FrameData[16] net55 VPWR VGND sg13g2_buf_1
XFILLER_8_50 VPWR VGND sg13g2_decap_8
XFILLER_7_178 VPWR VGND sg13g2_decap_8
X_036_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit20.Q net16 net28 net20 net24 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit21.Q
+ _000_ VPWR VGND sg13g2_mux4_1
XFILLER_3_373 VPWR VGND sg13g2_decap_8
XFILLER_0_310 VPWR VGND sg13g2_decap_8
XFILLER_8_454 VPWR VGND sg13g2_fill_1
XFILLER_8_410 VPWR VGND sg13g2_decap_8
XFILLER_0_387 VPWR VGND sg13g2_decap_8
XFILLER_0_184 VPWR VGND sg13g2_decap_8
XFILLER_8_262 VPWR VGND sg13g2_decap_8
XFILLER_5_84 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_2_449 VPWR VGND sg13g2_fill_2
Xinput8 FrameData[26] net10 VPWR VGND sg13g2_buf_1
XFILLER_5_287 VPWR VGND sg13g2_decap_8
XFILLER_5_210 VPWR VGND sg13g2_decap_8
XANTENNA_13 VPWR VGND FrameData[10] sg13g2_antennanp
XANTENNA_35 VPWR VGND FrameData[10] sg13g2_antennanp
Xoutput142 net144 NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput153 net155 NN4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput120 net122 N2BEGb[6] VPWR VGND sg13g2_buf_1
XANTENNA_46 VPWR VGND FrameData[11] sg13g2_antennanp
Xoutput131 net133 N4BEG[3] VPWR VGND sg13g2_buf_1
XANTENNA_24 VPWR VGND net64 sg13g2_antennanp
XFILLER_1_290 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_121_ net5 net80 VPWR VGND sg13g2_buf_1
XFILLER_7_338 VPWR VGND sg13g2_decap_8
X_052_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q VPWR _015_ VGND Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q
+ net41 sg13g2_o21ai_1
Xinput44 SS4END[6] net46 VPWR VGND sg13g2_buf_1
Xinput33 S4END[3] net35 VPWR VGND sg13g2_buf_1
Xinput22 S2END[4] net24 VPWR VGND sg13g2_buf_1
Xinput11 FrameData[29] net13 VPWR VGND sg13g2_buf_1
X_104_ FrameData[15] net54 VPWR VGND sg13g2_buf_1
XFILLER_3_352 VPWR VGND sg13g2_decap_8
XFILLER_4_105 VPWR VGND sg13g2_decap_8
XFILLER_0_366 VPWR VGND sg13g2_decap_8
XFILLER_5_436 VPWR VGND sg13g2_fill_1
XFILLER_0_163 VPWR VGND sg13g2_decap_8
XFILLER_8_241 VPWR VGND sg13g2_decap_8
XFILLER_5_63 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_fill_1
Xinput9 FrameData[27] net11 VPWR VGND sg13g2_buf_1
XFILLER_5_266 VPWR VGND sg13g2_decap_8
XANTENNA_25 VPWR VGND FrameData[10] sg13g2_antennanp
Xoutput143 net145 NN4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput132 net134 N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput121 net123 N2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput110 net112 N2BEG[4] VPWR VGND sg13g2_buf_1
XANTENNA_36 VPWR VGND FrameData[11] sg13g2_antennanp
XANTENNA_14 VPWR VGND FrameData[11] sg13g2_antennanp
XANTENNA_47 VPWR VGND FrameData[8] sg13g2_antennanp
XFILLER_2_42 VPWR VGND sg13g2_decap_8
Xoutput154 net156 UserCLKo VPWR VGND sg13g2_buf_1
X_120_ net15 net72 VPWR VGND sg13g2_buf_1
X_051_ net45 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q _014_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_390 VPWR VGND sg13g2_decap_8
Xinput45 SS4END[7] net47 VPWR VGND sg13g2_buf_1
Xinput34 S4END[4] net36 VPWR VGND sg13g2_buf_1
Xinput23 S2END[5] net25 VPWR VGND sg13g2_buf_1
Xinput12 FrameData[30] net14 VPWR VGND sg13g2_buf_1
XFILLER_6_372 VPWR VGND sg13g2_fill_1
X_103_ FrameData[14] net53 VPWR VGND sg13g2_buf_1
XFILLER_7_158 VPWR VGND sg13g2_fill_2
XFILLER_7_125 VPWR VGND sg13g2_decap_8
XFILLER_8_85 VPWR VGND sg13g2_decap_8
XFILLER_8_401 VPWR VGND sg13g2_fill_1
XFILLER_0_345 VPWR VGND sg13g2_decap_8
XFILLER_4_139 VPWR VGND sg13g2_decap_8
XFILLER_3_150 VPWR VGND sg13g2_decap_8
XFILLER_3_172 VPWR VGND sg13g2_fill_1
XFILLER_5_415 VPWR VGND sg13g2_decap_8
XFILLER_8_220 VPWR VGND sg13g2_decap_8
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_0_142 VPWR VGND sg13g2_decap_8
XFILLER_5_245 VPWR VGND sg13g2_decap_8
XANTENNA_48 VPWR VGND net63 sg13g2_antennanp
XANTENNA_26 VPWR VGND FrameData[11] sg13g2_antennanp
XANTENNA_37 VPWR VGND FrameData[8] sg13g2_antennanp
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XANTENNA_15 VPWR VGND FrameData[18] sg13g2_antennanp
Xoutput144 net146 NN4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput133 net135 N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput122 net124 N4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput111 net113 N2BEG[5] VPWR VGND sg13g2_buf_1
Xoutput100 net102 IRQ_top2 VPWR VGND sg13g2_buf_1
X_050_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q _011_ _012_ _013_ VPWR VGND sg13g2_nor3_1
X_179_ SS4END[13] net148 VPWR VGND sg13g2_buf_1
Xinput35 S4END[5] net37 VPWR VGND sg13g2_buf_1
Xinput24 S2END[6] net26 VPWR VGND sg13g2_buf_1
Xinput13 FrameData[31] net15 VPWR VGND sg13g2_buf_1
XFILLER_6_384 VPWR VGND sg13g2_decap_8
X_102_ FrameData[13] net52 VPWR VGND sg13g2_buf_1
XFILLER_7_148 VPWR VGND sg13g2_fill_1
XFILLER_0_0 VPWR VGND sg13g2_fill_2
XFILLER_3_398 VPWR VGND sg13g2_decap_8
XFILLER_8_64 VPWR VGND sg13g2_decap_8
XFILLER_0_324 VPWR VGND sg13g2_decap_8
XFILLER_8_424 VPWR VGND sg13g2_fill_2
XFILLER_3_140 VPWR VGND sg13g2_decap_4
XFILLER_8_276 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_0_198 VPWR VGND sg13g2_decap_8
XFILLER_0_121 VPWR VGND sg13g2_decap_8
XFILLER_5_98 VPWR VGND sg13g2_decap_8
XFILLER_5_224 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_4
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_fill_1
XANTENNA_38 VPWR VGND net63 sg13g2_antennanp
XFILLER_9_382 VPWR VGND sg13g2_fill_1
Xoutput145 net147 NN4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput123 net125 N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput134 net136 N4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput112 net114 N2BEG[6] VPWR VGND sg13g2_buf_1
XANTENNA_49 VPWR VGND net64 sg13g2_antennanp
Xoutput101 net103 IRQ_top3 VPWR VGND sg13g2_buf_1
XANTENNA_27 VPWR VGND FrameData[8] sg13g2_antennanp
XANTENNA_16 VPWR VGND FrameData[8] sg13g2_antennanp
Xinput36 S4END[6] net38 VPWR VGND sg13g2_buf_1
Xinput25 S2END[7] net27 VPWR VGND sg13g2_buf_1
Xinput14 S1END[0] net16 VPWR VGND sg13g2_buf_1
X_178_ SS4END[14] net147 VPWR VGND sg13g2_buf_1
XFILLER_6_363 VPWR VGND sg13g2_decap_8
XFILLER_6_352 VPWR VGND sg13g2_fill_2
X_101_ FrameData[12] net51 VPWR VGND sg13g2_buf_1
XFILLER_3_322 VPWR VGND sg13g2_decap_8
XFILLER_3_333 VPWR VGND sg13g2_fill_1
XFILLER_3_366 VPWR VGND sg13g2_decap_8
XFILLER_8_43 VPWR VGND sg13g2_decap_8
XFILLER_6_182 VPWR VGND sg13g2_decap_8
XFILLER_0_303 VPWR VGND sg13g2_decap_8
XFILLER_4_119 VPWR VGND sg13g2_fill_2
XFILLER_0_177 VPWR VGND sg13g2_decap_8
XFILLER_0_100 VPWR VGND sg13g2_decap_8
XFILLER_8_255 VPWR VGND sg13g2_fill_2
XFILLER_5_77 VPWR VGND sg13g2_decap_8
XFILLER_5_203 VPWR VGND sg13g2_decap_8
XFILLER_1_283 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XANTENNA_17 VPWR VGND net63 sg13g2_antennanp
XFILLER_9_361 VPWR VGND sg13g2_decap_8
Xoutput146 net148 NN4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput124 net126 N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput135 net137 N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput113 net115 N2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput102 net104 N1BEG[0] VPWR VGND sg13g2_buf_1
XANTENNA_28 VPWR VGND net63 sg13g2_antennanp
XANTENNA_39 VPWR VGND net64 sg13g2_antennanp
Xinput37 S4END[7] net39 VPWR VGND sg13g2_buf_1
Xinput26 S2MID[0] net28 VPWR VGND sg13g2_buf_1
Xinput15 S1END[1] net17 VPWR VGND sg13g2_buf_1
X_177_ SS4END[15] net140 VPWR VGND sg13g2_buf_1
XFILLER_6_342 VPWR VGND sg13g2_decap_4
X_100_ FrameData[11] net50 VPWR VGND sg13g2_buf_1
XFILLER_7_139 VPWR VGND sg13g2_decap_4
XFILLER_8_99 VPWR VGND sg13g2_fill_2
XFILLER_8_22 VPWR VGND sg13g2_decap_8
XFILLER_6_161 VPWR VGND sg13g2_decap_8
XFILLER_0_2 VPWR VGND sg13g2_fill_1
XFILLER_3_301 VPWR VGND sg13g2_decap_8
XFILLER_3_345 VPWR VGND sg13g2_decap_8
XFILLER_0_359 VPWR VGND sg13g2_decap_8
XFILLER_3_164 VPWR VGND sg13g2_decap_4
XFILLER_3_197 VPWR VGND sg13g2_decap_8
XFILLER_5_429 VPWR VGND sg13g2_decap_8
XFILLER_0_156 VPWR VGND sg13g2_decap_8
XFILLER_8_234 VPWR VGND sg13g2_decap_8
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_5_259 VPWR VGND sg13g2_decap_8
XFILLER_4_292 VPWR VGND sg13g2_decap_8
X_193_ UserCLK net156 VPWR VGND sg13g2_buf_1
XANTENNA_18 VPWR VGND net64 sg13g2_antennanp
XANTENNA_29 VPWR VGND net64 sg13g2_antennanp
XFILLER_9_351 VPWR VGND sg13g2_fill_2
Xoutput147 net149 NN4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput125 net127 N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput136 net138 N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput114 net116 N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput103 net105 N1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_1_262 VPWR VGND sg13g2_decap_8
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_10_383 VPWR VGND sg13g2_decap_8
Xinput38 SS4END[0] net40 VPWR VGND sg13g2_buf_1
Xinput16 S1END[2] net18 VPWR VGND sg13g2_buf_1
Xinput27 S2MID[1] net29 VPWR VGND sg13g2_buf_1
XFILLER_6_398 VPWR VGND sg13g2_decap_8
XFILLER_6_354 VPWR VGND sg13g2_fill_1
XFILLER_6_321 VPWR VGND sg13g2_decap_8
X_176_ net32 net130 VPWR VGND sg13g2_buf_1
XFILLER_8_78 VPWR VGND sg13g2_decap_8
XFILLER_6_140 VPWR VGND sg13g2_decap_8
X_159_ net21 net122 VPWR VGND sg13g2_buf_1
XFILLER_2_390 VPWR VGND sg13g2_fill_1
XFILLER_0_338 VPWR VGND sg13g2_decap_8
XFILLER_5_408 VPWR VGND sg13g2_decap_8
XFILLER_0_135 VPWR VGND sg13g2_decap_8
XFILLER_8_257 VPWR VGND sg13g2_fill_1
XFILLER_8_213 VPWR VGND sg13g2_decap_8
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_4_430 VPWR VGND sg13g2_decap_8
XFILLER_5_238 VPWR VGND sg13g2_decap_8
X_192_ net40 net146 VPWR VGND sg13g2_buf_1
XFILLER_2_208 VPWR VGND sg13g2_fill_1
XANTENNA_19 VPWR VGND FrameData[10] sg13g2_antennanp
Xoutput148 net150 NN4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput126 net128 N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput137 net139 N4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput115 net117 N2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput104 net106 N1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_1_241 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
Xinput39 SS4END[1] net41 VPWR VGND sg13g2_buf_1
Xinput28 S2MID[2] net30 VPWR VGND sg13g2_buf_1
Xinput17 S1END[3] net19 VPWR VGND sg13g2_buf_1
XFILLER_6_377 VPWR VGND sg13g2_decap_8
X_175_ net33 net129 VPWR VGND sg13g2_buf_1
XFILLER_8_57 VPWR VGND sg13g2_decap_8
X_158_ net22 net121 VPWR VGND sg13g2_buf_1
XFILLER_6_196 VPWR VGND sg13g2_decap_8
XFILLER_2_380 VPWR VGND sg13g2_fill_2
X_089_ FrameData[0] net48 VPWR VGND sg13g2_buf_1
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_0_317 VPWR VGND sg13g2_decap_8
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_fill_1
XFILLER_8_269 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_0_114 VPWR VGND sg13g2_decap_8
XFILLER_5_217 VPWR VGND sg13g2_decap_8
XFILLER_1_401 VPWR VGND sg13g2_fill_2
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_1_445 VPWR VGND sg13g2_fill_2
XFILLER_9_375 VPWR VGND sg13g2_decap_8
XFILLER_1_297 VPWR VGND sg13g2_decap_8
X_191_ net41 net145 VPWR VGND sg13g2_buf_1
Xoutput149 net151 NN4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput138 net140 NN4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput127 net129 N4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput116 net118 N2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput105 net107 N1BEG[3] VPWR VGND sg13g2_buf_1
Xinput18 S2END[0] net20 VPWR VGND sg13g2_buf_1
Xinput29 S2MID[3] net31 VPWR VGND sg13g2_buf_1
X_174_ net34 net128 VPWR VGND sg13g2_buf_1
XFILLER_3_91 VPWR VGND sg13g2_decap_8
XFILLER_3_315 VPWR VGND sg13g2_decap_8
XFILLER_3_359 VPWR VGND sg13g2_decap_8
X_157_ net23 net120 VPWR VGND sg13g2_buf_1
XFILLER_8_36 VPWR VGND sg13g2_decap_8
XFILLER_6_175 VPWR VGND sg13g2_decap_8
XFILLER_8_248 VPWR VGND sg13g2_decap_8
XFILLER_7_281 VPWR VGND sg13g2_fill_2
XFILLER_4_262 VPWR VGND sg13g2_decap_8
XFILLER_4_273 VPWR VGND sg13g2_fill_2
XFILLER_6_91 VPWR VGND sg13g2_decap_8
X_190_ net42 net144 VPWR VGND sg13g2_buf_1
XFILLER_1_276 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_9_321 VPWR VGND sg13g2_fill_2
Xoutput139 net141 NN4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput128 net130 N4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput117 net119 N2BEGb[3] VPWR VGND sg13g2_buf_1
Xoutput106 net108 N2BEG[0] VPWR VGND sg13g2_buf_1
X_173_ net35 net127 VPWR VGND sg13g2_buf_1
Xinput19 S2END[1] net21 VPWR VGND sg13g2_buf_1
XFILLER_6_335 VPWR VGND sg13g2_decap_8
XFILLER_6_302 VPWR VGND sg13g2_decap_8
XFILLER_10_397 VPWR VGND sg13g2_decap_8
XFILLER_9_162 VPWR VGND sg13g2_fill_2
XFILLER_6_346 VPWR VGND sg13g2_fill_2
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_3_338 VPWR VGND sg13g2_decap_8
XFILLER_8_15 VPWR VGND sg13g2_decap_8
X_087_ net15 net6 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_154 VPWR VGND sg13g2_decap_8
X_156_ net24 net119 VPWR VGND sg13g2_buf_1
XFILLER_3_157 VPWR VGND sg13g2_decap_8
X_139_ FrameStrobe[18] net89 VPWR VGND sg13g2_buf_1
XFILLER_0_93 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_fill_1
XFILLER_8_227 VPWR VGND sg13g2_decap_8
XFILLER_0_149 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_444 VPWR VGND sg13g2_decap_8
XFILLER_1_403 VPWR VGND sg13g2_fill_1
XFILLER_1_425 VPWR VGND sg13g2_fill_1
XFILLER_4_241 VPWR VGND sg13g2_decap_8
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_1_255 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_9_300 VPWR VGND sg13g2_decap_8
Xoutput129 net131 N4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput118 net120 N2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput107 net109 N2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_10_376 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_6_314 VPWR VGND sg13g2_decap_8
X_172_ net36 net126 VPWR VGND sg13g2_buf_1
XFILLER_5_380 VPWR VGND sg13g2_decap_8
XFILLER_6_133 VPWR VGND sg13g2_decap_8
X_155_ net25 net118 VPWR VGND sg13g2_buf_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
X_086_ net14 net6 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q VPWR VGND sg13g2_dlhq_1
X_138_ FrameStrobe[17] net88 VPWR VGND sg13g2_buf_1
XFILLER_7_431 VPWR VGND sg13g2_fill_1
X_069_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q net35 _030_ VPWR VGND sg13g2_nor2_1
XFILLER_2_180 VPWR VGND sg13g2_decap_8
XFILLER_0_128 VPWR VGND sg13g2_decap_8
XFILLER_0_61 VPWR VGND sg13g2_decap_8
XFILLER_0_50 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_4_423 VPWR VGND sg13g2_decap_8
XFILLER_7_283 VPWR VGND sg13g2_fill_1
XFILLER_7_250 VPWR VGND sg13g2_fill_2
Xoutput90 net92 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput119 net121 N2BEGb[5] VPWR VGND sg13g2_buf_1
Xoutput108 net110 N2BEG[2] VPWR VGND sg13g2_buf_1
X_171_ net37 net125 VPWR VGND sg13g2_buf_1
XFILLER_9_164 VPWR VGND sg13g2_fill_1
XFILLER_3_329 VPWR VGND sg13g2_decap_4
X_154_ net26 net117 VPWR VGND sg13g2_buf_1
X_085_ net13 net6 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_189 VPWR VGND sg13g2_decap_8
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_2_373 VPWR VGND sg13g2_decap_8
XFILLER_2_395 VPWR VGND sg13g2_fill_2
X_137_ FrameStrobe[16] net87 VPWR VGND sg13g2_buf_1
X_068_ net39 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q _029_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_82 VPWR VGND sg13g2_decap_8
XFILLER_0_107 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_9_368 VPWR VGND sg13g2_decap_8
Xoutput109 net111 N2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput80 net82 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput91 net93 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_170_ net38 net139 VPWR VGND sg13g2_buf_1
XFILLER_3_84 VPWR VGND sg13g2_decap_8
XFILLER_3_308 VPWR VGND sg13g2_decap_8
X_153_ net27 net116 VPWR VGND sg13g2_buf_1
X_084_ net12 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q VPWR VGND sg13g2_dlhq_1
XFILLER_8_29 VPWR VGND sg13g2_decap_8
XFILLER_6_168 VPWR VGND sg13g2_decap_8
XFILLER_2_352 VPWR VGND sg13g2_decap_8
XFILLER_7_422 VPWR VGND sg13g2_decap_8
X_136_ FrameStrobe[15] net86 VPWR VGND sg13g2_buf_1
XFILLER_3_105 VPWR VGND sg13g2_decap_4
XFILLER_9_61 VPWR VGND sg13g2_decap_8
X_067_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit31.Q _027_ _028_ VPWR VGND sg13g2_nor2_1
XFILLER_7_274 VPWR VGND sg13g2_decap_8
XFILLER_7_252 VPWR VGND sg13g2_fill_1
X_119_ net14 net71 VPWR VGND sg13g2_buf_1
XFILLER_4_255 VPWR VGND sg13g2_decap_8
XFILLER_4_299 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_9_314 VPWR VGND sg13g2_decap_8
XFILLER_1_269 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
Xoutput70 net72 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput81 net83 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput92 net94 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_391 VPWR VGND sg13g2_fill_2
XFILLER_6_328 VPWR VGND sg13g2_decap_8
XFILLER_5_394 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
X_083_ net11 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit27.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_147 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
X_152_ net28 net115 VPWR VGND sg13g2_buf_1
XFILLER_2_331 VPWR VGND sg13g2_decap_8
XFILLER_2_397 VPWR VGND sg13g2_fill_1
XFILLER_9_40 VPWR VGND sg13g2_decap_8
X_135_ FrameStrobe[14] net85 VPWR VGND sg13g2_buf_1
X_066_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit29.Q net19 net31 net23 net27 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit30.Q
+ _027_ VPWR VGND sg13g2_mux4_1
XFILLER_0_86 VPWR VGND sg13g2_decap_8
XFILLER_2_150 VPWR VGND sg13g2_fill_2
XFILLER_2_194 VPWR VGND sg13g2_decap_8
XFILLER_4_437 VPWR VGND sg13g2_decap_8
X_118_ net13 net69 VPWR VGND sg13g2_buf_1
X_049_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q net33 _012_ VPWR VGND sg13g2_nor2_1
XFILLER_4_234 VPWR VGND sg13g2_decap_8
XANTENNA_1 VPWR VGND FrameData[10] sg13g2_antennanp
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_1_248 VPWR VGND sg13g2_decap_8
Xoutput60 net62 FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput82 net84 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput93 net95 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput71 net73 FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_10_369 VPWR VGND sg13g2_decap_8
XFILLER_5_373 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
X_082_ net10 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit26.Q VPWR VGND sg13g2_dlhq_1
XFILLER_6_126 VPWR VGND sg13g2_decap_8
X_151_ net29 net114 VPWR VGND sg13g2_buf_1
XFILLER_2_310 VPWR VGND sg13g2_decap_8
X_065_ _019_ _026_ net102 VPWR VGND sg13g2_nor2_1
X_134_ FrameStrobe[13] net84 VPWR VGND sg13g2_buf_1
XFILLER_0_43 VPWR VGND sg13g2_decap_8
XFILLER_0_32 VPWR VGND sg13g2_decap_8
XFILLER_2_173 VPWR VGND sg13g2_decap_8
X_117_ net12 net68 VPWR VGND sg13g2_buf_1
XFILLER_7_243 VPWR VGND sg13g2_decap_8
XFILLER_4_416 VPWR VGND sg13g2_decap_8
X_048_ net37 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q _011_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_202 VPWR VGND sg13g2_fill_2
XANTENNA_2 VPWR VGND FrameData[11] sg13g2_antennanp
XFILLER_6_42 VPWR VGND sg13g2_decap_8
Xoutput61 net63 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput83 net85 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput94 net96 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
Xoutput50 net52 FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_0_282 VPWR VGND sg13g2_decap_8
Xoutput72 net74 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_360 VPWR VGND sg13g2_decap_8
XFILLER_9_179 VPWR VGND sg13g2_fill_1
XFILLER_5_352 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
X_150_ net30 net113 VPWR VGND sg13g2_buf_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
X_081_ net9 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_dlhq_1
XFILLER_5_182 VPWR VGND sg13g2_decap_8
XFILLER_2_366 VPWR VGND sg13g2_decap_8
X_133_ FrameStrobe[12] net83 VPWR VGND sg13g2_buf_1
X_064_ net1 VPWR _026_ VGND _022_ _025_ sg13g2_o21ai_1
XFILLER_7_447 VPWR VGND sg13g2_fill_1
XFILLER_9_75 VPWR VGND sg13g2_decap_8
X_116_ net11 net67 VPWR VGND sg13g2_buf_1
XFILLER_7_222 VPWR VGND sg13g2_decap_8
X_047_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit25.Q _009_ _010_ VPWR VGND sg13g2_nor2_1
Xfanout5 FrameStrobe[0] net5 VPWR VGND sg13g2_buf_1
XFILLER_6_98 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_4_225 VPWR VGND sg13g2_decap_4
XFILLER_4_269 VPWR VGND sg13g2_decap_4
XANTENNA_3 VPWR VGND FrameData[18] sg13g2_antennanp
XFILLER_1_217 VPWR VGND sg13g2_fill_2
XFILLER_3_280 VPWR VGND sg13g2_decap_8
Xoutput62 net64 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput84 net86 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
Xoutput95 net97 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
Xoutput51 net53 FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_0_261 VPWR VGND sg13g2_decap_8
Xoutput73 net75 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_6_309 VPWR VGND sg13g2_fill_1
XFILLER_9_169 VPWR VGND sg13g2_fill_2
XFILLER_3_77 VPWR VGND sg13g2_decap_8
X_080_ net8 net5 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q VPWR VGND sg13g2_dlhq_1
XFILLER_2_345 VPWR VGND sg13g2_decap_8
XFILLER_5_161 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_fill_2
X_132_ FrameStrobe[11] net82 VPWR VGND sg13g2_buf_1
XFILLER_7_415 VPWR VGND sg13g2_decap_8
X_063_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit28.Q VPWR _025_ VGND _023_ _024_ sg13g2_o21ai_1
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_9_54 VPWR VGND sg13g2_decap_8
X_115_ net10 net66 VPWR VGND sg13g2_buf_1
X_046_ Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit23.Q net17 net29 net21 net25 Inst_S_CPU_IRQ_ConfigMem.Inst_frame0_bit24.Q
+ _009_ VPWR VGND sg13g2_mux4_1
Xfanout6 FrameStrobe[0] net6 VPWR VGND sg13g2_buf_1
XFILLER_4_248 VPWR VGND sg13g2_decap_8
XFILLER_6_77 VPWR VGND sg13g2_decap_8
XANTENNA_4 VPWR VGND FrameData[8] sg13g2_antennanp
XFILLER_9_307 VPWR VGND sg13g2_decap_8
Xoutput52 net54 FrameData_O[15] VPWR VGND sg13g2_buf_1
Xoutput63 net65 FrameData_O[25] VPWR VGND sg13g2_buf_1
Xoutput85 net87 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
Xoutput96 net98 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
XFILLER_0_240 VPWR VGND sg13g2_decap_8
Xoutput74 net76 FrameData_O[6] VPWR VGND sg13g2_buf_1
.ends

