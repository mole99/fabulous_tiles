module DSP (Tile_X0Y0_UserCLKo,
    Tile_X0Y1_UserCLK,
    Tile_X0Y0_E1BEG,
    Tile_X0Y0_E1END,
    Tile_X0Y0_E2BEG,
    Tile_X0Y0_E2BEGb,
    Tile_X0Y0_E2END,
    Tile_X0Y0_E2MID,
    Tile_X0Y0_E6BEG,
    Tile_X0Y0_E6END,
    Tile_X0Y0_EE4BEG,
    Tile_X0Y0_EE4END,
    Tile_X0Y0_FrameData,
    Tile_X0Y0_FrameData_O,
    Tile_X0Y0_FrameStrobe_O,
    Tile_X0Y0_N1BEG,
    Tile_X0Y0_N2BEG,
    Tile_X0Y0_N2BEGb,
    Tile_X0Y0_N4BEG,
    Tile_X0Y0_NN4BEG,
    Tile_X0Y0_S1END,
    Tile_X0Y0_S2END,
    Tile_X0Y0_S2MID,
    Tile_X0Y0_S4END,
    Tile_X0Y0_SS4END,
    Tile_X0Y0_W1BEG,
    Tile_X0Y0_W1END,
    Tile_X0Y0_W2BEG,
    Tile_X0Y0_W2BEGb,
    Tile_X0Y0_W2END,
    Tile_X0Y0_W2MID,
    Tile_X0Y0_W6BEG,
    Tile_X0Y0_W6END,
    Tile_X0Y0_WW4BEG,
    Tile_X0Y0_WW4END,
    Tile_X0Y1_E1BEG,
    Tile_X0Y1_E1END,
    Tile_X0Y1_E2BEG,
    Tile_X0Y1_E2BEGb,
    Tile_X0Y1_E2END,
    Tile_X0Y1_E2MID,
    Tile_X0Y1_E6BEG,
    Tile_X0Y1_E6END,
    Tile_X0Y1_EE4BEG,
    Tile_X0Y1_EE4END,
    Tile_X0Y1_FrameData,
    Tile_X0Y1_FrameData_O,
    Tile_X0Y1_FrameStrobe,
    Tile_X0Y1_N1END,
    Tile_X0Y1_N2END,
    Tile_X0Y1_N2MID,
    Tile_X0Y1_N4END,
    Tile_X0Y1_NN4END,
    Tile_X0Y1_S1BEG,
    Tile_X0Y1_S2BEG,
    Tile_X0Y1_S2BEGb,
    Tile_X0Y1_S4BEG,
    Tile_X0Y1_SS4BEG,
    Tile_X0Y1_W1BEG,
    Tile_X0Y1_W1END,
    Tile_X0Y1_W2BEG,
    Tile_X0Y1_W2BEGb,
    Tile_X0Y1_W2END,
    Tile_X0Y1_W2MID,
    Tile_X0Y1_W6BEG,
    Tile_X0Y1_W6END,
    Tile_X0Y1_WW4BEG,
    Tile_X0Y1_WW4END);
 output Tile_X0Y0_UserCLKo;
 input Tile_X0Y1_UserCLK;
 output [3:0] Tile_X0Y0_E1BEG;
 input [3:0] Tile_X0Y0_E1END;
 output [7:0] Tile_X0Y0_E2BEG;
 output [7:0] Tile_X0Y0_E2BEGb;
 input [7:0] Tile_X0Y0_E2END;
 input [7:0] Tile_X0Y0_E2MID;
 output [11:0] Tile_X0Y0_E6BEG;
 input [11:0] Tile_X0Y0_E6END;
 output [15:0] Tile_X0Y0_EE4BEG;
 input [15:0] Tile_X0Y0_EE4END;
 input [31:0] Tile_X0Y0_FrameData;
 output [31:0] Tile_X0Y0_FrameData_O;
 output [19:0] Tile_X0Y0_FrameStrobe_O;
 output [3:0] Tile_X0Y0_N1BEG;
 output [7:0] Tile_X0Y0_N2BEG;
 output [7:0] Tile_X0Y0_N2BEGb;
 output [15:0] Tile_X0Y0_N4BEG;
 output [15:0] Tile_X0Y0_NN4BEG;
 input [3:0] Tile_X0Y0_S1END;
 input [7:0] Tile_X0Y0_S2END;
 input [7:0] Tile_X0Y0_S2MID;
 input [15:0] Tile_X0Y0_S4END;
 input [15:0] Tile_X0Y0_SS4END;
 output [3:0] Tile_X0Y0_W1BEG;
 input [3:0] Tile_X0Y0_W1END;
 output [7:0] Tile_X0Y0_W2BEG;
 output [7:0] Tile_X0Y0_W2BEGb;
 input [7:0] Tile_X0Y0_W2END;
 input [7:0] Tile_X0Y0_W2MID;
 output [11:0] Tile_X0Y0_W6BEG;
 input [11:0] Tile_X0Y0_W6END;
 output [15:0] Tile_X0Y0_WW4BEG;
 input [15:0] Tile_X0Y0_WW4END;
 output [3:0] Tile_X0Y1_E1BEG;
 input [3:0] Tile_X0Y1_E1END;
 output [7:0] Tile_X0Y1_E2BEG;
 output [7:0] Tile_X0Y1_E2BEGb;
 input [7:0] Tile_X0Y1_E2END;
 input [7:0] Tile_X0Y1_E2MID;
 output [11:0] Tile_X0Y1_E6BEG;
 input [11:0] Tile_X0Y1_E6END;
 output [15:0] Tile_X0Y1_EE4BEG;
 input [15:0] Tile_X0Y1_EE4END;
 input [31:0] Tile_X0Y1_FrameData;
 output [31:0] Tile_X0Y1_FrameData_O;
 input [19:0] Tile_X0Y1_FrameStrobe;
 input [3:0] Tile_X0Y1_N1END;
 input [7:0] Tile_X0Y1_N2END;
 input [7:0] Tile_X0Y1_N2MID;
 input [15:0] Tile_X0Y1_N4END;
 input [15:0] Tile_X0Y1_NN4END;
 output [3:0] Tile_X0Y1_S1BEG;
 output [7:0] Tile_X0Y1_S2BEG;
 output [7:0] Tile_X0Y1_S2BEGb;
 output [15:0] Tile_X0Y1_S4BEG;
 output [15:0] Tile_X0Y1_SS4BEG;
 output [3:0] Tile_X0Y1_W1BEG;
 input [3:0] Tile_X0Y1_W1END;
 output [7:0] Tile_X0Y1_W2BEG;
 output [7:0] Tile_X0Y1_W2BEGb;
 input [7:0] Tile_X0Y1_W2END;
 input [7:0] Tile_X0Y1_W2MID;
 output [11:0] Tile_X0Y1_W6BEG;
 input [11:0] Tile_X0Y1_W6END;
 output [15:0] Tile_X0Y1_WW4BEG;
 input [15:0] Tile_X0Y1_WW4END;

 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ;
 wire \Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ;
 wire \Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ;
 wire net728;
 wire net730;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net734;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net726;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net732;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net733;
 wire net736;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net648;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net731;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire \Tile_X0Y1_DSP_bot.A0 ;
 wire \Tile_X0Y1_DSP_bot.A1 ;
 wire \Tile_X0Y1_DSP_bot.A2 ;
 wire \Tile_X0Y1_DSP_bot.A3 ;
 wire \Tile_X0Y1_DSP_bot.B0 ;
 wire \Tile_X0Y1_DSP_bot.B1 ;
 wire \Tile_X0Y1_DSP_bot.B2 ;
 wire \Tile_X0Y1_DSP_bot.B3 ;
 wire \Tile_X0Y1_DSP_bot.C0 ;
 wire \Tile_X0Y1_DSP_bot.C1 ;
 wire \Tile_X0Y1_DSP_bot.C2 ;
 wire \Tile_X0Y1_DSP_bot.C3 ;
 wire \Tile_X0Y1_DSP_bot.C4 ;
 wire \Tile_X0Y1_DSP_bot.C5 ;
 wire \Tile_X0Y1_DSP_bot.C6 ;
 wire \Tile_X0Y1_DSP_bot.C7 ;
 wire \Tile_X0Y1_DSP_bot.C8 ;
 wire \Tile_X0Y1_DSP_bot.C9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ;
 wire \Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ;
 wire \Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ;
 wire net374;
 wire net375;
 wire net376;
 wire net727;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net729;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net735;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net649;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net617;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net687;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net554;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net667;
 wire net668;
 wire net669;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;

 sg13g2_o21ai_1 _2468_ (.B1(_0557_),
    .Y(_0558_),
    .A1(net1680),
    .A2(net1521));
 sg13g2_a21oi_1 _2469_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0558_),
    .Y(_0559_),
    .B1(_0108_));
 sg13g2_a21oi_1 _2470_ (.A1(_0556_),
    .A2(_0559_),
    .Y(_0560_),
    .B1(_0109_));
 sg13g2_mux2_1 _2471_ (.A0(net142),
    .A1(net53),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .X(_0561_));
 sg13g2_nor2b_1 _2472_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ),
    .B_N(net169),
    .Y(_0562_));
 sg13g2_a21oi_2 _2473_ (.B1(_0562_),
    .Y(_0563_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_nand2_2 _2474_ (.Y(_0564_),
    .A(_0563_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_o21ai_1 _2475_ (.B1(_0564_),
    .Y(_0565_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ),
    .A2(_0561_));
 sg13g2_inv_1 _2476_ (.Y(_0566_),
    .A(net684));
 sg13g2_mux4_1 _2477_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(net1529),
    .A1(net636),
    .A2(net1550),
    .A3(net1560),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0567_));
 sg13g2_mux4_1 _2478_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(net1565),
    .A1(net1572),
    .A2(net1579),
    .A3(net1618),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0568_));
 sg13g2_nand2b_1 _2479_ (.Y(_0569_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A_N(_0568_));
 sg13g2_o21ai_1 _2480_ (.B1(_0569_),
    .Y(_0570_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0567_));
 sg13g2_mux4_1 _2481_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(net1712),
    .A1(net118),
    .A2(net94),
    .A3(net1922),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0571_));
 sg13g2_nand2b_1 _2482_ (.Y(_0572_),
    .B(_0571_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_nand2b_1 _2483_ (.Y(_0573_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .A_N(net168));
 sg13g2_o21ai_1 _2484_ (.B1(_0573_),
    .Y(_0574_),
    .A1(net154),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_nand2_1 _2485_ (.Y(_0575_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ),
    .B(net53));
 sg13g2_o21ai_1 _2486_ (.B1(_0575_),
    .Y(_0576_),
    .A1(_0068_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_o21ai_1 _2487_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0577_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0576_));
 sg13g2_a21oi_1 _2488_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0574_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nor2_1 _2489_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ),
    .B(_0578_),
    .Y(_0579_));
 sg13g2_a22oi_1 _2490_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .B1(_0572_),
    .B2(_0579_),
    .A2(_0570_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_inv_1 _2491_ (.Y(_0580_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ));
 sg13g2_mux4_1 _2492_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net1632),
    .A1(net1585),
    .A2(net1522),
    .A3(net1520),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0581_));
 sg13g2_mux4_1 _2493_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net1597),
    .A1(net1610),
    .A2(net649),
    .A3(net1623),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_0582_));
 sg13g2_nand2b_1 _2494_ (.Y(_0583_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .A_N(_0581_));
 sg13g2_o21ai_1 _2495_ (.B1(_0583_),
    .Y(_0584_),
    .A1(_0582_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_mux4_1 _2496_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .A0(net1516),
    .A1(net2003),
    .A2(net129),
    .A3(net10),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_0585_));
 sg13g2_nor2b_1 _2497_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .B_N(_0585_),
    .Y(_0586_));
 sg13g2_nor2_1 _2498_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .B(net28),
    .Y(_0587_));
 sg13g2_a21oi_1 _2499_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0086_),
    .Y(_0588_),
    .B1(_0587_));
 sg13g2_nand2b_1 _2500_ (.Y(_0589_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ),
    .A_N(net1932));
 sg13g2_o21ai_1 _2501_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net62),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_o21ai_1 _2502_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ),
    .Y(_0591_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .A2(_0588_));
 sg13g2_a21oi_1 _2503_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ),
    .A2(_0590_),
    .Y(_0592_),
    .B1(_0591_));
 sg13g2_nor3_1 _2504_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .B(_0586_),
    .C(_0592_),
    .Y(_0593_));
 sg13g2_a21o_2 _2505_ (.A2(_0584_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ),
    .B1(_0593_),
    .X(_0594_));
 sg13g2_inv_8 _2506_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A(_0594_));
 sg13g2_mux4_1 _2507_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(_0083_),
    .A1(_0084_),
    .A2(_0594_),
    .A3(_0085_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0595_));
 sg13g2_inv_1 _2508_ (.Y(_0596_),
    .A(net643));
 sg13g2_mux4_1 _2509_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ),
    .A0(net1562),
    .A1(_0580_),
    .A2(_0595_),
    .A3(_0565_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ),
    .X(_0597_));
 sg13g2_inv_1 _2510_ (.Y(_0598_),
    .A(net621));
 sg13g2_a21oi_1 _2511_ (.A1(net124),
    .A2(net1680),
    .Y(_0599_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_o21ai_1 _2512_ (.B1(_0599_),
    .Y(_0600_),
    .A1(net1680),
    .A2(net610));
 sg13g2_nor2b_1 _2513_ (.A(net1680),
    .B_N(net136),
    .Y(_0601_));
 sg13g2_a21oi_1 _2514_ (.A1(net1680),
    .A2(net23),
    .Y(_0602_),
    .B1(_0601_));
 sg13g2_a21oi_1 _2515_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0602_),
    .Y(_0603_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_a21oi_1 _2516_ (.A1(net31),
    .A2(net1681),
    .Y(_0604_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_o21ai_1 _2517_ (.B1(_0604_),
    .Y(_0605_),
    .A1(_0075_),
    .A2(net1680));
 sg13g2_nand2_1 _2518_ (.Y(_0606_),
    .A(_0076_),
    .B(net1681));
 sg13g2_o21ai_1 _2519_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net66),
    .A2(net1681));
 sg13g2_a21oi_1 _2520_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0607_),
    .Y(_0608_),
    .B1(_0108_));
 sg13g2_a221oi_1 _2521_ (.B2(_0608_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ),
    .B1(_0605_),
    .A1(_0600_),
    .Y(_0609_),
    .A2(_0603_));
 sg13g2_a21oi_2 _2522_ (.B1(_0609_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .A2(_0560_),
    .A1(_0554_));
 sg13g2_inv_2 _2523_ (.Y(_0610_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ));
 sg13g2_mux4_1 _2524_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net136),
    .A1(net55),
    .A2(net69),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0611_));
 sg13g2_inv_1 _2525_ (.Y(_0612_),
    .A(_0611_));
 sg13g2_mux4_1 _2526_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .A0(_0435_),
    .A1(_0081_),
    .A2(_0080_),
    .A3(_0082_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0613_));
 sg13g2_mux4_1 _2527_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ),
    .A0(net723),
    .A1(net45),
    .A2(net19),
    .A3(net80),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0614_));
 sg13g2_mux4_1 _2528_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ),
    .A0(net1590),
    .A1(_0610_),
    .A2(_0613_),
    .A3(_0612_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ),
    .X(_0615_));
 sg13g2_inv_4 _2529_ (.A(_0615_),
    .Y(_0616_));
 sg13g2_a21o_1 _2530_ (.A2(net1660),
    .A1(_0099_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0617_));
 sg13g2_a21oi_1 _2531_ (.A1(_0107_),
    .A2(_0615_),
    .Y(_0618_),
    .B1(_0617_));
 sg13g2_o21ai_1 _2532_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0619_),
    .A1(net148),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_a21oi_1 _2533_ (.A1(_0104_),
    .A2(net1660),
    .Y(_0620_),
    .B1(_0619_));
 sg13g2_nor2b_1 _2534_ (.A(_0620_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0621_));
 sg13g2_inv_1 _2535_ (.Y(_0622_),
    .A(_0621_));
 sg13g2_mux4_1 _2536_ (.S0(net1660),
    .A0(net1712),
    .A1(net120),
    .A2(net1927),
    .A3(net96),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0623_));
 sg13g2_nor2_1 _2537_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_nor2_1 _2538_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_o21ai_1 _2539_ (.B1(_0625_),
    .Y(_0626_),
    .A1(_0618_),
    .A2(_0622_));
 sg13g2_nor2b_2 _2540_ (.A(_0552_),
    .B_N(_0626_),
    .Y(_0627_));
 sg13g2_inv_8 _2541_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A(_0627_));
 sg13g2_a21oi_1 _2542_ (.A1(net16),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .Y(_0628_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_o21ai_1 _2543_ (.B1(_0628_),
    .Y(_0629_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .A2(_0627_));
 sg13g2_nand2b_2 _2544_ (.Y(_0630_),
    .B(_0629_),
    .A_N(_0544_));
 sg13g2_a21oi_1 _2545_ (.A1(_0083_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .Y(_0631_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_o21ai_1 _2546_ (.B1(_0631_),
    .Y(_0632_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(net1527));
 sg13g2_mux2_1 _2547_ (.A0(net2),
    .A1(net9),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0633_));
 sg13g2_a21oi_1 _2548_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0633_),
    .Y(_0634_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_mux4_1 _2549_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A0(net27),
    .A1(net35),
    .A2(net29),
    .A3(net1933),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0635_));
 sg13g2_o21ai_1 _2550_ (.B1(_0093_),
    .Y(_0636_),
    .A1(_0092_),
    .A2(_0635_));
 sg13g2_a21oi_1 _2551_ (.A1(_0632_),
    .A2(_0634_),
    .Y(_0637_),
    .B1(_0636_));
 sg13g2_nand2b_1 _2552_ (.Y(_0638_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A_N(net1588));
 sg13g2_o21ai_1 _2553_ (.B1(_0638_),
    .Y(_0639_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(net1593));
 sg13g2_mux2_1 _2554_ (.A0(net1524),
    .A1(net1520),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0640_));
 sg13g2_a21oi_1 _2555_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0640_),
    .Y(_0641_),
    .B1(_0092_));
 sg13g2_o21ai_1 _2556_ (.B1(_0641_),
    .Y(_0642_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0639_));
 sg13g2_mux4_1 _2557_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(net1599),
    .A1(net1613),
    .A2(net1606),
    .A3(net1626),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0643_));
 sg13g2_o21ai_1 _2558_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ),
    .Y(_0644_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0643_));
 sg13g2_nand2b_1 _2559_ (.Y(_0645_),
    .B(_0642_),
    .A_N(_0644_));
 sg13g2_nand2b_2 _2560_ (.Y(_0646_),
    .B(_0645_),
    .A_N(_0637_));
 sg13g2_mux4_1 _2561_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ),
    .A0(net143),
    .A1(net65),
    .A2(net20),
    .A3(_0646_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_0647_));
 sg13g2_mux4_1 _2562_ (.S0(net1682),
    .A0(net1596),
    .A1(net1602),
    .A2(net1621),
    .A3(net1630),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0648_));
 sg13g2_inv_4 _2563_ (.A(_0648_),
    .Y(_0649_));
 sg13g2_mux4_1 _2564_ (.S0(net1682),
    .A0(net1592),
    .A1(net1583),
    .A2(net1521),
    .A3(net699),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0650_));
 sg13g2_o21ai_1 _2565_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .Y(_0651_),
    .A1(_0649_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_a21oi_2 _2566_ (.B1(_0651_),
    .Y(_0652_),
    .A2(_0650_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_a21oi_1 _2567_ (.A1(net125),
    .A2(net1682),
    .Y(_0653_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_o21ai_1 _2568_ (.B1(_0653_),
    .Y(_0654_),
    .A1(net1682),
    .A2(net687));
 sg13g2_nor2b_1 _2569_ (.A(net1682),
    .B_N(net137),
    .Y(_0655_));
 sg13g2_a21oi_1 _2570_ (.A1(net6),
    .A2(net1682),
    .Y(_0656_),
    .B1(_0655_));
 sg13g2_a21oi_1 _2571_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .A2(_0656_),
    .Y(_0657_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_a21oi_1 _2572_ (.A1(net32),
    .A2(net1682),
    .Y(_0658_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_o21ai_1 _2573_ (.B1(_0658_),
    .Y(_0659_),
    .A1(_0059_),
    .A2(net1682));
 sg13g2_nand2b_1 _2574_ (.Y(_0660_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .A_N(net86));
 sg13g2_o21ai_1 _2575_ (.B1(_0660_),
    .Y(_0661_),
    .A1(net67),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_a21oi_1 _2576_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ),
    .A2(_0661_),
    .Y(_0662_),
    .B1(_0094_));
 sg13g2_a221oi_1 _2577_ (.B2(_0662_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ),
    .B1(_0659_),
    .A1(_0654_),
    .Y(_0663_),
    .A2(_0657_));
 sg13g2_nor2_2 _2578_ (.A(_0663_),
    .B(_0652_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ));
 sg13g2_mux4_1 _2579_ (.S0(net1659),
    .A0(net1528),
    .A1(net1534),
    .A2(net1543),
    .A3(net1558),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0664_));
 sg13g2_nand2_2 _2580_ (.Y(_0665_),
    .A(_0664_),
    .B(_0089_));
 sg13g2_nor2_1 _2581_ (.A(net1658),
    .B(net1564),
    .Y(_0666_));
 sg13g2_a21oi_1 _2582_ (.A1(net1658),
    .A2(net1569),
    .Y(_0667_),
    .B1(_0666_));
 sg13g2_nand2b_1 _2583_ (.Y(_0668_),
    .B(net1658),
    .A_N(net1617));
 sg13g2_o21ai_1 _2584_ (.B1(_0668_),
    .Y(_0669_),
    .A1(net1658),
    .A2(net1578));
 sg13g2_a21oi_1 _2585_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0669_),
    .Y(_0670_),
    .B1(_0089_));
 sg13g2_o21ai_1 _2586_ (.B1(_0670_),
    .Y(_0671_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0667_));
 sg13g2_nand3_1 _2587_ (.B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .C(_0671_),
    .A(_0665_),
    .Y(_0672_));
 sg13g2_nor2_1 _2588_ (.A(net1924),
    .B(net1659),
    .Y(_0673_));
 sg13g2_a21oi_1 _2589_ (.A1(_0066_),
    .A2(net1658),
    .Y(_0674_),
    .B1(_0673_));
 sg13g2_nor2_1 _2590_ (.A(net155),
    .B(net1658),
    .Y(_0675_));
 sg13g2_a21oi_1 _2591_ (.A1(_0058_),
    .A2(net1658),
    .Y(_0676_),
    .B1(_0675_));
 sg13g2_mux2_1 _2592_ (.A0(net1926),
    .A1(net95),
    .S(net1659),
    .X(_0677_));
 sg13g2_mux2_1 _2593_ (.A0(net119),
    .A1(net131),
    .S(net1658),
    .X(_0678_));
 sg13g2_mux4_1 _2594_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ),
    .A0(_0674_),
    .A1(_0676_),
    .A2(_0678_),
    .A3(_0677_),
    .S1(_0089_),
    .X(_0679_));
 sg13g2_o21ai_1 _2595_ (.B1(_0672_),
    .Y(_0680_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ),
    .A2(_0679_));
 sg13g2_inv_16 _2596_ (.A(net633),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ));
 sg13g2_mux4_1 _2597_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net15),
    .A2(net41),
    .A3(net76),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_0681_));
 sg13g2_mux4_1 _2598_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ),
    .A0(net1584),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .A2(net1576),
    .A3(_0647_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ),
    .X(_0682_));
 sg13g2_a21oi_1 _2599_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0095_),
    .Y(_0683_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_o21ai_1 _2600_ (.B1(_0683_),
    .Y(_0684_),
    .A1(_0682_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_mux2_1 _2601_ (.A0(net147),
    .A1(net1705),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0685_));
 sg13g2_a21oi_1 _2602_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_0685_),
    .Y(_0686_),
    .B1(_0096_));
 sg13g2_mux4_1 _2603_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A0(net1711),
    .A1(net1926),
    .A2(net121),
    .A3(net97),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0687_));
 sg13g2_o21ai_1 _2604_ (.B1(_0097_),
    .Y(_0688_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0687_));
 sg13g2_a21oi_2 _2605_ (.B1(_0688_),
    .Y(_0689_),
    .A2(_0684_),
    .A1(_0686_));
 sg13g2_mux2_1 _2606_ (.A0(net1555),
    .A1(net1571),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0690_));
 sg13g2_mux2_1 _2607_ (.A0(net1581),
    .A1(net1619),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_0691_));
 sg13g2_o21ai_1 _2608_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0692_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_0690_));
 sg13g2_a21o_1 _2609_ (.A2(_0691_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .B1(_0692_),
    .X(_0693_));
 sg13g2_mux4_1 _2610_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(net1531),
    .A1(net1537),
    .A2(net1545),
    .A3(net1552),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0694_));
 sg13g2_nor2_2 _2611_ (.A(_0694_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0695_));
 sg13g2_nor2_2 _2612_ (.A(_0695_),
    .B(_0097_),
    .Y(_0696_));
 sg13g2_a21oi_2 _2613_ (.B1(_0689_),
    .Y(_0697_),
    .A2(_0696_),
    .A1(_0693_));
 sg13g2_inv_8 _2614_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .A(_0697_));
 sg13g2_mux4_1 _2615_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .A0(_0697_),
    .A1(_0099_),
    .A2(_0098_),
    .A3(_0100_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(_0698_));
 sg13g2_mux4_1 _2616_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .A1(net43),
    .A2(net17),
    .A3(net78),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ),
    .X(_0699_));
 sg13g2_mux2_1 _2617_ (.A0(_0630_),
    .A1(_0698_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .X(_0700_));
 sg13g2_o21ai_1 _2618_ (.B1(_0527_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0700_));
 sg13g2_nand2b_1 _2619_ (.Y(_0701_),
    .B(net1642),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ));
 sg13g2_mux2_2 _2620_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ),
    .S(net1642),
    .X(_0702_));
 sg13g2_o21ai_1 _2621_ (.B1(_0701_),
    .Y(_0703_),
    .A1(net1642),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ));
 sg13g2_mux4_1 _2622_ (.S0(net1675),
    .A0(net1598),
    .A1(net1603),
    .A2(net1623),
    .A3(net1633),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0704_));
 sg13g2_nand2b_1 _2623_ (.Y(_0705_),
    .B(_0704_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_mux2_1 _2624_ (.A0(net690),
    .A1(net1587),
    .S(net1674),
    .X(_0706_));
 sg13g2_nand2b_1 _2625_ (.Y(_0707_),
    .B(net1675),
    .A_N(net1520));
 sg13g2_o21ai_1 _2626_ (.B1(_0707_),
    .Y(_0708_),
    .A1(net1675),
    .A2(net1522));
 sg13g2_o21ai_1 _2627_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0709_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0706_));
 sg13g2_a21oi_1 _2628_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0708_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_nor2_1 _2629_ (.A(_0101_),
    .B(_0710_),
    .Y(_0711_));
 sg13g2_nand2b_1 _2630_ (.Y(_0712_),
    .B(net1674),
    .A_N(net32));
 sg13g2_o21ai_1 _2631_ (.B1(_0712_),
    .Y(_0713_),
    .A1(net20),
    .A2(net1674));
 sg13g2_nand2b_1 _2632_ (.Y(_0714_),
    .B(net1674),
    .A_N(net81));
 sg13g2_o21ai_1 _2633_ (.B1(_0714_),
    .Y(_0715_),
    .A1(net67),
    .A2(net1674));
 sg13g2_nand2b_1 _2634_ (.Y(_0716_),
    .B(net1674),
    .A_N(net6));
 sg13g2_o21ai_1 _2635_ (.B1(_0716_),
    .Y(_0717_),
    .A1(net1),
    .A2(net1674));
 sg13g2_nand2b_1 _2636_ (.Y(_0718_),
    .B(net1675),
    .A_N(net137));
 sg13g2_o21ai_1 _2637_ (.B1(_0718_),
    .Y(_0719_),
    .A1(net125),
    .A2(net1674));
 sg13g2_mux4_1 _2638_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ),
    .A0(_0719_),
    .A1(_0717_),
    .A2(_0713_),
    .A3(_0715_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ),
    .X(_0720_));
 sg13g2_a22oi_1 _2639_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .B1(_0720_),
    .B2(_0101_),
    .A2(_0711_),
    .A1(_0705_));
 sg13g2_mux4_1 _2640_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ),
    .A0(net146),
    .A1(net83),
    .A2(net49),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ),
    .X(_0721_));
 sg13g2_inv_2 _2641_ (.Y(_0722_),
    .A(_0721_));
 sg13g2_mux4_1 _2642_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .A0(net1521),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .A2(_0699_),
    .A3(_0721_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .X(_0723_));
 sg13g2_mux4_1 _2643_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ),
    .A0(_0175_),
    .A1(_0384_),
    .A2(_0698_),
    .A3(_0722_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ),
    .X(_0724_));
 sg13g2_mux4_1 _2644_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(net645),
    .A1(_0724_),
    .A2(_0099_),
    .A3(_0105_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0725_));
 sg13g2_mux4_1 _2645_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(net1712),
    .A1(net120),
    .A2(net88),
    .A3(net96),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0726_));
 sg13g2_nor2_1 _2646_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .B(_0726_),
    .Y(_0727_));
 sg13g2_nor2_1 _2647_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .B(_0727_),
    .Y(_0728_));
 sg13g2_inv_1 _2648_ (.Y(_0729_),
    .A(_0728_));
 sg13g2_a21oi_2 _2649_ (.B1(_0729_),
    .Y(_0730_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .A1(_0725_));
 sg13g2_mux2_1 _2650_ (.A0(net1562),
    .A1(net1571),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0731_));
 sg13g2_mux2_1 _2651_ (.A0(net1582),
    .A1(net1619),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0732_));
 sg13g2_o21ai_1 _2652_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0733_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0731_));
 sg13g2_a21o_1 _2653_ (.A2(_0732_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .B1(_0733_),
    .X(_0734_));
 sg13g2_nand2_1 _2654_ (.Y(_0735_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .B(_0180_));
 sg13g2_o21ai_1 _2655_ (.B1(_0735_),
    .Y(_0736_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(net1531));
 sg13g2_mux2_1 _2656_ (.A0(net1545),
    .A1(net1552),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ),
    .X(_0737_));
 sg13g2_a21oi_1 _2657_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0737_),
    .Y(_0738_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_o21ai_1 _2658_ (.B1(_0738_),
    .Y(_0739_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ),
    .A2(_0736_));
 sg13g2_and3_1 _2659_ (.X(_0740_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ),
    .B(_0734_),
    .C(_0739_));
 sg13g2_or2_1 _2660_ (.X(_0741_),
    .B(_0740_),
    .A(_0730_));
 sg13g2_nor3_1 _2661_ (.A(_0124_),
    .B(_0730_),
    .C(_0740_),
    .Y(_0742_));
 sg13g2_o21ai_1 _2662_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ),
    .Y(_0743_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .A2(net159));
 sg13g2_mux4_1 _2663_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net1609),
    .A1(net1602),
    .A2(net1621),
    .A3(net1629),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0744_));
 sg13g2_nand2b_1 _2664_ (.Y(_0745_),
    .B(_0744_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_mux4_1 _2665_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net1592),
    .A1(net1583),
    .A2(net1521),
    .A3(net699),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0746_));
 sg13g2_a21oi_2 _2666_ (.B1(_0103_),
    .Y(_0747_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .A1(_0746_));
 sg13g2_mux4_1 _2667_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net144),
    .A1(net2002),
    .A2(net5),
    .A3(net21),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0748_));
 sg13g2_nand2b_1 _2668_ (.Y(_0749_),
    .B(_0748_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_mux4_1 _2669_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net31),
    .A1(net47),
    .A2(net66),
    .A3(net82),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_0750_));
 sg13g2_a21oi_1 _2670_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0750_),
    .Y(_0751_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_a22oi_1 _2671_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .B1(_0749_),
    .B2(_0751_),
    .A2(_0747_),
    .A1(_0745_));
 sg13g2_nand2_1 _2672_ (.Y(_0752_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ));
 sg13g2_o21ai_1 _2673_ (.B1(_0752_),
    .Y(_0753_),
    .A1(_0069_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_a21oi_1 _2674_ (.A1(_0125_),
    .A2(_0753_),
    .Y(_0754_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_o21ai_1 _2675_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0742_),
    .A2(_0743_));
 sg13g2_a21oi_1 _2676_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0290_),
    .Y(_0756_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_o21ai_1 _2677_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .Y(_0757_),
    .A1(net167),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_a21oi_1 _2678_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .A2(_0580_),
    .Y(_0758_),
    .B1(_0757_));
 sg13g2_nor2b_1 _2679_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .B_N(net131),
    .Y(_0759_));
 sg13g2_a21oi_1 _2680_ (.A1(net58),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ),
    .Y(_0760_),
    .B1(_0759_));
 sg13g2_o21ai_1 _2681_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .Y(_0761_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_0760_));
 sg13g2_nor2_1 _2682_ (.A(_0758_),
    .B(_0761_),
    .Y(_0762_));
 sg13g2_mux4_1 _2683_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ),
    .A0(net115),
    .A1(net38),
    .A2(net108),
    .A3(net151),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0763_));
 sg13g2_o21ai_1 _2684_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_0764_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0763_));
 sg13g2_nor2_1 _2685_ (.A(_0762_),
    .B(_0764_),
    .Y(_0765_));
 sg13g2_a21oi_2 _2686_ (.B1(_0765_),
    .Y(_0766_),
    .A2(_0756_),
    .A1(_0755_));
 sg13g2_inv_1 _2687_ (.Y(\Tile_X0Y1_DSP_bot.B3 ),
    .A(_0766_));
 sg13g2_nor2_1 _2688_ (.A(net1640),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ),
    .Y(_0767_));
 sg13g2_a21o_1 _2689_ (.A2(_0766_),
    .A1(net1640),
    .B1(_0767_),
    .X(_0768_));
 sg13g2_nor2_2 _2690_ (.A(_0703_),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_nor2_1 _2691_ (.A(_0462_),
    .B(_0703_),
    .Y(_0770_));
 sg13g2_nor2_1 _2692_ (.A(net1515),
    .B(net1608),
    .Y(_0771_));
 sg13g2_nand2_1 _2693_ (.Y(_0772_),
    .A(_0519_),
    .B(_0769_));
 sg13g2_o21ai_1 _2694_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0773_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(net642));
 sg13g2_a21oi_2 _2695_ (.B1(_0773_),
    .Y(_0774_),
    .A2(net712),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_nor2b_1 _2696_ (.A(net99),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .Y(_0775_));
 sg13g2_nor2_1 _2697_ (.A(net1709),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ),
    .Y(_0776_));
 sg13g2_nor3_1 _2698_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_0775_),
    .C(_0776_),
    .Y(_0777_));
 sg13g2_nor3_2 _2699_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .B(_0777_),
    .C(_0774_),
    .Y(_0778_));
 sg13g2_nand2_1 _2700_ (.Y(_0779_),
    .A(net160),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_o21ai_1 _2701_ (.B1(_0779_),
    .Y(_0780_),
    .A1(net696),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_nand2b_1 _2702_ (.Y(_0781_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ),
    .A_N(net100));
 sg13g2_o21ai_1 _2703_ (.B1(_0781_),
    .Y(_0782_),
    .A1(net124),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_o21ai_1 _2704_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .Y(_0783_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0782_));
 sg13g2_a21oi_1 _2705_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0780_),
    .Y(_0784_),
    .B1(_0783_));
 sg13g2_or3_1 _2706_ (.A(_0778_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .C(_0784_),
    .X(_0785_));
 sg13g2_mux4_1 _2707_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(net1528),
    .A1(net1542),
    .A2(net1549),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0786_));
 sg13g2_mux2_1 _2708_ (.A0(net1561),
    .A1(net1569),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0787_));
 sg13g2_mux2_1 _2709_ (.A0(net1577),
    .A1(net1615),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0788_));
 sg13g2_o21ai_1 _2710_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0789_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0787_));
 sg13g2_a21oi_2 _2711_ (.B1(_0789_),
    .Y(_0790_),
    .A2(_0788_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_nor2b_1 _2712_ (.A(_0790_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0791_));
 sg13g2_o21ai_1 _2713_ (.B1(_0791_),
    .Y(_0792_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0786_));
 sg13g2_mux4_1 _2714_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(net1713),
    .A1(net117),
    .A2(net93),
    .A3(net1923),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0793_));
 sg13g2_mux2_1 _2715_ (.A0(net153),
    .A1(net167),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0794_));
 sg13g2_nor2b_1 _2716_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .B_N(net1935),
    .Y(_0795_));
 sg13g2_a21oi_1 _2717_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(net52),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_o21ai_1 _2718_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0797_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0796_));
 sg13g2_a21o_1 _2719_ (.A2(_0794_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ),
    .B1(_0797_),
    .X(_0798_));
 sg13g2_o21ai_1 _2720_ (.B1(_0798_),
    .Y(_0799_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0793_));
 sg13g2_o21ai_1 _2721_ (.B1(_0792_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0799_));
 sg13g2_mux2_1 _2722_ (.A0(net50),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0800_));
 sg13g2_nor2b_1 _2723_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .B_N(net131),
    .Y(_0801_));
 sg13g2_a21oi_1 _2724_ (.A1(net1924),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_o21ai_1 _2725_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .Y(_0803_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0802_));
 sg13g2_a21oi_1 _2726_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_0800_),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_mux4_1 _2727_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ),
    .A0(net115),
    .A1(net38),
    .A2(net91),
    .A3(net172),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0805_));
 sg13g2_o21ai_1 _2728_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ),
    .Y(_0806_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0805_));
 sg13g2_o21ai_1 _2729_ (.B1(_0785_),
    .Y(\Tile_X0Y1_DSP_bot.A3 ),
    .A1(_0804_),
    .A2(_0806_));
 sg13g2_mux2_2 _2730_ (.A0(\Tile_X0Y1_DSP_bot.A3 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ),
    .S(net1641),
    .X(_0807_));
 sg13g2_inv_8 _2731_ (.Y(_0808_),
    .A(_0807_));
 sg13g2_mux4_1 _2732_ (.S0(net1697),
    .A0(net1596),
    .A1(net1609),
    .A2(net1621),
    .A3(net1629),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0809_));
 sg13g2_nand2b_1 _2733_ (.Y(_0810_),
    .B(net1697),
    .A_N(net1583));
 sg13g2_o21ai_1 _2734_ (.B1(_0810_),
    .Y(_0811_),
    .A1(net1697),
    .A2(net1592));
 sg13g2_nand2_1 _2735_ (.Y(_0812_),
    .A(net1698),
    .B(net1518));
 sg13g2_o21ai_1 _2736_ (.B1(_0812_),
    .Y(_0813_),
    .A1(net1698),
    .A2(_0175_));
 sg13g2_o21ai_1 _2737_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0814_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0811_));
 sg13g2_a21oi_1 _2738_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0813_),
    .Y(_0815_),
    .B1(_0814_));
 sg13g2_o21ai_1 _2739_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0816_),
    .A1(_0809_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_a21oi_1 _2740_ (.A1(_0074_),
    .A2(net1697),
    .Y(_0817_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_o21ai_1 _2741_ (.B1(_0817_),
    .Y(_0818_),
    .A1(net1697),
    .A2(net1527));
 sg13g2_o21ai_1 _2742_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Y(_0819_),
    .A1(net7),
    .A2(net1697));
 sg13g2_a21oi_1 _2743_ (.A1(_0075_),
    .A2(net1697),
    .Y(_0820_),
    .B1(_0819_));
 sg13g2_nor2_1 _2744_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_nand2_1 _2745_ (.Y(_0822_),
    .A(_0818_),
    .B(_0821_));
 sg13g2_nand2b_1 _2746_ (.Y(_0823_),
    .B(net1698),
    .A_N(net49));
 sg13g2_o21ai_1 _2747_ (.B1(_0823_),
    .Y(_0824_),
    .A1(net33),
    .A2(net1698));
 sg13g2_o21ai_1 _2748_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .Y(_0825_),
    .A1(net68),
    .A2(net1697));
 sg13g2_a21oi_1 _2749_ (.A1(_0076_),
    .A2(net1698),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_nor2b_1 _2750_ (.A(_0826_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ),
    .Y(_0827_));
 sg13g2_o21ai_1 _2751_ (.B1(_0827_),
    .Y(_0828_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0824_));
 sg13g2_nand3b_1 _2752_ (.B(_0822_),
    .C(_0828_),
    .Y(_0829_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_o21ai_1 _2753_ (.B1(_0829_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .A1(_0816_),
    .A2(_0815_));
 sg13g2_mux2_1 _2754_ (.A0(net1929),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0830_));
 sg13g2_nor2b_1 _2755_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .B_N(net135),
    .Y(_0831_));
 sg13g2_a21oi_1 _2756_ (.A1(net54),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ),
    .Y(_0832_),
    .B1(_0831_));
 sg13g2_o21ai_1 _2757_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .Y(_0833_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_0832_));
 sg13g2_a21oi_2 _2758_ (.B1(_0833_),
    .Y(_0834_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ),
    .A1(_0830_));
 sg13g2_mux4_1 _2759_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ),
    .A0(net123),
    .A1(net30),
    .A2(net23),
    .A3(net65),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0835_));
 sg13g2_o21ai_1 _2760_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_0836_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0835_));
 sg13g2_nor2_2 _2761_ (.A(_0836_),
    .B(_0834_),
    .Y(_0837_));
 sg13g2_or2_1 _2762_ (.X(_0838_),
    .B(_0646_),
    .A(_0115_));
 sg13g2_nor2_1 _2763_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .B(net73),
    .Y(_0839_));
 sg13g2_nor2b_1 _2764_ (.A(_0839_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ),
    .Y(_0840_));
 sg13g2_a21oi_1 _2765_ (.A1(_0077_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .Y(_0841_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_o21ai_1 _2766_ (.B1(_0841_),
    .Y(_0842_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ));
 sg13g2_nand2b_1 _2767_ (.Y(_0843_),
    .B(_0842_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_a21o_1 _2768_ (.A2(_0840_),
    .A1(_0838_),
    .B1(_0843_),
    .X(_0844_));
 sg13g2_a21oi_1 _2769_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0412_),
    .Y(_0845_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_a21oi_2 _2770_ (.B1(_0837_),
    .Y(_0846_),
    .A2(_0845_),
    .A1(_0844_));
 sg13g2_inv_1 _2771_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .A(_0846_));
 sg13g2_nor2_2 _2772_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_a21oi_2 _2773_ (.B1(_0847_),
    .Y(_0848_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ));
 sg13g2_inv_8 _2774_ (.Y(_0849_),
    .A(_0848_));
 sg13g2_nand2_2 _2775_ (.Y(_0850_),
    .A(_0807_),
    .B(_0849_));
 sg13g2_mux4_1 _2776_ (.S0(net1690),
    .A0(net1599),
    .A1(net1612),
    .A2(net1605),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0851_));
 sg13g2_inv_1 _2777_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_mux4_1 _2778_ (.S0(net1690),
    .A0(net1594),
    .A1(net1588),
    .A2(net1523),
    .A3(net1541),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0853_));
 sg13g2_o21ai_1 _2779_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .Y(_0854_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0852_));
 sg13g2_a21oi_1 _2780_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0853_),
    .Y(_0855_),
    .B1(_0854_));
 sg13g2_nand2b_1 _2781_ (.Y(_0856_),
    .B(net1527),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_a21oi_1 _2782_ (.A1(net128),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .Y(_0857_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_nor2b_1 _2783_ (.A(net1690),
    .B_N(net2004),
    .Y(_0858_));
 sg13g2_a21oi_1 _2784_ (.A1(net9),
    .A2(net1690),
    .Y(_0859_),
    .B1(_0858_));
 sg13g2_a221oi_1 _2785_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ),
    .B1(_0859_),
    .A1(_0856_),
    .Y(_0860_),
    .A2(_0857_));
 sg13g2_nand2b_1 _2786_ (.Y(_0861_),
    .B(net27),
    .A_N(net1690));
 sg13g2_a21oi_1 _2787_ (.A1(net35),
    .A2(net1690),
    .Y(_0862_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_nand2b_1 _2788_ (.Y(_0863_),
    .B(net1690),
    .A_N(net1930));
 sg13g2_o21ai_1 _2789_ (.B1(_0863_),
    .Y(_0864_),
    .A1(net1933),
    .A2(net1690));
 sg13g2_a221oi_1 _2790_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ),
    .C1(_0114_),
    .B1(_0864_),
    .A1(_0861_),
    .Y(_0865_),
    .A2(_0862_));
 sg13g2_nor3_1 _2791_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ),
    .B(_0860_),
    .C(_0865_),
    .Y(_0866_));
 sg13g2_nor2_2 _2792_ (.A(_0866_),
    .B(_0855_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ));
 sg13g2_inv_1 _2793_ (.Y(_0867_),
    .A(net615));
 sg13g2_mux4_1 _2794_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(_0627_),
    .A1(_0110_),
    .A2(_0066_),
    .A3(_0867_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_0868_));
 sg13g2_mux4_1 _2795_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .A1(net43),
    .A2(net17),
    .A3(net78),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ),
    .X(_0869_));
 sg13g2_inv_1 _2796_ (.Y(_0870_),
    .A(_0869_));
 sg13g2_nand2b_1 _2797_ (.Y(_0871_),
    .B(net1688),
    .A_N(net1629));
 sg13g2_o21ai_1 _2798_ (.B1(_0871_),
    .Y(_0872_),
    .A1(net1688),
    .A2(net1621));
 sg13g2_mux2_1 _2799_ (.A0(net1596),
    .A1(net1609),
    .S(net1688),
    .X(_0873_));
 sg13g2_a21oi_1 _2800_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_0872_),
    .Y(_0874_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_o21ai_1 _2801_ (.B1(_0874_),
    .Y(_0875_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_0873_));
 sg13g2_nand2_1 _2802_ (.Y(_0876_),
    .A(net1688),
    .B(net1583));
 sg13g2_o21ai_1 _2803_ (.B1(_0876_),
    .Y(_0877_),
    .A1(net1688),
    .A2(net1590));
 sg13g2_o21ai_1 _2804_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .Y(_0878_),
    .A1(net1688),
    .A2(_0175_));
 sg13g2_a21oi_1 _2805_ (.A1(net1688),
    .A2(net699),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_o21ai_1 _2806_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_0880_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_0877_));
 sg13g2_nor2_1 _2807_ (.A(_0879_),
    .B(_0880_),
    .Y(_0881_));
 sg13g2_nor2b_1 _2808_ (.A(_0881_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_0882_));
 sg13g2_mux4_1 _2809_ (.S0(net1688),
    .A0(net146),
    .A1(net2004),
    .A2(net7),
    .A3(net21),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0883_));
 sg13g2_nand2b_1 _2810_ (.Y(_0884_),
    .B(_0883_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_nand2_1 _2811_ (.Y(_0885_),
    .A(_0076_),
    .B(net1689));
 sg13g2_o21ai_1 _2812_ (.B1(_0885_),
    .Y(_0886_),
    .A1(net68),
    .A2(net1689));
 sg13g2_mux2_1 _2813_ (.A0(net33),
    .A1(net49),
    .S(net1689),
    .X(_0887_));
 sg13g2_o21ai_1 _2814_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_0888_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_0887_));
 sg13g2_a21oi_1 _2815_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_0886_),
    .Y(_0889_),
    .B1(_0888_));
 sg13g2_nor2_1 _2816_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ),
    .B(_0889_),
    .Y(_0890_));
 sg13g2_a22oi_1 _2817_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .B1(_0884_),
    .B2(_0890_),
    .A2(_0875_),
    .A1(_0882_));
 sg13g2_o21ai_1 _2818_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .Y(_0891_),
    .A1(_0087_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_a21o_1 _2819_ (.A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .B1(_0891_),
    .X(_0892_));
 sg13g2_mux2_1 _2820_ (.A0(net144),
    .A1(net23),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0893_));
 sg13g2_o21ai_1 _2821_ (.B1(_0892_),
    .Y(_0894_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_0893_));
 sg13g2_mux4_1 _2822_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(net127),
    .A1(net8),
    .A2(net56),
    .A3(net69),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0895_));
 sg13g2_inv_1 _2823_ (.Y(_0896_),
    .A(_0895_));
 sg13g2_mux4_1 _2824_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ),
    .A0(_0868_),
    .A1(_0870_),
    .A2(_0896_),
    .A3(_0894_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_0897_));
 sg13g2_inv_1 _2825_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ),
    .A(_0897_));
 sg13g2_nor2_1 _2826_ (.A(net1640),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ),
    .Y(_0898_));
 sg13g2_a21oi_2 _2827_ (.B1(_0898_),
    .Y(_0899_),
    .A2(_0123_),
    .A1(_0897_));
 sg13g2_mux2_1 _2828_ (.A0(net1708),
    .A1(net103),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0900_));
 sg13g2_nand2_1 _2829_ (.Y(_0901_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ));
 sg13g2_nand2b_1 _2830_ (.Y(_0902_),
    .B(net163),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_nand3_1 _2831_ (.B(_0901_),
    .C(_0902_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .Y(_0903_));
 sg13g2_o21ai_1 _2832_ (.B1(_0903_),
    .Y(_0904_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ),
    .A2(_0900_));
 sg13g2_inv_1 _2833_ (.Y(_0905_),
    .A(_0904_));
 sg13g2_mux4_1 _2834_ (.S0(net1667),
    .A0(net1528),
    .A1(net1542),
    .A2(net1549),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0906_));
 sg13g2_or2_1 _2835_ (.X(_0907_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .A(_0906_));
 sg13g2_a21oi_1 _2836_ (.A1(net1667),
    .A2(net1569),
    .Y(_0908_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_o21ai_1 _2837_ (.B1(_0908_),
    .Y(_0909_),
    .A1(net1667),
    .A2(net1563));
 sg13g2_mux2_1 _2838_ (.A0(net1577),
    .A1(net1617),
    .S(net1667),
    .X(_0910_));
 sg13g2_nand2_1 _2839_ (.Y(_0911_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .B(_0910_));
 sg13g2_nand3_1 _2840_ (.B(_0909_),
    .C(_0911_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0912_));
 sg13g2_nand3_1 _2841_ (.B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .C(_0912_),
    .A(_0907_),
    .Y(_0913_));
 sg13g2_mux2_1 _2842_ (.A0(net109),
    .A1(net1923),
    .S(net1667),
    .X(_0914_));
 sg13g2_nor2b_1 _2843_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .B_N(net141),
    .Y(_0915_));
 sg13g2_a21oi_1 _2844_ (.A1(net1928),
    .A2(net1667),
    .Y(_0916_),
    .B1(_0915_));
 sg13g2_a21oi_1 _2845_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0914_),
    .Y(_0917_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_o21ai_1 _2846_ (.B1(_0917_),
    .Y(_0918_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0916_));
 sg13g2_o21ai_1 _2847_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .Y(_0919_),
    .A1(net153),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_a21oi_1 _2848_ (.A1(_0058_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .Y(_0920_),
    .B1(_0919_));
 sg13g2_nor2b_1 _2849_ (.A(net1667),
    .B_N(net52),
    .Y(_0921_));
 sg13g2_a21oi_1 _2850_ (.A1(net1667),
    .A2(net60),
    .Y(_0922_),
    .B1(_0921_));
 sg13g2_o21ai_1 _2851_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ),
    .Y(_0923_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0922_));
 sg13g2_o21ai_1 _2852_ (.B1(_0918_),
    .Y(_0924_),
    .A1(_0920_),
    .A2(_0923_));
 sg13g2_o21ai_1 _2853_ (.B1(_0913_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_0924_));
 sg13g2_mux4_1 _2854_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ),
    .A0(net132),
    .A1(net1703),
    .A2(net1921),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_0925_));
 sg13g2_mux4_1 _2855_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(net119),
    .A1(net42),
    .A2(net107),
    .A3(net155),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0926_));
 sg13g2_mux4_1 _2856_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ),
    .A0(_0905_),
    .A1(_0926_),
    .A2(_0596_),
    .A3(_0925_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ),
    .X(\Tile_X0Y1_DSP_bot.A2 ));
 sg13g2_nand2b_1 _2857_ (.Y(_0927_),
    .B(net1641),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ));
 sg13g2_o21ai_1 _2858_ (.B1(_0927_),
    .Y(_0928_),
    .A1(\Tile_X0Y1_DSP_bot.A2 ),
    .A2(net1641));
 sg13g2_inv_4 _2859_ (.A(_0928_),
    .Y(_0929_));
 sg13g2_nand2_1 _2860_ (.Y(_0930_),
    .A(_0899_),
    .B(net714));
 sg13g2_nand2_1 _2861_ (.Y(_0931_),
    .A(_0807_),
    .B(_0899_));
 sg13g2_nand2_1 _2862_ (.Y(_0932_),
    .A(_0849_),
    .B(net714));
 sg13g2_nor2_1 _2863_ (.A(_0850_),
    .B(_0930_),
    .Y(_0933_));
 sg13g2_mux4_1 _2864_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ),
    .A0(net125),
    .A1(net32),
    .A2(net6),
    .A3(net85),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0934_));
 sg13g2_nor2b_1 _2865_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .B_N(_0934_),
    .Y(_0935_));
 sg13g2_a21oi_1 _2866_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0385_),
    .Y(_0936_),
    .B1(_0935_));
 sg13g2_mux4_1 _2867_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net1599),
    .A1(net1612),
    .A2(net1605),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0937_));
 sg13g2_inv_1 _2868_ (.Y(_0938_),
    .A(_0937_));
 sg13g2_mux4_1 _2869_ (.S0(net1686),
    .A0(net1593),
    .A1(net1588),
    .A2(net1524),
    .A3(net1519),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0939_));
 sg13g2_o21ai_1 _2870_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .Y(_0940_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0938_));
 sg13g2_a21oi_1 _2871_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0939_),
    .Y(_0941_),
    .B1(_0940_));
 sg13g2_nand2_1 _2872_ (.Y(_0942_),
    .A(_0083_),
    .B(net1686));
 sg13g2_o21ai_1 _2873_ (.B1(_0942_),
    .Y(_0943_),
    .A1(_0376_),
    .A2(net1686));
 sg13g2_nand2b_1 _2874_ (.Y(_0944_),
    .B(net2004),
    .A_N(net1686));
 sg13g2_a21oi_1 _2875_ (.A1(net9),
    .A2(net1686),
    .Y(_0945_),
    .B1(_0113_));
 sg13g2_a221oi_1 _2876_ (.B2(_0945_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .B1(_0944_),
    .A1(_0113_),
    .Y(_0946_),
    .A2(_0943_));
 sg13g2_a21oi_1 _2877_ (.A1(net29),
    .A2(net1686),
    .Y(_0947_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_o21ai_1 _2878_ (.B1(_0947_),
    .Y(_0948_),
    .A1(_0091_),
    .A2(net1686));
 sg13g2_mux2_1 _2879_ (.A0(net35),
    .A1(net1933),
    .S(net1686),
    .X(_0949_));
 sg13g2_o21ai_1 _2880_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_0950_),
    .A1(_0113_),
    .A2(_0949_));
 sg13g2_nor2b_1 _2881_ (.A(_0950_),
    .B_N(_0948_),
    .Y(_0951_));
 sg13g2_nor3_2 _2882_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ),
    .B(_0946_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_nor2_2 _2883_ (.A(_0952_),
    .B(_0941_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ));
 sg13g2_mux4_1 _2884_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(net1565),
    .A1(net1572),
    .A2(net1579),
    .A3(net1616),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0953_));
 sg13g2_mux4_1 _2885_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(net1529),
    .A1(net1535),
    .A2(net1550),
    .A3(net1559),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0954_));
 sg13g2_nand2b_1 _2886_ (.Y(_0955_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .A_N(_0953_));
 sg13g2_o21ai_1 _2887_ (.B1(_0955_),
    .Y(_0956_),
    .A1(_0954_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_mux4_1 _2888_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(net118),
    .A1(net134),
    .A2(net1927),
    .A3(net94),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0957_));
 sg13g2_nor2b_1 _2889_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .B_N(_0957_),
    .Y(_0958_));
 sg13g2_nor2_1 _2890_ (.A(net1922),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .Y(_0959_));
 sg13g2_a21oi_1 _2891_ (.A1(_0068_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .Y(_0960_),
    .B1(_0959_));
 sg13g2_nand2b_1 _2892_ (.Y(_0961_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ),
    .A_N(net170));
 sg13g2_o21ai_1 _2893_ (.B1(_0961_),
    .Y(_0962_),
    .A1(net154),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_o21ai_1 _2894_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0963_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0960_));
 sg13g2_a21oi_1 _2895_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0962_),
    .Y(_0964_),
    .B1(_0963_));
 sg13g2_nor3_1 _2896_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .B(_0958_),
    .C(_0964_),
    .Y(_0965_));
 sg13g2_a21o_2 _2897_ (.A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ),
    .A1(_0956_),
    .B1(_0965_),
    .X(_0966_));
 sg13g2_inv_4 _2898_ (.A(_0966_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ));
 sg13g2_mux4_1 _2899_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net75),
    .A2(net14),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_0967_));
 sg13g2_nor2b_1 _2900_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ),
    .B_N(_0967_),
    .Y(_0968_));
 sg13g2_mux4_1 _2901_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net15),
    .A2(net41),
    .A3(net76),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0969_));
 sg13g2_a21oi_2 _2902_ (.B1(_0968_),
    .Y(_0970_),
    .A2(_0969_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_mux2_1 _2903_ (.A0(_0970_),
    .A1(_0936_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ),
    .X(_0971_));
 sg13g2_inv_1 _2904_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .A(_0971_));
 sg13g2_nand2_1 _2905_ (.Y(_0972_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ));
 sg13g2_o21ai_1 _2906_ (.B1(_0972_),
    .Y(_0973_),
    .A1(_0971_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ));
 sg13g2_mux4_1 _2907_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(net1707),
    .A1(net10),
    .A2(net57),
    .A3(net71),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0974_));
 sg13g2_mux4_1 _2908_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A0(net1597),
    .A1(net1610),
    .A2(net649),
    .A3(net1632),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0975_));
 sg13g2_mux4_1 _2909_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A0(net1591),
    .A1(net1585),
    .A2(net1522),
    .A3(net1520),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0976_));
 sg13g2_nand2b_1 _2910_ (.Y(_0977_),
    .B(_0102_),
    .A_N(_0975_));
 sg13g2_o21ai_1 _2911_ (.B1(_0977_),
    .Y(_0978_),
    .A1(_0976_),
    .A2(_0102_));
 sg13g2_mux4_1 _2912_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A0(net1708),
    .A1(net135),
    .A2(net2003),
    .A3(net8),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0979_));
 sg13g2_nand2_1 _2913_ (.Y(_0980_),
    .A(_0102_),
    .B(_0979_));
 sg13g2_nand2_1 _2914_ (.Y(_0981_),
    .A(net34),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_o21ai_1 _2915_ (.B1(_0981_),
    .Y(_0982_),
    .A1(_0059_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_or2_1 _2916_ (.X(_0983_),
    .B(_0982_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_nand2b_1 _2917_ (.Y(_0984_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ),
    .A_N(net1929));
 sg13g2_o21ai_1 _2918_ (.B1(_0984_),
    .Y(_0985_),
    .A1(net69),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_a21oi_1 _2919_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0985_),
    .Y(_0986_),
    .B1(_0102_));
 sg13g2_a21oi_1 _2920_ (.A1(_0983_),
    .A2(_0986_),
    .Y(_0987_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_a22oi_1 _2921_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .B1(_0980_),
    .B2(_0987_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ),
    .A1(_0978_));
 sg13g2_mux4_1 _2922_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .A0(net1531),
    .A1(net1537),
    .A2(net1545),
    .A3(net1552),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0988_));
 sg13g2_nor2_2 _2923_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_mux2_1 _2924_ (.A0(net1555),
    .A1(net1562),
    .S(net1661),
    .X(_0990_));
 sg13g2_o21ai_1 _2925_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0991_),
    .A1(net1661),
    .A2(net1581));
 sg13g2_a21oi_1 _2926_ (.A1(net1661),
    .A2(_0178_),
    .Y(_0992_),
    .B1(_0991_));
 sg13g2_o21ai_1 _2927_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_0993_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0990_));
 sg13g2_nor2_2 _2928_ (.A(_0106_),
    .B(_0989_),
    .Y(_0994_));
 sg13g2_o21ai_1 _2929_ (.B1(_0994_),
    .Y(_0995_),
    .A1(_0992_),
    .A2(_0993_));
 sg13g2_a21oi_1 _2930_ (.A1(_0081_),
    .A2(net1661),
    .Y(_0996_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_o21ai_1 _2931_ (.B1(_0996_),
    .Y(_0997_),
    .A1(net1661),
    .A2(_0723_));
 sg13g2_nor2b_1 _2932_ (.A(net150),
    .B_N(net1661),
    .Y(_0998_));
 sg13g2_o21ai_1 _2933_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .Y(_0999_),
    .A1(net1661),
    .A2(net148));
 sg13g2_o21ai_1 _2934_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .Y(_1000_),
    .A1(_0998_),
    .A2(_0999_));
 sg13g2_nor2b_1 _2935_ (.A(_1000_),
    .B_N(_0997_),
    .Y(_1001_));
 sg13g2_mux4_1 _2936_ (.S0(net1661),
    .A0(net1710),
    .A1(net122),
    .A2(net1925),
    .A3(net98),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_1002_));
 sg13g2_o21ai_1 _2937_ (.B1(_0106_),
    .Y(_1003_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_1002_));
 sg13g2_o21ai_1 _2938_ (.B1(_0995_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(_1003_),
    .A2(_1001_));
 sg13g2_mux4_1 _2939_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(net79),
    .A2(net44),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ),
    .X(_1004_));
 sg13g2_mux4_1 _2940_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .A1(net45),
    .A2(net19),
    .A3(net80),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ),
    .X(_1005_));
 sg13g2_mux4_1 _2941_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ),
    .A0(_1004_),
    .A1(_1005_),
    .A2(_0974_),
    .A3(_0721_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ));
 sg13g2_mux2_2 _2942_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ),
    .S(net1642),
    .X(_1006_));
 sg13g2_inv_1 _2943_ (.Y(_1007_),
    .A(_1006_));
 sg13g2_nand2_2 _2944_ (.Y(_1008_),
    .A(_0973_),
    .B(_1006_));
 sg13g2_xnor2_1 _2945_ (.Y(_1009_),
    .A(_0931_),
    .B(_0932_));
 sg13g2_nor2_2 _2946_ (.A(_1009_),
    .B(_1008_),
    .Y(_1010_));
 sg13g2_mux4_1 _2947_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A1(net15),
    .A2(net41),
    .A3(net76),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_1011_));
 sg13g2_mux4_1 _2948_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ),
    .A0(net14),
    .A1(net75),
    .A2(net40),
    .A3(net705),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_1012_));
 sg13g2_nor2b_1 _2949_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .B_N(_1012_),
    .Y(_1013_));
 sg13g2_a21oi_1 _2950_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_1011_),
    .Y(_1014_),
    .B1(_1013_));
 sg13g2_mux2_1 _2951_ (.A0(net72),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_1015_));
 sg13g2_nand2_1 _2952_ (.Y(_1016_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ),
    .B(_1015_));
 sg13g2_a21oi_1 _2953_ (.A1(_0062_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ),
    .Y(_1017_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_o21ai_1 _2954_ (.B1(_1017_),
    .Y(_1018_),
    .A1(net24),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_nand3_1 _2955_ (.B(_1016_),
    .C(_1018_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .Y(_1019_));
 sg13g2_mux4_1 _2956_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(net143),
    .A1(net32),
    .A2(net6),
    .A3(net67),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_1020_));
 sg13g2_o21ai_1 _2957_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ),
    .Y(_1021_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_1020_));
 sg13g2_nand2b_1 _2958_ (.Y(_1022_),
    .B(_1019_),
    .A_N(_1021_));
 sg13g2_o21ai_1 _2959_ (.B1(_1022_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .A1(_1014_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_mux2_2 _2960_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ),
    .S(net1642),
    .X(_1023_));
 sg13g2_inv_1 _2961_ (.Y(_1024_),
    .A(_1023_));
 sg13g2_nand2_1 _2962_ (.Y(_1025_),
    .A(net1575),
    .B(_1023_));
 sg13g2_nand2_1 _2963_ (.Y(_1026_),
    .A(_0849_),
    .B(_1006_));
 sg13g2_nand2_2 _2964_ (.Y(_1027_),
    .A(_1006_),
    .B(_0899_));
 sg13g2_or2_1 _2965_ (.X(_1028_),
    .B(_1026_),
    .A(_0931_));
 sg13g2_xnor2_1 _2966_ (.Y(_1029_),
    .A(_1027_),
    .B(_0850_));
 sg13g2_xor2_1 _2967_ (.B(_1029_),
    .A(_1025_),
    .X(_1030_));
 sg13g2_o21ai_1 _2968_ (.B1(_1030_),
    .Y(_1031_),
    .A1(_1010_),
    .A2(_0933_));
 sg13g2_xnor2_1 _2969_ (.Y(_1032_),
    .A(_0770_),
    .B(_0771_));
 sg13g2_or3_1 _2970_ (.A(_0933_),
    .B(_1010_),
    .C(_1030_),
    .X(_1033_));
 sg13g2_nand2_2 _2971_ (.Y(_1034_),
    .A(_1033_),
    .B(_1031_));
 sg13g2_or2_1 _2972_ (.X(_1035_),
    .B(_1032_),
    .A(_1034_));
 sg13g2_o21ai_1 _2973_ (.B1(_1028_),
    .Y(_1036_),
    .A1(_1025_),
    .A2(_1029_));
 sg13g2_nand2_1 _2974_ (.Y(_1037_),
    .A(_0702_),
    .B(net1575));
 sg13g2_nand2_1 _2975_ (.Y(_1038_),
    .A(_0849_),
    .B(_1023_));
 sg13g2_nand2_1 _2976_ (.Y(_1039_),
    .A(_0899_),
    .B(_1023_));
 sg13g2_nor2_2 _2977_ (.A(_1038_),
    .B(_1027_),
    .Y(_1040_));
 sg13g2_xor2_1 _2978_ (.B(_1039_),
    .A(_1026_),
    .X(_1041_));
 sg13g2_nor2b_1 _2979_ (.A(_1037_),
    .B_N(_1041_),
    .Y(_1042_));
 sg13g2_xnor2_1 _2980_ (.Y(_1043_),
    .A(_1037_),
    .B(_1041_));
 sg13g2_and2_1 _2981_ (.A(_1043_),
    .B(_1036_),
    .X(_1044_));
 sg13g2_xnor2_1 _2982_ (.Y(_1045_),
    .A(_1036_),
    .B(_1043_));
 sg13g2_nor3_1 _2983_ (.A(net1511),
    .B(net1515),
    .C(_1045_),
    .Y(_1046_));
 sg13g2_xor2_1 _2984_ (.B(_1045_),
    .A(_0519_),
    .X(_1047_));
 sg13g2_a21oi_2 _2985_ (.B1(_1047_),
    .Y(_1048_),
    .A2(_1035_),
    .A1(_1031_));
 sg13g2_nand3_1 _2986_ (.B(_1035_),
    .C(_1047_),
    .A(_1031_),
    .Y(_1049_));
 sg13g2_nand2b_1 _2987_ (.Y(_1050_),
    .B(_1049_),
    .A_N(_1048_));
 sg13g2_nor2_1 _2988_ (.A(_0772_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_xnor2_1 _2989_ (.Y(_1052_),
    .A(_1050_),
    .B(_0772_));
 sg13g2_a21oi_1 _2990_ (.A1(net102),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .Y(_1053_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_o21ai_1 _2991_ (.B1(_1053_),
    .Y(_1054_),
    .A1(_0074_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_nor2b_1 _2992_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .B_N(net638),
    .Y(_1055_));
 sg13g2_nand2_1 _2993_ (.Y(_1056_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ),
    .B(net162));
 sg13g2_nand2_1 _2994_ (.Y(_1057_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ),
    .B(_1056_));
 sg13g2_o21ai_1 _2995_ (.B1(_1054_),
    .Y(_1058_),
    .A1(_1055_),
    .A2(_1057_));
 sg13g2_mux4_1 _2996_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net1530),
    .A1(net1534),
    .A2(net1543),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1059_));
 sg13g2_mux4_1 _2997_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net1563),
    .A1(net1573),
    .A2(net1578),
    .A3(net1615),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1060_));
 sg13g2_nand2b_1 _2998_ (.Y(_1061_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A_N(_1060_));
 sg13g2_o21ai_1 _2999_ (.B1(_1061_),
    .Y(_1062_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_1059_));
 sg13g2_mux4_1 _3000_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net1711),
    .A1(net119),
    .A2(net131),
    .A3(net95),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1063_));
 sg13g2_nand2b_1 _3001_ (.Y(_1064_),
    .B(_1063_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_nand2_1 _3002_ (.Y(_1065_),
    .A(_0058_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_o21ai_1 _3003_ (.B1(_1065_),
    .Y(_1066_),
    .A1(net155),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_nor2_1 _3004_ (.A(net1924),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .Y(_1067_));
 sg13g2_a21oi_1 _3005_ (.A1(_0066_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ),
    .Y(_1068_),
    .B1(_1067_));
 sg13g2_o21ai_1 _3006_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ),
    .Y(_1069_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_1068_));
 sg13g2_a21oi_1 _3007_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_1066_),
    .Y(_1070_),
    .B1(_1069_));
 sg13g2_nor2_1 _3008_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .B(_1070_),
    .Y(_1071_));
 sg13g2_a22oi_1 _3009_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .B1(_1064_),
    .B2(_1071_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ),
    .A1(_1062_));
 sg13g2_mux2_1 _3010_ (.A0(net1550),
    .A1(net1559),
    .S(net1665),
    .X(_1072_));
 sg13g2_or2_1 _3011_ (.X(_1073_),
    .B(net1529),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_a21oi_1 _3012_ (.A1(net1665),
    .A2(_0176_),
    .Y(_1074_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_a221oi_1 _3013_ (.B2(_1074_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .B1(_1073_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_1075_),
    .A2(_1072_));
 sg13g2_o21ai_1 _3014_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_1076_),
    .A1(net1665),
    .A2(net1579));
 sg13g2_a21oi_1 _3015_ (.A1(net1665),
    .A2(_0178_),
    .Y(_1077_),
    .B1(_1076_));
 sg13g2_a21oi_1 _3016_ (.A1(net1665),
    .A2(net1570),
    .Y(_1078_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_o21ai_1 _3017_ (.B1(_1078_),
    .Y(_1079_),
    .A1(net1665),
    .A2(net1565));
 sg13g2_nand2_1 _3018_ (.Y(_1080_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .B(_1079_));
 sg13g2_o21ai_1 _3019_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ),
    .Y(_1081_),
    .A1(_1077_),
    .A2(_1080_));
 sg13g2_nor2_1 _3020_ (.A(_1075_),
    .B(_1081_),
    .Y(_1082_));
 sg13g2_mux4_1 _3021_ (.S0(net1665),
    .A0(net1713),
    .A1(net117),
    .A2(net133),
    .A3(net93),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_1083_));
 sg13g2_mux4_1 _3022_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ),
    .A0(net1924),
    .A1(net153),
    .A2(net1935),
    .A3(net172),
    .S1(net1665),
    .X(_1084_));
 sg13g2_mux2_1 _3023_ (.A0(_1083_),
    .A1(_1084_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_1085_));
 sg13g2_a21oi_2 _3024_ (.B1(_1082_),
    .Y(_1086_),
    .A2(_1085_),
    .A1(_0126_));
 sg13g2_inv_1 _3025_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .A(_1086_));
 sg13g2_o21ai_1 _3026_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .Y(_1087_),
    .A1(net158),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_a21oi_1 _3027_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .A2(_1086_),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_nand2b_1 _3028_ (.Y(_1089_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ),
    .A_N(net52));
 sg13g2_o21ai_1 _3029_ (.B1(_1089_),
    .Y(_1090_),
    .A1(net109),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_mux4_1 _3030_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(net139),
    .A1(net1935),
    .A2(net93),
    .A3(net153),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_1091_));
 sg13g2_nand2b_1 _3031_ (.Y(_1092_),
    .B(_1058_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_o21ai_1 _3032_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_1093_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ),
    .A2(_1090_));
 sg13g2_o21ai_1 _3033_ (.B1(_1092_),
    .Y(_1094_),
    .A1(_1088_),
    .A2(_1093_));
 sg13g2_nor2b_1 _3034_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .B_N(net161),
    .Y(_1095_));
 sg13g2_a21oi_2 _3035_ (.B1(_1095_),
    .Y(_1096_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ));
 sg13g2_a21oi_2 _3036_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_1097_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .A1(_1096_));
 sg13g2_mux2_1 _3037_ (.A0(net101),
    .A1(net715),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_1098_));
 sg13g2_o21ai_1 _3038_ (.B1(_1097_),
    .Y(_1099_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ),
    .A2(_1098_));
 sg13g2_a21oi_1 _3039_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ),
    .A2(_1091_),
    .Y(_1100_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_a22oi_1 _3040_ (.Y(\Tile_X0Y1_DSP_bot.A1 ),
    .B1(_1099_),
    .B2(_1100_),
    .A2(_1094_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_nand2_1 _3041_ (.Y(_1101_),
    .A(net1641),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ));
 sg13g2_nand2b_1 _3042_ (.Y(_1102_),
    .B(\Tile_X0Y1_DSP_bot.A1 ),
    .A_N(net1641));
 sg13g2_nand2_2 _3043_ (.Y(_1103_),
    .A(_1101_),
    .B(_1102_));
 sg13g2_inv_2 _3044_ (.Y(_1104_),
    .A(_1103_));
 sg13g2_a221oi_1 _3045_ (.B2(_1102_),
    .C1(_0898_),
    .B1(_1101_),
    .A1(_0123_),
    .Y(_1105_),
    .A2(_0897_));
 sg13g2_nand2_2 _3046_ (.Y(_1106_),
    .A(_1103_),
    .B(_0899_));
 sg13g2_nand2_1 _3047_ (.Y(_1107_),
    .A(_0849_),
    .B(_1103_));
 sg13g2_nand2_1 _3048_ (.Y(_1108_),
    .A(_0807_),
    .B(net1575));
 sg13g2_xnor2_1 _3049_ (.Y(_1109_),
    .A(_0930_),
    .B(_1107_));
 sg13g2_or2_1 _3050_ (.X(_1110_),
    .B(_1109_),
    .A(_1108_));
 sg13g2_o21ai_1 _3051_ (.B1(_1110_),
    .Y(_1111_),
    .A1(_0932_),
    .A2(_1106_));
 sg13g2_xor2_1 _3052_ (.B(_1009_),
    .A(_1008_),
    .X(_1112_));
 sg13g2_xnor2_1 _3053_ (.Y(_1113_),
    .A(_1111_),
    .B(_1112_));
 sg13g2_mux4_1 _3054_ (.S0(net1668),
    .A0(net1531),
    .A1(net1536),
    .A2(net1545),
    .A3(net1552),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_1114_));
 sg13g2_nor2_2 _3055_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .B(_1114_),
    .Y(_1115_));
 sg13g2_mux2_1 _3056_ (.A0(net1562),
    .A1(net1571),
    .S(net1668),
    .X(_1116_));
 sg13g2_o21ai_1 _3057_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_1117_),
    .A1(net1668),
    .A2(net1582));
 sg13g2_a21oi_1 _3058_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0178_),
    .Y(_1118_),
    .B1(_1117_));
 sg13g2_o21ai_1 _3059_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_1119_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_1116_));
 sg13g2_nor2_2 _3060_ (.A(_0127_),
    .B(_1115_),
    .Y(_1120_));
 sg13g2_o21ai_1 _3061_ (.B1(_1120_),
    .Y(_1121_),
    .A1(_1118_),
    .A2(_1119_));
 sg13g2_nand2b_1 _3062_ (.Y(_1122_),
    .B(_0615_),
    .A_N(net1668));
 sg13g2_a21oi_1 _3063_ (.A1(_0099_),
    .A2(net1668),
    .Y(_1123_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_nor2b_1 _3064_ (.A(net150),
    .B_N(net1668),
    .Y(_1124_));
 sg13g2_o21ai_1 _3065_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_1125_),
    .A1(net148),
    .A2(net1668));
 sg13g2_o21ai_1 _3066_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_1126_),
    .A1(_1124_),
    .A2(_1125_));
 sg13g2_a21oi_1 _3067_ (.A1(_1122_),
    .A2(_1123_),
    .Y(_1127_),
    .B1(_1126_));
 sg13g2_mux4_1 _3068_ (.S0(net1668),
    .A0(net112),
    .A1(net120),
    .A2(net1927),
    .A3(net96),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_1128_));
 sg13g2_o21ai_1 _3069_ (.B1(_0127_),
    .Y(_1129_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_1128_));
 sg13g2_o21ai_1 _3070_ (.B1(_1121_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .A1(_1127_),
    .A2(_1129_));
 sg13g2_mux4_1 _3071_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(net1708),
    .A1(net103),
    .A2(net615),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ),
    .X(_1130_));
 sg13g2_mux4_1 _3072_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(net128),
    .A1(net104),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net164),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_1131_));
 sg13g2_mux2_1 _3073_ (.A0(net1579),
    .A1(net1616),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_1132_));
 sg13g2_mux2_1 _3074_ (.A0(net1561),
    .A1(net1570),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_1133_));
 sg13g2_o21ai_1 _3075_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_1134_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_1133_));
 sg13g2_a21oi_1 _3076_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_1132_),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_mux4_1 _3077_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net1529),
    .A1(net1535),
    .A2(net1550),
    .A3(net1559),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_1136_));
 sg13g2_o21ai_1 _3078_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_1137_),
    .A1(_1136_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_nor2_1 _3079_ (.A(_0068_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .Y(_1138_));
 sg13g2_a21oi_1 _3080_ (.A1(net53),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .Y(_1139_),
    .B1(_1138_));
 sg13g2_mux2_1 _3081_ (.A0(net154),
    .A1(net168),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_1140_));
 sg13g2_o21ai_1 _3082_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_1141_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_1139_));
 sg13g2_a21oi_1 _3083_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .A2(_1140_),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_mux4_1 _3084_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net142),
    .A1(net1927),
    .A2(net94),
    .A3(net1922),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_1143_));
 sg13g2_nor2_1 _3085_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ),
    .B(_1142_),
    .Y(_1144_));
 sg13g2_o21ai_1 _3086_ (.B1(_1144_),
    .Y(_1145_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_1143_));
 sg13g2_o21ai_1 _3087_ (.B1(_1145_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .A1(_1137_),
    .A2(_1135_));
 sg13g2_mux4_1 _3088_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(net140),
    .A1(net108),
    .A2(net51),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_1146_));
 sg13g2_mux4_1 _3089_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(net119),
    .A1(net95),
    .A2(net60),
    .A3(net155),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_1147_));
 sg13g2_mux4_1 _3090_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ),
    .A0(_1130_),
    .A1(_1131_),
    .A2(_1147_),
    .A3(_1146_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.B2 ));
 sg13g2_mux2_1 _3091_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ),
    .A1(\Tile_X0Y1_DSP_bot.B2 ),
    .S(net1640),
    .X(_1148_));
 sg13g2_nand2b_1 _3092_ (.Y(_1149_),
    .B(_1148_),
    .A_N(_0518_));
 sg13g2_nor2_1 _3093_ (.A(net1608),
    .B(_1024_),
    .Y(_1150_));
 sg13g2_inv_1 _3094_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_nor2_1 _3095_ (.A(net1511),
    .B(_1024_),
    .Y(_1152_));
 sg13g2_xor2_1 _3096_ (.B(_1152_),
    .A(_0769_),
    .X(_1153_));
 sg13g2_nor2b_1 _3097_ (.A(_1149_),
    .B_N(_1153_),
    .Y(_1154_));
 sg13g2_xnor2_1 _3098_ (.Y(_1155_),
    .A(_1149_),
    .B(_1153_));
 sg13g2_nor2b_1 _3099_ (.A(_1113_),
    .B_N(_1155_),
    .Y(_1156_));
 sg13g2_a21o_1 _3100_ (.A2(_1112_),
    .A1(_1111_),
    .B1(_1156_),
    .X(_1157_));
 sg13g2_xnor2_1 _3101_ (.Y(_1158_),
    .A(_1032_),
    .B(_1034_));
 sg13g2_nand2b_1 _3102_ (.Y(_1159_),
    .B(_1157_),
    .A_N(_1158_));
 sg13g2_a21o_1 _3103_ (.A2(_1152_),
    .A1(_0769_),
    .B1(_1154_),
    .X(_1160_));
 sg13g2_xor2_1 _3104_ (.B(_1158_),
    .A(_1157_),
    .X(_1161_));
 sg13g2_nand2b_1 _3105_ (.Y(_1162_),
    .B(_1160_),
    .A_N(_1161_));
 sg13g2_a21o_1 _3106_ (.A2(_1162_),
    .A1(_1159_),
    .B1(_1052_),
    .X(_1163_));
 sg13g2_nand2b_1 _3107_ (.Y(_1164_),
    .B(net1575),
    .A_N(net1515));
 sg13g2_nor2_1 _3108_ (.A(_0703_),
    .B(_0848_),
    .Y(_1165_));
 sg13g2_nand2_2 _3109_ (.Y(_1166_),
    .A(_0702_),
    .B(_0899_));
 sg13g2_or2_1 _3110_ (.X(_1167_),
    .B(_1166_),
    .A(_1038_));
 sg13g2_xnor2_1 _3111_ (.Y(_1168_),
    .A(_1038_),
    .B(_1166_));
 sg13g2_xor2_1 _3112_ (.B(_1168_),
    .A(_1164_),
    .X(_1169_));
 sg13g2_nor2_2 _3113_ (.A(_1042_),
    .B(_1040_),
    .Y(_1170_));
 sg13g2_nand2b_1 _3114_ (.Y(_1171_),
    .B(_1169_),
    .A_N(_1170_));
 sg13g2_xnor2_1 _3115_ (.Y(_1172_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_o21ai_1 _3116_ (.B1(_1172_),
    .Y(_1173_),
    .A1(_1046_),
    .A2(_1044_));
 sg13g2_or3_1 _3117_ (.A(_1044_),
    .B(_1046_),
    .C(_1172_),
    .X(_1174_));
 sg13g2_and2_1 _3118_ (.A(_1174_),
    .B(_1173_),
    .X(_1175_));
 sg13g2_o21ai_1 _3119_ (.B1(_1175_),
    .Y(_1176_),
    .A1(_1048_),
    .A2(_1051_));
 sg13g2_or3_1 _3120_ (.A(_1048_),
    .B(_1051_),
    .C(_1175_),
    .X(_1177_));
 sg13g2_and2_1 _3121_ (.A(_1177_),
    .B(_1176_),
    .X(_1178_));
 sg13g2_nor2b_1 _3122_ (.A(_1163_),
    .B_N(_1178_),
    .Y(_1179_));
 sg13g2_xnor2_1 _3123_ (.Y(_1180_),
    .A(_1178_),
    .B(_1163_));
 sg13g2_mux4_1 _3124_ (.S0(net1691),
    .A0(net1599),
    .A1(net1612),
    .A2(net1605),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1181_));
 sg13g2_inv_1 _3125_ (.Y(_1182_),
    .A(_1181_));
 sg13g2_mux4_1 _3126_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(net1634),
    .A1(net1523),
    .A2(net1593),
    .A3(net1540),
    .S1(net1691),
    .X(_1183_));
 sg13g2_o21ai_1 _3127_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .Y(_1184_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1182_));
 sg13g2_a21oi_1 _3128_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_1183_),
    .Y(_1185_),
    .B1(_1184_));
 sg13g2_a21oi_1 _3129_ (.A1(net130),
    .A2(net1691),
    .Y(_1186_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_o21ai_1 _3130_ (.B1(_1186_),
    .Y(_1187_),
    .A1(net1691),
    .A2(net622));
 sg13g2_nor2b_1 _3131_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .B_N(net2001),
    .Y(_1188_));
 sg13g2_a21oi_1 _3132_ (.A1(net11),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .Y(_1189_),
    .B1(_1188_));
 sg13g2_a21oi_1 _3133_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_1189_),
    .Y(_1190_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_a21oi_1 _3134_ (.A1(net37),
    .A2(net1691),
    .Y(_1191_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_o21ai_1 _3135_ (.B1(_1191_),
    .Y(_1192_),
    .A1(_0090_),
    .A2(net1691));
 sg13g2_nand2b_1 _3136_ (.Y(_1193_),
    .B(net1691),
    .A_N(net1930));
 sg13g2_o21ai_1 _3137_ (.B1(_1193_),
    .Y(_1194_),
    .A1(net1933),
    .A2(net1691));
 sg13g2_a21oi_1 _3138_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_1194_),
    .Y(_1195_),
    .B1(_0120_));
 sg13g2_a221oi_1 _3139_ (.B2(_1195_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ),
    .B1(_1192_),
    .A1(_1190_),
    .Y(_1196_),
    .A2(_1187_));
 sg13g2_nor2_2 _3140_ (.A(_1196_),
    .B(_1185_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ));
 sg13g2_nor2b_1 _3141_ (.A(net624),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .Y(_1197_));
 sg13g2_nor2_1 _3142_ (.A(net1707),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .Y(_1198_));
 sg13g2_nor3_1 _3143_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .B(_1197_),
    .C(_1198_),
    .Y(_1199_));
 sg13g2_o21ai_1 _3144_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ),
    .Y(_1200_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(net165));
 sg13g2_a21oi_1 _3145_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ),
    .A2(net633),
    .Y(_1201_),
    .B1(_1200_));
 sg13g2_nor3_1 _3146_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .B(_1199_),
    .C(_1201_),
    .Y(_1202_));
 sg13g2_nand2_1 _3147_ (.Y(_1203_),
    .A(net166),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_o21ai_1 _3148_ (.B1(_1203_),
    .Y(_1204_),
    .A1(_0347_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_nand2b_1 _3149_ (.Y(_1205_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ),
    .A_N(net106));
 sg13g2_o21ai_1 _3150_ (.B1(_1205_),
    .Y(_1206_),
    .A1(net1706),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_o21ai_1 _3151_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .Y(_1207_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .A2(_1206_));
 sg13g2_a21oi_2 _3152_ (.B1(_1207_),
    .Y(_1208_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ),
    .A1(_1204_));
 sg13g2_nor3_2 _3153_ (.A(_1208_),
    .B(_1202_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .Y(_1209_));
 sg13g2_mux4_1 _3154_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(net121),
    .A1(net97),
    .A2(net61),
    .A3(net157),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_1210_));
 sg13g2_o21ai_1 _3155_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ),
    .Y(_1211_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_1210_));
 sg13g2_a21oi_1 _3156_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(net668),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_or2_1 _3157_ (.X(\Tile_X0Y1_DSP_bot.A0 ),
    .B(_1209_),
    .A(_1212_));
 sg13g2_mux2_2 _3158_ (.A0(\Tile_X0Y1_DSP_bot.A0 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ),
    .S(net1641),
    .X(_1213_));
 sg13g2_inv_8 _3159_ (.Y(_1214_),
    .A(_1213_));
 sg13g2_nor2_1 _3160_ (.A(_0848_),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_nand2_1 _3161_ (.Y(_1216_),
    .A(_1105_),
    .B(_1215_));
 sg13g2_nand2_1 _3162_ (.Y(_1217_),
    .A(net714),
    .B(net1575));
 sg13g2_xnor2_1 _3163_ (.Y(_1218_),
    .A(_1105_),
    .B(_1215_));
 sg13g2_o21ai_1 _3164_ (.B1(_1216_),
    .Y(_1219_),
    .A1(_1217_),
    .A2(_1218_));
 sg13g2_xor2_1 _3165_ (.B(_1109_),
    .A(_1108_),
    .X(_1220_));
 sg13g2_xnor2_1 _3166_ (.Y(_1221_),
    .A(_1219_),
    .B(_1220_));
 sg13g2_nand2b_1 _3167_ (.Y(_1222_),
    .B(_1006_),
    .A_N(net1608));
 sg13g2_nand2b_1 _3168_ (.Y(_1223_),
    .B(_1006_),
    .A_N(net1511));
 sg13g2_xnor2_1 _3169_ (.Y(_1224_),
    .A(_1150_),
    .B(_1223_));
 sg13g2_nand3_1 _3170_ (.B(net1628),
    .C(_1224_),
    .A(_0702_),
    .Y(_1225_));
 sg13g2_a21o_1 _3171_ (.A2(net1628),
    .A1(_0702_),
    .B1(_1224_),
    .X(_1226_));
 sg13g2_and2_1 _3172_ (.A(_1225_),
    .B(_1226_),
    .X(_1227_));
 sg13g2_nor2b_1 _3173_ (.A(_1221_),
    .B_N(_1227_),
    .Y(_1228_));
 sg13g2_a21o_1 _3174_ (.A2(_1220_),
    .A1(_1219_),
    .B1(_1228_),
    .X(_1229_));
 sg13g2_xnor2_1 _3175_ (.Y(_1230_),
    .A(_1113_),
    .B(_1155_));
 sg13g2_o21ai_1 _3176_ (.B1(_1225_),
    .Y(_1231_),
    .A1(_1151_),
    .A2(_1223_));
 sg13g2_xnor2_1 _3177_ (.Y(_1232_),
    .A(_1229_),
    .B(_1230_));
 sg13g2_nor2b_1 _3178_ (.A(_1232_),
    .B_N(_1231_),
    .Y(_1233_));
 sg13g2_a21o_1 _3179_ (.A2(_1230_),
    .A1(_1229_),
    .B1(_1233_),
    .X(_1234_));
 sg13g2_xnor2_1 _3180_ (.Y(_1235_),
    .A(_1160_),
    .B(_1161_));
 sg13g2_nand3_1 _3181_ (.B(_1159_),
    .C(_1162_),
    .A(_1052_),
    .Y(_1236_));
 sg13g2_and2_1 _3182_ (.A(_1236_),
    .B(_1163_),
    .X(_1237_));
 sg13g2_a21o_1 _3183_ (.A2(_1235_),
    .A1(_1234_),
    .B1(_1237_),
    .X(_1238_));
 sg13g2_and3_1 _3184_ (.X(_1239_),
    .A(_1234_),
    .B(_1235_),
    .C(_1237_));
 sg13g2_inv_1 _3185_ (.Y(_1240_),
    .A(_1239_));
 sg13g2_xnor2_1 _3186_ (.Y(_1241_),
    .A(_1234_),
    .B(_1235_));
 sg13g2_nand2_1 _3187_ (.Y(_1242_),
    .A(net1575),
    .B(_1213_));
 sg13g2_nor2_2 _3188_ (.A(_1106_),
    .B(_1242_),
    .Y(_1243_));
 sg13g2_nand3_1 _3189_ (.B(_1105_),
    .C(_1213_),
    .A(net1575),
    .Y(_1244_));
 sg13g2_xnor2_1 _3190_ (.Y(_1245_),
    .A(_1217_),
    .B(_1218_));
 sg13g2_nand2_1 _3191_ (.Y(_1246_),
    .A(_1023_),
    .B(net1628));
 sg13g2_nor2_2 _3192_ (.A(net1608),
    .B(_0808_),
    .Y(_1247_));
 sg13g2_nor2_1 _3193_ (.A(net1511),
    .B(_0808_),
    .Y(_1248_));
 sg13g2_nand2b_1 _3194_ (.Y(_1249_),
    .B(_1247_),
    .A_N(_1223_));
 sg13g2_xnor2_1 _3195_ (.Y(_1250_),
    .A(_1222_),
    .B(_1248_));
 sg13g2_inv_1 _3196_ (.Y(_1251_),
    .A(_1250_));
 sg13g2_xnor2_1 _3197_ (.Y(_1252_),
    .A(_1246_),
    .B(_1250_));
 sg13g2_xnor2_1 _3198_ (.Y(_1253_),
    .A(_1243_),
    .B(_1245_));
 sg13g2_nand2_1 _3199_ (.Y(_1254_),
    .A(_1252_),
    .B(_1253_));
 sg13g2_o21ai_1 _3200_ (.B1(_1254_),
    .Y(_1255_),
    .A1(_1244_),
    .A2(_1245_));
 sg13g2_xor2_1 _3201_ (.B(_1227_),
    .A(_1221_),
    .X(_1256_));
 sg13g2_nor2b_1 _3202_ (.A(_1256_),
    .B_N(_1255_),
    .Y(_1257_));
 sg13g2_o21ai_1 _3203_ (.B1(_1249_),
    .Y(_1258_),
    .A1(_1246_),
    .A2(_1251_));
 sg13g2_mux4_1 _3204_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(net117),
    .A1(net93),
    .A2(net1935),
    .A3(net171),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ),
    .X(_1259_));
 sg13g2_mux2_1 _3205_ (.A0(_1259_),
    .A1(_0308_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .X(_1260_));
 sg13g2_mux4_1 _3206_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net645),
    .A1(_0724_),
    .A2(_0099_),
    .A3(_0105_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_1261_));
 sg13g2_mux4_1 _3207_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net1712),
    .A1(net120),
    .A2(net1927),
    .A3(net96),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_1262_));
 sg13g2_o21ai_1 _3208_ (.B1(_0128_),
    .Y(_1263_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_1262_));
 sg13g2_a21o_1 _3209_ (.A2(_1261_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .B1(_1263_),
    .X(_1264_));
 sg13g2_mux2_1 _3210_ (.A0(net1562),
    .A1(net1571),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_1265_));
 sg13g2_mux2_1 _3211_ (.A0(net1582),
    .A1(net1619),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_1266_));
 sg13g2_o21ai_1 _3212_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .Y(_1267_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .A2(_1265_));
 sg13g2_a21o_1 _3213_ (.A2(_1266_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .B1(_1267_),
    .X(_1268_));
 sg13g2_mux4_1 _3214_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net1533),
    .A1(net635),
    .A2(net1547),
    .A3(net1554),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_1269_));
 sg13g2_o21ai_1 _3215_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ),
    .Y(_1270_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_1269_));
 sg13g2_nand2b_1 _3216_ (.Y(_1271_),
    .B(_1268_),
    .A_N(_1270_));
 sg13g2_nand2_2 _3217_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .A(_1264_),
    .B(_1271_));
 sg13g2_and3_1 _3218_ (.X(_1272_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .B(_1264_),
    .C(_1271_));
 sg13g2_o21ai_1 _3219_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ),
    .Y(_1273_),
    .A1(net161),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_mux2_1 _3220_ (.A0(net125),
    .A1(net101),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_1274_));
 sg13g2_a21oi_1 _3221_ (.A1(_0129_),
    .A2(_1274_),
    .Y(_1275_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_o21ai_1 _3222_ (.B1(_1275_),
    .Y(_1276_),
    .A1(_1272_),
    .A2(_1273_));
 sg13g2_mux4_1 _3223_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(net126),
    .A1(net102),
    .A2(net639),
    .A3(net162),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_1277_));
 sg13g2_inv_4 _3224_ (.A(_1277_),
    .Y(_1278_));
 sg13g2_a21oi_2 _3225_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_1279_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ),
    .A1(_1278_));
 sg13g2_a22oi_1 _3226_ (.Y(_1280_),
    .B1(_1276_),
    .B2(_1279_),
    .A2(_1260_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_inv_1 _3227_ (.Y(\Tile_X0Y1_DSP_bot.B1 ),
    .A(_1280_));
 sg13g2_nor2_1 _3228_ (.A(net1640),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ),
    .Y(_1281_));
 sg13g2_a21o_2 _3229_ (.A2(net1640),
    .A1(_1280_),
    .B1(_1281_),
    .X(_1282_));
 sg13g2_nor2_2 _3230_ (.A(_1282_),
    .B(net1515),
    .Y(_1283_));
 sg13g2_nand2_2 _3231_ (.Y(_1284_),
    .A(_1258_),
    .B(_1283_));
 sg13g2_xnor2_1 _3232_ (.Y(_1285_),
    .A(_1258_),
    .B(_1283_));
 sg13g2_xnor2_1 _3233_ (.Y(_1286_),
    .A(_1255_),
    .B(_1256_));
 sg13g2_nand2b_1 _3234_ (.Y(_1287_),
    .B(_1286_),
    .A_N(_1285_));
 sg13g2_nand2b_1 _3235_ (.Y(_1288_),
    .B(_1287_),
    .A_N(_1257_));
 sg13g2_xor2_1 _3236_ (.B(_1232_),
    .A(_1231_),
    .X(_1289_));
 sg13g2_nand2b_1 _3237_ (.Y(_1290_),
    .B(_1288_),
    .A_N(_1289_));
 sg13g2_xor2_1 _3238_ (.B(_1289_),
    .A(_1288_),
    .X(_1291_));
 sg13g2_or2_1 _3239_ (.X(_1292_),
    .B(_1291_),
    .A(_1284_));
 sg13g2_a21oi_2 _3240_ (.B1(_1241_),
    .Y(_1293_),
    .A2(_1292_),
    .A1(_1290_));
 sg13g2_nand3_1 _3241_ (.B(_1290_),
    .C(_1292_),
    .A(_1241_),
    .Y(_1294_));
 sg13g2_nand2b_1 _3242_ (.Y(_1295_),
    .B(_1294_),
    .A_N(_1293_));
 sg13g2_a22oi_1 _3243_ (.Y(_1296_),
    .B1(_1213_),
    .B2(_0899_),
    .A2(_1103_),
    .A1(net1575));
 sg13g2_nor2_1 _3244_ (.A(_1243_),
    .B(_1296_),
    .Y(_1297_));
 sg13g2_nand2_1 _3245_ (.Y(_1298_),
    .A(_1006_),
    .B(net1628));
 sg13g2_nor2_1 _3246_ (.A(net1608),
    .B(net625),
    .Y(_1299_));
 sg13g2_nor2_1 _3247_ (.A(net1511),
    .B(net625),
    .Y(_1300_));
 sg13g2_nand2_1 _3248_ (.Y(_1301_),
    .A(_1248_),
    .B(_1299_));
 sg13g2_nor2_1 _3249_ (.A(_1247_),
    .B(_1300_),
    .Y(_1302_));
 sg13g2_xor2_1 _3250_ (.B(_1300_),
    .A(_1247_),
    .X(_1303_));
 sg13g2_xnor2_1 _3251_ (.Y(_1304_),
    .A(_1303_),
    .B(_1298_));
 sg13g2_nand2_1 _3252_ (.Y(_1305_),
    .A(_1297_),
    .B(_1304_));
 sg13g2_xnor2_1 _3253_ (.Y(_1306_),
    .A(_1252_),
    .B(_1253_));
 sg13g2_nor2_1 _3254_ (.A(_1305_),
    .B(_1306_),
    .Y(_1307_));
 sg13g2_or2_1 _3255_ (.X(_1308_),
    .B(net1548),
    .A(_0703_));
 sg13g2_o21ai_1 _3256_ (.B1(_1301_),
    .Y(_1309_),
    .A1(_1298_),
    .A2(_1302_));
 sg13g2_o21ai_1 _3257_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .Y(_1310_),
    .A1(net171),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_a21oi_1 _3258_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .A2(_0966_),
    .Y(_1311_),
    .B1(_1310_));
 sg13g2_nor2b_1 _3259_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .B_N(net94),
    .Y(_1312_));
 sg13g2_a21oi_1 _3260_ (.A1(net61),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ),
    .Y(_1313_),
    .B1(_1312_));
 sg13g2_o21ai_1 _3261_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .Y(_1314_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_1313_));
 sg13g2_mux4_1 _3262_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(net142),
    .A1(net97),
    .A2(net44),
    .A3(net157),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_1315_));
 sg13g2_inv_1 _3263_ (.Y(_1316_),
    .A(_1315_));
 sg13g2_o21ai_1 _3264_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_1317_),
    .A1(_1311_),
    .A2(_1314_));
 sg13g2_inv_1 _3265_ (.Y(_1318_),
    .A(_1317_));
 sg13g2_o21ai_1 _3266_ (.B1(_1318_),
    .Y(_1319_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_1315_));
 sg13g2_nand3b_1 _3267_ (.B(_0626_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .Y(_1320_),
    .A_N(_0552_));
 sg13g2_o21ai_1 _3268_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ),
    .Y(_1321_),
    .A1(net165),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_inv_1 _3269_ (.Y(_1322_),
    .A(_1321_));
 sg13g2_mux2_1 _3270_ (.A0(net105),
    .A1(net624),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_1323_));
 sg13g2_a221oi_1 _3271_ (.B2(_1323_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .B1(_0130_),
    .A1(_1320_),
    .Y(_1324_),
    .A2(_1322_));
 sg13g2_o21ai_1 _3272_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .Y(_1325_),
    .A1(net166),
    .A2(_0131_));
 sg13g2_a21oi_1 _3273_ (.A1(_0131_),
    .A2(_0347_),
    .Y(_1326_),
    .B1(_1325_));
 sg13g2_nand2b_1 _3274_ (.Y(_1327_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ),
    .A_N(net106));
 sg13g2_o21ai_1 _3275_ (.B1(_1327_),
    .Y(_1328_),
    .A1(net1706),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_o21ai_1 _3276_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ),
    .Y(_1329_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ),
    .A2(_1328_));
 sg13g2_o21ai_1 _3277_ (.B1(_0132_),
    .Y(_1330_),
    .A1(_1326_),
    .A2(_1329_));
 sg13g2_o21ai_1 _3278_ (.B1(_1319_),
    .Y(\Tile_X0Y1_DSP_bot.B0 ),
    .A1(_1324_),
    .A2(_1330_));
 sg13g2_mux2_1 _3279_ (.A0(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ),
    .A1(\Tile_X0Y1_DSP_bot.B0 ),
    .S(net1640),
    .X(_1331_));
 sg13g2_nor2b_1 _3280_ (.A(net1515),
    .B_N(_1331_),
    .Y(_1332_));
 sg13g2_xnor2_1 _3281_ (.Y(_1333_),
    .A(_1309_),
    .B(_1332_));
 sg13g2_nor2_1 _3282_ (.A(_1308_),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_xor2_1 _3283_ (.B(_1333_),
    .A(_1308_),
    .X(_1335_));
 sg13g2_xor2_1 _3284_ (.B(_1306_),
    .A(_1305_),
    .X(_1336_));
 sg13g2_a21oi_1 _3285_ (.A1(_1335_),
    .A2(_1336_),
    .Y(_1337_),
    .B1(_1307_));
 sg13g2_xnor2_1 _3286_ (.Y(_1338_),
    .A(_1285_),
    .B(_1286_));
 sg13g2_nor2b_1 _3287_ (.A(_1337_),
    .B_N(_1338_),
    .Y(_1339_));
 sg13g2_a21o_1 _3288_ (.A2(_1332_),
    .A1(_1309_),
    .B1(_1334_),
    .X(_1340_));
 sg13g2_xnor2_1 _3289_ (.Y(_1341_),
    .A(_1337_),
    .B(_1338_));
 sg13g2_a21o_1 _3290_ (.A2(_1341_),
    .A1(_1340_),
    .B1(_1339_),
    .X(_1342_));
 sg13g2_xnor2_1 _3291_ (.Y(_1343_),
    .A(_1284_),
    .B(_1291_));
 sg13g2_inv_4 _3292_ (.A(_1343_),
    .Y(_1344_));
 sg13g2_nor2_2 _3293_ (.A(_1344_),
    .B(_1342_),
    .Y(_1345_));
 sg13g2_nand2_1 _3294_ (.Y(_1346_),
    .A(_0807_),
    .B(net1628));
 sg13g2_nor2_1 _3295_ (.A(net1511),
    .B(_1104_),
    .Y(_1347_));
 sg13g2_nand2_1 _3296_ (.Y(_1348_),
    .A(_1299_),
    .B(_1347_));
 sg13g2_xnor2_1 _3297_ (.Y(_1349_),
    .A(_1299_),
    .B(_1347_));
 sg13g2_xor2_1 _3298_ (.B(_1346_),
    .A(_1349_),
    .X(_1350_));
 sg13g2_nand2b_1 _3299_ (.Y(_1351_),
    .B(_1350_),
    .A_N(_1242_));
 sg13g2_xnor2_1 _3300_ (.Y(_1352_),
    .A(_1297_),
    .B(_1304_));
 sg13g2_nor2_1 _3301_ (.A(_1351_),
    .B(_1352_),
    .Y(_1353_));
 sg13g2_nor2_1 _3302_ (.A(_1024_),
    .B(_1282_),
    .Y(_1354_));
 sg13g2_inv_1 _3303_ (.Y(_1355_),
    .A(_1354_));
 sg13g2_o21ai_1 _3304_ (.B1(_1348_),
    .Y(_1356_),
    .A1(_1346_),
    .A2(_1349_));
 sg13g2_nand2_1 _3305_ (.Y(_1357_),
    .A(_0702_),
    .B(net1568));
 sg13g2_nand2b_1 _3306_ (.Y(_1358_),
    .B(_1356_),
    .A_N(_1357_));
 sg13g2_xor2_1 _3307_ (.B(_1357_),
    .A(_1356_),
    .X(_1359_));
 sg13g2_xnor2_1 _3308_ (.Y(_1360_),
    .A(_1355_),
    .B(_1359_));
 sg13g2_xor2_1 _3309_ (.B(_1352_),
    .A(_1351_),
    .X(_1361_));
 sg13g2_nor2b_1 _3310_ (.A(_1360_),
    .B_N(_1361_),
    .Y(_1362_));
 sg13g2_nor2_1 _3311_ (.A(_1353_),
    .B(_1362_),
    .Y(_1363_));
 sg13g2_xnor2_1 _3312_ (.Y(_1364_),
    .A(_1335_),
    .B(_1336_));
 sg13g2_nor2_1 _3313_ (.A(_1363_),
    .B(_1364_),
    .Y(_1365_));
 sg13g2_o21ai_1 _3314_ (.B1(_1358_),
    .Y(_1366_),
    .A1(_1355_),
    .A2(_1359_));
 sg13g2_xor2_1 _3315_ (.B(_1363_),
    .A(_1364_),
    .X(_1367_));
 sg13g2_a21oi_1 _3316_ (.A1(_1366_),
    .A2(_1367_),
    .Y(_1368_),
    .B1(_1365_));
 sg13g2_xnor2_1 _3317_ (.Y(_1369_),
    .A(_1340_),
    .B(_1341_));
 sg13g2_nor2_1 _3318_ (.A(_1368_),
    .B(_1369_),
    .Y(_1370_));
 sg13g2_xnor2_1 _3319_ (.Y(_1371_),
    .A(_1242_),
    .B(_1350_));
 sg13g2_nor2_1 _3320_ (.A(_1007_),
    .B(net1548),
    .Y(_1372_));
 sg13g2_nand2b_1 _3321_ (.Y(_1373_),
    .B(_1213_),
    .A_N(net1608));
 sg13g2_nor2_1 _3322_ (.A(net1511),
    .B(_1214_),
    .Y(_1374_));
 sg13g2_inv_1 _3323_ (.Y(_1375_),
    .A(_1374_));
 sg13g2_nor3_2 _3324_ (.A(net1608),
    .B(_1104_),
    .C(_1375_),
    .Y(_1376_));
 sg13g2_and2_1 _3325_ (.A(net714),
    .B(net1628),
    .X(_1377_));
 sg13g2_o21ai_1 _3326_ (.B1(_1375_),
    .Y(_1378_),
    .A1(net1608),
    .A2(_1104_));
 sg13g2_nand2b_1 _3327_ (.Y(_1379_),
    .B(_1378_),
    .A_N(_1376_));
 sg13g2_a21o_1 _3328_ (.A2(_1378_),
    .A1(_1377_),
    .B1(_1376_),
    .X(_1380_));
 sg13g2_nand2_1 _3329_ (.Y(_1381_),
    .A(_1023_),
    .B(net1568));
 sg13g2_inv_1 _3330_ (.Y(_1382_),
    .A(_1381_));
 sg13g2_xnor2_1 _3331_ (.Y(_1383_),
    .A(_1380_),
    .B(_1382_));
 sg13g2_nor3_1 _3332_ (.A(_1007_),
    .B(net1548),
    .C(_1383_),
    .Y(_1384_));
 sg13g2_xnor2_1 _3333_ (.Y(_1385_),
    .A(_1372_),
    .B(_1383_));
 sg13g2_nand2_2 _3334_ (.Y(_1386_),
    .A(_1371_),
    .B(_1385_));
 sg13g2_xnor2_1 _3335_ (.Y(_1387_),
    .A(_1360_),
    .B(_1361_));
 sg13g2_nand2b_1 _3336_ (.Y(_1388_),
    .B(_1387_),
    .A_N(_1386_));
 sg13g2_a21oi_1 _3337_ (.A1(_1380_),
    .A2(_1382_),
    .Y(_1389_),
    .B1(_1384_));
 sg13g2_xnor2_1 _3338_ (.Y(_1390_),
    .A(_1386_),
    .B(_1387_));
 sg13g2_nand2b_1 _3339_ (.Y(_1391_),
    .B(_1390_),
    .A_N(_1389_));
 sg13g2_nand2_1 _3340_ (.Y(_1392_),
    .A(_1388_),
    .B(_1391_));
 sg13g2_xnor2_1 _3341_ (.Y(_1393_),
    .A(_1366_),
    .B(_1367_));
 sg13g2_nand2b_1 _3342_ (.Y(_1394_),
    .B(_1392_),
    .A_N(_1393_));
 sg13g2_xnor2_1 _3343_ (.Y(_1395_),
    .A(_1379_),
    .B(_1377_));
 sg13g2_nor2_2 _3344_ (.A(net1548),
    .B(_0808_),
    .Y(_1396_));
 sg13g2_nand2_1 _3345_ (.Y(_1397_),
    .A(net1628),
    .B(_1213_));
 sg13g2_nand2_2 _3346_ (.Y(_1398_),
    .A(_1103_),
    .B(net1628));
 sg13g2_or2_1 _3347_ (.X(_1399_),
    .B(_1373_),
    .A(_1398_));
 sg13g2_nand2_1 _3348_ (.Y(_1400_),
    .A(_1006_),
    .B(net1568));
 sg13g2_nor2_2 _3349_ (.A(_1400_),
    .B(_1399_),
    .Y(_1401_));
 sg13g2_xor2_1 _3350_ (.B(_1400_),
    .A(_1399_),
    .X(_1402_));
 sg13g2_xor2_1 _3351_ (.B(_1402_),
    .A(_1396_),
    .X(_1403_));
 sg13g2_nand2_2 _3352_ (.Y(_1404_),
    .A(_1395_),
    .B(_1403_));
 sg13g2_xnor2_1 _3353_ (.Y(_1405_),
    .A(_1371_),
    .B(_1385_));
 sg13g2_nor2_1 _3354_ (.A(_1404_),
    .B(_1405_),
    .Y(_1406_));
 sg13g2_a21oi_2 _3355_ (.B1(_1401_),
    .Y(_1407_),
    .A2(_1402_),
    .A1(_1396_));
 sg13g2_xor2_1 _3356_ (.B(_1404_),
    .A(_1405_),
    .X(_1408_));
 sg13g2_nor2b_1 _3357_ (.A(_1407_),
    .B_N(_1408_),
    .Y(_1409_));
 sg13g2_nor2_2 _3358_ (.A(_1406_),
    .B(_1409_),
    .Y(_1410_));
 sg13g2_xnor2_1 _3359_ (.Y(_1411_),
    .A(_1389_),
    .B(_1390_));
 sg13g2_nor2b_1 _3360_ (.A(_1410_),
    .B_N(_1411_),
    .Y(_1412_));
 sg13g2_xnor2_1 _3361_ (.Y(_1413_),
    .A(_1373_),
    .B(_1398_));
 sg13g2_and2_1 _3362_ (.A(_0929_),
    .B(net1568),
    .X(_1414_));
 sg13g2_nor2_1 _3363_ (.A(net625),
    .B(net1548),
    .Y(_1415_));
 sg13g2_nand2_2 _3364_ (.Y(_1416_),
    .A(_1396_),
    .B(_1414_));
 sg13g2_a21o_1 _3365_ (.A2(net1568),
    .A1(_0807_),
    .B1(_1415_),
    .X(_1417_));
 sg13g2_nand2_1 _3366_ (.Y(_1418_),
    .A(_1416_),
    .B(_1417_));
 sg13g2_nor2_1 _3367_ (.A(_1413_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_xor2_1 _3368_ (.B(_1403_),
    .A(_1395_),
    .X(_1420_));
 sg13g2_xnor2_1 _3369_ (.Y(_1421_),
    .A(_1419_),
    .B(_1420_));
 sg13g2_and4_1 _3370_ (.A(_0807_),
    .B(net1568),
    .C(_1415_),
    .D(_1420_),
    .X(_1422_));
 sg13g2_a21oi_1 _3371_ (.A1(_1419_),
    .A2(_1420_),
    .Y(_1423_),
    .B1(_1422_));
 sg13g2_xnor2_1 _3372_ (.Y(_1424_),
    .A(_1407_),
    .B(_1408_));
 sg13g2_nand2b_1 _3373_ (.Y(_1425_),
    .B(_1424_),
    .A_N(_1423_));
 sg13g2_xor2_1 _3374_ (.B(_1418_),
    .A(_1413_),
    .X(_1426_));
 sg13g2_nand2_2 _3375_ (.Y(_1427_),
    .A(_1103_),
    .B(net1568));
 sg13g2_nor2_2 _3376_ (.A(_1104_),
    .B(net1548),
    .Y(_1428_));
 sg13g2_nand2_1 _3377_ (.Y(_1429_),
    .A(_1414_),
    .B(_1428_));
 sg13g2_xnor2_1 _3378_ (.Y(_1430_),
    .A(_1428_),
    .B(_1414_));
 sg13g2_o21ai_1 _3379_ (.B1(_1429_),
    .Y(_1431_),
    .A1(_1397_),
    .A2(_1430_));
 sg13g2_nand2_1 _3380_ (.Y(_1432_),
    .A(_1426_),
    .B(_1431_));
 sg13g2_xor2_1 _3381_ (.B(_1430_),
    .A(_1397_),
    .X(_1433_));
 sg13g2_nand2_2 _3382_ (.Y(_1434_),
    .A(_1213_),
    .B(net1568));
 sg13g2_nor3_2 _3383_ (.A(_1214_),
    .B(net1548),
    .C(_1427_),
    .Y(_1435_));
 sg13g2_nand2_2 _3384_ (.Y(_1436_),
    .A(net682),
    .B(_1435_));
 sg13g2_nor2_1 _3385_ (.A(_1426_),
    .B(_1431_),
    .Y(_1437_));
 sg13g2_xor2_1 _3386_ (.B(_1431_),
    .A(_1426_),
    .X(_1438_));
 sg13g2_o21ai_1 _3387_ (.B1(_1432_),
    .Y(_1439_),
    .A1(_1437_),
    .A2(_1436_));
 sg13g2_xnor2_1 _3388_ (.Y(_1440_),
    .A(_1416_),
    .B(_1421_));
 sg13g2_nand2b_1 _3389_ (.Y(_1441_),
    .B(_1439_),
    .A_N(_1440_));
 sg13g2_nor2b_1 _3390_ (.A(_1424_),
    .B_N(_1423_),
    .Y(_1442_));
 sg13g2_xnor2_1 _3391_ (.Y(_1443_),
    .A(_1423_),
    .B(_1424_));
 sg13g2_o21ai_1 _3392_ (.B1(_1425_),
    .Y(_1444_),
    .A1(_1441_),
    .A2(_1442_));
 sg13g2_xnor2_1 _3393_ (.Y(_1445_),
    .A(_1410_),
    .B(_1411_));
 sg13g2_a21oi_2 _3394_ (.B1(_1412_),
    .Y(_1446_),
    .A2(_1445_),
    .A1(_1444_));
 sg13g2_nor2b_1 _3395_ (.A(_1392_),
    .B_N(_1393_),
    .Y(_1447_));
 sg13g2_xnor2_1 _3396_ (.Y(_1448_),
    .A(_1392_),
    .B(_1393_));
 sg13g2_o21ai_1 _3397_ (.B1(_1394_),
    .Y(_1449_),
    .A1(_1446_),
    .A2(_1447_));
 sg13g2_xor2_1 _3398_ (.B(_1369_),
    .A(_1368_),
    .X(_1450_));
 sg13g2_a21oi_2 _3399_ (.B1(_1370_),
    .Y(_1451_),
    .A2(_1450_),
    .A1(_1449_));
 sg13g2_a221oi_1 _3400_ (.B2(_1450_),
    .C1(_1370_),
    .B1(_1449_),
    .A1(_1342_),
    .Y(_1452_),
    .A2(_1344_));
 sg13g2_nor3_2 _3401_ (.A(_1345_),
    .B(_1295_),
    .C(_1452_),
    .Y(_1453_));
 sg13g2_nor2_2 _3402_ (.A(_1453_),
    .B(_1293_),
    .Y(_1454_));
 sg13g2_or3_1 _3403_ (.A(_1239_),
    .B(_1293_),
    .C(_1453_),
    .X(_1455_));
 sg13g2_and3_1 _3404_ (.X(_1456_),
    .A(_1455_),
    .B(_1238_),
    .C(_1180_));
 sg13g2_nand2_1 _3405_ (.Y(_1457_),
    .A(_1173_),
    .B(_1176_));
 sg13g2_o21ai_1 _3406_ (.B1(_1167_),
    .Y(_1458_),
    .A1(_1164_),
    .A2(_1168_));
 sg13g2_nor2b_1 _3407_ (.A(net1515),
    .B_N(_0899_),
    .Y(_1459_));
 sg13g2_xnor2_1 _3408_ (.Y(_1460_),
    .A(_1165_),
    .B(_1459_));
 sg13g2_nand2b_1 _3409_ (.Y(_1461_),
    .B(_1458_),
    .A_N(_1460_));
 sg13g2_xor2_1 _3410_ (.B(_1458_),
    .A(_1460_),
    .X(_1462_));
 sg13g2_xor2_1 _3411_ (.B(_1462_),
    .A(_1171_),
    .X(_1463_));
 sg13g2_xor2_1 _3412_ (.B(_1463_),
    .A(_1457_),
    .X(_1464_));
 sg13g2_o21ai_1 _3413_ (.B1(_1464_),
    .Y(_1465_),
    .A1(_1456_),
    .A2(_1179_));
 sg13g2_or3_1 _3414_ (.A(_1179_),
    .B(_1456_),
    .C(_1464_),
    .X(_1466_));
 sg13g2_nand2_2 _3415_ (.Y(_1467_),
    .A(_1466_),
    .B(_1465_));
 sg13g2_or2_1 _3416_ (.X(_1468_),
    .B(_0235_),
    .A(_1467_));
 sg13g2_mux4_1 _3417_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ),
    .A0(net128),
    .A1(net55),
    .A2(net9),
    .A3(net70),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ),
    .X(_1469_));
 sg13g2_mux4_1 _3418_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A1(net77),
    .A2(net42),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1470_));
 sg13g2_mux4_1 _3419_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .A1(net43),
    .A2(net17),
    .A3(net78),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ),
    .X(_1471_));
 sg13g2_mux4_1 _3420_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(_1470_),
    .A1(_1471_),
    .A2(_1469_),
    .A3(_0611_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ));
 sg13g2_nand2_1 _3421_ (.Y(_1472_),
    .A(net1638),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ));
 sg13g2_a21oi_1 _3422_ (.A1(_0133_),
    .A2(net1645),
    .Y(_1473_),
    .B1(net1650));
 sg13g2_a22oi_1 _3423_ (.Y(_1474_),
    .B1(_1472_),
    .B2(_1473_),
    .A2(net1650),
    .A1(_0000_));
 sg13g2_a21o_1 _3424_ (.A2(_1238_),
    .A1(_1455_),
    .B1(_1180_),
    .X(_1475_));
 sg13g2_nand2b_1 _3425_ (.Y(_1476_),
    .B(_1475_),
    .A_N(_1456_));
 sg13g2_a221oi_1 _3426_ (.B2(_1473_),
    .C1(_1476_),
    .B1(_1472_),
    .A1(_0000_),
    .Y(_1477_),
    .A2(net1650));
 sg13g2_o21ai_1 _3427_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ),
    .Y(_1478_),
    .A1(_0068_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_a21oi_1 _3428_ (.A1(net76),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ),
    .Y(_1479_),
    .B1(_1478_));
 sg13g2_a21oi_1 _3429_ (.A1(net15),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ),
    .Y(_1480_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_o21ai_1 _3430_ (.B1(_1480_),
    .Y(_1481_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ),
    .A2(net616));
 sg13g2_nand2b_1 _3431_ (.Y(_1482_),
    .B(_1481_),
    .A_N(_1479_));
 sg13g2_inv_1 _3432_ (.Y(_1483_),
    .A(_1482_));
 sg13g2_o21ai_1 _3433_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_1484_),
    .A1(net1687),
    .A2(_0175_));
 sg13g2_a21oi_1 _3434_ (.A1(net1687),
    .A2(net1539),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_mux2_1 _3435_ (.A0(net1635),
    .A1(net1586),
    .S(net1687),
    .X(_1486_));
 sg13g2_o21ai_1 _3436_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .Y(_1487_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .A2(_1486_));
 sg13g2_mux4_1 _3437_ (.S0(net1687),
    .A0(net1598),
    .A1(net1611),
    .A2(net1603),
    .A3(net1623),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1488_));
 sg13g2_o21ai_1 _3438_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ),
    .Y(_1489_),
    .A1(_1485_),
    .A2(_1487_));
 sg13g2_a21oi_1 _3439_ (.A1(_0116_),
    .A2(_1488_),
    .Y(_1490_),
    .B1(_1489_));
 sg13g2_mux4_1 _3440_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .A0(net1516),
    .A1(net2003),
    .A2(net1707),
    .A3(net10),
    .S1(net1687),
    .X(_1491_));
 sg13g2_o21ai_1 _3441_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_1492_),
    .A1(_0086_),
    .A2(net1687));
 sg13g2_a21oi_1 _3442_ (.A1(net64),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .Y(_1493_),
    .B1(_1492_));
 sg13g2_nand2_1 _3443_ (.Y(_1494_),
    .A(net28),
    .B(net1687));
 sg13g2_o21ai_1 _3444_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_0070_),
    .A2(net1687));
 sg13g2_o21ai_1 _3445_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ),
    .Y(_1496_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ),
    .A2(_1495_));
 sg13g2_nor2_1 _3446_ (.A(_1493_),
    .B(_1496_),
    .Y(_1497_));
 sg13g2_a21oi_1 _3447_ (.A1(_0116_),
    .A2(_1491_),
    .Y(_1498_),
    .B1(_1497_));
 sg13g2_a21oi_1 _3448_ (.A1(_0117_),
    .A2(_1498_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .B1(_1490_));
 sg13g2_mux4_1 _3449_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(net126),
    .A1(net7),
    .A2(net33),
    .A3(net84),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1499_));
 sg13g2_mux4_1 _3450_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net14),
    .A2(net1935),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1500_));
 sg13g2_mux4_1 _3451_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ),
    .A0(net145),
    .A1(net48),
    .A2(net6),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1501_));
 sg13g2_mux4_1 _3452_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ),
    .A0(_1500_),
    .A1(_1499_),
    .A2(_1483_),
    .A3(_1501_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ));
 sg13g2_nand2_1 _3453_ (.Y(_1502_),
    .A(net1638),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ));
 sg13g2_a21oi_1 _3454_ (.A1(net1645),
    .A2(_0136_),
    .Y(_1503_),
    .B1(net1650));
 sg13g2_a22oi_1 _3455_ (.Y(_1504_),
    .B1(_1502_),
    .B2(_1503_),
    .A2(_0002_),
    .A1(net1650));
 sg13g2_nand2_1 _3456_ (.Y(_1505_),
    .A(_1238_),
    .B(_1240_));
 sg13g2_xor2_1 _3457_ (.B(_1505_),
    .A(_1454_),
    .X(_1506_));
 sg13g2_nand2_2 _3458_ (.Y(_1507_),
    .A(_1506_),
    .B(_1504_));
 sg13g2_o21ai_1 _3459_ (.B1(_1295_),
    .Y(_1508_),
    .A1(_1345_),
    .A2(_1452_));
 sg13g2_nor2b_2 _3460_ (.A(_1453_),
    .B_N(_1508_),
    .Y(_1509_));
 sg13g2_mux4_1 _3461_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(net138),
    .A1(net7),
    .A2(net68),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_1510_));
 sg13g2_inv_1 _3462_ (.Y(_1511_),
    .A(_1510_));
 sg13g2_mux4_1 _3463_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(net130),
    .A1(net24),
    .A2(net37),
    .A3(net72),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_1512_));
 sg13g2_nand2_1 _3464_ (.Y(_1513_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .B(_1511_));
 sg13g2_o21ai_1 _3465_ (.B1(_1513_),
    .Y(_1514_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_1512_));
 sg13g2_mux2_1 _3466_ (.A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(net18),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .X(_1515_));
 sg13g2_mux4_1 _3467_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(net1597),
    .A1(net1610),
    .A2(net649),
    .A3(net1624),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_1516_));
 sg13g2_mux4_1 _3468_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .A0(net1632),
    .A1(net1585),
    .A2(net1525),
    .A3(net1520),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_1517_));
 sg13g2_nand2b_1 _3469_ (.Y(_1518_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .A_N(_1517_));
 sg13g2_o21ai_1 _3470_ (.B1(_1518_),
    .Y(_1519_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_1516_));
 sg13g2_nor2_1 _3471_ (.A(net28),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_1520_));
 sg13g2_a21oi_1 _3472_ (.A1(_0086_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .Y(_1521_),
    .B1(_1520_));
 sg13g2_nand2b_1 _3473_ (.Y(_1522_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .A_N(net1932));
 sg13g2_o21ai_1 _3474_ (.B1(_1522_),
    .Y(_1523_),
    .A1(net62),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_o21ai_1 _3475_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_1524_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_1521_));
 sg13g2_a21oi_1 _3476_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .A2(_1523_),
    .Y(_1525_),
    .B1(_1524_));
 sg13g2_mux4_1 _3477_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ),
    .A0(net1516),
    .A1(net2003),
    .A2(net1707),
    .A3(net10),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ),
    .X(_1526_));
 sg13g2_nand2b_1 _3478_ (.Y(_1527_),
    .B(_1526_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_nor2_1 _3479_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .B(_1525_),
    .Y(_1528_));
 sg13g2_a22oi_1 _3480_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .B1(_1527_),
    .B2(_1528_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ),
    .A1(_1519_));
 sg13g2_nor2b_1 _3481_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .B_N(net79),
    .Y(_1529_));
 sg13g2_a21oi_1 _3482_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ),
    .A2(net729),
    .Y(_1530_),
    .B1(_1529_));
 sg13g2_a21oi_1 _3483_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .A2(_1530_),
    .Y(_1531_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_o21ai_1 _3484_ (.B1(_1531_),
    .Y(_1532_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ),
    .A2(_1515_));
 sg13g2_a21oi_1 _3485_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0614_),
    .Y(_1533_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_a22oi_1 _3486_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .B1(_1532_),
    .B2(_1533_),
    .A2(_1514_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_o21ai_1 _3487_ (.B1(_0135_),
    .Y(_1534_),
    .A1(net1638),
    .A2(_0005_));
 sg13g2_a21oi_1 _3488_ (.A1(net1638),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .Y(_1535_),
    .B1(_1534_));
 sg13g2_a21o_1 _3489_ (.A2(_0004_),
    .A1(net1650),
    .B1(_1535_),
    .X(_1536_));
 sg13g2_inv_1 _3490_ (.Y(_1537_),
    .A(_1536_));
 sg13g2_and2_1 _3491_ (.A(_1509_),
    .B(_1537_),
    .X(_1538_));
 sg13g2_nand2b_1 _3492_ (.Y(_1539_),
    .B(net1531),
    .A_N(net1669));
 sg13g2_a21oi_1 _3493_ (.A1(net1670),
    .A2(net1536),
    .Y(_1540_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_nand2b_1 _3494_ (.Y(_1541_),
    .B(net1669),
    .A_N(net1552));
 sg13g2_o21ai_1 _3495_ (.B1(_1541_),
    .Y(_1542_),
    .A1(net1669),
    .A2(net1545));
 sg13g2_a221oi_1 _3496_ (.B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .B1(_1542_),
    .A1(_1539_),
    .Y(_1543_),
    .A2(_1540_));
 sg13g2_a21oi_1 _3497_ (.A1(net1669),
    .A2(net1574),
    .Y(_1544_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_o21ai_1 _3498_ (.B1(_1544_),
    .Y(_1545_),
    .A1(net1669),
    .A2(net1555));
 sg13g2_nand2b_1 _3499_ (.Y(_1546_),
    .B(net1581),
    .A_N(net1669));
 sg13g2_nand2_1 _3500_ (.Y(_1547_),
    .A(net1670),
    .B(net1616));
 sg13g2_nand3_1 _3501_ (.B(_1546_),
    .C(_1547_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .Y(_1548_));
 sg13g2_nand3_1 _3502_ (.B(_1545_),
    .C(_1548_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ),
    .Y(_1549_));
 sg13g2_nor2b_1 _3503_ (.A(_1543_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ),
    .Y(_1550_));
 sg13g2_nand2_1 _3504_ (.Y(_1551_),
    .A(net1670),
    .B(_0682_));
 sg13g2_o21ai_1 _3505_ (.B1(_1551_),
    .Y(_1552_),
    .A1(_0416_),
    .A2(net1670));
 sg13g2_o21ai_1 _3506_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .Y(_1553_),
    .A1(_0095_),
    .A2(net1669));
 sg13g2_a21oi_1 _3507_ (.A1(net1705),
    .A2(net1670),
    .Y(_1554_),
    .B1(_1553_));
 sg13g2_nor2_1 _3508_ (.A(_0142_),
    .B(_1554_),
    .Y(_1555_));
 sg13g2_o21ai_1 _3509_ (.B1(_1555_),
    .Y(_1556_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_1552_));
 sg13g2_mux4_1 _3510_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ),
    .A0(net1711),
    .A1(net1926),
    .A2(net121),
    .A3(net97),
    .S1(net1669),
    .X(_1557_));
 sg13g2_a21oi_1 _3511_ (.A1(_0142_),
    .A2(_1557_),
    .Y(_1558_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_a22oi_1 _3512_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .B1(_1558_),
    .B2(_1556_),
    .A2(_1550_),
    .A1(_1549_));
 sg13g2_inv_1 _3513_ (.Y(_1559_),
    .A(net717));
 sg13g2_nand2_1 _3514_ (.Y(_1560_),
    .A(net1671),
    .B(_0682_));
 sg13g2_o21ai_1 _3515_ (.B1(_1560_),
    .Y(_1561_),
    .A1(net1671),
    .A2(_0416_));
 sg13g2_o21ai_1 _3516_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_1562_),
    .A1(_0077_),
    .A2(net1671));
 sg13g2_a21oi_1 _3517_ (.A1(net147),
    .A2(net1671),
    .Y(_1563_),
    .B1(_1562_));
 sg13g2_nor2_1 _3518_ (.A(_0143_),
    .B(_1563_),
    .Y(_1564_));
 sg13g2_o21ai_1 _3519_ (.B1(_1564_),
    .Y(_1565_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_1561_));
 sg13g2_mux4_1 _3520_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .A0(net111),
    .A1(net87),
    .A2(net115),
    .A3(net91),
    .S1(net1671),
    .X(_1566_));
 sg13g2_a21oi_1 _3521_ (.A1(_0143_),
    .A2(_1566_),
    .Y(_1567_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_mux4_1 _3522_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(net1532),
    .A1(net1537),
    .A2(net1546),
    .A3(net1553),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1568_));
 sg13g2_and2_1 _3523_ (.A(_0143_),
    .B(_1568_),
    .X(_1569_));
 sg13g2_o21ai_1 _3524_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_1570_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .A2(net1571));
 sg13g2_a21oi_1 _3525_ (.A1(net1671),
    .A2(net1616),
    .Y(_1571_),
    .B1(_1570_));
 sg13g2_nor2_1 _3526_ (.A(net1671),
    .B(net1558),
    .Y(_1572_));
 sg13g2_a21oi_1 _3527_ (.A1(net1671),
    .A2(net1561),
    .Y(_1573_),
    .B1(_1572_));
 sg13g2_o21ai_1 _3528_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_1574_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_1573_));
 sg13g2_o21ai_1 _3529_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ),
    .Y(_1575_),
    .A1(_1571_),
    .A2(_1574_));
 sg13g2_o21ai_1 _3530_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .Y(_1576_),
    .A1(_1569_),
    .A2(_1575_));
 sg13g2_a21oi_1 _3531_ (.A1(_1565_),
    .A2(_1567_),
    .Y(_1577_),
    .B1(_1576_));
 sg13g2_mux4_1 _3532_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(net1532),
    .A1(net1536),
    .A2(net1546),
    .A3(net1553),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_1578_));
 sg13g2_mux4_1 _3533_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(net1558),
    .A1(net1564),
    .A2(net1574),
    .A3(net1619),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_1579_));
 sg13g2_mux4_1 _3534_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(net708),
    .A1(net147),
    .A2(net38),
    .A3(net1705),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1580_));
 sg13g2_mux4_1 _3535_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(net111),
    .A1(net1928),
    .A2(net115),
    .A3(net91),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_1581_));
 sg13g2_mux4_1 _3536_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(_1581_),
    .A1(_1580_),
    .A2(_1578_),
    .A3(_1579_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ));
 sg13g2_mux4_1 _3537_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net1531),
    .A1(net1537),
    .A2(net1545),
    .A3(net1552),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1582_));
 sg13g2_nand2_1 _3538_ (.Y(_1583_),
    .A(_0140_),
    .B(_1582_));
 sg13g2_a21oi_1 _3539_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(net1574),
    .Y(_1584_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_o21ai_1 _3540_ (.B1(_1584_),
    .Y(_1585_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(net1555));
 sg13g2_nand2b_1 _3541_ (.Y(_1586_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A_N(net1619));
 sg13g2_o21ai_1 _3542_ (.B1(_1586_),
    .Y(_1587_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(net1581));
 sg13g2_a21oi_1 _3543_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .A2(_1587_),
    .Y(_1588_),
    .B1(_0140_));
 sg13g2_a21oi_1 _3544_ (.A1(_1585_),
    .A2(_1588_),
    .Y(_1589_),
    .B1(_0141_));
 sg13g2_mux4_1 _3545_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(_0682_),
    .A1(net44),
    .A2(net147),
    .A3(net1705),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1590_));
 sg13g2_nand2_1 _3546_ (.Y(_1591_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_1590_));
 sg13g2_mux4_1 _3547_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ),
    .A0(net1711),
    .A1(net1926),
    .A2(net121),
    .A3(net97),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1592_));
 sg13g2_a21oi_1 _3548_ (.A1(_0140_),
    .A2(_1592_),
    .Y(_1593_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_a22oi_1 _3549_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .B1(_1591_),
    .B2(_1593_),
    .A2(_1589_),
    .A1(_1583_));
 sg13g2_mux4_1 _3550_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net703),
    .A1(_0682_),
    .A2(net58),
    .A3(net169),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1594_));
 sg13g2_mux4_1 _3551_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .A0(net1713),
    .A1(net1928),
    .A2(net115),
    .A3(net91),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_1595_));
 sg13g2_mux4_1 _3552_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net1560),
    .A1(net1566),
    .A2(net1574),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1596_));
 sg13g2_mux4_1 _3553_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net1533),
    .A1(net635),
    .A2(net1547),
    .A3(net1554),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_1597_));
 sg13g2_mux4_1 _3554_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(_1595_),
    .A1(_1597_),
    .A2(_1594_),
    .A3(_1596_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ));
 sg13g2_a21oi_2 _3555_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_1598_),
    .A2(net720),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_o21ai_1 _3556_ (.B1(_1598_),
    .Y(_1599_),
    .A1(net718),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_o21ai_1 _3557_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_1600_),
    .A1(_0095_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_a21oi_1 _3558_ (.A1(net1705),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .Y(_1601_),
    .B1(_1600_));
 sg13g2_nor2_1 _3559_ (.A(_0138_),
    .B(_1601_),
    .Y(_1602_));
 sg13g2_mux4_1 _3560_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .A0(net1711),
    .A1(net1926),
    .A2(net121),
    .A3(net97),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .X(_1603_));
 sg13g2_a221oi_1 _3561_ (.B2(_0138_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ),
    .B1(_1603_),
    .A1(_1599_),
    .Y(_1604_),
    .A2(_1602_));
 sg13g2_mux4_1 _3562_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net1558),
    .A1(net1574),
    .A2(net1582),
    .A3(net1616),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1605_));
 sg13g2_mux4_1 _3563_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net1531),
    .A1(net1536),
    .A2(net1545),
    .A3(net1552),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1606_));
 sg13g2_nand2_1 _3564_ (.Y(_1607_),
    .A(_0138_),
    .B(_1606_));
 sg13g2_a21oi_1 _3565_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1605_),
    .Y(_1608_),
    .B1(_0139_));
 sg13g2_a21oi_2 _3566_ (.B1(_1604_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .A2(_1608_),
    .A1(_1607_));
 sg13g2_nand2_2 _3567_ (.Y(_1609_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .B(_0137_));
 sg13g2_mux4_1 _3568_ (.S0(_0137_),
    .A0(net725),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1610_));
 sg13g2_a21oi_1 _3569_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .Y(_1611_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_a21oi_1 _3570_ (.A1(_0137_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .Y(_1612_),
    .B1(_1577_));
 sg13g2_a22oi_1 _3571_ (.Y(_1613_),
    .B1(_1612_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ),
    .A2(_1611_),
    .A1(_1609_));
 sg13g2_mux2_1 _3572_ (.A0(_1610_),
    .A1(_1613_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ),
    .X(\Tile_X0Y1_DSP_bot.C9 ));
 sg13g2_o21ai_1 _3573_ (.B1(net1636),
    .Y(_1614_),
    .A1(net1637),
    .A2(_0007_));
 sg13g2_a21oi_2 _3574_ (.B1(_1614_),
    .Y(_1615_),
    .A2(\Tile_X0Y1_DSP_bot.C9 ),
    .A1(net1637));
 sg13g2_a21o_1 _3575_ (.A2(_0006_),
    .A1(net1651),
    .B1(_1615_),
    .X(_1616_));
 sg13g2_xor2_1 _3576_ (.B(_1343_),
    .A(_1342_),
    .X(_1617_));
 sg13g2_xor2_1 _3577_ (.B(_1617_),
    .A(_1451_),
    .X(_1618_));
 sg13g2_nand2b_1 _3578_ (.Y(_1619_),
    .B(_1618_),
    .A_N(_1616_));
 sg13g2_nand2_1 _3579_ (.Y(_1620_),
    .A(net1648),
    .B(_0008_));
 sg13g2_mux2_1 _3580_ (.A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .A1(_0741_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .X(_1621_));
 sg13g2_mux4_1 _3581_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(_0616_),
    .A1(_0723_),
    .A2(net1934),
    .A3(net1704),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1622_));
 sg13g2_nand2_1 _3582_ (.Y(_1623_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ),
    .B(_1622_));
 sg13g2_mux4_1 _3583_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net114),
    .A1(net122),
    .A2(net1925),
    .A3(net98),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1624_));
 sg13g2_a21oi_1 _3584_ (.A1(_0148_),
    .A2(_1624_),
    .Y(_1625_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_a21oi_1 _3585_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(net1567),
    .Y(_1626_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_o21ai_1 _3586_ (.B1(_1626_),
    .Y(_1627_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(net1555));
 sg13g2_nand2b_1 _3587_ (.Y(_1628_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A_N(net1619));
 sg13g2_o21ai_1 _3588_ (.B1(_1628_),
    .Y(_1629_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(net1581));
 sg13g2_a21oi_1 _3589_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_1629_),
    .Y(_1630_),
    .B1(_0148_));
 sg13g2_mux4_1 _3590_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net1532),
    .A1(net1536),
    .A2(net1546),
    .A3(net1553),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1631_));
 sg13g2_nand2_2 _3591_ (.Y(_1632_),
    .A(_0148_),
    .B(_1631_));
 sg13g2_a21oi_1 _3592_ (.A1(_1627_),
    .A2(_1630_),
    .Y(_1633_),
    .B1(_0149_));
 sg13g2_a22oi_1 _3593_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .B1(_1632_),
    .B2(_1633_),
    .A2(_1625_),
    .A1(_1623_));
 sg13g2_mux4_1 _3594_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(_0616_),
    .A1(_0723_),
    .A2(net1934),
    .A3(net1704),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1634_));
 sg13g2_nand2_1 _3595_ (.Y(_1635_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ),
    .B(_1634_));
 sg13g2_mux4_1 _3596_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(net114),
    .A1(net122),
    .A2(net90),
    .A3(net98),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1636_));
 sg13g2_a21oi_1 _3597_ (.A1(_0144_),
    .A2(_1636_),
    .Y(_1637_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_a21oi_1 _3598_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(net1566),
    .Y(_1638_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_o21ai_1 _3599_ (.B1(_1638_),
    .Y(_1639_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0171_));
 sg13g2_nand2b_1 _3600_ (.Y(_1640_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A_N(net1620));
 sg13g2_o21ai_1 _3601_ (.B1(_1640_),
    .Y(_1641_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(net1582));
 sg13g2_a21oi_1 _3602_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1641_),
    .Y(_1642_),
    .B1(_0144_));
 sg13g2_mux4_1 _3603_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(net1532),
    .A1(net1536),
    .A2(net1547),
    .A3(net1554),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1643_));
 sg13g2_nand2_2 _3604_ (.Y(_1644_),
    .A(_0144_),
    .B(_1643_));
 sg13g2_a21oi_1 _3605_ (.A1(_1639_),
    .A2(_1642_),
    .Y(_1645_),
    .B1(_0145_));
 sg13g2_a22oi_1 _3606_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .B1(_1644_),
    .B2(_1645_),
    .A2(_1637_),
    .A1(_1635_));
 sg13g2_nor2b_1 _3607_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .Y(_1646_));
 sg13g2_a21oi_1 _3608_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .Y(_1647_),
    .B1(_1646_));
 sg13g2_o21ai_1 _3609_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .Y(_1648_),
    .A1(_1621_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_a21oi_2 _3610_ (.B1(_1648_),
    .Y(_1649_),
    .A2(_1647_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_mux4_1 _3611_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net1532),
    .A1(net1536),
    .A2(net1546),
    .A3(net1553),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1650_));
 sg13g2_nand2_1 _3612_ (.Y(_1651_),
    .A(_0146_),
    .B(_1650_));
 sg13g2_a21oi_1 _3613_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(net1564),
    .Y(_1652_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_o21ai_1 _3614_ (.B1(_1652_),
    .Y(_1653_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(net1555));
 sg13g2_nand2_1 _3615_ (.Y(_1654_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .B(_0178_));
 sg13g2_o21ai_1 _3616_ (.B1(_1654_),
    .Y(_1655_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(net1581));
 sg13g2_a21oi_1 _3617_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_1655_),
    .Y(_1656_),
    .B1(_0146_));
 sg13g2_a21oi_1 _3618_ (.A1(_1653_),
    .A2(_1656_),
    .Y(_1657_),
    .B1(_0147_));
 sg13g2_mux4_1 _3619_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(_0723_),
    .A1(net148),
    .A2(net1934),
    .A3(net1704),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_1658_));
 sg13g2_nand2_1 _3620_ (.Y(_1659_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_1658_));
 sg13g2_mux4_1 _3621_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net1710),
    .A1(net122),
    .A2(net1925),
    .A3(net98),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_1660_));
 sg13g2_a21oi_1 _3622_ (.A1(_0146_),
    .A2(_1660_),
    .Y(_1661_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_a22oi_1 _3623_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .B1(_1659_),
    .B2(_1661_),
    .A2(_1657_),
    .A1(_1651_));
 sg13g2_nor2b_1 _3624_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .Y(_1662_));
 sg13g2_a21oi_1 _3625_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_nand2b_1 _3626_ (.Y(_1664_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_a21oi_1 _3627_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .Y(_1665_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_a221oi_1 _3628_ (.B2(_1665_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ),
    .B1(_1664_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ),
    .Y(_1666_),
    .A2(_1663_));
 sg13g2_or2_1 _3629_ (.X(\Tile_X0Y1_DSP_bot.C8 ),
    .B(_1666_),
    .A(_1649_));
 sg13g2_nor2_2 _3630_ (.A(net1643),
    .B(\Tile_X0Y1_DSP_bot.C8 ),
    .Y(_1667_));
 sg13g2_a21oi_2 _3631_ (.B1(_1667_),
    .Y(_1668_),
    .A2(_0009_),
    .A1(net1646));
 sg13g2_o21ai_1 _3632_ (.B1(_1620_),
    .Y(_1669_),
    .A1(_1668_),
    .A2(net1648));
 sg13g2_xor2_1 _3633_ (.B(_1449_),
    .A(_1450_),
    .X(_1670_));
 sg13g2_nor2b_1 _3634_ (.A(_1669_),
    .B_N(_1670_),
    .Y(_1671_));
 sg13g2_nand2_1 _3635_ (.Y(_1672_),
    .A(net1651),
    .B(_0010_));
 sg13g2_mux4_1 _3636_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ),
    .A0(net139),
    .A1(net151),
    .A2(net1923),
    .A3(_0741_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_1673_));
 sg13g2_mux4_1 _3637_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(net116),
    .A1(net110),
    .A2(net1936),
    .A3(net152),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ),
    .X(_1674_));
 sg13g2_nor2b_1 _3638_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .B_N(_1674_),
    .Y(_1675_));
 sg13g2_a21oi_1 _3639_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_1673_),
    .Y(_1676_),
    .B1(_1675_));
 sg13g2_nand2_1 _3640_ (.Y(_1677_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ),
    .B(_1676_));
 sg13g2_nand2b_1 _3641_ (.Y(_1678_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ));
 sg13g2_o21ai_1 _3642_ (.B1(_1678_),
    .Y(_1679_),
    .A1(net159),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_nand2b_1 _3643_ (.Y(_1680_),
    .B(net1709),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_a21oi_1 _3644_ (.A1(net99),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ),
    .Y(_1681_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_a221oi_1 _3645_ (.B2(_1681_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .B1(_1680_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ),
    .Y(_1682_),
    .A2(_1679_));
 sg13g2_a21oi_1 _3646_ (.A1(net160),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .Y(_1683_),
    .B1(_0150_));
 sg13g2_o21ai_1 _3647_ (.B1(_1683_),
    .Y(_1684_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .A2(net696));
 sg13g2_a21oi_1 _3648_ (.A1(net100),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ),
    .Y(_1685_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_o21ai_1 _3649_ (.B1(_1685_),
    .Y(_1686_),
    .A1(_0060_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_nand3_1 _3650_ (.B(_1684_),
    .C(_1686_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ),
    .Y(_1687_));
 sg13g2_nand2b_1 _3651_ (.Y(_1688_),
    .B(_1687_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_o21ai_1 _3652_ (.B1(_1677_),
    .Y(_1689_),
    .A1(_1688_),
    .A2(_1682_));
 sg13g2_inv_1 _3653_ (.Y(\Tile_X0Y1_DSP_bot.C7 ),
    .A(_1689_));
 sg13g2_nor2_1 _3654_ (.A(net1646),
    .B(_1689_),
    .Y(_1690_));
 sg13g2_o21ai_1 _3655_ (.B1(net1636),
    .Y(_1691_),
    .A1(net1639),
    .A2(_0011_));
 sg13g2_o21ai_1 _3656_ (.B1(_1672_),
    .Y(_1692_),
    .A1(_1691_),
    .A2(_1690_));
 sg13g2_xnor2_1 _3657_ (.Y(_1693_),
    .A(_1446_),
    .B(_1448_));
 sg13g2_nand2b_1 _3658_ (.Y(_1694_),
    .B(_1693_),
    .A_N(_1692_));
 sg13g2_mux4_1 _3659_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(net140),
    .A1(net96),
    .A2(net43),
    .A3(net156),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_1695_));
 sg13g2_mux4_1 _3660_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ),
    .A0(net1922),
    .A1(net51),
    .A2(net172),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_1696_));
 sg13g2_nand2b_1 _3661_ (.Y(_1697_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A_N(_1696_));
 sg13g2_o21ai_1 _3662_ (.B1(_1697_),
    .Y(_1698_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1695_));
 sg13g2_mux4_1 _3663_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ),
    .A0(net103),
    .A1(net163),
    .A2(net615),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_1699_));
 sg13g2_nand2b_1 _3664_ (.Y(_1700_),
    .B(_1699_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_a21oi_1 _3665_ (.A1(net164),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .Y(_1701_),
    .B1(_0151_));
 sg13g2_o21ai_1 _3666_ (.B1(_1701_),
    .Y(_1702_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .A2(_0594_));
 sg13g2_a21oi_1 _3667_ (.A1(net104),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ),
    .Y(_1703_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_o21ai_1 _3668_ (.B1(_1703_),
    .Y(_1704_),
    .A1(_0083_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_nand3_1 _3669_ (.B(_1702_),
    .C(_1704_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_1705_));
 sg13g2_nor2b_1 _3670_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ),
    .B_N(_1705_),
    .Y(_1706_));
 sg13g2_a22oi_1 _3671_ (.Y(\Tile_X0Y1_DSP_bot.C6 ),
    .B1(_1700_),
    .B2(_1706_),
    .A2(_1698_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_nand2_1 _3672_ (.Y(_1707_),
    .A(net1637),
    .B(\Tile_X0Y1_DSP_bot.C6 ));
 sg13g2_a21oi_1 _3673_ (.A1(net1643),
    .A2(_0152_),
    .Y(_1708_),
    .B1(net1648));
 sg13g2_a22oi_1 _3674_ (.Y(_1709_),
    .B1(_1707_),
    .B2(_1708_),
    .A2(_0012_),
    .A1(net1648));
 sg13g2_inv_1 _3675_ (.Y(_1710_),
    .A(_1709_));
 sg13g2_xnor2_1 _3676_ (.Y(_1711_),
    .A(_1444_),
    .B(_1445_));
 sg13g2_nor2_1 _3677_ (.A(_1710_),
    .B(_1711_),
    .Y(_1712_));
 sg13g2_nand2_1 _3678_ (.Y(_1713_),
    .A(net1647),
    .B(_0014_));
 sg13g2_mux4_1 _3679_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(net118),
    .A1(net94),
    .A2(net58),
    .A3(net154),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_1714_));
 sg13g2_mux4_1 _3680_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ),
    .A0(net133),
    .A1(net153),
    .A2(net60),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_1715_));
 sg13g2_nand2b_1 _3681_ (.Y(_1716_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .A_N(_1715_));
 sg13g2_o21ai_1 _3682_ (.B1(_1716_),
    .Y(_1717_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_1714_));
 sg13g2_nor2b_1 _3683_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .B_N(net161),
    .Y(_1718_));
 sg13g2_a21oi_1 _3684_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .Y(_1719_),
    .B1(_1718_));
 sg13g2_nand2_1 _3685_ (.Y(_1720_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ),
    .B(_1719_));
 sg13g2_nand2_1 _3686_ (.Y(_1721_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ),
    .B(net715));
 sg13g2_a21oi_1 _3687_ (.A1(net125),
    .A2(_0153_),
    .Y(_1722_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_a21oi_1 _3688_ (.A1(_1721_),
    .A2(_1722_),
    .Y(_1723_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_mux4_1 _3689_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(net126),
    .A1(net102),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(net162),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_1724_));
 sg13g2_a221oi_1 _3690_ (.B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .B1(_1724_),
    .A1(_1720_),
    .Y(_1725_),
    .A2(_1723_));
 sg13g2_a21oi_2 _3691_ (.B1(_1725_),
    .Y(\Tile_X0Y1_DSP_bot.C5 ),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ),
    .A1(_1717_));
 sg13g2_nor2_2 _3692_ (.A(net1643),
    .B(\Tile_X0Y1_DSP_bot.C5 ),
    .Y(_1726_));
 sg13g2_a21oi_2 _3693_ (.B1(_1726_),
    .Y(_1727_),
    .A2(_0015_),
    .A1(net1643));
 sg13g2_o21ai_1 _3694_ (.B1(_1713_),
    .Y(_1728_),
    .A1(_1727_),
    .A2(net1647));
 sg13g2_inv_4 _3695_ (.A(_1728_),
    .Y(_1729_));
 sg13g2_xnor2_1 _3696_ (.Y(_1730_),
    .A(_1441_),
    .B(_1443_));
 sg13g2_nand2_2 _3697_ (.Y(_1731_),
    .A(_1729_),
    .B(_1730_));
 sg13g2_xor2_1 _3698_ (.B(_1440_),
    .A(_1439_),
    .X(_1732_));
 sg13g2_mux4_1 _3699_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(net134),
    .A1(net53),
    .A2(net107),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_1733_));
 sg13g2_mux4_1 _3700_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(net122),
    .A1(net98),
    .A2(net1934),
    .A3(net169),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ),
    .X(_1734_));
 sg13g2_mux4_1 _3701_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ),
    .A0(net1707),
    .A1(net105),
    .A2(net619),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_1735_));
 sg13g2_mux4_1 _3702_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(net1706),
    .A1(net106),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .A3(net166),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_1736_));
 sg13g2_mux4_1 _3703_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(_1735_),
    .A1(_1736_),
    .A2(_1734_),
    .A3(_1733_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Tile_X0Y1_DSP_bot.C4 ));
 sg13g2_o21ai_1 _3704_ (.B1(net1636),
    .Y(_1737_),
    .A1(net1639),
    .A2(_0017_));
 sg13g2_a21oi_1 _3705_ (.A1(net1637),
    .A2(\Tile_X0Y1_DSP_bot.C4 ),
    .Y(_1738_),
    .B1(_1737_));
 sg13g2_a21o_1 _3706_ (.A2(_0016_),
    .A1(net1648),
    .B1(_1738_),
    .X(_1739_));
 sg13g2_nor2_1 _3707_ (.A(_1732_),
    .B(_1739_),
    .Y(_1740_));
 sg13g2_mux4_1 _3708_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ),
    .A0(net99),
    .A1(net159),
    .A2(net642),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_1741_));
 sg13g2_mux4_1 _3709_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(net124),
    .A1(net100),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A3(net160),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ),
    .X(_1742_));
 sg13g2_mux4_1 _3710_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(net110),
    .A1(net170),
    .A2(net50),
    .A3(_0323_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_1743_));
 sg13g2_mux4_1 _3711_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(net141),
    .A1(net92),
    .A2(net1936),
    .A3(net152),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_1744_));
 sg13g2_mux4_1 _3712_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(_1741_),
    .A1(_1742_),
    .A2(_1744_),
    .A3(_1743_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Tile_X0Y1_DSP_bot.C3 ));
 sg13g2_o21ai_1 _3713_ (.B1(net1636),
    .Y(_1745_),
    .A1(net1637),
    .A2(_0019_));
 sg13g2_a21oi_2 _3714_ (.B1(_1745_),
    .Y(_1746_),
    .A2(\Tile_X0Y1_DSP_bot.C3 ),
    .A1(net1637));
 sg13g2_a21o_1 _3715_ (.A2(_0018_),
    .A1(net1648),
    .B1(_1746_),
    .X(_1747_));
 sg13g2_xnor2_1 _3716_ (.Y(_1748_),
    .A(_1436_),
    .B(_1438_));
 sg13g2_inv_2 _3717_ (.Y(_1749_),
    .A(_1748_));
 sg13g2_nand2_1 _3718_ (.Y(_1750_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .B(_0362_));
 sg13g2_mux4_1 _3719_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(net120),
    .A1(net96),
    .A2(net59),
    .A3(net156),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_1751_));
 sg13g2_nand2b_1 _3720_ (.Y(_1752_),
    .B(_1751_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_nand3_1 _3721_ (.B(_1750_),
    .C(_1752_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ),
    .Y(_1753_));
 sg13g2_nand2_1 _3722_ (.Y(_1754_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .B(_0867_));
 sg13g2_nor2_1 _3723_ (.A(net1708),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .Y(_1755_));
 sg13g2_nor2_1 _3724_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .B(_1755_),
    .Y(_1756_));
 sg13g2_mux2_1 _3725_ (.A0(net163),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1757_));
 sg13g2_a22oi_1 _3726_ (.Y(_1758_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ),
    .B2(_1757_),
    .A2(_1756_),
    .A1(_1754_));
 sg13g2_inv_4 _3727_ (.A(_1758_),
    .Y(_1759_));
 sg13g2_mux4_1 _3728_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(net128),
    .A1(net104),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .A3(net164),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_1760_));
 sg13g2_a21oi_1 _3729_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_1760_),
    .Y(_1761_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_o21ai_1 _3730_ (.B1(_1761_),
    .Y(_1762_),
    .A1(_1758_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_nand2_2 _3731_ (.Y(_1763_),
    .A(_1762_),
    .B(_1753_));
 sg13g2_inv_2 _3732_ (.Y(\Tile_X0Y1_DSP_bot.C2 ),
    .A(_1763_));
 sg13g2_nand2_2 _3733_ (.Y(_1764_),
    .A(net1637),
    .B(\Tile_X0Y1_DSP_bot.C2 ));
 sg13g2_a21oi_1 _3734_ (.A1(net1643),
    .A2(_0154_),
    .Y(_1765_),
    .B1(net1647));
 sg13g2_a22oi_1 _3735_ (.Y(_1766_),
    .B1(_1764_),
    .B2(_1765_),
    .A2(_0020_),
    .A1(net1647));
 sg13g2_xnor2_1 _3736_ (.Y(_1767_),
    .A(net685),
    .B(_1435_));
 sg13g2_a221oi_1 _3737_ (.B2(_1765_),
    .C1(_1767_),
    .B1(_1764_),
    .A1(net1647),
    .Y(_1768_),
    .A2(_0020_));
 sg13g2_nand2_1 _3738_ (.Y(_1769_),
    .A(net1647),
    .B(_0022_));
 sg13g2_mux4_1 _3739_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ),
    .A0(net141),
    .A1(net52),
    .A2(net93),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1770_));
 sg13g2_nor2b_1 _3740_ (.A(_1770_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .Y(_1771_));
 sg13g2_mux4_1 _3741_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(net118),
    .A1(net94),
    .A2(net41),
    .A3(net170),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1772_));
 sg13g2_o21ai_1 _3742_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ),
    .Y(_1773_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1772_));
 sg13g2_mux4_1 _3743_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(net125),
    .A1(net101),
    .A2(net715),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ),
    .X(_1774_));
 sg13g2_nand2b_1 _3744_ (.Y(_1775_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .A_N(net162));
 sg13g2_o21ai_1 _3745_ (.B1(_1775_),
    .Y(_1776_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ));
 sg13g2_nand2_1 _3746_ (.Y(_1777_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .B(_1776_));
 sg13g2_nand2_1 _3747_ (.Y(_1778_),
    .A(net102),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_o21ai_1 _3748_ (.B1(_1778_),
    .Y(_1779_),
    .A1(_0074_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_o21ai_1 _3749_ (.B1(_1777_),
    .Y(_1780_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ),
    .A2(_1779_));
 sg13g2_a21oi_1 _3750_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_1780_),
    .Y(_1781_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_o21ai_1 _3751_ (.B1(_1781_),
    .Y(_1782_),
    .A1(_1774_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_o21ai_1 _3752_ (.B1(_1782_),
    .Y(\Tile_X0Y1_DSP_bot.C1 ),
    .A1(_1771_),
    .A2(_1773_));
 sg13g2_nor2_2 _3753_ (.A(net1643),
    .B(\Tile_X0Y1_DSP_bot.C1 ),
    .Y(_1783_));
 sg13g2_a21oi_2 _3754_ (.B1(_1783_),
    .Y(_1784_),
    .A2(_0023_),
    .A1(net1643));
 sg13g2_o21ai_1 _3755_ (.B1(_1769_),
    .Y(_1785_),
    .A1(_1784_),
    .A2(net1647));
 sg13g2_o21ai_1 _3756_ (.B1(_1427_),
    .Y(_1786_),
    .A1(_1214_),
    .A2(net1548));
 sg13g2_nand2b_1 _3757_ (.Y(_1787_),
    .B(_1786_),
    .A_N(_1435_));
 sg13g2_nor2_1 _3758_ (.A(_1785_),
    .B(_1787_),
    .Y(_1788_));
 sg13g2_nand2_1 _3759_ (.Y(_1789_),
    .A(net1647),
    .B(net745));
 sg13g2_mux4_1 _3760_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(net134),
    .A1(net94),
    .A2(net154),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_1790_));
 sg13g2_nand2_1 _3761_ (.Y(_1791_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .B(_1790_));
 sg13g2_mux4_1 _3762_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(net122),
    .A1(net109),
    .A2(net1934),
    .A3(net158),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_1792_));
 sg13g2_nand2b_1 _3763_ (.Y(_1793_),
    .B(_1792_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_nand3_1 _3764_ (.B(_1791_),
    .C(_1793_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_1794_));
 sg13g2_nor2b_1 _3765_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .B_N(net165),
    .Y(_1795_));
 sg13g2_a21oi_2 _3766_ (.B1(_1795_),
    .Y(_1796_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ));
 sg13g2_nand2b_1 _3767_ (.Y(_1797_),
    .B(net1707),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_a21oi_1 _3768_ (.A1(net105),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ),
    .Y(_1798_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_a221oi_1 _3769_ (.B2(_1798_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .B1(_1797_),
    .A1(_1796_),
    .Y(_1799_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_a21o_1 _3770_ (.A2(_0348_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_1800_));
 sg13g2_o21ai_1 _3771_ (.B1(_1794_),
    .Y(_1801_),
    .A1(_1799_),
    .A2(_1800_));
 sg13g2_inv_1 _3772_ (.Y(\Tile_X0Y1_DSP_bot.C0 ),
    .A(net704));
 sg13g2_nor2_2 _3773_ (.A(net1643),
    .B(_1801_),
    .Y(_1802_));
 sg13g2_o21ai_1 _3774_ (.B1(net1636),
    .Y(_1803_),
    .A1(net1637),
    .A2(_0025_));
 sg13g2_o21ai_1 _3775_ (.B1(_1789_),
    .Y(_1804_),
    .A1(_1803_),
    .A2(_1802_));
 sg13g2_nor2_2 _3776_ (.A(net686),
    .B(_1434_),
    .Y(_1805_));
 sg13g2_xor2_1 _3777_ (.B(_1785_),
    .A(_1787_),
    .X(_1806_));
 sg13g2_a21oi_2 _3778_ (.B1(_1788_),
    .Y(_1807_),
    .A2(_1805_),
    .A1(_1806_));
 sg13g2_xnor2_1 _3779_ (.Y(_1808_),
    .A(_1767_),
    .B(_1766_));
 sg13g2_nor2b_1 _3780_ (.A(_1807_),
    .B_N(_1808_),
    .Y(_1809_));
 sg13g2_nor2_2 _3781_ (.A(_1768_),
    .B(_1809_),
    .Y(_1810_));
 sg13g2_xnor2_1 _3782_ (.Y(_1811_),
    .A(_1747_),
    .B(_1748_));
 sg13g2_nand2b_1 _3783_ (.Y(_1812_),
    .B(_1811_),
    .A_N(_1810_));
 sg13g2_o21ai_1 _3784_ (.B1(_1812_),
    .Y(_1813_),
    .A1(_1747_),
    .A2(_1749_));
 sg13g2_xor2_1 _3785_ (.B(_1739_),
    .A(_1732_),
    .X(_1814_));
 sg13g2_a21oi_2 _3786_ (.B1(_1740_),
    .Y(_1815_),
    .A2(_1813_),
    .A1(_1814_));
 sg13g2_nor2_1 _3787_ (.A(_1729_),
    .B(_1730_),
    .Y(_1816_));
 sg13g2_xnor2_1 _3788_ (.Y(_1817_),
    .A(_1728_),
    .B(_1730_));
 sg13g2_o21ai_1 _3789_ (.B1(_1731_),
    .Y(_1818_),
    .A1(_1815_),
    .A2(_1816_));
 sg13g2_xnor2_1 _3790_ (.Y(_1819_),
    .A(_1709_),
    .B(_1711_));
 sg13g2_a21oi_2 _3791_ (.B1(_1712_),
    .Y(_1820_),
    .A2(_1818_),
    .A1(_1819_));
 sg13g2_xor2_1 _3792_ (.B(_1692_),
    .A(_1693_),
    .X(_1821_));
 sg13g2_o21ai_1 _3793_ (.B1(_1694_),
    .Y(_1822_),
    .A1(_1821_),
    .A2(_1820_));
 sg13g2_xnor2_1 _3794_ (.Y(_1823_),
    .A(_1669_),
    .B(_1670_));
 sg13g2_a21oi_2 _3795_ (.B1(_1671_),
    .Y(_1824_),
    .A2(_1823_),
    .A1(_1822_));
 sg13g2_xor2_1 _3796_ (.B(_1616_),
    .A(_1618_),
    .X(_1825_));
 sg13g2_o21ai_1 _3797_ (.B1(_1619_),
    .Y(_1826_),
    .A1(_1825_),
    .A2(_1824_));
 sg13g2_xnor2_1 _3798_ (.Y(_1827_),
    .A(_1536_),
    .B(_1509_));
 sg13g2_a21oi_2 _3799_ (.B1(_1538_),
    .Y(_1828_),
    .A2(_1826_),
    .A1(_1827_));
 sg13g2_xnor2_1 _3800_ (.Y(_1829_),
    .A(_1504_),
    .B(_1506_));
 sg13g2_o21ai_1 _3801_ (.B1(_1507_),
    .Y(_1830_),
    .A1(_1829_),
    .A2(_1828_));
 sg13g2_xnor2_1 _3802_ (.Y(_1831_),
    .A(_1474_),
    .B(_1476_));
 sg13g2_a21oi_2 _3803_ (.B1(_1477_),
    .Y(_1832_),
    .A2(_1831_),
    .A1(_1830_));
 sg13g2_and2_1 _3804_ (.A(_0235_),
    .B(_1467_),
    .X(_1833_));
 sg13g2_xor2_1 _3805_ (.B(_1467_),
    .A(_0235_),
    .X(_1834_));
 sg13g2_o21ai_1 _3806_ (.B1(_1468_),
    .Y(_1835_),
    .A1(_1832_),
    .A2(_1833_));
 sg13g2_o21ai_1 _3807_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_1836_),
    .A1(_0445_),
    .A2(_0456_));
 sg13g2_o21ai_1 _3808_ (.B1(_1836_),
    .Y(_1837_),
    .A1(net49),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_mux2_1 _3809_ (.A0(net138),
    .A1(net22),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_1838_));
 sg13g2_o21ai_1 _3810_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_1839_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_1838_));
 sg13g2_a21oi_1 _3811_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_1837_),
    .Y(_1840_),
    .B1(_1839_));
 sg13g2_mux4_1 _3812_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ),
    .A0(net1706),
    .A1(net37),
    .A2(net11),
    .A3(net83),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_1841_));
 sg13g2_nand2b_1 _3813_ (.Y(_1842_),
    .B(_1841_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_nor2b_1 _3814_ (.A(_1840_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_1843_));
 sg13g2_mux4_1 _3815_ (.S0(net1678),
    .A0(net1600),
    .A1(net1612),
    .A2(net1605),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_1844_));
 sg13g2_inv_1 _3816_ (.Y(_1845_),
    .A(_1844_));
 sg13g2_mux4_1 _3817_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A0(net1634),
    .A1(net1523),
    .A2(net1593),
    .A3(net1540),
    .S1(net1678),
    .X(_1846_));
 sg13g2_o21ai_1 _3818_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .Y(_1847_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_1845_));
 sg13g2_a21oi_1 _3819_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_1846_),
    .Y(_1848_),
    .B1(_1847_));
 sg13g2_a21oi_1 _3820_ (.A1(net1706),
    .A2(net1678),
    .Y(_1849_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_o21ai_1 _3821_ (.B1(_1849_),
    .Y(_1850_),
    .A1(net1678),
    .A2(net622));
 sg13g2_nor2b_1 _3822_ (.A(net1678),
    .B_N(net2001),
    .Y(_1851_));
 sg13g2_a21oi_1 _3823_ (.A1(net1678),
    .A2(net11),
    .Y(_1852_),
    .B1(_1851_));
 sg13g2_a21oi_1 _3824_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_1852_),
    .Y(_1853_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_a21oi_1 _3825_ (.A1(net37),
    .A2(net1678),
    .Y(_1854_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_o21ai_1 _3826_ (.B1(_1854_),
    .Y(_1855_),
    .A1(_0090_),
    .A2(net1678));
 sg13g2_nand2b_1 _3827_ (.Y(_1856_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .A_N(net1930));
 sg13g2_o21ai_1 _3828_ (.B1(_1856_),
    .Y(_1857_),
    .A1(net1933),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_a21oi_1 _3829_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_1857_),
    .Y(_1858_),
    .B1(_0118_));
 sg13g2_a221oi_1 _3830_ (.B2(_1858_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ),
    .B1(_1855_),
    .A1(_1850_),
    .Y(_1859_),
    .A2(_1853_));
 sg13g2_nor2_2 _3831_ (.A(_1848_),
    .B(_1859_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ));
 sg13g2_mux4_1 _3832_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .A1(net18),
    .A2(net44),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ),
    .X(_1860_));
 sg13g2_nand2b_1 _3833_ (.Y(_1861_),
    .B(_1860_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_mux4_1 _3834_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ),
    .A0(net724),
    .A1(net1934),
    .A2(net19),
    .A3(net80),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_1862_));
 sg13g2_a21oi_1 _3835_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1862_),
    .Y(_1863_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_a22oi_1 _3836_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .B1(_1861_),
    .B2(_1863_),
    .A2(_1843_),
    .A1(_1842_));
 sg13g2_o21ai_1 _3837_ (.B1(net1636),
    .Y(_1864_),
    .A1(net1639),
    .A2(_0029_));
 sg13g2_a21oi_1 _3838_ (.A1(net1638),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .Y(_1865_),
    .B1(_1864_));
 sg13g2_a21oi_1 _3839_ (.A1(net1649),
    .A2(_0028_),
    .Y(_1866_),
    .B1(_1865_));
 sg13g2_inv_1 _3840_ (.Y(_1867_),
    .A(_1866_));
 sg13g2_nand2b_1 _3841_ (.Y(_1868_),
    .B(_1463_),
    .A_N(_1176_));
 sg13g2_nor2_2 _3842_ (.A(_1173_),
    .B(net697),
    .Y(_1869_));
 sg13g2_nor2_2 _3843_ (.A(net1515),
    .B(_0848_),
    .Y(_1870_));
 sg13g2_nand2_2 _3844_ (.Y(_1871_),
    .A(_1870_),
    .B(_1166_));
 sg13g2_o21ai_1 _3845_ (.B1(_1461_),
    .Y(_1872_),
    .A1(_1462_),
    .A2(_1171_));
 sg13g2_xor2_1 _3846_ (.B(_1872_),
    .A(_1871_),
    .X(_1873_));
 sg13g2_nor2b_1 _3847_ (.A(_1873_),
    .B_N(_1869_),
    .Y(_1874_));
 sg13g2_xor2_1 _3848_ (.B(_1869_),
    .A(_1873_),
    .X(_1875_));
 sg13g2_a21oi_2 _3849_ (.B1(_1875_),
    .Y(_1876_),
    .A2(_1868_),
    .A1(_1465_));
 sg13g2_nand3_1 _3850_ (.B(_1868_),
    .C(_1875_),
    .A(_1465_),
    .Y(_1877_));
 sg13g2_nand2b_1 _3851_ (.Y(_1878_),
    .B(_1877_),
    .A_N(_1876_));
 sg13g2_nor2_2 _3852_ (.A(_1878_),
    .B(_1867_),
    .Y(_1879_));
 sg13g2_xnor2_1 _3853_ (.Y(_1880_),
    .A(_1866_),
    .B(_1878_));
 sg13g2_xnor2_1 _3854_ (.Y(_1881_),
    .A(_1835_),
    .B(_1880_));
 sg13g2_nand2_1 _3855_ (.Y(_1882_),
    .A(net1655),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ));
 sg13g2_o21ai_1 _3856_ (.B1(_1882_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .A1(net1655),
    .A2(_1881_));
 sg13g2_xnor2_1 _3857_ (.Y(_1883_),
    .A(_1808_),
    .B(_1807_));
 sg13g2_mux2_1 _3858_ (.A0(_1883_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ),
    .S(net1652),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ));
 sg13g2_xnor2_1 _3859_ (.Y(_1884_),
    .A(_1434_),
    .B(net644));
 sg13g2_nand2_1 _3860_ (.Y(_1885_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ),
    .B(net1652));
 sg13g2_o21ai_1 _3861_ (.B1(_1885_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .A1(net1652),
    .A2(_1884_));
 sg13g2_xnor2_1 _3862_ (.Y(_1886_),
    .A(_1813_),
    .B(_1814_));
 sg13g2_nand2_1 _3863_ (.Y(_1887_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ),
    .B(net1653));
 sg13g2_o21ai_1 _3864_ (.B1(_1887_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .A1(_1886_),
    .A2(net1652));
 sg13g2_xnor2_1 _3865_ (.Y(_1888_),
    .A(_1811_),
    .B(_1810_));
 sg13g2_mux2_2 _3866_ (.A0(_1888_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ),
    .S(net1652),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ));
 sg13g2_xnor2_1 _3867_ (.Y(_1889_),
    .A(_1815_),
    .B(_1817_));
 sg13g2_mux2_1 _3868_ (.A0(_1889_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ),
    .S(net1652),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ));
 sg13g2_xnor2_1 _3869_ (.Y(_1890_),
    .A(_1818_),
    .B(_1819_));
 sg13g2_nand2_1 _3870_ (.Y(_1891_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ),
    .B(net1653));
 sg13g2_o21ai_1 _3871_ (.B1(_1891_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .A1(net1653),
    .A2(_1890_));
 sg13g2_xor2_1 _3872_ (.B(_1820_),
    .A(_1821_),
    .X(_1892_));
 sg13g2_mux2_1 _3873_ (.A0(_1892_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ),
    .S(net1654),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ));
 sg13g2_xnor2_1 _3874_ (.Y(_1893_),
    .A(_1824_),
    .B(_1825_));
 sg13g2_nand2_1 _3875_ (.Y(_1894_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ),
    .B(net1654));
 sg13g2_o21ai_1 _3876_ (.B1(_1894_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .A1(net1654),
    .A2(_1893_));
 sg13g2_mux4_1 _3877_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ),
    .A0(net1558),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .A2(net1517),
    .A3(_1673_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ));
 sg13g2_xnor2_1 _3878_ (.Y(_1895_),
    .A(_1826_),
    .B(_1827_));
 sg13g2_nand2_1 _3879_ (.Y(_1896_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ),
    .B(net1656));
 sg13g2_o21ai_1 _3880_ (.B1(_1896_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .A1(_1895_),
    .A2(net1656));
 sg13g2_xor2_1 _3881_ (.B(_1829_),
    .A(_1828_),
    .X(_1897_));
 sg13g2_mux2_1 _3882_ (.A0(_1897_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ),
    .S(net1656),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ));
 sg13g2_xnor2_1 _3883_ (.Y(_1898_),
    .A(_1830_),
    .B(_1831_));
 sg13g2_nand2_1 _3884_ (.Y(_1899_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ),
    .B(net1656));
 sg13g2_o21ai_1 _3885_ (.B1(_1899_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .A1(_1898_),
    .A2(net1656));
 sg13g2_a21oi_2 _3886_ (.B1(_1879_),
    .Y(_1900_),
    .A2(_1880_),
    .A1(_1835_));
 sg13g2_nand2b_1 _3887_ (.Y(_1901_),
    .B(_1166_),
    .A_N(_1872_));
 sg13g2_and2_1 _3888_ (.A(_1870_),
    .B(_1901_),
    .X(_1902_));
 sg13g2_nor3_2 _3889_ (.A(_1902_),
    .B(_1876_),
    .C(_1874_),
    .Y(_1903_));
 sg13g2_nand2_1 _3890_ (.Y(_1904_),
    .A(net1649),
    .B(_0030_));
 sg13g2_mux4_1 _3891_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(net1599),
    .A1(net1612),
    .A2(net1605),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_1905_));
 sg13g2_inv_1 _3892_ (.Y(_1906_),
    .A(_1905_));
 sg13g2_mux4_1 _3893_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .A0(net1634),
    .A1(net1523),
    .A2(net1593),
    .A3(net1519),
    .S1(net2005),
    .X(_1907_));
 sg13g2_o21ai_1 _3894_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_1908_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1906_));
 sg13g2_a21oi_1 _3895_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_1907_),
    .Y(_1909_),
    .B1(_1908_));
 sg13g2_a21oi_1 _3896_ (.A1(net1706),
    .A2(net2005),
    .Y(_1910_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_o21ai_1 _3897_ (.B1(_1910_),
    .Y(_1911_),
    .A1(_0597_),
    .A2(net2005));
 sg13g2_nor2b_1 _3898_ (.A(net2005),
    .B_N(net2001),
    .Y(_1912_));
 sg13g2_a21oi_1 _3899_ (.A1(net11),
    .A2(net2005),
    .Y(_1913_),
    .B1(_1912_));
 sg13g2_a21oi_1 _3900_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1913_),
    .Y(_1914_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_a21oi_1 _3901_ (.A1(net29),
    .A2(net2005),
    .Y(_1915_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_o21ai_1 _3902_ (.B1(_1915_),
    .Y(_1916_),
    .A1(_0091_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_nand2b_1 _3903_ (.Y(_1917_),
    .B(net2005),
    .A_N(net1930));
 sg13g2_o21ai_1 _3904_ (.B1(_1917_),
    .Y(_1918_),
    .A1(net37),
    .A2(net2005));
 sg13g2_a21oi_1 _3905_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_1918_),
    .Y(_1919_),
    .B1(_0119_));
 sg13g2_a221oi_1 _3906_ (.B2(_1919_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ),
    .B1(_1916_),
    .A1(_1914_),
    .Y(_1920_),
    .A2(_1911_));
 sg13g2_nor2_2 _3907_ (.A(_1920_),
    .B(_1909_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ));
 sg13g2_mux4_1 _3908_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A1(net75),
    .A2(net1935),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_1921_));
 sg13g2_mux4_1 _3909_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(net126),
    .A1(net7),
    .A2(net54),
    .A3(net68),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_1922_));
 sg13g2_mux4_1 _3910_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ),
    .A0(net137),
    .A1(net56),
    .A2(net67),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_1923_));
 sg13g2_mux4_1 _3911_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ),
    .A0(_1921_),
    .A1(_1922_),
    .A2(net1576),
    .A3(_1923_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ));
 sg13g2_nor2_2 _3912_ (.A(net1645),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .Y(_1924_));
 sg13g2_a21oi_2 _3913_ (.B1(_1924_),
    .Y(_1925_),
    .A2(_0031_),
    .A1(net1644));
 sg13g2_o21ai_1 _3914_ (.B1(_1904_),
    .Y(_1926_),
    .A1(net1649),
    .A2(_1925_));
 sg13g2_and2_1 _3915_ (.A(_1903_),
    .B(_1926_),
    .X(_1927_));
 sg13g2_or2_1 _3916_ (.X(_1928_),
    .B(_1926_),
    .A(_1903_));
 sg13g2_nor2b_1 _3917_ (.A(_1927_),
    .B_N(_1928_),
    .Y(_1929_));
 sg13g2_xnor2_1 _3918_ (.Y(_1930_),
    .A(_1929_),
    .B(_1900_));
 sg13g2_mux2_2 _3919_ (.A0(_1930_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ),
    .S(net1655),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ));
 sg13g2_nand2b_2 _3920_ (.Y(_1931_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ),
    .A_N(_1903_));
 sg13g2_inv_1 _3921_ (.Y(_1932_),
    .A(_1931_));
 sg13g2_nand2_1 _3922_ (.Y(_1933_),
    .A(net1649),
    .B(_0032_));
 sg13g2_mux4_1 _3923_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ),
    .A0(net21),
    .A1(net47),
    .A2(net86),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_1934_));
 sg13g2_mux4_1 _3924_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ),
    .A0(net144),
    .A1(net35),
    .A2(net9),
    .A3(net70),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ),
    .X(_1935_));
 sg13g2_nand2b_1 _3925_ (.Y(_1936_),
    .B(_0121_),
    .A_N(_1935_));
 sg13g2_o21ai_1 _3926_ (.B1(_1936_),
    .Y(_1937_),
    .A1(_0121_),
    .A2(_1934_));
 sg13g2_a21oi_1 _3927_ (.A1(net17),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .Y(_1938_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_o21ai_1 _3928_ (.B1(_1938_),
    .Y(_1939_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .A2(_0697_));
 sg13g2_o21ai_1 _3929_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ),
    .Y(_1940_),
    .A1(_0099_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_a21oi_1 _3930_ (.A1(net78),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ),
    .Y(_1941_),
    .B1(_1940_));
 sg13g2_nor2_1 _3931_ (.A(_0121_),
    .B(_1941_),
    .Y(_1942_));
 sg13g2_mux4_1 _3932_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ),
    .A0(net16),
    .A1(net77),
    .A2(net42),
    .A3(net618),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ),
    .X(_1943_));
 sg13g2_a221oi_1 _3933_ (.B2(_0121_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .B1(_1943_),
    .A1(_1939_),
    .Y(_1944_),
    .A2(_1942_));
 sg13g2_a21oi_1 _3934_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_1937_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .B1(_1944_));
 sg13g2_nor2_1 _3935_ (.A(net1644),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .Y(_1945_));
 sg13g2_a21oi_1 _3936_ (.A1(net1644),
    .A2(_0033_),
    .Y(_1946_),
    .B1(_1945_));
 sg13g2_o21ai_1 _3937_ (.B1(_1933_),
    .Y(_1947_),
    .A1(_1946_),
    .A2(net1649));
 sg13g2_nor2_2 _3938_ (.A(_1931_),
    .B(_1947_),
    .Y(_1948_));
 sg13g2_nand2_2 _3939_ (.Y(_1949_),
    .A(_1931_),
    .B(_1947_));
 sg13g2_nand2b_1 _3940_ (.Y(_1950_),
    .B(_1949_),
    .A_N(_1948_));
 sg13g2_a21oi_2 _3941_ (.B1(_1927_),
    .Y(_1951_),
    .A2(_1900_),
    .A1(_1928_));
 sg13g2_xnor2_1 _3942_ (.Y(_1952_),
    .A(_1950_),
    .B(_1951_));
 sg13g2_mux2_1 _3943_ (.A0(_1952_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ),
    .S(net1656),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ));
 sg13g2_a21oi_2 _3944_ (.B1(_1948_),
    .Y(_1953_),
    .A2(_1951_),
    .A1(_1949_));
 sg13g2_mux4_1 _3945_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(net124),
    .A1(net31),
    .A2(net25),
    .A3(net66),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_1954_));
 sg13g2_mux4_1 _3946_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net1600),
    .A1(net1612),
    .A2(net1606),
    .A3(net1626),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_1955_));
 sg13g2_inv_1 _3947_ (.Y(_1956_),
    .A(_1955_));
 sg13g2_mux4_1 _3948_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .A0(net1634),
    .A1(net1524),
    .A2(net1594),
    .A3(net1519),
    .S1(net1700),
    .X(_1957_));
 sg13g2_o21ai_1 _3949_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .Y(_1958_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1956_));
 sg13g2_a21oi_1 _3950_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_1957_),
    .Y(_1959_),
    .B1(_1958_));
 sg13g2_a21oi_1 _3951_ (.A1(net1706),
    .A2(net1700),
    .Y(_1960_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_o21ai_1 _3952_ (.B1(_1960_),
    .Y(_1961_),
    .A1(net1700),
    .A2(net620));
 sg13g2_nor2b_1 _3953_ (.A(net1700),
    .B_N(net2001),
    .Y(_1962_));
 sg13g2_a21oi_1 _3954_ (.A1(net11),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .Y(_1963_),
    .B1(_1962_));
 sg13g2_a21oi_1 _3955_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_1963_),
    .Y(_1964_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_a21oi_1 _3956_ (.A1(net29),
    .A2(net1700),
    .Y(_1965_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_o21ai_1 _3957_ (.B1(_1965_),
    .Y(_1966_),
    .A1(_0091_),
    .A2(net1700));
 sg13g2_nand2b_1 _3958_ (.Y(_1967_),
    .B(net1700),
    .A_N(net1930));
 sg13g2_o21ai_1 _3959_ (.B1(_1967_),
    .Y(_1968_),
    .A1(net37),
    .A2(net1700));
 sg13g2_a21oi_1 _3960_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_1968_),
    .Y(_1969_),
    .B1(_0122_));
 sg13g2_a221oi_1 _3961_ (.B2(_1969_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ),
    .B1(_1966_),
    .A1(_1961_),
    .Y(_1970_),
    .A2(_1964_));
 sg13g2_nor2_2 _3962_ (.A(_1970_),
    .B(_1959_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ));
 sg13g2_mux4_1 _3963_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(net611),
    .A1(net39),
    .A2(net13),
    .A3(net74),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_1971_));
 sg13g2_mux4_1 _3964_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A1(net73),
    .A2(net12),
    .A3(net727),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ),
    .X(_1972_));
 sg13g2_mux4_1 _3965_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ),
    .A0(_1972_),
    .A1(_1971_),
    .A2(_1954_),
    .A3(_0647_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ));
 sg13g2_nor2_2 _3966_ (.A(net1644),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .Y(_1973_));
 sg13g2_a21oi_2 _3967_ (.B1(_1973_),
    .Y(_1974_),
    .A2(_0035_),
    .A1(net1645));
 sg13g2_nor2_2 _3968_ (.A(net1651),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_a21oi_2 _3969_ (.B1(_1975_),
    .Y(_1976_),
    .A2(_0034_),
    .A1(net1651));
 sg13g2_nor2_2 _3970_ (.A(_1976_),
    .B(_1932_),
    .Y(_1977_));
 sg13g2_nand2_2 _3971_ (.Y(_1978_),
    .A(_1932_),
    .B(_1976_));
 sg13g2_nor2b_1 _3972_ (.A(_1977_),
    .B_N(_1978_),
    .Y(_1979_));
 sg13g2_xnor2_1 _3973_ (.Y(_1980_),
    .A(_1953_),
    .B(_1979_));
 sg13g2_mux2_1 _3974_ (.A0(_1980_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ),
    .S(net1655),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ));
 sg13g2_mux4_1 _3975_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .A2(_0646_),
    .A3(net727),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .X(_1981_));
 sg13g2_mux4_1 _3976_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1982_));
 sg13g2_mux2_1 _3977_ (.A0(_1982_),
    .A1(_1981_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ));
 sg13g2_nand2_1 _3978_ (.Y(_1983_),
    .A(net1638),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ));
 sg13g2_a21oi_1 _3979_ (.A1(net1644),
    .A2(_0155_),
    .Y(_1984_),
    .B1(net1651));
 sg13g2_a22oi_1 _3980_ (.Y(_1985_),
    .B1(_1983_),
    .B2(_1984_),
    .A2(_0036_),
    .A1(net1649));
 sg13g2_nor2b_1 _3981_ (.A(net700),
    .B_N(_1985_),
    .Y(_1986_));
 sg13g2_or2_1 _3982_ (.X(_1987_),
    .B(_1985_),
    .A(_1932_));
 sg13g2_nand2b_1 _3983_ (.Y(_1988_),
    .B(_1987_),
    .A_N(_1986_));
 sg13g2_a21oi_2 _3984_ (.B1(_1977_),
    .Y(_1989_),
    .A2(_1978_),
    .A1(_1953_));
 sg13g2_a21oi_1 _3985_ (.A1(_1987_),
    .A2(_1989_),
    .Y(_1990_),
    .B1(_1986_));
 sg13g2_a21oi_1 _3986_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .Y(_1991_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_o21ai_1 _3987_ (.B1(_1991_),
    .Y(_1992_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_0594_));
 sg13g2_mux4_1 _3988_ (.S0(net1701),
    .A0(net681),
    .A1(net1709),
    .A2(net1),
    .A3(net4),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_1993_));
 sg13g2_a21oi_1 _3989_ (.A1(net28),
    .A2(net1701),
    .Y(_1994_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_o21ai_1 _3990_ (.B1(_1994_),
    .Y(_1995_),
    .A1(_0070_),
    .A2(net1701));
 sg13g2_nor2b_1 _3991_ (.A(net1701),
    .B_N(net30),
    .Y(_1996_));
 sg13g2_a21oi_1 _3992_ (.A1(net62),
    .A2(net1701),
    .Y(_1997_),
    .B1(_1996_));
 sg13g2_a21oi_1 _3993_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_1997_),
    .Y(_1998_),
    .B1(_0158_));
 sg13g2_a221oi_1 _3994_ (.B2(_1998_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .B1(_1995_),
    .A1(_0158_),
    .Y(_1999_),
    .A2(_1993_));
 sg13g2_o21ai_1 _3995_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_2000_),
    .A1(net1702),
    .A2(_0177_));
 sg13g2_a21oi_1 _3996_ (.A1(net1701),
    .A2(net1623),
    .Y(_2001_),
    .B1(_2000_));
 sg13g2_mux2_1 _3997_ (.A0(net1598),
    .A1(net1611),
    .S(net1701),
    .X(_2002_));
 sg13g2_o21ai_1 _3998_ (.B1(_0158_),
    .Y(_2003_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_2002_));
 sg13g2_nand2_1 _3999_ (.Y(_2004_),
    .A(net1702),
    .B(_0179_));
 sg13g2_o21ai_1 _4000_ (.B1(_2004_),
    .Y(_2005_),
    .A1(net1702),
    .A2(net1586));
 sg13g2_nor2_1 _4001_ (.A(net1701),
    .B(net1633),
    .Y(_2006_));
 sg13g2_a21oi_1 _4002_ (.A1(net1702),
    .A2(_0174_),
    .Y(_2007_),
    .B1(_2006_));
 sg13g2_o21ai_1 _4003_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_2008_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_2007_));
 sg13g2_a21oi_1 _4004_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ),
    .A2(_2005_),
    .Y(_2009_),
    .B1(_2008_));
 sg13g2_o21ai_1 _4005_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ),
    .Y(_2010_),
    .A1(_2001_),
    .A2(_2003_));
 sg13g2_o21ai_1 _4006_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .Y(_2011_),
    .A1(_2009_),
    .A2(_2010_));
 sg13g2_nor2_2 _4007_ (.A(_0230_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .Y(_2012_));
 sg13g2_o21ai_1 _4008_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .Y(_2013_),
    .A1(_1999_),
    .A2(_2011_));
 sg13g2_or2_1 _4009_ (.X(_2014_),
    .B(_2012_),
    .A(_2013_));
 sg13g2_nand3_1 _4010_ (.B(_1992_),
    .C(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ),
    .A(_2014_),
    .Y(_2015_));
 sg13g2_mux4_1 _4011_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net1598),
    .A1(net1610),
    .A2(net649),
    .A3(net1623),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_2016_));
 sg13g2_inv_1 _4012_ (.Y(_2017_),
    .A(_2016_));
 sg13g2_mux4_1 _4013_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .A0(net1632),
    .A1(net1586),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .A3(net1539),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_2018_));
 sg13g2_o21ai_1 _4014_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_2019_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_2017_));
 sg13g2_a21oi_1 _4015_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_2018_),
    .Y(_2020_),
    .B1(_2019_));
 sg13g2_a21oi_1 _4016_ (.A1(net1709),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_2021_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_o21ai_1 _4017_ (.B1(_2021_),
    .Y(_2022_),
    .A1(net688),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_o21ai_1 _4018_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .Y(_2023_),
    .A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_a21oi_1 _4019_ (.A1(net4),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_2024_),
    .B1(_2023_));
 sg13g2_nor2_1 _4020_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .B(_2024_),
    .Y(_2025_));
 sg13g2_mux4_1 _4021_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net26),
    .A1(net28),
    .A2(net54),
    .A3(net83),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_2026_));
 sg13g2_a221oi_1 _4022_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ),
    .B1(_2026_),
    .A1(_2022_),
    .Y(_2027_),
    .A2(_2025_));
 sg13g2_nor2_2 _4023_ (.A(_2027_),
    .B(_2020_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ));
 sg13g2_nor2b_1 _4024_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .Y(_2028_));
 sg13g2_a21oi_1 _4025_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .Y(_2029_),
    .B1(_2028_));
 sg13g2_nand2_1 _4026_ (.Y(_2030_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .B(_2029_));
 sg13g2_mux4_1 _4027_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(net1597),
    .A1(net1610),
    .A2(net1603),
    .A3(net1624),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_2031_));
 sg13g2_inv_1 _4028_ (.Y(_2032_),
    .A(_2031_));
 sg13g2_mux4_1 _4029_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .A0(net1632),
    .A1(net1585),
    .A2(net1591),
    .A3(net1520),
    .S1(net1679),
    .X(_2033_));
 sg13g2_o21ai_1 _4030_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .Y(_2034_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_2032_));
 sg13g2_a21oi_1 _4031_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_2033_),
    .Y(_2035_),
    .B1(_2034_));
 sg13g2_a21oi_1 _4032_ (.A1(net1709),
    .A2(net1679),
    .Y(_2036_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_o21ai_1 _4033_ (.B1(_2036_),
    .Y(_2037_),
    .A1(net1679),
    .A2(net687));
 sg13g2_o21ai_1 _4034_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .Y(_2038_),
    .A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_a21oi_1 _4035_ (.A1(net22),
    .A2(net1679),
    .Y(_2039_),
    .B1(_2038_));
 sg13g2_nor2_1 _4036_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ),
    .B(_2039_),
    .Y(_2040_));
 sg13g2_a21oi_1 _4037_ (.A1(net30),
    .A2(net1679),
    .Y(_2041_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_o21ai_1 _4038_ (.B1(_2041_),
    .Y(_2042_),
    .A1(_0070_),
    .A2(net1679));
 sg13g2_nand2b_1 _4039_ (.Y(_2043_),
    .B(net1679),
    .A_N(net1932));
 sg13g2_o21ai_1 _4040_ (.B1(_2043_),
    .Y(_2044_),
    .A1(net62),
    .A2(net1679));
 sg13g2_a21oi_1 _4041_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_2044_),
    .Y(_2045_),
    .B1(_0157_));
 sg13g2_a221oi_1 _4042_ (.B2(_2045_),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ),
    .B1(_2042_),
    .A1(_2037_),
    .Y(_2046_),
    .A2(_2040_));
 sg13g2_nor2_2 _4043_ (.A(_2046_),
    .B(_2035_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ));
 sg13g2_mux2_1 _4044_ (.A0(net729),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_2047_));
 sg13g2_o21ai_1 _4045_ (.B1(_2030_),
    .Y(_2048_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_2047_));
 sg13g2_o21ai_1 _4046_ (.B1(_2015_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .A1(_2048_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_a21oi_1 _4047_ (.A1(net1644),
    .A2(_0159_),
    .Y(_2049_),
    .B1(net1649));
 sg13g2_o21ai_1 _4048_ (.B1(_2049_),
    .Y(_2050_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .A2(net1644));
 sg13g2_o21ai_1 _4049_ (.B1(_2050_),
    .Y(_2051_),
    .A1(net1636),
    .A2(_0160_));
 sg13g2_xnor2_1 _4050_ (.Y(_2052_),
    .A(net700),
    .B(_2051_));
 sg13g2_xor2_1 _4051_ (.B(_2052_),
    .A(_1990_),
    .X(_2053_));
 sg13g2_nand2_1 _4052_ (.Y(_2054_),
    .A(net1655),
    .B(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ));
 sg13g2_o21ai_1 _4053_ (.B1(_2054_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .A1(net1655),
    .A2(_2053_));
 sg13g2_xnor2_1 _4054_ (.Y(_2055_),
    .A(_1834_),
    .B(_1832_));
 sg13g2_mux2_1 _4055_ (.A0(_2055_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ),
    .S(net1655),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ));
 sg13g2_xnor2_1 _4056_ (.Y(_2056_),
    .A(_1989_),
    .B(_1988_));
 sg13g2_mux2_2 _4057_ (.A0(_2056_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ),
    .S(net1655),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ));
 sg13g2_xnor2_1 _4058_ (.Y(_2057_),
    .A(_1805_),
    .B(_1806_));
 sg13g2_nand2_1 _4059_ (.Y(_2058_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ),
    .B(net1652));
 sg13g2_o21ai_1 _4060_ (.B1(_2058_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .A1(_2057_),
    .A2(net1652));
 sg13g2_xnor2_1 _4061_ (.Y(_2059_),
    .A(_1822_),
    .B(_1823_));
 sg13g2_nand2_1 _4062_ (.Y(_2060_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ),
    .B(net1653));
 sg13g2_o21ai_1 _4063_ (.B1(_2060_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .A1(_2059_),
    .A2(net1653));
 sg13g2_nand2b_1 _4064_ (.Y(_2061_),
    .B(net610),
    .A_N(net1694));
 sg13g2_a21oi_1 _4065_ (.A1(_0060_),
    .A2(net1694),
    .Y(_2062_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_nor2_1 _4066_ (.A(net1694),
    .B(net5),
    .Y(_2063_));
 sg13g2_a21oi_1 _4067_ (.A1(_0075_),
    .A2(net1694),
    .Y(_2064_),
    .B1(_2063_));
 sg13g2_a221oi_1 _4068_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .B1(_2064_),
    .A1(_2061_),
    .Y(_2065_),
    .A2(_2062_));
 sg13g2_nand2_1 _4069_ (.Y(_2066_),
    .A(net1694),
    .B(_0087_));
 sg13g2_o21ai_1 _4070_ (.B1(_2066_),
    .Y(_2067_),
    .A1(net1694),
    .A2(net31));
 sg13g2_o21ai_1 _4071_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_2068_),
    .A1(net1693),
    .A2(net66));
 sg13g2_a21oi_1 _4072_ (.A1(_0076_),
    .A2(net1694),
    .Y(_2069_),
    .B1(_2068_));
 sg13g2_o21ai_1 _4073_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_2070_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_2067_));
 sg13g2_o21ai_1 _4074_ (.B1(_0088_),
    .Y(_2071_),
    .A1(_2069_),
    .A2(_2070_));
 sg13g2_mux2_1 _4075_ (.A0(net1621),
    .A1(net1629),
    .S(net1693),
    .X(_2072_));
 sg13g2_nor2b_1 _4076_ (.A(net1693),
    .B_N(net1609),
    .Y(_2073_));
 sg13g2_a21oi_1 _4077_ (.A1(net1693),
    .A2(net1602),
    .Y(_2074_),
    .B1(_2073_));
 sg13g2_a21oi_1 _4078_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_2072_),
    .Y(_2075_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_o21ai_1 _4079_ (.B1(_2075_),
    .Y(_2076_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_2074_));
 sg13g2_nand2_1 _4080_ (.Y(_2077_),
    .A(net1693),
    .B(net1518));
 sg13g2_o21ai_1 _4081_ (.B1(_2077_),
    .Y(_2078_),
    .A1(net1693),
    .A2(_0175_));
 sg13g2_nor2_1 _4082_ (.A(net1693),
    .B(net1590),
    .Y(_2079_));
 sg13g2_a21oi_1 _4083_ (.A1(net1693),
    .A2(net1584),
    .Y(_2080_),
    .B1(_2079_));
 sg13g2_o21ai_1 _4084_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_2081_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .A2(_2080_));
 sg13g2_a21o_1 _4085_ (.A2(_2078_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ),
    .B1(_2081_),
    .X(_2082_));
 sg13g2_nand3_1 _4086_ (.B(_2076_),
    .C(_2082_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_2083_));
 sg13g2_o21ai_1 _4087_ (.B1(_2083_),
    .Y(_2084_),
    .A1(_2065_),
    .A2(_2071_));
 sg13g2_mux4_1 _4088_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ),
    .A0(net1622),
    .A1(_0614_),
    .A2(_2084_),
    .A3(_0611_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ));
 sg13g2_mux4_1 _4089_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ),
    .A0(net1633),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .A2(net694),
    .A3(_0647_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ));
 sg13g2_mux4_1 _4090_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ),
    .A0(net1592),
    .A1(_0699_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .A3(_0721_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _4091_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ),
    .A0(net125),
    .A1(net136),
    .A2(net21),
    .A3(net1633),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ));
 sg13g2_mux4_1 _4092_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ),
    .A0(net126),
    .A1(net137),
    .A2(net20),
    .A3(net1591),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ));
 sg13g2_mux4_1 _4093_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ),
    .A0(net1709),
    .A1(net138),
    .A2(net82),
    .A3(net1586),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ));
 sg13g2_mux4_1 _4094_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ),
    .A0(net124),
    .A1(net1929),
    .A2(net135),
    .A3(net1522),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ));
 sg13g2_mux4_1 _4095_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ),
    .A0(net1621),
    .A1(net701),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .A3(_0385_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ));
 sg13g2_mux4_1 _4096_ (.S0(net1673),
    .A0(net1611),
    .A1(net1603),
    .A2(net1623),
    .A3(net1633),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_2085_));
 sg13g2_nor2_1 _4097_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .B(_2085_),
    .Y(_2086_));
 sg13g2_nor2_1 _4098_ (.A(net1672),
    .B(net1590),
    .Y(_2087_));
 sg13g2_a21oi_1 _4099_ (.A1(net1673),
    .A2(net1587),
    .Y(_2088_),
    .B1(_2087_));
 sg13g2_o21ai_1 _4100_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_2089_),
    .A1(net1673),
    .A2(net1522));
 sg13g2_a21oi_1 _4101_ (.A1(net1673),
    .A2(_0179_),
    .Y(_2090_),
    .B1(_2089_));
 sg13g2_o21ai_1 _4102_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .Y(_2091_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .A2(_2088_));
 sg13g2_o21ai_1 _4103_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_2092_),
    .A1(_2090_),
    .A2(_2091_));
 sg13g2_or2_1 _4104_ (.X(_2093_),
    .B(_2092_),
    .A(_2086_));
 sg13g2_nor2_1 _4105_ (.A(_0075_),
    .B(net1673),
    .Y(_2094_));
 sg13g2_a21oi_1 _4106_ (.A1(net55),
    .A2(net1672),
    .Y(_2095_),
    .B1(_2094_));
 sg13g2_nor2b_1 _4107_ (.A(net1672),
    .B_N(net66),
    .Y(_2096_));
 sg13g2_a21oi_1 _4108_ (.A1(net82),
    .A2(net1672),
    .Y(_2097_),
    .B1(_2096_));
 sg13g2_nor2b_1 _4109_ (.A(net1672),
    .B_N(net2002),
    .Y(_2098_));
 sg13g2_a21oi_1 _4110_ (.A1(net5),
    .A2(net1672),
    .Y(_2099_),
    .B1(_2098_));
 sg13g2_nor2_1 _4111_ (.A(_0060_),
    .B(net1672),
    .Y(_2100_));
 sg13g2_a21oi_1 _4112_ (.A1(net136),
    .A2(net1672),
    .Y(_2101_),
    .B1(_2100_));
 sg13g2_mux4_1 _4113_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ),
    .A0(_2101_),
    .A1(_2099_),
    .A2(_2095_),
    .A3(_2097_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ),
    .X(_2102_));
 sg13g2_o21ai_1 _4114_ (.B1(_2093_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ),
    .A2(_2102_));
 sg13g2_mux4_1 _4115_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ),
    .A0(net1630),
    .A1(_0614_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .A3(_0611_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ));
 sg13g2_mux4_1 _4116_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ),
    .A0(net690),
    .A1(net694),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .A3(_0647_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ));
 sg13g2_mux4_1 _4117_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ),
    .A0(net1583),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .A2(_0699_),
    .A3(_0721_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ));
 sg13g2_mux4_1 _4118_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ),
    .A0(net21),
    .A1(net47),
    .A2(net32),
    .A3(net1596),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ));
 sg13g2_mux4_1 _4119_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ),
    .A0(net20),
    .A1(net48),
    .A2(net33),
    .A3(net1609),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ));
 sg13g2_mux4_1 _4120_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ),
    .A0(net30),
    .A1(net82),
    .A2(net49),
    .A3(net648),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ));
 sg13g2_mux4_1 _4121_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ),
    .A0(net31),
    .A1(net46),
    .A2(net1929),
    .A3(net1622),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _4122_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ),
    .A0(net1592),
    .A1(net701),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .A3(_0385_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _4123_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ),
    .A0(net1583),
    .A1(_0614_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .A3(_0611_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _4124_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ),
    .A0(net1521),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A2(net1576),
    .A3(_0647_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _4125_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ),
    .A0(net1596),
    .A1(_0699_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .A3(_0721_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _4126_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .A0(net1588),
    .A1(_0969_),
    .A2(_1011_),
    .A3(_1922_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .X(_2103_));
 sg13g2_mux4_1 _4127_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ),
    .A0(net1516),
    .A1(net3),
    .A2(net1932),
    .A3(net1605),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_2104_));
 sg13g2_mux2_1 _4128_ (.A0(_2104_),
    .A1(_2103_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ));
 sg13g2_mux4_1 _4129_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .A0(_0598_),
    .A1(net1930),
    .A2(net2001),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_2105_));
 sg13g2_nor2_1 _4130_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .B(_2105_),
    .Y(_2106_));
 sg13g2_nand2_1 _4131_ (.Y(_2107_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .B(_1499_));
 sg13g2_o21ai_1 _4132_ (.B1(_2107_),
    .Y(_2108_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_0868_));
 sg13g2_nand2_1 _4133_ (.Y(_2109_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .B(_0630_));
 sg13g2_o21ai_1 _4134_ (.B1(_2109_),
    .Y(_2110_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(net1523));
 sg13g2_o21ai_1 _4135_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ),
    .Y(_2111_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_2110_));
 sg13g2_a21oi_1 _4136_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ),
    .A2(_2108_),
    .Y(_2112_),
    .B1(_2111_));
 sg13g2_nor2_1 _4137_ (.A(_2106_),
    .B(_2112_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ));
 sg13g2_a21oi_1 _4138_ (.A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .Y(_2113_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ));
 sg13g2_o21ai_1 _4139_ (.B1(_2113_),
    .Y(_2114_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(net681));
 sg13g2_mux2_1 _4140_ (.A0(net62),
    .A1(net1634),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_2115_));
 sg13g2_a21oi_1 _4141_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .A2(_2115_),
    .Y(_2116_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ));
 sg13g2_o21ai_1 _4142_ (.B1(_0156_),
    .Y(_2117_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(net1519));
 sg13g2_a21oi_1 _4143_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_1482_),
    .Y(_2118_),
    .B1(_2117_));
 sg13g2_mux2_1 _4144_ (.A0(net1576),
    .A1(_0934_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ),
    .X(_2119_));
 sg13g2_nand2_1 _4145_ (.Y(_2120_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ),
    .B(_2119_));
 sg13g2_nor2b_1 _4146_ (.A(_2118_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ),
    .Y(_2121_));
 sg13g2_a22oi_1 _4147_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ),
    .B1(_2120_),
    .B2(_2121_),
    .A2(_2114_),
    .A1(_2116_));
 sg13g2_mux4_1 _4148_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .A0(net1527),
    .A1(net1933),
    .A2(net2004),
    .A3(net1594),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .X(_2122_));
 sg13g2_mux4_1 _4149_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ),
    .A0(net1539),
    .A1(_1470_),
    .A2(net623),
    .A3(_1020_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ),
    .X(_2123_));
 sg13g2_mux2_1 _4150_ (.A0(_2122_),
    .A1(_2123_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ));
 sg13g2_mux4_1 _4151_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .A0(net1588),
    .A1(_0969_),
    .A2(_1011_),
    .A3(_1841_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_2124_));
 sg13g2_mux4_1 _4152_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ),
    .A0(net1516),
    .A1(net28),
    .A2(net3),
    .A3(net1606),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_2125_));
 sg13g2_mux2_1 _4153_ (.A0(_2125_),
    .A1(_2124_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ));
 sg13g2_mux4_1 _4154_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(_0598_),
    .A1(net2001),
    .A2(net29),
    .A3(net1626),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_2126_));
 sg13g2_nand2_1 _4155_ (.Y(_2127_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .B(_0630_));
 sg13g2_o21ai_1 _4156_ (.B1(_2127_),
    .Y(_2128_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(net1524));
 sg13g2_nand2_1 _4157_ (.Y(_2129_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .B(_1512_));
 sg13g2_o21ai_1 _4158_ (.B1(_2129_),
    .Y(_2130_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_0868_));
 sg13g2_a21oi_1 _4159_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .A2(_2130_),
    .Y(_2131_),
    .B1(_0161_));
 sg13g2_o21ai_1 _4160_ (.B1(_2131_),
    .Y(_2132_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ),
    .A2(_2128_));
 sg13g2_o21ai_1 _4161_ (.B1(_2132_),
    .Y(_2133_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ),
    .A2(_2126_));
 sg13g2_inv_1 _4162_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ),
    .A(_2133_));
 sg13g2_a21oi_1 _4163_ (.A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .Y(_2134_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_o21ai_1 _4164_ (.B1(_2134_),
    .Y(_2135_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(net681));
 sg13g2_mux2_1 _4165_ (.A0(net26),
    .A1(net1634),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_2136_));
 sg13g2_a21oi_1 _4166_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_2136_),
    .Y(_2137_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_o21ai_1 _4167_ (.B1(_0163_),
    .Y(_2138_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(net1519));
 sg13g2_a21oi_1 _4168_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_1482_),
    .Y(_2139_),
    .B1(_2138_));
 sg13g2_nor2_1 _4169_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ),
    .B(net1576),
    .Y(_2140_));
 sg13g2_o21ai_1 _4170_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ),
    .Y(_2141_),
    .A1(_0162_),
    .A2(_0257_));
 sg13g2_o21ai_1 _4171_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ),
    .Y(_2142_),
    .A1(_2140_),
    .A2(_2141_));
 sg13g2_nor2_1 _4172_ (.A(_2139_),
    .B(_2142_),
    .Y(_2143_));
 sg13g2_a21oi_2 _4173_ (.B1(_2143_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ),
    .A2(_2137_),
    .A1(_2135_));
 sg13g2_mux4_1 _4174_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .A0(net1527),
    .A1(net27),
    .A2(net2004),
    .A3(net1593),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_2144_));
 sg13g2_mux4_1 _4175_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ),
    .A0(net1540),
    .A1(_1470_),
    .A2(net623),
    .A3(_0974_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_2145_));
 sg13g2_mux2_1 _4176_ (.A0(_2144_),
    .A1(_2145_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ));
 sg13g2_mux4_1 _4177_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net2001),
    .A1(net1930),
    .A2(net1599),
    .A3(net1613),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_2146_));
 sg13g2_mux4_1 _4178_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .A0(net1606),
    .A1(net1634),
    .A2(net1626),
    .A3(net1593),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_2147_));
 sg13g2_inv_1 _4179_ (.Y(_2148_),
    .A(_2147_));
 sg13g2_a21oi_1 _4180_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2148_),
    .Y(_2149_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ));
 sg13g2_o21ai_1 _4181_ (.B1(_2149_),
    .Y(_2150_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2146_));
 sg13g2_mux4_1 _4182_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .A0(_1011_),
    .A1(_1483_),
    .A2(_0969_),
    .A3(net1576),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .X(_2151_));
 sg13g2_nor2b_1 _4183_ (.A(_2151_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .Y(_2152_));
 sg13g2_mux4_1 _4184_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net1588),
    .A1(net1523),
    .A2(net1519),
    .A3(net1540),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_2153_));
 sg13g2_o21ai_1 _4185_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ),
    .Y(_2154_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_2153_));
 sg13g2_o21ai_1 _4186_ (.B1(_2150_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ),
    .A1(_2152_),
    .A2(_2154_));
 sg13g2_mux4_1 _4187_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .A0(net3),
    .A1(net1600),
    .A2(net1932),
    .A3(net1613),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_2155_));
 sg13g2_mux4_1 _4188_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .A0(net1606),
    .A1(net1634),
    .A2(net1626),
    .A3(net1593),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_2156_));
 sg13g2_inv_1 _4189_ (.Y(_2157_),
    .A(_2156_));
 sg13g2_a21oi_1 _4190_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_2157_),
    .Y(_2158_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_o21ai_1 _4191_ (.B1(_2158_),
    .Y(_2159_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_2155_));
 sg13g2_mux2_1 _4192_ (.A0(_0630_),
    .A1(_0868_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_2160_));
 sg13g2_mux2_1 _4193_ (.A0(_1470_),
    .A1(net623),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .X(_2161_));
 sg13g2_o21ai_1 _4194_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .Y(_2162_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_2160_));
 sg13g2_a21oi_1 _4195_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_2161_),
    .Y(_2163_),
    .B1(_2162_));
 sg13g2_mux4_1 _4196_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(net1588),
    .A1(net1524),
    .A2(net1519),
    .A3(net1540),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ),
    .X(_2164_));
 sg13g2_o21ai_1 _4197_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ),
    .Y(_2165_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_2164_));
 sg13g2_o21ai_1 _4198_ (.B1(_2159_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ),
    .A1(_2163_),
    .A2(_2165_));
 sg13g2_mux4_1 _4199_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .A0(net1584),
    .A1(_0969_),
    .A2(_1011_),
    .A3(_1954_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_2166_));
 sg13g2_mux4_1 _4200_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net2003),
    .A2(net1932),
    .A3(net1602),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_2167_));
 sg13g2_mux2_1 _4201_ (.A0(_2167_),
    .A1(_2166_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ));
 sg13g2_nand2_1 _4202_ (.Y(_2168_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .B(_0232_));
 sg13g2_o21ai_1 _4203_ (.B1(_2168_),
    .Y(_2169_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_0868_));
 sg13g2_nand2_2 _4204_ (.Y(_2170_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .B(_0630_));
 sg13g2_o21ai_1 _4205_ (.B1(_2170_),
    .Y(_2171_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(net1526));
 sg13g2_o21ai_1 _4206_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ),
    .Y(_2172_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_2171_));
 sg13g2_a21oi_2 _4207_ (.B1(_2172_),
    .Y(_2173_),
    .A2(_2169_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ));
 sg13g2_mux4_1 _4208_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ),
    .A0(_0598_),
    .A1(net1931),
    .A2(net2001),
    .A3(net1622),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_2174_));
 sg13g2_nor2_1 _4209_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ),
    .B(_2174_),
    .Y(_2175_));
 sg13g2_nor2_2 _4210_ (.A(_2173_),
    .B(_2175_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ));
 sg13g2_a21oi_1 _4211_ (.A1(_0061_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .Y(_2176_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ));
 sg13g2_o21ai_1 _4212_ (.B1(_2176_),
    .Y(_2177_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(net681));
 sg13g2_mux2_1 _4213_ (.A0(net62),
    .A1(net1631),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_2178_));
 sg13g2_a21oi_1 _4214_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .A2(_2178_),
    .Y(_2179_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ));
 sg13g2_nand2_1 _4215_ (.Y(_2180_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .B(_1482_));
 sg13g2_o21ai_1 _4216_ (.B1(_2180_),
    .Y(_2181_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(net1518));
 sg13g2_mux2_1 _4217_ (.A0(net1576),
    .A1(_0835_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ),
    .X(_2182_));
 sg13g2_o21ai_1 _4218_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ),
    .Y(_2183_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .A2(_2181_));
 sg13g2_a21oi_1 _4219_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ),
    .A2(_2182_),
    .Y(_2184_),
    .B1(_2183_));
 sg13g2_a21oi_2 _4220_ (.B1(_2184_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ),
    .A2(_2179_),
    .A1(_2177_));
 sg13g2_mux4_1 _4221_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .A0(net1527),
    .A1(net1933),
    .A2(net2004),
    .A3(net691),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .X(_2185_));
 sg13g2_mux4_1 _4222_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ),
    .A0(net699),
    .A1(_1470_),
    .A2(net623),
    .A3(_0513_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ),
    .X(_2186_));
 sg13g2_mux2_1 _4223_ (.A0(_2185_),
    .A1(_2186_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ));
 sg13g2_mux4_1 _4224_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .A0(net1584),
    .A1(_0969_),
    .A2(_1011_),
    .A3(_1935_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_2187_));
 sg13g2_mux4_1 _4225_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ),
    .A0(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .A1(net28),
    .A2(net1932),
    .A3(net1607),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_2188_));
 sg13g2_mux2_1 _4226_ (.A0(_2188_),
    .A1(_2187_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _4227_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .A0(_0598_),
    .A1(net1931),
    .A2(net29),
    .A3(net1622),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_2189_));
 sg13g2_nand2_1 _4228_ (.Y(_2190_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .B(_0630_));
 sg13g2_o21ai_1 _4229_ (.B1(_2190_),
    .Y(_2191_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(net1526));
 sg13g2_nand2_1 _4230_ (.Y(_2192_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .B(_1469_));
 sg13g2_o21ai_1 _4231_ (.B1(_2192_),
    .Y(_2193_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_0868_));
 sg13g2_a21oi_1 _4232_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .A2(_2193_),
    .Y(_2194_),
    .B1(_0164_));
 sg13g2_o21ai_1 _4233_ (.B1(_2194_),
    .Y(_2195_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ),
    .A2(_2191_));
 sg13g2_o21ai_1 _4234_ (.B1(_2195_),
    .Y(_2196_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ),
    .A2(_2189_));
 sg13g2_inv_1 _4235_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ),
    .A(_2196_));
 sg13g2_a21oi_1 _4236_ (.A1(_0070_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .Y(_2197_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_o21ai_1 _4237_ (.B1(_2197_),
    .Y(_2198_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(net681));
 sg13g2_mux2_1 _4238_ (.A0(net62),
    .A1(net1630),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .X(_2199_));
 sg13g2_a21oi_1 _4239_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_2199_),
    .Y(_2200_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_o21ai_1 _4240_ (.B1(_0165_),
    .Y(_2201_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(net1518));
 sg13g2_a21o_1 _4241_ (.A2(_1482_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .B1(_2201_),
    .X(_2202_));
 sg13g2_o21ai_1 _4242_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ),
    .Y(_2203_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(net694));
 sg13g2_a21oi_1 _4243_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0896_),
    .Y(_2204_),
    .B1(_2203_));
 sg13g2_nor2b_1 _4244_ (.A(_2204_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ),
    .Y(_2205_));
 sg13g2_a22oi_1 _4245_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ),
    .B1(_2202_),
    .B2(_2205_),
    .A2(_2198_),
    .A1(_2200_));
 sg13g2_mux4_1 _4246_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .A0(_0376_),
    .A1(net63),
    .A2(net27),
    .A3(net1591),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2206_));
 sg13g2_mux4_1 _4247_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ),
    .A0(net1539),
    .A1(_1470_),
    .A2(net623),
    .A3(_0525_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_2207_));
 sg13g2_mux2_1 _4248_ (.A0(_2206_),
    .A1(_2207_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _4249_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(net2002),
    .A1(net1931),
    .A2(net1599),
    .A3(net1612),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2208_));
 sg13g2_mux4_1 _4250_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .A0(net1605),
    .A1(net1635),
    .A2(net1625),
    .A3(net1594),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_2209_));
 sg13g2_inv_1 _4251_ (.Y(_2210_),
    .A(_2209_));
 sg13g2_a21oi_1 _4252_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2210_),
    .Y(_2211_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_o21ai_1 _4253_ (.B1(_2211_),
    .Y(_2212_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2208_));
 sg13g2_mux4_1 _4254_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .A0(_1011_),
    .A1(_1483_),
    .A2(_0969_),
    .A3(net1576),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .X(_2213_));
 sg13g2_nor2b_1 _4255_ (.A(_2213_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .Y(_2214_));
 sg13g2_mux4_1 _4256_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(net1589),
    .A1(net1523),
    .A2(net1519),
    .A3(net1541),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2215_));
 sg13g2_o21ai_1 _4257_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ),
    .Y(_2216_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2215_));
 sg13g2_o21ai_1 _4258_ (.B1(_2212_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ),
    .A1(_2214_),
    .A2(_2216_));
 sg13g2_mux4_1 _4259_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(net2003),
    .A1(net1597),
    .A2(net64),
    .A3(net1610),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_2217_));
 sg13g2_mux4_1 _4260_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A0(net649),
    .A1(net1632),
    .A2(net1624),
    .A3(net1591),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_2218_));
 sg13g2_inv_1 _4261_ (.Y(_2219_),
    .A(_2218_));
 sg13g2_a21oi_1 _4262_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_2219_),
    .Y(_2220_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_o21ai_1 _4263_ (.B1(_2220_),
    .Y(_2221_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_2217_));
 sg13g2_mux2_1 _4264_ (.A0(_0630_),
    .A1(_0868_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_2222_));
 sg13g2_mux2_1 _4265_ (.A0(_1470_),
    .A1(net623),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .X(_2223_));
 sg13g2_o21ai_1 _4266_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .Y(_2224_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_2222_));
 sg13g2_a21oi_1 _4267_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .A2(_2223_),
    .Y(_2225_),
    .B1(_2224_));
 sg13g2_mux4_1 _4268_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ),
    .A0(net1585),
    .A1(net1522),
    .A2(net1520),
    .A3(net1540),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ),
    .X(_2226_));
 sg13g2_o21ai_1 _4269_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_2227_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_2226_));
 sg13g2_o21ai_1 _4270_ (.B1(_2221_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ),
    .A1(_2227_),
    .A2(_2225_));
 sg13g2_mux4_1 _4271_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ),
    .A0(net1602),
    .A1(_0194_),
    .A2(net701),
    .A3(_0385_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ));
 sg13g2_mux4_1 _4272_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ),
    .A0(net117),
    .A1(net1921),
    .A2(net132),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ));
 sg13g2_mux4_1 _4273_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ),
    .A0(net118),
    .A1(net1923),
    .A2(net133),
    .A3(net1563),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ));
 sg13g2_mux4_1 _4274_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ),
    .A0(net115),
    .A1(net134),
    .A2(net1703),
    .A3(net1573),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ));
 sg13g2_mux4_1 _4275_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ),
    .A0(net116),
    .A1(net131),
    .A2(net167),
    .A3(net1577),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ),
    .X(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ));
 sg13g2_mux4_1 _4276_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ),
    .A0(net1551),
    .A1(net693),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A3(_0308_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ));
 sg13g2_mux4_1 _4277_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ),
    .A0(net1559),
    .A1(net689),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .A3(_0362_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ));
 sg13g2_mux4_1 _4278_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ),
    .A0(net1565),
    .A1(net613),
    .A2(_1724_),
    .A3(_1673_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ));
 sg13g2_mux4_1 _4279_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ),
    .A0(net1570),
    .A1(net643),
    .A2(_0966_),
    .A3(net669),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ),
    .X(_2228_));
 sg13g2_inv_2 _4280_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ),
    .A(_2228_));
 sg13g2_mux4_1 _4281_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(net1557),
    .A1(net693),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .A3(_0308_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ));
 sg13g2_mux2_1 _4282_ (.A0(net1579),
    .A1(net1617),
    .S(net1663),
    .X(_2229_));
 sg13g2_mux2_1 _4283_ (.A0(net1561),
    .A1(net1570),
    .S(net1663),
    .X(_2230_));
 sg13g2_o21ai_1 _4284_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_2231_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_2230_));
 sg13g2_a21o_1 _4285_ (.A2(_2229_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .B1(_2231_),
    .X(_2232_));
 sg13g2_mux2_1 _4286_ (.A0(net1550),
    .A1(net1557),
    .S(net1663),
    .X(_2233_));
 sg13g2_mux2_1 _4287_ (.A0(_0180_),
    .A1(_0176_),
    .S(net1664),
    .X(_2234_));
 sg13g2_a21oi_1 _4288_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_2233_),
    .Y(_2235_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_o21ai_1 _4289_ (.B1(_2235_),
    .Y(_2236_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_2234_));
 sg13g2_nand3_1 _4290_ (.B(_2232_),
    .C(_2236_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_2237_));
 sg13g2_nor2b_1 _4291_ (.A(net1664),
    .B_N(net132),
    .Y(_2238_));
 sg13g2_a21oi_1 _4292_ (.A1(net108),
    .A2(net1664),
    .Y(_2239_),
    .B1(_2238_));
 sg13g2_nor2b_1 _4293_ (.A(net1663),
    .B_N(net1710),
    .Y(_2240_));
 sg13g2_a21oi_1 _4294_ (.A1(net116),
    .A2(net1663),
    .Y(_2241_),
    .B1(_2240_));
 sg13g2_nor2b_1 _4295_ (.A(net1664),
    .B_N(net152),
    .Y(_2242_));
 sg13g2_a21oi_1 _4296_ (.A1(net1703),
    .A2(net1663),
    .Y(_2243_),
    .B1(_2242_));
 sg13g2_nor2b_1 _4297_ (.A(net1663),
    .B_N(net1921),
    .Y(_2244_));
 sg13g2_a21oi_1 _4298_ (.A1(net1936),
    .A2(net1663),
    .Y(_2245_),
    .B1(_2244_));
 sg13g2_mux4_1 _4299_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ),
    .A0(_2241_),
    .A1(_2245_),
    .A2(_2239_),
    .A3(_2243_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_2246_));
 sg13g2_o21ai_1 _4300_ (.B1(_2237_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_2246_));
 sg13g2_mux4_1 _4301_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ),
    .A0(net1565),
    .A1(net689),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .A3(_0362_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _4302_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ),
    .A0(net1572),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .A2(net1517),
    .A3(_1673_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _4303_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ),
    .A0(net1579),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .A2(_0596_),
    .A3(_0566_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _4304_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ),
    .A0(net1921),
    .A1(net51),
    .A2(net1935),
    .A3(net1529),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ));
 sg13g2_mux4_1 _4305_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ),
    .A0(net1923),
    .A1(net41),
    .A2(net52),
    .A3(net1535),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ));
 sg13g2_mux4_1 _4306_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ),
    .A0(net38),
    .A1(net53),
    .A2(net1703),
    .A3(net1544),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ));
 sg13g2_mux4_1 _4307_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ),
    .A0(net1936),
    .A1(net50),
    .A2(net167),
    .A3(net1551),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _4308_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ),
    .A0(net1564),
    .A1(net693),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .A3(_0308_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ));
 sg13g2_o21ai_1 _4309_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_2247_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(net1577));
 sg13g2_a21oi_1 _4310_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(_0178_),
    .Y(_2248_),
    .B1(_2247_));
 sg13g2_a21oi_1 _4311_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(net1569),
    .Y(_2249_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_o21ai_1 _4312_ (.B1(_2249_),
    .Y(_2250_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(net1564));
 sg13g2_nand2_1 _4313_ (.Y(_2251_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_2250_));
 sg13g2_mux4_1 _4314_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net1534),
    .A1(net1542),
    .A2(net1549),
    .A3(net1557),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_2252_));
 sg13g2_nor2_1 _4315_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_2252_),
    .Y(_2253_));
 sg13g2_o21ai_1 _4316_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ),
    .Y(_2254_),
    .A1(_2248_),
    .A2(_2251_));
 sg13g2_mux4_1 _4317_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net1936),
    .A1(net51),
    .A2(net152),
    .A3(net1703),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_2255_));
 sg13g2_mux4_1 _4318_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(net140),
    .A1(net1925),
    .A2(net92),
    .A3(net1921),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_2256_));
 sg13g2_mux2_1 _4319_ (.A0(_2256_),
    .A1(_2255_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_2257_));
 sg13g2_nand2b_1 _4320_ (.Y(_2258_),
    .B(_2257_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_o21ai_1 _4321_ (.B1(_2258_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .A1(_2253_),
    .A2(_2254_));
 sg13g2_mux4_1 _4322_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ),
    .A0(net1573),
    .A1(net689),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .A3(_0362_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _4323_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ),
    .A0(net1577),
    .A1(net683),
    .A2(net1517),
    .A3(_1673_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _4324_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ),
    .A0(net1529),
    .A1(_0596_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .A3(_0566_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _4325_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A0(net1711),
    .A1(net89),
    .A2(net149),
    .A3(net1544),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_2259_));
 sg13g2_nor2_1 _4326_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ),
    .B(_2259_),
    .Y(_2260_));
 sg13g2_o21ai_1 _4327_ (.B1(_0166_),
    .Y(_2261_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(net1572));
 sg13g2_a21oi_1 _4328_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_1058_),
    .Y(_2262_),
    .B1(_2261_));
 sg13g2_nor2b_1 _4329_ (.A(_1714_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .Y(_2263_));
 sg13g2_nor2_1 _4330_ (.A(_0166_),
    .B(_2263_),
    .Y(_2264_));
 sg13g2_o21ai_1 _4331_ (.B1(_2264_),
    .Y(_2265_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_1277_));
 sg13g2_nor2b_1 _4332_ (.A(_2262_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ),
    .Y(_2266_));
 sg13g2_a21oi_1 _4333_ (.A1(_2265_),
    .A2(_2266_),
    .Y(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ),
    .B1(_2260_));
 sg13g2_nand2_1 _4334_ (.Y(_2267_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .B(net1553));
 sg13g2_o21ai_1 _4335_ (.B1(_2267_),
    .Y(_2268_),
    .A1(_0104_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ));
 sg13g2_mux2_1 _4336_ (.A0(net1710),
    .A1(net1925),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .X(_2269_));
 sg13g2_mux2_1 _4337_ (.A0(_1130_),
    .A1(_1772_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .X(_2270_));
 sg13g2_mux2_1 _4338_ (.A0(net1581),
    .A1(_0905_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ),
    .X(_2271_));
 sg13g2_mux4_1 _4339_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ),
    .A0(_2269_),
    .A1(_2271_),
    .A2(_2268_),
    .A3(_2270_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ));
 sg13g2_mux4_1 _4340_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .A0(net1713),
    .A1(net1928),
    .A2(net147),
    .A3(net1559),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .X(_2272_));
 sg13g2_nor2_1 _4341_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ),
    .B(_2272_),
    .Y(_2273_));
 sg13g2_mux2_1 _4342_ (.A0(_1724_),
    .A1(_1259_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .X(_2274_));
 sg13g2_nand2_1 _4343_ (.Y(_2275_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .B(_1780_));
 sg13g2_o21ai_1 _4344_ (.B1(_2275_),
    .Y(_2276_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(net1615));
 sg13g2_o21ai_1 _4345_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ),
    .Y(_2277_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_2276_));
 sg13g2_a21oi_1 _4346_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ),
    .A2(_2274_),
    .Y(_2278_),
    .B1(_2277_));
 sg13g2_nor2_1 _4347_ (.A(_2273_),
    .B(_2278_),
    .Y(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ));
 sg13g2_mux4_1 _4348_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .A0(net1619),
    .A1(_1699_),
    .A2(_1759_),
    .A3(_1091_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_2279_));
 sg13g2_mux4_1 _4349_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ),
    .A0(net1712),
    .A1(net148),
    .A2(net1927),
    .A3(net1566),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ),
    .X(_2280_));
 sg13g2_mux2_1 _4350_ (.A0(_2280_),
    .A1(_2279_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ),
    .X(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ));
 sg13g2_nor2_1 _4351_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .B(_0682_),
    .Y(_2281_));
 sg13g2_a21oi_1 _4352_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(_0176_),
    .Y(_2282_),
    .B1(_2281_));
 sg13g2_or2_1 _4353_ (.X(_2283_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A(net1711));
 sg13g2_a21oi_1 _4354_ (.A1(_0073_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .Y(_2284_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ));
 sg13g2_a221oi_1 _4355_ (.B2(_2284_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ),
    .B1(_2283_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .Y(_2285_),
    .A2(_2282_));
 sg13g2_nand2_1 _4356_ (.Y(_2286_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .B(_1058_));
 sg13g2_o21ai_1 _4357_ (.B1(_2286_),
    .Y(_2287_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(net1573));
 sg13g2_nand2_1 _4358_ (.Y(_2288_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .B(_1734_));
 sg13g2_o21ai_1 _4359_ (.B1(_2288_),
    .Y(_2289_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ),
    .A2(_1278_));
 sg13g2_o21ai_1 _4360_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ),
    .Y(_2290_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_2287_));
 sg13g2_a21oi_1 _4361_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_2289_),
    .Y(_2291_),
    .B1(_2290_));
 sg13g2_nor2_1 _4362_ (.A(_2285_),
    .B(_2291_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ));
 sg13g2_mux4_1 _4363_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A0(net1710),
    .A1(net1925),
    .A2(_0723_),
    .A3(net1554),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_2292_));
 sg13g2_mux4_1 _4364_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ),
    .A0(net1582),
    .A1(_0905_),
    .A2(_1130_),
    .A3(_1792_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ),
    .X(_2293_));
 sg13g2_mux2_1 _4365_ (.A0(_2292_),
    .A1(_2293_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ));
 sg13g2_a21oi_1 _4366_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(net1555),
    .Y(_2294_),
    .B1(_0167_));
 sg13g2_o21ai_1 _4367_ (.B1(_2294_),
    .Y(_2295_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(net703));
 sg13g2_mux2_1 _4368_ (.A0(net1713),
    .A1(net1928),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .X(_2296_));
 sg13g2_a21oi_1 _4369_ (.A1(_0167_),
    .A2(_2296_),
    .Y(_2297_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ));
 sg13g2_a21oi_1 _4370_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(_1316_),
    .Y(_2298_),
    .B1(_0167_));
 sg13g2_o21ai_1 _4371_ (.B1(_2298_),
    .Y(_2299_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(net1517));
 sg13g2_nand2_1 _4372_ (.Y(_2300_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .B(_1780_));
 sg13g2_o21ai_1 _4373_ (.B1(_2300_),
    .Y(_2301_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(net1616));
 sg13g2_o21ai_1 _4374_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ),
    .Y(_2302_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ),
    .A2(_2301_));
 sg13g2_inv_1 _4375_ (.Y(_2303_),
    .A(_2302_));
 sg13g2_a22oi_1 _4376_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ),
    .B1(_2299_),
    .B2(_2303_),
    .A2(_2297_),
    .A1(_2295_));
 sg13g2_mux4_1 _4377_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .A0(net1712),
    .A1(net1927),
    .A2(_0616_),
    .A3(net1566),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .X(_2304_));
 sg13g2_mux4_1 _4378_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ),
    .A0(net1620),
    .A1(_1699_),
    .A2(_1759_),
    .A3(_1210_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ),
    .X(_2305_));
 sg13g2_mux2_1 _4379_ (.A0(_2304_),
    .A1(_2305_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ));
 sg13g2_mux4_1 _4380_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .A0(net90),
    .A1(net1704),
    .A2(net1529),
    .A3(net1535),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_2306_));
 sg13g2_mux4_1 _4381_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .A0(net1544),
    .A1(net1550),
    .A2(net1559),
    .A3(net1565),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_2307_));
 sg13g2_or2_1 _4382_ (.X(_2308_),
    .B(_1058_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_a21oi_1 _4383_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .A2(_1277_),
    .Y(_2309_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ));
 sg13g2_nor2_1 _4384_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .B(_1780_),
    .Y(_2310_));
 sg13g2_a21oi_1 _4385_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .A2(net1517),
    .Y(_2311_),
    .B1(_2310_));
 sg13g2_a22oi_1 _4386_ (.Y(_2312_),
    .B1(_2311_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .A2(_2309_),
    .A1(_2308_));
 sg13g2_mux4_1 _4387_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ),
    .A0(net1572),
    .A1(net1579),
    .A2(net1615),
    .A3(net1618),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ),
    .X(_2313_));
 sg13g2_mux4_1 _4388_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ),
    .A0(_2306_),
    .A1(_2307_),
    .A2(_2313_),
    .A3(_2312_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ));
 sg13g2_mux4_1 _4389_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(_0905_),
    .A1(_1130_),
    .A2(_1759_),
    .A3(_1699_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_2314_));
 sg13g2_mux4_1 _4390_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net1574),
    .A1(net1580),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .A3(net1618),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_2315_));
 sg13g2_mux2_1 _4391_ (.A0(_2315_),
    .A1(_2314_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_2316_));
 sg13g2_mux4_1 _4392_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net89),
    .A1(net149),
    .A2(net1530),
    .A3(net1535),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_2317_));
 sg13g2_mux4_1 _4393_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(net1544),
    .A1(net1551),
    .A2(net1560),
    .A3(net1566),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ),
    .X(_2318_));
 sg13g2_mux2_1 _4394_ (.A0(_2317_),
    .A1(_2318_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ),
    .X(_2319_));
 sg13g2_mux2_1 _4395_ (.A0(_2319_),
    .A1(_2316_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ));
 sg13g2_mux4_1 _4396_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A0(net113),
    .A1(net1926),
    .A2(net149),
    .A3(net1544),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_2320_));
 sg13g2_nor2_1 _4397_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ),
    .B(_2320_),
    .Y(_2321_));
 sg13g2_o21ai_1 _4398_ (.B1(_0168_),
    .Y(_2322_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(net1572));
 sg13g2_a21oi_1 _4399_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(_1058_),
    .Y(_2323_),
    .B1(_2322_));
 sg13g2_nand2_1 _4400_ (.Y(_2324_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .B(_1674_));
 sg13g2_o21ai_1 _4401_ (.B1(_2324_),
    .Y(_2325_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ),
    .A2(_1278_));
 sg13g2_nand2_1 _4402_ (.Y(_2326_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ),
    .B(_2325_));
 sg13g2_nor2b_1 _4403_ (.A(_2323_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ),
    .Y(_2327_));
 sg13g2_a21oi_1 _4404_ (.A1(_2326_),
    .A2(_2327_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ),
    .B1(_2321_));
 sg13g2_mux4_1 _4405_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A0(net1580),
    .A1(_0905_),
    .A2(_1130_),
    .A3(_1744_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_2328_));
 sg13g2_mux4_1 _4406_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ),
    .A0(net1710),
    .A1(net90),
    .A2(net1704),
    .A3(net1550),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ),
    .X(_2329_));
 sg13g2_mux2_1 _4407_ (.A0(_2329_),
    .A1(_2328_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ));
 sg13g2_mux4_1 _4408_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .A0(net1713),
    .A1(net1928),
    .A2(net147),
    .A3(net1559),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .X(_2330_));
 sg13g2_nor2_1 _4409_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ),
    .B(_2330_),
    .Y(_2331_));
 sg13g2_nand2_1 _4410_ (.Y(_2332_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .B(_1780_));
 sg13g2_o21ai_1 _4411_ (.B1(_2332_),
    .Y(_2333_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(net1615));
 sg13g2_mux2_1 _4412_ (.A0(net1517),
    .A1(_0763_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ),
    .X(_2334_));
 sg13g2_o21ai_1 _4413_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ),
    .Y(_2335_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_2333_));
 sg13g2_a21oi_1 _4414_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_2334_),
    .Y(_2336_),
    .B1(_2335_));
 sg13g2_nor2_1 _4415_ (.A(_2331_),
    .B(_2336_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ));
 sg13g2_mux4_1 _4416_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .A0(net1618),
    .A1(_1699_),
    .A2(_1759_),
    .A3(_0805_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_2337_));
 sg13g2_mux4_1 _4417_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ),
    .A0(net1712),
    .A1(net148),
    .A2(net1927),
    .A3(net1565),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ),
    .X(_2338_));
 sg13g2_mux2_1 _4418_ (.A0(_2338_),
    .A1(_2337_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ));
 sg13g2_a21oi_1 _4419_ (.A1(_0065_),
    .A2(_0169_),
    .Y(_2339_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ));
 sg13g2_o21ai_1 _4420_ (.B1(_2339_),
    .Y(_2340_),
    .A1(_0169_),
    .A2(_0682_));
 sg13g2_o21ai_1 _4421_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .Y(_2341_),
    .A1(net1705),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_a21oi_1 _4422_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(_0176_),
    .Y(_2342_),
    .B1(_2341_));
 sg13g2_nor2_1 _4423_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ),
    .B(_2342_),
    .Y(_2343_));
 sg13g2_a21o_1 _4424_ (.A2(net1570),
    .A1(_0169_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .X(_2344_));
 sg13g2_a21oi_1 _4425_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .A2(_1058_),
    .Y(_2345_),
    .B1(_2344_));
 sg13g2_nor2_1 _4426_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ),
    .B(_1277_),
    .Y(_2346_));
 sg13g2_o21ai_1 _4427_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ),
    .Y(_2347_),
    .A1(_0169_),
    .A2(_1695_));
 sg13g2_o21ai_1 _4428_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ),
    .Y(_2348_),
    .A1(_2346_),
    .A2(_2347_));
 sg13g2_nor2_1 _4429_ (.A(_2345_),
    .B(_2348_),
    .Y(_2349_));
 sg13g2_a21oi_1 _4430_ (.A1(_2340_),
    .A2(_2343_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ),
    .B1(_2349_));
 sg13g2_mux4_1 _4431_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .A0(net1710),
    .A1(net1704),
    .A2(_0723_),
    .A3(net1551),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .X(_2350_));
 sg13g2_mux4_1 _4432_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ),
    .A0(net1578),
    .A1(_0905_),
    .A2(_1130_),
    .A3(_1751_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ),
    .X(_2351_));
 sg13g2_mux2_1 _4433_ (.A0(_2350_),
    .A1(_2351_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ));
 sg13g2_nand2_1 _4434_ (.Y(_2352_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .B(net718));
 sg13g2_o21ai_1 _4435_ (.B1(_2352_),
    .Y(_2353_),
    .A1(net1713),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_o21ai_1 _4436_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .Y(_2354_),
    .A1(net147),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_a21oi_1 _4437_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(net1555),
    .Y(_2355_),
    .B1(_2354_));
 sg13g2_nor2_1 _4438_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .B(_2355_),
    .Y(_2356_));
 sg13g2_o21ai_1 _4439_ (.B1(_2356_),
    .Y(_2357_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_2353_));
 sg13g2_a21o_1 _4440_ (.A2(_0178_),
    .A1(_0170_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .X(_2358_));
 sg13g2_a21oi_1 _4441_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_1780_),
    .Y(_2359_),
    .B1(_2358_));
 sg13g2_nor2_1 _4442_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ),
    .B(net1517),
    .Y(_2360_));
 sg13g2_o21ai_1 _4443_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ),
    .Y(_2361_),
    .A1(_0170_),
    .A2(_1147_));
 sg13g2_o21ai_1 _4444_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ),
    .Y(_2362_),
    .A1(_2360_),
    .A2(_2361_));
 sg13g2_o21ai_1 _4445_ (.B1(_2357_),
    .Y(_2363_),
    .A1(_2359_),
    .A2(_2362_));
 sg13g2_inv_1 _4446_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ),
    .A(_2363_));
 sg13g2_mux4_1 _4447_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .A0(net112),
    .A1(net148),
    .A2(_0616_),
    .A3(net1564),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_2364_));
 sg13g2_mux4_1 _4448_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ),
    .A0(net1618),
    .A1(_1699_),
    .A2(_1759_),
    .A3(_0926_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ),
    .X(_2365_));
 sg13g2_mux2_1 _4449_ (.A0(_2364_),
    .A1(_2365_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _4450_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .A0(net1925),
    .A1(net1704),
    .A2(net1528),
    .A3(net1534),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2366_));
 sg13g2_mux4_1 _4451_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .A0(net1542),
    .A1(net1549),
    .A2(net1556),
    .A3(net1563),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2367_));
 sg13g2_or2_1 _4452_ (.X(_2368_),
    .B(_1058_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_a21oi_1 _4453_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(_1277_),
    .Y(_2369_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_nor2_1 _4454_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .B(_1780_),
    .Y(_2370_));
 sg13g2_a21oi_1 _4455_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .A2(net1517),
    .Y(_2371_),
    .B1(_2370_));
 sg13g2_a22oi_1 _4456_ (.Y(_2372_),
    .B1(_2371_),
    .B2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .A2(_2369_),
    .A1(_2368_));
 sg13g2_mux4_1 _4457_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ),
    .A0(net1573),
    .A1(net1577),
    .A2(net1615),
    .A3(net1617),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ),
    .X(_2373_));
 sg13g2_mux4_1 _4458_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ),
    .A0(_2366_),
    .A1(_2367_),
    .A2(_2373_),
    .A3(_2372_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ),
    .X(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ));
 sg13g2_mux4_1 _4459_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(net1926),
    .A1(net1705),
    .A2(net1528),
    .A3(net1535),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2374_));
 sg13g2_mux4_1 _4460_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(net1543),
    .A1(net1551),
    .A2(net1558),
    .A3(net1564),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2375_));
 sg13g2_inv_1 _4461_ (.Y(_2376_),
    .A(_2375_));
 sg13g2_a21oi_1 _4462_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2376_),
    .Y(_2377_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_o21ai_1 _4463_ (.B1(_2377_),
    .Y(_2378_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2374_));
 sg13g2_mux4_1 _4464_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(_0905_),
    .A1(_1130_),
    .A2(_1759_),
    .A3(_1699_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2379_));
 sg13g2_nor2b_1 _4465_ (.A(_2379_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .Y(_2380_));
 sg13g2_mux4_1 _4466_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(net1573),
    .A1(net1578),
    .A2(net1615),
    .A3(net1617),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ),
    .X(_2381_));
 sg13g2_o21ai_1 _4467_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ),
    .Y(_2382_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_2381_));
 sg13g2_o21ai_1 _4468_ (.B1(_2378_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ),
    .A1(_2380_),
    .A2(_2382_));
 sg13g2_nor2b_1 _4469_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .Y(_2383_));
 sg13g2_mux4_1 _4470_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .A1(net617),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_2384_));
 sg13g2_nor2b_1 _4471_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .B_N(_2384_),
    .Y(_2385_));
 sg13g2_nor2_1 _4472_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .B(net712),
    .Y(_2386_));
 sg13g2_o21ai_1 _4473_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .Y(_2387_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(_2386_));
 sg13g2_a21oi_1 _4474_ (.A1(_1559_),
    .A2(_2383_),
    .Y(_2388_),
    .B1(_2387_));
 sg13g2_o21ai_1 _4475_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .Y(_2389_),
    .A1(_2385_),
    .A2(_2388_));
 sg13g2_mux4_1 _4476_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(net1707),
    .A1(net99),
    .A2(net105),
    .A3(net642),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .X(_2390_));
 sg13g2_nor2b_1 _4477_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .B_N(_2390_),
    .Y(_2391_));
 sg13g2_mux4_1 _4478_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ),
    .A0(net159),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .A3(net614),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ),
    .X(_2392_));
 sg13g2_a21oi_1 _4479_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_2392_),
    .Y(_2393_),
    .B1(_2391_));
 sg13g2_o21ai_1 _4480_ (.B1(_2389_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ),
    .A2(_2393_));
 sg13g2_nor2_1 _4481_ (.A(net1512),
    .B(_1884_),
    .Y(_0038_));
 sg13g2_nor2_1 _4482_ (.A(net1512),
    .B(_2057_),
    .Y(_0039_));
 sg13g2_nor2b_1 _4483_ (.A(net1512),
    .B_N(_1883_),
    .Y(_0040_));
 sg13g2_nor2b_1 _4484_ (.A(net1512),
    .B_N(_1888_),
    .Y(_0041_));
 sg13g2_nor2_1 _4485_ (.A(net1512),
    .B(_1886_),
    .Y(_0042_));
 sg13g2_nor2b_1 _4486_ (.A(net1512),
    .B_N(_1889_),
    .Y(_0043_));
 sg13g2_nor2_1 _4487_ (.A(net1512),
    .B(_1890_),
    .Y(_0044_));
 sg13g2_nor2b_1 _4488_ (.A(net1514),
    .B_N(_1892_),
    .Y(_0045_));
 sg13g2_nor2_1 _4489_ (.A(net1512),
    .B(_2059_),
    .Y(_0046_));
 sg13g2_nor2_1 _4490_ (.A(net1514),
    .B(_1893_),
    .Y(_0047_));
 sg13g2_nor2_1 _4491_ (.A(net1513),
    .B(_1895_),
    .Y(_0048_));
 sg13g2_nor2b_1 _4492_ (.A(net1513),
    .B_N(_1897_),
    .Y(_0049_));
 sg13g2_nor2_1 _4493_ (.A(net1513),
    .B(_1898_),
    .Y(_0050_));
 sg13g2_nor2b_1 _4494_ (.A(net1514),
    .B_N(_2055_),
    .Y(_0051_));
 sg13g2_nor2_1 _4495_ (.A(net1513),
    .B(_1881_),
    .Y(_0052_));
 sg13g2_nor2b_1 _4496_ (.A(net1513),
    .B_N(_1930_),
    .Y(_0053_));
 sg13g2_nor2b_1 _4497_ (.A(net1514),
    .B_N(_1952_),
    .Y(_0054_));
 sg13g2_nor2b_1 _4498_ (.A(net1513),
    .B_N(_1980_),
    .Y(_0055_));
 sg13g2_nor2b_1 _4499_ (.A(net1513),
    .B_N(_2056_),
    .Y(_0056_));
 sg13g2_nor2_1 _4500_ (.A(net1513),
    .B(net711),
    .Y(_0057_));
 sg13g2_inv_1 _4501_ (.Y(_0058_),
    .A(net167));
 sg13g2_inv_1 _4502_ (.Y(_0059_),
    .A(net20));
 sg13g2_inv_1 _4503_ (.Y(_0060_),
    .A(net124));
 sg13g2_inv_1 _4504_ (.Y(_0061_),
    .A(net1));
 sg13g2_inv_1 _4505_ (.Y(_0062_),
    .A(net48));
 sg13g2_inv_1 _4506_ (.Y(_0063_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_inv_1 _4507_ (.Y(_0064_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_inv_1 _4508_ (.Y(_0065_),
    .A(net113));
 sg13g2_inv_1 _4509_ (.Y(_0066_),
    .A(net42));
 sg13g2_inv_1 _4510_ (.Y(_0067_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_inv_1 _4511_ (.Y(_0068_),
    .A(net41));
 sg13g2_inv_1 _4512_ (.Y(_0069_),
    .A(net1709));
 sg13g2_inv_1 _4513_ (.Y(_0070_),
    .A(net26));
 sg13g2_inv_1 _4514_ (.Y(_0071_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_inv_1 _4515_ (.Y(_0072_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_inv_1 _4516_ (.Y(_0073_),
    .A(net89));
 sg13g2_inv_1 _4517_ (.Y(_0074_),
    .A(net126));
 sg13g2_inv_1 _4518_ (.Y(_0075_),
    .A(net21));
 sg13g2_inv_1 _4519_ (.Y(_0076_),
    .A(net82));
 sg13g2_inv_1 _4520_ (.Y(_0077_),
    .A(net38));
 sg13g2_inv_1 _4521_ (.Y(_0078_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_inv_1 _4522_ (.Y(_0079_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_inv_1 _4523_ (.Y(_0080_),
    .A(net19));
 sg13g2_inv_1 _4524_ (.Y(_0081_),
    .A(net1934));
 sg13g2_inv_1 _4525_ (.Y(_0082_),
    .A(net80));
 sg13g2_inv_1 _4526_ (.Y(_0083_),
    .A(net128));
 sg13g2_inv_1 _4527_ (.Y(_0084_),
    .A(net104));
 sg13g2_inv_1 _4528_ (.Y(_0085_),
    .A(net164));
 sg13g2_inv_1 _4529_ (.Y(_0086_),
    .A(net36));
 sg13g2_inv_1 _4530_ (.Y(_0087_),
    .A(net47));
 sg13g2_inv_1 _4531_ (.Y(_0088_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_inv_1 _4532_ (.Y(_0089_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_inv_1 _4533_ (.Y(_0090_),
    .A(net29));
 sg13g2_inv_1 _4534_ (.Y(_0091_),
    .A(net27));
 sg13g2_inv_1 _4535_ (.Y(_0092_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_inv_1 _4536_ (.Y(_0093_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_inv_1 _4537_ (.Y(_0094_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_inv_1 _4538_ (.Y(_0095_),
    .A(net44));
 sg13g2_inv_1 _4539_ (.Y(_0096_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_inv_1 _4540_ (.Y(_0097_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_inv_1 _4541_ (.Y(_0098_),
    .A(net17));
 sg13g2_inv_1 _4542_ (.Y(_0099_),
    .A(net43));
 sg13g2_inv_1 _4543_ (.Y(_0100_),
    .A(net78));
 sg13g2_inv_1 _4544_ (.Y(_0101_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_inv_1 _4545_ (.Y(_0102_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_inv_1 _4546_ (.Y(_0103_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_inv_1 _4547_ (.Y(_0104_),
    .A(net1704));
 sg13g2_inv_1 _4548_ (.Y(_0105_),
    .A(net148));
 sg13g2_inv_1 _4549_ (.Y(_0106_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_inv_1 _4550_ (.Y(_0107_),
    .A(net1660));
 sg13g2_inv_1 _4551_ (.Y(_0108_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_inv_1 _4552_ (.Y(_0109_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_inv_1 _4553_ (.Y(_0110_),
    .A(net16));
 sg13g2_inv_1 _4554_ (.Y(_0111_),
    .A(net77));
 sg13g2_inv_1 _4555_ (.Y(_0112_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_inv_1 _4556_ (.Y(_0113_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_inv_1 _4557_ (.Y(_0114_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_inv_1 _4558_ (.Y(_0115_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_inv_1 _4559_ (.Y(_0116_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_inv_1 _4560_ (.Y(_0117_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_inv_1 _4561_ (.Y(_0118_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_inv_1 _4562_ (.Y(_0119_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_inv_1 _4563_ (.Y(_0120_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_inv_1 _4564_ (.Y(_0121_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_inv_1 _4565_ (.Y(_0122_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_inv_1 _4566_ (.Y(_0123_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ));
 sg13g2_inv_1 _4567_ (.Y(_0124_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_inv_1 _4568_ (.Y(_0125_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_inv_1 _4569_ (.Y(_0126_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_inv_1 _4570_ (.Y(_0127_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_inv_1 _4571_ (.Y(_0128_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_inv_1 _4572_ (.Y(_0129_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_inv_1 _4573_ (.Y(_0130_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_inv_1 _4574_ (.Y(_0131_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_inv_1 _4575_ (.Y(_0132_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_inv_1 _4576_ (.Y(_0133_),
    .A(_0001_));
 sg13g2_inv_1 _4577_ (.Y(_0134_),
    .A(net1644));
 sg13g2_inv_1 _4578_ (.Y(_0135_),
    .A(net1649));
 sg13g2_inv_1 _4579_ (.Y(_0136_),
    .A(_0003_));
 sg13g2_inv_1 _4580_ (.Y(_0137_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_inv_1 _4581_ (.Y(_0138_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_inv_1 _4582_ (.Y(_0139_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_inv_1 _4583_ (.Y(_0140_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_inv_1 _4584_ (.Y(_0141_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_inv_1 _4585_ (.Y(_0142_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_inv_1 _4586_ (.Y(_0143_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_inv_1 _4587_ (.Y(_0144_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_inv_1 _4588_ (.Y(_0145_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_inv_1 _4589_ (.Y(_0146_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_inv_1 _4590_ (.Y(_0147_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_inv_1 _4591_ (.Y(_0148_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_inv_1 _4592_ (.Y(_0149_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_inv_1 _4593_ (.Y(_0150_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_inv_1 _4594_ (.Y(_0151_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_inv_1 _4595_ (.Y(_0152_),
    .A(_0013_));
 sg13g2_inv_1 _4596_ (.Y(_0153_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_inv_1 _4597_ (.Y(_0154_),
    .A(_0021_));
 sg13g2_inv_1 _4598_ (.Y(_0155_),
    .A(_0037_));
 sg13g2_inv_1 _4599_ (.Y(_0156_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ));
 sg13g2_inv_1 _4600_ (.Y(_0157_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_inv_1 _4601_ (.Y(_0158_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_inv_1 _4602_ (.Y(_0159_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ));
 sg13g2_inv_1 _4603_ (.Y(_0160_),
    .A(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ));
 sg13g2_inv_1 _4604_ (.Y(_0161_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ));
 sg13g2_inv_1 _4605_ (.Y(_0162_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ));
 sg13g2_inv_1 _4606_ (.Y(_0163_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_inv_1 _4607_ (.Y(_0164_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_inv_1 _4608_ (.Y(_0165_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_inv_1 _4609_ (.Y(_0166_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ));
 sg13g2_inv_1 _4610_ (.Y(_0167_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ));
 sg13g2_inv_1 _4611_ (.Y(_0168_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ));
 sg13g2_inv_1 _4612_ (.Y(_0169_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_inv_1 _4613_ (.Y(_0170_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_inv_1 _4614_ (.Y(_0171_),
    .A(net1558));
 sg13g2_inv_8 _4615_ (.Y(_0172_),
    .A(net1563));
 sg13g2_inv_1 _4616_ (.Y(_0173_),
    .A(net1572));
 sg13g2_inv_1 _4617_ (.Y(_0174_),
    .A(net1591));
 sg13g2_inv_1 _4618_ (.Y(_0175_),
    .A(net1525));
 sg13g2_inv_1 _4619_ (.Y(_0176_),
    .A(net1544));
 sg13g2_inv_1 _4620_ (.Y(_0177_),
    .A(net1603));
 sg13g2_inv_1 _4621_ (.Y(_0178_),
    .A(net1616));
 sg13g2_inv_1 _4622_ (.Y(_0179_),
    .A(net1539));
 sg13g2_inv_4 _4623_ (.A(net1535),
    .Y(_0180_));
 sg13g2_mux4_1 _4624_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(net1598),
    .A1(net1611),
    .A2(net1603),
    .A3(net1633),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0181_));
 sg13g2_mux4_1 _4625_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(net1591),
    .A1(net1587),
    .A2(net1522),
    .A3(net1539),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0182_));
 sg13g2_nand2b_1 _4626_ (.Y(_0183_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A_N(_0182_));
 sg13g2_o21ai_1 _4627_ (.B1(_0183_),
    .Y(_0184_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0181_));
 sg13g2_mux4_1 _4628_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .A0(net1516),
    .A1(net8),
    .A2(net1708),
    .A3(net20),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0185_));
 sg13g2_nor2b_1 _4629_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .B_N(_0185_),
    .Y(_0186_));
 sg13g2_mux2_1 _4630_ (.A0(net34),
    .A1(net46),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0187_));
 sg13g2_nand2b_1 _4631_ (.Y(_0188_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ),
    .A_N(net1929));
 sg13g2_o21ai_1 _4632_ (.B1(_0188_),
    .Y(_0189_),
    .A1(net69),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_o21ai_1 _4633_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0190_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .A2(_0187_));
 sg13g2_a21oi_1 _4634_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ),
    .A2(_0189_),
    .Y(_0191_),
    .B1(_0190_));
 sg13g2_nor3_1 _4635_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .B(_0186_),
    .C(_0191_),
    .Y(_0192_));
 sg13g2_a21o_1 _4636_ (.A2(_0184_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ),
    .B1(_0192_),
    .X(_0193_));
 sg13g2_inv_1 _4637_ (.Y(_0194_),
    .A(_0193_));
 sg13g2_mux4_1 _4638_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ),
    .A0(net25),
    .A1(net84),
    .A2(net46),
    .A3(_0194_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0195_));
 sg13g2_mux4_1 _4639_ (.S0(net1657),
    .A0(net1528),
    .A1(net1542),
    .A2(net1549),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0196_));
 sg13g2_nand2b_1 _4640_ (.Y(_0197_),
    .B(_0196_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_nor2_1 _4641_ (.A(net1657),
    .B(net1563),
    .Y(_0198_));
 sg13g2_a21oi_1 _4642_ (.A1(net1657),
    .A2(net1569),
    .Y(_0199_),
    .B1(_0198_));
 sg13g2_nand2b_1 _4643_ (.Y(_0200_),
    .B(net1657),
    .A_N(net1617));
 sg13g2_o21ai_1 _4644_ (.B1(_0200_),
    .Y(_0201_),
    .A1(net1657),
    .A2(net1577));
 sg13g2_o21ai_1 _4645_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0202_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0199_));
 sg13g2_a21oi_1 _4646_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0201_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_nor2b_1 _4647_ (.A(_0203_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_0204_));
 sg13g2_mux4_1 _4648_ (.S0(net1657),
    .A0(net117),
    .A1(net133),
    .A2(net1928),
    .A3(net93),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0205_));
 sg13g2_nand2b_1 _4649_ (.Y(_0206_),
    .B(_0205_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_nand2_1 _4650_ (.Y(_0207_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .B(_0058_));
 sg13g2_o21ai_1 _4651_ (.B1(_0207_),
    .Y(_0208_),
    .A1(net1657),
    .A2(net153));
 sg13g2_mux2_1 _4652_ (.A0(net1923),
    .A1(net1935),
    .S(net1657),
    .X(_0209_));
 sg13g2_o21ai_1 _4653_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ),
    .Y(_0210_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0209_));
 sg13g2_a21oi_1 _4654_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ),
    .A2(_0208_),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_nor2_1 _4655_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_a22oi_1 _4656_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .B1(_0206_),
    .B2(_0212_),
    .A2(_0204_),
    .A1(_0197_));
 sg13g2_mux4_1 _4657_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ),
    .A0(net611),
    .A1(net39),
    .A2(net13),
    .A3(net74),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0213_));
 sg13g2_o21ai_1 _4658_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .Y(_0214_),
    .A1(net1699),
    .A2(_0175_));
 sg13g2_a21oi_1 _4659_ (.A1(net1699),
    .A2(net1539),
    .Y(_0215_),
    .B1(_0214_));
 sg13g2_mux2_1 _4660_ (.A0(net1632),
    .A1(net1585),
    .S(net1699),
    .X(_0216_));
 sg13g2_o21ai_1 _4661_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .Y(_0217_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_0216_));
 sg13g2_mux4_1 _4662_ (.S0(net1699),
    .A0(net1597),
    .A1(net1610),
    .A2(net1603),
    .A3(net1623),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0218_));
 sg13g2_nand2b_1 _4663_ (.Y(_0219_),
    .B(_0218_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_and2_1 _4664_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ),
    .B(_0219_),
    .X(_0220_));
 sg13g2_o21ai_1 _4665_ (.B1(_0220_),
    .Y(_0221_),
    .A1(_0215_),
    .A2(_0217_));
 sg13g2_mux4_1 _4666_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .A0(net1516),
    .A1(net2003),
    .A2(net1707),
    .A3(net10),
    .S1(net1699),
    .X(_0222_));
 sg13g2_nand2b_1 _4667_ (.Y(_0223_),
    .B(_0222_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_o21ai_1 _4668_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .Y(_0224_),
    .A1(_0086_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_a21oi_1 _4669_ (.A1(net64),
    .A2(net1699),
    .Y(_0225_),
    .B1(_0224_));
 sg13g2_nand2_1 _4670_ (.Y(_0226_),
    .A(net28),
    .B(net1699));
 sg13g2_o21ai_1 _4671_ (.B1(_0226_),
    .Y(_0227_),
    .A1(_0070_),
    .A2(net1699));
 sg13g2_o21ai_1 _4672_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ),
    .Y(_0228_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_0227_));
 sg13g2_o21ai_1 _4673_ (.B1(_0223_),
    .Y(_0229_),
    .A1(_0225_),
    .A2(_0228_));
 sg13g2_o21ai_1 _4674_ (.B1(_0221_),
    .Y(_0230_),
    .A1(_0229_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_inv_1 _4675_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .A(net722));
 sg13g2_mux4_1 _4676_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ),
    .A0(net12),
    .A1(net73),
    .A2(net38),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0231_));
 sg13g2_mux4_1 _4677_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(net145),
    .A1(net5),
    .A2(net31),
    .A3(net66),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_0232_));
 sg13g2_mux4_1 _4678_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ),
    .A0(_0231_),
    .A1(_0232_),
    .A2(_0213_),
    .A3(_0195_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ));
 sg13g2_o21ai_1 _4679_ (.B1(net1636),
    .Y(_0233_),
    .A1(net1638),
    .A2(_0027_));
 sg13g2_a21oi_1 _4680_ (.A1(net1638),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .Y(_0234_),
    .B1(_0233_));
 sg13g2_a21o_1 _4681_ (.A2(_0026_),
    .A1(net1650),
    .B1(_0234_),
    .X(_0235_));
 sg13g2_mux4_1 _4682_ (.S0(net1676),
    .A0(net1597),
    .A1(net1610),
    .A2(net1624),
    .A3(net1632),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0236_));
 sg13g2_nor2_1 _4683_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_nor2_1 _4684_ (.A(net1676),
    .B(net1590),
    .Y(_0238_));
 sg13g2_a21oi_1 _4685_ (.A1(net1676),
    .A2(net1585),
    .Y(_0239_),
    .B1(_0238_));
 sg13g2_o21ai_1 _4686_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .Y(_0240_),
    .A1(net1676),
    .A2(net1525));
 sg13g2_a21oi_1 _4687_ (.A1(net1676),
    .A2(_0179_),
    .Y(_0241_),
    .B1(_0240_));
 sg13g2_o21ai_1 _4688_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0242_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0239_));
 sg13g2_o21ai_1 _4689_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .Y(_0243_),
    .A1(_0241_),
    .A2(_0242_));
 sg13g2_mux4_1 _4690_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(net126),
    .A1(net138),
    .A2(net2004),
    .A3(net7),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .X(_0244_));
 sg13g2_mux2_1 _4691_ (.A0(net68),
    .A1(net84),
    .S(net1676),
    .X(_0245_));
 sg13g2_nor2_1 _4692_ (.A(_0075_),
    .B(net1676),
    .Y(_0246_));
 sg13g2_a21oi_1 _4693_ (.A1(net33),
    .A2(net1676),
    .Y(_0247_),
    .B1(_0246_));
 sg13g2_o21ai_1 _4694_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0248_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0247_));
 sg13g2_a21oi_1 _4695_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0245_),
    .Y(_0249_),
    .B1(_0248_));
 sg13g2_nor2_1 _4696_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ),
    .B(_0249_),
    .Y(_0250_));
 sg13g2_o21ai_1 _4697_ (.B1(_0250_),
    .Y(_0251_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0244_));
 sg13g2_o21ai_1 _4698_ (.B1(_0251_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .A1(_0237_),
    .A2(_0243_));
 sg13g2_mux2_1 _4699_ (.A0(net85),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_0252_));
 sg13g2_nor2b_1 _4700_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .B_N(net7),
    .Y(_0253_));
 sg13g2_a21oi_1 _4701_ (.A1(net57),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_o21ai_1 _4702_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .Y(_0255_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_0254_));
 sg13g2_a21oi_1 _4703_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_0252_),
    .Y(_0256_),
    .B1(_0255_));
 sg13g2_mux4_1 _4704_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ),
    .A0(net146),
    .A1(net36),
    .A2(net10),
    .A3(net71),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ),
    .X(_0257_));
 sg13g2_o21ai_1 _4705_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .Y(_0258_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0257_));
 sg13g2_nor2_1 _4706_ (.A(_0256_),
    .B(_0258_),
    .Y(_0259_));
 sg13g2_nand2b_1 _4707_ (.Y(_0260_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A_N(net1609));
 sg13g2_o21ai_1 _4708_ (.B1(_0260_),
    .Y(_0261_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(net1596));
 sg13g2_mux2_1 _4709_ (.A0(net1622),
    .A1(net1630),
    .S(net1683),
    .X(_0262_));
 sg13g2_a21oi_1 _4710_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0262_),
    .Y(_0263_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_o21ai_1 _4711_ (.B1(_0263_),
    .Y(_0264_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0261_));
 sg13g2_nand2b_1 _4712_ (.Y(_0265_),
    .B(net1683),
    .A_N(net1584));
 sg13g2_o21ai_1 _4713_ (.B1(_0265_),
    .Y(_0266_),
    .A1(net1683),
    .A2(net1592));
 sg13g2_mux2_1 _4714_ (.A0(net1521),
    .A1(net1518),
    .S(net1683),
    .X(_0267_));
 sg13g2_o21ai_1 _4715_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0268_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0266_));
 sg13g2_a21oi_1 _4716_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0267_),
    .Y(_0269_),
    .B1(_0268_));
 sg13g2_nor2b_1 _4717_ (.A(_0269_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .Y(_0270_));
 sg13g2_mux4_1 _4718_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(net1596),
    .A1(net1602),
    .A2(net1621),
    .A3(net1629),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0271_));
 sg13g2_inv_1 _4719_ (.Y(_0272_),
    .A(_0271_));
 sg13g2_mux2_1 _4720_ (.A0(net1592),
    .A1(net1583),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0273_));
 sg13g2_nand2b_1 _4721_ (.Y(_0274_),
    .B(_0273_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_mux2_1 _4722_ (.A0(net1521),
    .A1(net1518),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0275_));
 sg13g2_a21oi_1 _4723_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0275_),
    .Y(_0276_),
    .B1(_0063_));
 sg13g2_a221oi_1 _4724_ (.B2(_0274_),
    .C1(_0064_),
    .B1(_0276_),
    .A1(_0063_),
    .Y(_0277_),
    .A2(_0272_));
 sg13g2_nor2b_1 _4725_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .B_N(net48),
    .Y(_0278_));
 sg13g2_a21oi_1 _4726_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(net56),
    .Y(_0279_),
    .B1(_0278_));
 sg13g2_mux2_1 _4727_ (.A0(net67),
    .A1(net1929),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0280_));
 sg13g2_a21oi_1 _4728_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0280_),
    .Y(_0281_),
    .B1(_0063_));
 sg13g2_o21ai_1 _4729_ (.B1(_0281_),
    .Y(_0282_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0279_));
 sg13g2_mux2_1 _4730_ (.A0(net24),
    .A1(net20),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0283_));
 sg13g2_mux2_1 _4731_ (.A0(net145),
    .A1(net1),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0284_));
 sg13g2_nand2b_1 _4732_ (.Y(_0285_),
    .B(_0284_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_a21oi_1 _4733_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_0283_),
    .Y(_0286_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_a21oi_1 _4734_ (.A1(_0285_),
    .A2(_0286_),
    .Y(_0287_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_a21oi_2 _4735_ (.B1(_0277_),
    .Y(_0288_),
    .A2(_0287_),
    .A1(_0282_));
 sg13g2_inv_2 _4736_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A(_0288_));
 sg13g2_mux4_1 _4737_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(net124),
    .A1(net100),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .A3(net160),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_0289_));
 sg13g2_inv_1 _4738_ (.Y(_0290_),
    .A(net692));
 sg13g2_nand2_1 _4739_ (.Y(_0291_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .B(_0289_));
 sg13g2_o21ai_1 _4740_ (.B1(_0291_),
    .Y(_0292_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(_0176_));
 sg13g2_mux2_1 _4741_ (.A0(net1550),
    .A1(net1559),
    .S(net1666),
    .X(_0293_));
 sg13g2_or2_1 _4742_ (.X(_0294_),
    .B(net1529),
    .A(net1666));
 sg13g2_a21oi_1 _4743_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0180_),
    .Y(_0295_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_a221oi_1 _4744_ (.B2(_0295_),
    .C1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .B1(_0294_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Y(_0296_),
    .A2(_0293_));
 sg13g2_nand2_1 _4745_ (.Y(_0297_),
    .A(net1666),
    .B(net1572));
 sg13g2_nand2b_1 _4746_ (.Y(_0298_),
    .B(net1565),
    .A_N(net1666));
 sg13g2_a21oi_1 _4747_ (.A1(_0297_),
    .A2(_0298_),
    .Y(_0299_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_nor2b_1 _4748_ (.A(net1618),
    .B_N(net1666),
    .Y(_0300_));
 sg13g2_o21ai_1 _4749_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .Y(_0301_),
    .A1(net1666),
    .A2(net1579));
 sg13g2_o21ai_1 _4750_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0302_),
    .A1(_0300_),
    .A2(_0301_));
 sg13g2_o21ai_1 _4751_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ),
    .Y(_0303_),
    .A1(_0299_),
    .A2(_0302_));
 sg13g2_mux4_1 _4752_ (.S0(net1666),
    .A0(net1921),
    .A1(net41),
    .A2(net154),
    .A3(net1703),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0304_));
 sg13g2_mux4_1 _4753_ (.S0(net1666),
    .A0(net1712),
    .A1(net118),
    .A2(net134),
    .A3(net94),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0305_));
 sg13g2_mux2_1 _4754_ (.A0(_0305_),
    .A1(_0304_),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ),
    .X(_0306_));
 sg13g2_nand2b_1 _4755_ (.Y(_0307_),
    .B(_0306_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_o21ai_1 _4756_ (.B1(_0307_),
    .Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .A1(_0303_),
    .A2(_0296_));
 sg13g2_mux4_1 _4757_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net133),
    .A1(net93),
    .A2(net158),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0308_));
 sg13g2_mux4_1 _4758_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(net1528),
    .A1(net1534),
    .A2(net1543),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0309_));
 sg13g2_nand2b_1 _4759_ (.Y(_0310_),
    .B(_0067_),
    .A_N(_0309_));
 sg13g2_mux2_1 _4760_ (.A0(net1561),
    .A1(net1569),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0311_));
 sg13g2_mux2_1 _4761_ (.A0(net1578),
    .A1(net1615),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0312_));
 sg13g2_a21oi_2 _4762_ (.B1(_0067_),
    .Y(_0313_),
    .A2(_0312_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_o21ai_1 _4763_ (.B1(_0313_),
    .Y(_0314_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .A2(_0311_));
 sg13g2_nand3_1 _4764_ (.B(_0310_),
    .C(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .A(_0314_),
    .Y(_0315_));
 sg13g2_mux4_1 _4765_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(net1711),
    .A1(net119),
    .A2(net95),
    .A3(net1923),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0316_));
 sg13g2_mux2_1 _4766_ (.A0(net155),
    .A1(net167),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .X(_0317_));
 sg13g2_nor2b_1 _4767_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .B_N(net42),
    .Y(_0318_));
 sg13g2_a21oi_1 _4768_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ),
    .A2(net50),
    .Y(_0319_),
    .B1(_0318_));
 sg13g2_a21oi_1 _4769_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .A2(_0317_),
    .Y(_0320_),
    .B1(_0067_));
 sg13g2_o21ai_1 _4770_ (.B1(_0320_),
    .Y(_0321_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ),
    .A2(_0319_));
 sg13g2_o21ai_1 _4771_ (.B1(_0321_),
    .Y(_0322_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0316_));
 sg13g2_o21ai_1 _4772_ (.B1(_0315_),
    .Y(_0323_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0322_));
 sg13g2_inv_4 _4773_ (.A(net713),
    .Y(_0324_));
 sg13g2_o21ai_1 _4774_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .Y(_0325_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(_0324_));
 sg13g2_a21o_1 _4775_ (.A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A1(_0308_),
    .B1(_0325_),
    .X(_0326_));
 sg13g2_mux4_1 _4776_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(net1543),
    .A1(_0289_),
    .A2(net710),
    .A3(_0308_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .X(_0327_));
 sg13g2_o21ai_1 _4777_ (.B1(_0326_),
    .Y(_0328_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ),
    .A2(_0292_));
 sg13g2_a21oi_1 _4778_ (.A1(_0069_),
    .A2(net1692),
    .Y(_0329_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_o21ai_1 _4779_ (.B1(_0329_),
    .Y(_0330_),
    .A1(net1692),
    .A2(_0327_));
 sg13g2_mux2_1 _4780_ (.A0(net1),
    .A1(net4),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0331_));
 sg13g2_a21oi_1 _4781_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0331_),
    .Y(_0332_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_mux4_1 _4782_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .A0(net26),
    .A1(net30),
    .A2(net62),
    .A3(net1932),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0333_));
 sg13g2_inv_1 _4783_ (.Y(_0334_),
    .A(_0333_));
 sg13g2_a221oi_1 _4784_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .B1(_0334_),
    .A1(_0330_),
    .Y(_0335_),
    .A2(_0332_));
 sg13g2_nand2_1 _4785_ (.Y(_0336_),
    .A(net1692),
    .B(net1590));
 sg13g2_o21ai_1 _4786_ (.B1(_0336_),
    .Y(_0337_),
    .A1(net1692),
    .A2(net1631));
 sg13g2_mux2_1 _4787_ (.A0(net1584),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .S(net1692),
    .X(_0338_));
 sg13g2_o21ai_1 _4788_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ),
    .Y(_0339_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0337_));
 sg13g2_a21o_1 _4789_ (.A2(_0338_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .B1(_0339_),
    .X(_0340_));
 sg13g2_nand2b_1 _4790_ (.Y(_0341_),
    .B(net1692),
    .A_N(net1614));
 sg13g2_o21ai_1 _4791_ (.B1(_0341_),
    .Y(_0342_),
    .A1(net1692),
    .A2(net1601));
 sg13g2_mux2_1 _4792_ (.A0(net1607),
    .A1(net1622),
    .S(net1692),
    .X(_0343_));
 sg13g2_a21oi_1 _4793_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0343_),
    .Y(_0344_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_o21ai_1 _4794_ (.B1(_0344_),
    .Y(_0345_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0342_));
 sg13g2_nand3_1 _4795_ (.B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ),
    .C(_0345_),
    .A(_0340_),
    .Y(_0346_));
 sg13g2_nor2b_2 _4796_ (.A(_0335_),
    .B_N(_0346_),
    .Y(_0347_));
 sg13g2_inv_4 _4797_ (.A(_0347_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ));
 sg13g2_mux4_1 _4798_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(net1706),
    .A1(net106),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .A3(net166),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0348_));
 sg13g2_mux4_1 _4799_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net1528),
    .A1(net1534),
    .A2(net1542),
    .A3(net1557),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0349_));
 sg13g2_nand2b_1 _4800_ (.Y(_0350_),
    .B(_0349_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_nor2_1 _4801_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .B(net1563),
    .Y(_0351_));
 sg13g2_a21oi_1 _4802_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(net1569),
    .Y(_0352_),
    .B1(_0351_));
 sg13g2_nand2b_1 _4803_ (.Y(_0353_),
    .B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A_N(net1617));
 sg13g2_o21ai_1 _4804_ (.B1(_0353_),
    .Y(_0354_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(net1578));
 sg13g2_o21ai_1 _4805_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0355_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0352_));
 sg13g2_a21oi_1 _4806_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0354_),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_nor2b_1 _4807_ (.A(_0356_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0357_));
 sg13g2_mux4_1 _4808_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net42),
    .A1(net50),
    .A2(net155),
    .A3(net171),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0358_));
 sg13g2_mux4_1 _4809_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ),
    .A0(net119),
    .A1(net95),
    .A2(net1926),
    .A3(net1923),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0359_));
 sg13g2_nand2b_1 _4810_ (.Y(_0360_),
    .B(_0359_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_a21oi_1 _4811_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0358_),
    .Y(_0361_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_a22oi_1 _4812_ (.Y(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .B1(_0360_),
    .B2(_0361_),
    .A2(_0357_),
    .A1(_0350_));
 sg13g2_mux4_1 _4813_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net132),
    .A1(net59),
    .A2(net155),
    .A3(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0362_));
 sg13g2_nand2b_1 _4814_ (.Y(_0363_),
    .B(net1578),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_nand2_2 _4815_ (.Y(_0364_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .B(net1617));
 sg13g2_nand3_1 _4816_ (.B(_0364_),
    .C(_0363_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0365_));
 sg13g2_a21oi_1 _4817_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(net1573),
    .Y(_0366_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_o21ai_1 _4818_ (.B1(_0366_),
    .Y(_0367_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(net1561));
 sg13g2_nand3_1 _4819_ (.B(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .C(_0367_),
    .A(_0365_),
    .Y(_0368_));
 sg13g2_mux4_1 _4820_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(net1534),
    .A1(net1542),
    .A2(net1549),
    .A3(net1557),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0369_));
 sg13g2_a21oi_1 _4821_ (.A1(_0071_),
    .A2(_0369_),
    .Y(_0370_),
    .B1(_0072_));
 sg13g2_mux4_1 _4822_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(net1936),
    .A1(net51),
    .A2(net152),
    .A3(net1703),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0371_));
 sg13g2_nand2_1 _4823_ (.Y(_0372_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ),
    .B(_0371_));
 sg13g2_mux4_1 _4824_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ),
    .A0(net1710),
    .A1(net92),
    .A2(net116),
    .A3(net1921),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0373_));
 sg13g2_a21oi_1 _4825_ (.A1(_0071_),
    .A2(_0373_),
    .Y(_0374_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_a22oi_1 _4826_ (.Y(_0375_),
    .B1(_0372_),
    .B2(_0374_),
    .A2(_0370_),
    .A1(_0368_));
 sg13g2_mux4_1 _4827_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ),
    .A0(net1549),
    .A1(net689),
    .A2(_0375_),
    .A3(_0362_),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ),
    .X(_0376_));
 sg13g2_a21oi_1 _4828_ (.A1(_0074_),
    .A2(net1683),
    .Y(_0377_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_o21ai_1 _4829_ (.B1(_0377_),
    .Y(_0378_),
    .A1(net1683),
    .A2(net1527));
 sg13g2_mux2_1 _4830_ (.A0(net138),
    .A1(net7),
    .S(net1683),
    .X(_0379_));
 sg13g2_a21oi_1 _4831_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0379_),
    .Y(_0380_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_mux4_1 _4832_ (.S0(net1683),
    .A0(net21),
    .A1(net33),
    .A2(net68),
    .A3(net82),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0381_));
 sg13g2_inv_1 _4833_ (.Y(_0382_),
    .A(_0381_));
 sg13g2_a221oi_1 _4834_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ),
    .B1(_0382_),
    .A1(_0378_),
    .Y(_0383_),
    .A2(_0380_));
 sg13g2_a21o_2 _4835_ (.A2(_0270_),
    .A1(_0264_),
    .B1(_0383_),
    .X(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ));
 sg13g2_inv_1 _4836_ (.Y(_0384_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ));
 sg13g2_mux4_1 _4837_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net137),
    .A1(net6),
    .A2(net72),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0385_));
 sg13g2_o21ai_1 _4838_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_0386_),
    .A1(net1684),
    .A2(_0175_));
 sg13g2_a21oi_2 _4839_ (.B1(_0386_),
    .Y(_0387_),
    .A2(net1539),
    .A1(net1685));
 sg13g2_nand2_1 _4840_ (.Y(_0388_),
    .A(net1684),
    .B(net1585));
 sg13g2_o21ai_1 _4841_ (.B1(_0388_),
    .Y(_0389_),
    .A1(net1684),
    .A2(net1590));
 sg13g2_o21ai_1 _4842_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .Y(_0390_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_0389_));
 sg13g2_or2_1 _4843_ (.X(_0391_),
    .B(_0387_),
    .A(_0390_));
 sg13g2_o21ai_1 _4844_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_0392_),
    .A1(net1685),
    .A2(_0177_));
 sg13g2_a21oi_1 _4845_ (.A1(net1685),
    .A2(net1633),
    .Y(_0393_),
    .B1(_0392_));
 sg13g2_mux2_1 _4846_ (.A0(net1597),
    .A1(net1611),
    .S(net1685),
    .X(_0394_));
 sg13g2_nor2_1 _4847_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_nor3_1 _4848_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .B(_0393_),
    .C(_0395_),
    .Y(_0396_));
 sg13g2_nor2b_1 _4849_ (.A(_0396_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .Y(_0397_));
 sg13g2_nand2b_1 _4850_ (.Y(_0398_),
    .B(net1684),
    .A_N(net8));
 sg13g2_o21ai_1 _4851_ (.B1(_0398_),
    .Y(_0399_),
    .A1(net1684),
    .A2(net135));
 sg13g2_mux2_1 _4852_ (.A0(net1516),
    .A1(net1708),
    .S(net1684),
    .X(_0400_));
 sg13g2_a21oi_1 _4853_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_0399_),
    .Y(_0401_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_o21ai_1 _4854_ (.B1(_0401_),
    .Y(_0402_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_0400_));
 sg13g2_nand2b_1 _4855_ (.Y(_0403_),
    .B(net1684),
    .A_N(net1929));
 sg13g2_o21ai_1 _4856_ (.B1(_0403_),
    .Y(_0404_),
    .A1(net1684),
    .A2(net69));
 sg13g2_nand2_1 _4857_ (.Y(_0405_),
    .A(net1685),
    .B(net34));
 sg13g2_o21ai_1 _4858_ (.B1(_0405_),
    .Y(_0406_),
    .A1(net1685),
    .A2(_0059_));
 sg13g2_o21ai_1 _4859_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ),
    .Y(_0407_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_0406_));
 sg13g2_a21oi_1 _4860_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ),
    .A2(_0404_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_nor2_1 _4861_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ),
    .B(_0408_),
    .Y(_0409_));
 sg13g2_a22oi_1 _4862_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .B1(_0409_),
    .B2(_0402_),
    .A2(_0397_),
    .A1(_0391_));
 sg13g2_mux2_1 _4863_ (.A0(net647),
    .A1(_0385_),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_0410_));
 sg13g2_mux4_1 _4864_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ),
    .A0(net611),
    .A1(net1936),
    .A2(net13),
    .A3(net74),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ),
    .X(_0411_));
 sg13g2_inv_1 _4865_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_nand2_1 _4866_ (.Y(_0413_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .B(_0412_));
 sg13g2_nor2_1 _4867_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .B(net1629),
    .Y(_0414_));
 sg13g2_nor2_1 _4868_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_a22oi_1 _4869_ (.Y(_0416_),
    .B1(_0413_),
    .B2(_0415_),
    .A2(_0410_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ));
 sg13g2_mux4_1 _4870_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ),
    .A0(net1629),
    .A1(net647),
    .A2(_0411_),
    .A3(_0385_),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ),
    .X(_0417_));
 sg13g2_a21oi_1 _4871_ (.A1(net1662),
    .A2(_0077_),
    .Y(_0418_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_o21ai_1 _4872_ (.B1(_0418_),
    .Y(_0419_),
    .A1(net1662),
    .A2(_0417_));
 sg13g2_mux2_1 _4873_ (.A0(net147),
    .A1(net1705),
    .S(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0420_));
 sg13g2_a21oi_1 _4874_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0420_),
    .Y(_0421_),
    .B1(_0078_));
 sg13g2_mux4_1 _4875_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A0(net1713),
    .A1(net1928),
    .A2(net115),
    .A3(net107),
    .S1(net1662),
    .X(_0422_));
 sg13g2_o21ai_1 _4876_ (.B1(_0079_),
    .Y(_0423_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0422_));
 sg13g2_a21oi_2 _4877_ (.B1(_0423_),
    .Y(_0424_),
    .A2(_0419_),
    .A1(_0421_));
 sg13g2_mux2_1 _4878_ (.A0(_0171_),
    .A1(net1561),
    .S(net1662),
    .X(_0425_));
 sg13g2_mux2_1 _4879_ (.A0(net1574),
    .A1(net1619),
    .S(net1662),
    .X(_0426_));
 sg13g2_a21oi_1 _4880_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0426_),
    .Y(_0427_),
    .B1(_0078_));
 sg13g2_o21ai_1 _4881_ (.B1(_0427_),
    .Y(_0428_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0425_));
 sg13g2_nand2_1 _4882_ (.Y(_0429_),
    .A(net1662),
    .B(_0180_));
 sg13g2_o21ai_1 _4883_ (.B1(_0429_),
    .Y(_0430_),
    .A1(net1662),
    .A2(net1531));
 sg13g2_mux2_1 _4884_ (.A0(net1546),
    .A1(net1553),
    .S(net1662),
    .X(_0431_));
 sg13g2_a21oi_1 _4885_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0431_),
    .Y(_0432_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_o21ai_1 _4886_ (.B1(_0432_),
    .Y(_0433_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0430_));
 sg13g2_nand3_1 _4887_ (.B(_0428_),
    .C(_0433_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ),
    .Y(_0434_));
 sg13g2_nor2b_2 _4888_ (.A(_0424_),
    .B_N(_0434_),
    .Y(_0435_));
 sg13g2_inv_8 _4889_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .A(_0435_));
 sg13g2_a21oi_1 _4890_ (.A1(_0080_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .Y(_0436_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_o21ai_1 _4891_ (.B1(_0436_),
    .Y(_0437_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ));
 sg13g2_o21ai_1 _4892_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ),
    .Y(_0438_),
    .A1(net1934),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_a21o_1 _4893_ (.A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ),
    .A1(_0082_),
    .B1(_0438_),
    .X(_0439_));
 sg13g2_nand3_1 _4894_ (.B(_0437_),
    .C(_0439_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .Y(_0440_));
 sg13g2_mux4_1 _4895_ (.S0(net1677),
    .A0(net1599),
    .A1(net1612),
    .A2(net1605),
    .A3(net1625),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0441_));
 sg13g2_inv_1 _4896_ (.Y(_0442_),
    .A(_0441_));
 sg13g2_mux4_1 _4897_ (.S0(net1677),
    .A0(net1594),
    .A1(net1588),
    .A2(net1523),
    .A3(net1540),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0443_));
 sg13g2_o21ai_1 _4898_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .Y(_0444_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0442_));
 sg13g2_a21oi_1 _4899_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0443_),
    .Y(_0445_),
    .B1(_0444_));
 sg13g2_nand2b_1 _4900_ (.Y(_0446_),
    .B(net1527),
    .A_N(net1677));
 sg13g2_a21oi_1 _4901_ (.A1(net128),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .Y(_0447_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_nor2b_1 _4902_ (.A(net1677),
    .B_N(net2004),
    .Y(_0448_));
 sg13g2_a21oi_1 _4903_ (.A1(net9),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_a221oi_1 _4904_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .C1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ),
    .B1(_0449_),
    .A1(_0446_),
    .Y(_0450_),
    .A2(_0447_));
 sg13g2_nand2b_1 _4905_ (.Y(_0451_),
    .B(net27),
    .A_N(net1677));
 sg13g2_a21oi_1 _4906_ (.A1(net35),
    .A2(net1677),
    .Y(_0452_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_nand2b_1 _4907_ (.Y(_0453_),
    .B(net1677),
    .A_N(net1930));
 sg13g2_o21ai_1 _4908_ (.B1(_0453_),
    .Y(_0454_),
    .A1(net1933),
    .A2(net1677));
 sg13g2_a221oi_1 _4909_ (.B2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ),
    .C1(_0112_),
    .B1(_0454_),
    .A1(_0451_),
    .Y(_0455_),
    .A2(_0452_));
 sg13g2_nor3_1 _4910_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ),
    .B(_0450_),
    .C(_0455_),
    .Y(_0456_));
 sg13g2_nor2_1 _4911_ (.A(_0445_),
    .B(_0456_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ));
 sg13g2_mux4_1 _4912_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ),
    .A0(net18),
    .A1(net79),
    .A2(net44),
    .A3(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ),
    .X(_0457_));
 sg13g2_nor2_1 _4913_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_nor2_1 _4914_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_a21oi_2 _4915_ (.B1(_0259_),
    .Y(_0460_),
    .A2(_0440_),
    .A1(_0459_));
 sg13g2_inv_1 _4916_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .A(net707));
 sg13g2_nand2_2 _4917_ (.Y(_0461_),
    .A(net1640),
    .B(_0460_));
 sg13g2_o21ai_1 _4918_ (.B1(_0461_),
    .Y(_0462_),
    .A1(_0123_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ));
 sg13g2_o21ai_1 _4919_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_0463_),
    .A1(net38),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_a21oi_1 _4920_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .A2(_0193_),
    .Y(_0464_),
    .B1(_0463_));
 sg13g2_mux4_1 _4921_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(net1534),
    .A1(net1542),
    .A2(net1549),
    .A3(net1556),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0465_));
 sg13g2_nand2b_1 _4922_ (.Y(_0466_),
    .B(_0465_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_nor2_1 _4923_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .B(net1563),
    .Y(_0467_));
 sg13g2_a21oi_1 _4924_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(net1569),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_nand2_1 _4925_ (.Y(_0469_),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .B(_0178_));
 sg13g2_o21ai_1 _4926_ (.B1(_0469_),
    .Y(_0470_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(net1577));
 sg13g2_o21ai_1 _4927_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .Y(_0471_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .A2(_0468_));
 sg13g2_a21oi_2 _4928_ (.B1(_0471_),
    .Y(_0472_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .A1(_0470_));
 sg13g2_nor2b_1 _4929_ (.A(_0472_),
    .B_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ),
    .Y(_0473_));
 sg13g2_mux4_1 _4930_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(net116),
    .A1(net132),
    .A2(net1925),
    .A3(net92),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0474_));
 sg13g2_nand2b_1 _4931_ (.Y(_0475_),
    .B(_0474_),
    .A_N(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_mux4_1 _4932_ (.S0(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ),
    .A0(net1921),
    .A1(net152),
    .A2(net59),
    .A3(net1703),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ),
    .X(_0476_));
 sg13g2_a21oi_1 _4933_ (.A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_0476_),
    .Y(_0477_),
    .B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_a22oi_1 _4934_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .B1(_0475_),
    .B2(_0477_),
    .A2(_0466_),
    .A1(_0473_));
 sg13g2_nor2_1 _4935_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .Y(_0478_));
 sg13g2_nor2b_1 _4936_ (.A(net12),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ),
    .Y(_0479_));
 sg13g2_nor3_1 _4937_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_0478_),
    .C(_0479_),
    .Y(_0480_));
 sg13g2_nor3_1 _4938_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .B(_0464_),
    .C(_0480_),
    .Y(_0481_));
 sg13g2_nand2b_1 _4939_ (.Y(_0482_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A_N(net13));
 sg13g2_o21ai_1 _4940_ (.B1(_0482_),
    .Y(_0483_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .A2(net612));
 sg13g2_mux2_1 _4941_ (.A0(net1936),
    .A1(net74),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_0484_));
 sg13g2_o21ai_1 _4942_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .Y(_0485_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0483_));
 sg13g2_a21oi_1 _4943_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_0484_),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_nor3_1 _4944_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .B(_0481_),
    .C(_0486_),
    .Y(_0487_));
 sg13g2_mux4_1 _4945_ (.S0(net1695),
    .A0(net1598),
    .A1(net1603),
    .A2(net1623),
    .A3(net1633),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0488_));
 sg13g2_nor2_1 _4946_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0488_),
    .Y(_0489_));
 sg13g2_nand2b_1 _4947_ (.Y(_0490_),
    .B(net1695),
    .A_N(net1587));
 sg13g2_o21ai_1 _4948_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net1695),
    .A2(net1591));
 sg13g2_o21ai_1 _4949_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0492_),
    .A1(net1695),
    .A2(net1522));
 sg13g2_a21oi_1 _4950_ (.A1(net1695),
    .A2(_0179_),
    .Y(_0493_),
    .B1(_0492_));
 sg13g2_o21ai_1 _4951_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0494_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0491_));
 sg13g2_o21ai_1 _4952_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ),
    .Y(_0495_),
    .A1(_0494_),
    .A2(_0493_));
 sg13g2_nor2_1 _4953_ (.A(net1696),
    .B(net687),
    .Y(_0496_));
 sg13g2_a21oi_1 _4954_ (.A1(net125),
    .A2(net1696),
    .Y(_0497_),
    .B1(_0496_));
 sg13g2_o21ai_1 _4955_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0498_),
    .A1(net6),
    .A2(net1695));
 sg13g2_a21oi_1 _4956_ (.A1(_0059_),
    .A2(net1696),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_nor2_1 _4957_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_o21ai_1 _4958_ (.B1(_0500_),
    .Y(_0501_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0497_));
 sg13g2_a21oi_1 _4959_ (.A1(_0062_),
    .A2(net1696),
    .Y(_0502_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_o21ai_1 _4960_ (.B1(_0502_),
    .Y(_0503_),
    .A1(net1695),
    .A2(net32));
 sg13g2_mux2_1 _4961_ (.A0(net67),
    .A1(net1929),
    .S(net1695),
    .X(_0504_));
 sg13g2_nand2_1 _4962_ (.Y(_0505_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_0504_));
 sg13g2_nand3_1 _4963_ (.B(_0503_),
    .C(_0505_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0506_));
 sg13g2_nand3b_1 _4964_ (.B(_0501_),
    .C(_0506_),
    .Y(_0507_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_o21ai_1 _4965_ (.B1(_0507_),
    .Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .A1(_0489_),
    .A2(_0495_));
 sg13g2_mux2_1 _4966_ (.A0(net46),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_0508_));
 sg13g2_a21oi_1 _4967_ (.A1(_0059_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ),
    .Y(_0509_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_o21ai_1 _4968_ (.B1(_0509_),
    .Y(_0510_),
    .A1(net135),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_nand2_1 _4969_ (.Y(_0511_),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .B(_0510_));
 sg13g2_a21oi_2 _4970_ (.B1(_0511_),
    .Y(_0512_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ),
    .A1(_0508_));
 sg13g2_mux4_1 _4971_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ),
    .A0(net1709),
    .A1(net4),
    .A2(net30),
    .A3(net86),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ),
    .X(_0513_));
 sg13g2_o21ai_1 _4972_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_0514_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0513_));
 sg13g2_nor2_2 _4973_ (.A(_0514_),
    .B(_0512_),
    .Y(_0515_));
 sg13g2_nor2_2 _4974_ (.A(_0487_),
    .B(_0515_),
    .Y(_0516_));
 sg13g2_inv_1 _4975_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .A(_0516_));
 sg13g2_nor2_2 _4976_ (.A(net1641),
    .B(_0516_),
    .Y(_0517_));
 sg13g2_a21oi_2 _4977_ (.B1(_0517_),
    .Y(_0518_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ),
    .A1(net1641));
 sg13g2_nor2_1 _4978_ (.A(net1511),
    .B(net1515),
    .Y(_0519_));
 sg13g2_o21ai_1 _4979_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ),
    .Y(_0520_),
    .A1(net82),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_a21o_1 _4980_ (.A2(net695),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .B1(_0520_),
    .X(_0521_));
 sg13g2_a21oi_1 _4981_ (.A1(_0075_),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ),
    .Y(_0522_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_o21ai_1 _4982_ (.B1(_0522_),
    .Y(_0523_),
    .A1(net136),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_and2_1 _4983_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_0523_),
    .X(_0524_));
 sg13g2_mux4_1 _4984_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(net1708),
    .A1(net34),
    .A2(net22),
    .A3(net69),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0525_));
 sg13g2_o21ai_1 _4985_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_0526_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0525_));
 sg13g2_a21o_1 _4986_ (.A2(_0524_),
    .A1(_0521_),
    .B1(_0526_),
    .X(_0527_));
 sg13g2_mux4_1 _4987_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net1596),
    .A1(net1609),
    .A2(net1602),
    .A3(net1630),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0528_));
 sg13g2_nand2b_1 _4988_ (.Y(_0529_),
    .B(_0528_),
    .A_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_mux2_1 _4989_ (.A0(net1592),
    .A1(net1584),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0530_));
 sg13g2_nand2b_1 _4990_ (.Y(_0531_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .A_N(net1518));
 sg13g2_o21ai_1 _4991_ (.B1(_0531_),
    .Y(_0532_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(net1521));
 sg13g2_o21ai_1 _4992_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0533_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0530_));
 sg13g2_a21oi_2 _4993_ (.B1(_0533_),
    .Y(_0534_),
    .A2(_0532_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_nor2b_1 _4994_ (.A(_0534_),
    .B_N(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0535_));
 sg13g2_nand2_1 _4995_ (.Y(_0536_),
    .A(_0059_),
    .B(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_o21ai_1 _4996_ (.B1(_0536_),
    .Y(_0537_),
    .A1(net8),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_mux2_1 _4997_ (.A0(net1708),
    .A1(net2003),
    .S(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0538_));
 sg13g2_a21oi_1 _4998_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0537_),
    .Y(_0539_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_o21ai_1 _4999_ (.B1(_0539_),
    .Y(_0540_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0538_));
 sg13g2_mux4_1 _5000_ (.S0(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ),
    .A0(net34),
    .A1(net69),
    .A2(net46),
    .A3(net85),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0541_));
 sg13g2_a21oi_1 _5001_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0541_),
    .Y(_0542_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_a22oi_1 _5002_ (.Y(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .B1(_0540_),
    .B2(_0542_),
    .A2(_0529_),
    .A1(_0535_));
 sg13g2_o21ai_1 _5003_ (.B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ),
    .Y(_0543_),
    .A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .A2(_0111_));
 sg13g2_a21oi_1 _5004_ (.A1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ),
    .A2(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .Y(_0544_),
    .B1(_0543_));
 sg13g2_mux4_1 _5005_ (.S0(net1660),
    .A0(net1532),
    .A1(net1536),
    .A2(net1545),
    .A3(net1552),
    .S1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0545_));
 sg13g2_mux2_1 _5006_ (.A0(net1561),
    .A1(net1571),
    .S(net1660),
    .X(_0546_));
 sg13g2_o21ai_1 _5007_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0547_),
    .A1(net1660),
    .A2(net1581));
 sg13g2_a21oi_1 _5008_ (.A1(net1660),
    .A2(_0178_),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_o21ai_1 _5009_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0549_),
    .A1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ),
    .A2(_0546_));
 sg13g2_nor2_1 _5010_ (.A(_0548_),
    .B(_0549_),
    .Y(_0550_));
 sg13g2_o21ai_1 _5011_ (.B1(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ),
    .Y(_0551_),
    .A1(_0545_),
    .A2(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_nor2_2 _5012_ (.A(_0550_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_mux4_1 _5013_ (.S0(net1681),
    .A0(net1609),
    .A1(net1602),
    .A2(net1621),
    .A3(net1629),
    .S1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0553_));
 sg13g2_nand2_2 _5014_ (.Y(_0554_),
    .A(_0553_),
    .B(_0108_));
 sg13g2_a21oi_1 _5015_ (.A1(net1680),
    .A2(net1583),
    .Y(_0555_),
    .B1(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_o21ai_1 _5016_ (.B1(_0555_),
    .Y(_0556_),
    .A1(net1680),
    .A2(net1590));
 sg13g2_nand2b_1 _5017_ (.Y(_0557_),
    .B(net1681),
    .A_N(net1518));
 sg13g2_dlhq_1 _5018_ (.D(net1951),
    .GATE(net1852),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dlhq_1 _5019_ (.D(net1953),
    .GATE(net1853),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _5020_ (.D(net1957),
    .GATE(net1853),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _5021_ (.D(net1959),
    .GATE(net1853),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _5022_ (.D(net1962),
    .GATE(net1855),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _5023_ (.D(net1963),
    .GATE(net1855),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _5024_ (.D(net1965),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _5025_ (.D(net1968),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _5026_ (.D(net1969),
    .GATE(net1852),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _5027_ (.D(net1971),
    .GATE(net1852),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _5028_ (.D(net1974),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _5029_ (.D(net1976),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _5030_ (.D(net1980),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _5031_ (.D(net1982),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _5032_ (.D(net1983),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _5033_ (.D(net1985),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _5034_ (.D(net1987),
    .GATE(net1853),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _5035_ (.D(net1989),
    .GATE(net1852),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _5036_ (.D(net1992),
    .GATE(net1849),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _5037_ (.D(net1994),
    .GATE(net1849),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _5038_ (.D(net1995),
    .GATE(net1852),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _5039_ (.D(net1997),
    .GATE(net1852),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _5040_ (.D(net1938),
    .GATE(net1855),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _5041_ (.D(net1939),
    .GATE(net1854),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _5042_ (.D(net1941),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _5043_ (.D(net1943),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _5044_ (.D(net1945),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _5045_ (.D(net1947),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _5046_ (.D(net1949),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _5047_ (.D(net1955),
    .GATE(net1851),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _5048_ (.D(net1977),
    .GATE(net1853),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _5049_ (.D(net1999),
    .GATE(net1853),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _5050_ (.D(net1952),
    .GATE(net1807),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _5051_ (.D(net1954),
    .GATE(net1807),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _5052_ (.D(net1958),
    .GATE(net1807),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _5053_ (.D(net1960),
    .GATE(net1807),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _5054_ (.D(net1961),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _5055_ (.D(net1964),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _5056_ (.D(net1965),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _5057_ (.D(net1967),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _5058_ (.D(net1970),
    .GATE(net1808),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _5059_ (.D(net1972),
    .GATE(net1808),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _5060_ (.D(net1973),
    .GATE(net1808),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _5061_ (.D(net1975),
    .GATE(net1808),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _5062_ (.D(net1980),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _5063_ (.D(net1982),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _5064_ (.D(net1984),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _5065_ (.D(net1986),
    .GATE(net1809),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _5066_ (.D(net1988),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _5067_ (.D(net1990),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _5068_ (.D(net1991),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _5069_ (.D(net1993),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _5070_ (.D(net1995),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _5071_ (.D(net1997),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _5072_ (.D(net1937),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _5073_ (.D(net1939),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _5074_ (.D(net1942),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _5075_ (.D(net1944),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _5076_ (.D(net1946),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _5077_ (.D(net1948),
    .GATE(net1806),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _5078_ (.D(net1949),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _5079_ (.D(net1955),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _5080_ (.D(net1977),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _5081_ (.D(net1999),
    .GATE(net1810),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _5082_ (.D(net1951),
    .GATE(net1797),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _5083_ (.D(net1953),
    .GATE(net1797),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _5084_ (.D(net1957),
    .GATE(net1797),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _5085_ (.D(net1959),
    .GATE(net1797),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _5086_ (.D(net1961),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _5087_ (.D(net1963),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _5088_ (.D(net1965),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _5089_ (.D(net1967),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _5090_ (.D(net1970),
    .GATE(net1799),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _5091_ (.D(net1971),
    .GATE(net1799),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _5092_ (.D(net1973),
    .GATE(net1799),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _5093_ (.D(net1975),
    .GATE(net1799),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _5094_ (.D(net1979),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _5095_ (.D(net1981),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _5096_ (.D(net1983),
    .GATE(net1799),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _5097_ (.D(net1986),
    .GATE(net1798),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _5098_ (.D(net1987),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _5099_ (.D(net1989),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _5100_ (.D(net1991),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _5101_ (.D(net1993),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _5102_ (.D(net1995),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _5103_ (.D(net1997),
    .GATE(net1797),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _5104_ (.D(net1937),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _5105_ (.D(net1939),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _5106_ (.D(net1941),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _5107_ (.D(net1943),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _5108_ (.D(net1945),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _5109_ (.D(net1947),
    .GATE(net1795),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _5110_ (.D(net1949),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _5111_ (.D(net1955),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _5112_ (.D(net1977),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _5113_ (.D(net1999),
    .GATE(net1796),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _5114_ (.D(net1952),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _5115_ (.D(net1954),
    .GATE(net1788),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _5116_ (.D(net1958),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _5117_ (.D(net1960),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _5118_ (.D(net1962),
    .GATE(net1788),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _5119_ (.D(net1964),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _5120_ (.D(net1966),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _5121_ (.D(net1967),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _5122_ (.D(net1970),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _5123_ (.D(net1972),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _5124_ (.D(net1973),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _5125_ (.D(net1975),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _5126_ (.D(net1979),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _5127_ (.D(net1981),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _5128_ (.D(net1984),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _5129_ (.D(net1985),
    .GATE(net1787),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _5130_ (.D(net1987),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _5131_ (.D(net1989),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _5132_ (.D(net1991),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _5133_ (.D(net1993),
    .GATE(net1785),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _5134_ (.D(net1995),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _5135_ (.D(net1997),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _5136_ (.D(net1938),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _5137_ (.D(net1939),
    .GATE(net1786),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _5138_ (.D(net1941),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _5139_ (.D(net1943),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _5140_ (.D(net1945),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _5141_ (.D(net1947),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _5142_ (.D(net1949),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _5143_ (.D(net1955),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _5144_ (.D(net1977),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _5145_ (.D(net1999),
    .GATE(net1789),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _5146_ (.D(net1952),
    .GATE(net1779),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _5147_ (.D(net1954),
    .GATE(net1779),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _5148_ (.D(net1958),
    .GATE(net1776),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _5149_ (.D(net1960),
    .GATE(net1776),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _5150_ (.D(net1961),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _5151_ (.D(net1964),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _5152_ (.D(net1965),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _5153_ (.D(net1967),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _5154_ (.D(net1970),
    .GATE(net1776),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _5155_ (.D(net1972),
    .GATE(net1776),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _5156_ (.D(net1973),
    .GATE(net1776),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _5157_ (.D(net1975),
    .GATE(net1776),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _5158_ (.D(net1980),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _5159_ (.D(net1982),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _5160_ (.D(net1983),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _5161_ (.D(net1985),
    .GATE(net1778),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _5162_ (.D(net1987),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _5163_ (.D(net1989),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _5164_ (.D(net1991),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _5165_ (.D(net1993),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _5166_ (.D(net1996),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _5167_ (.D(net1997),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _5168_ (.D(net1938),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _5169_ (.D(net1940),
    .GATE(net1775),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _5170_ (.D(net1942),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _5171_ (.D(net1944),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _5172_ (.D(net1946),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _5173_ (.D(net1948),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _5174_ (.D(net1950),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _5175_ (.D(net1956),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _5176_ (.D(net1978),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _5177_ (.D(net1999),
    .GATE(net1777),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _5178_ (.D(net1951),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _5179_ (.D(net1953),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _5180_ (.D(net1957),
    .GATE(net1768),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _5181_ (.D(net1959),
    .GATE(net1768),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _5182_ (.D(net1961),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _5183_ (.D(net1964),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _5184_ (.D(net1965),
    .GATE(net1767),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _5185_ (.D(net1967),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _5186_ (.D(net1969),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _5187_ (.D(net1971),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _5188_ (.D(net1974),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _5189_ (.D(net1976),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _5190_ (.D(net1980),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _5191_ (.D(net1982),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _5192_ (.D(net1983),
    .GATE(net1767),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _5193_ (.D(net1985),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _5194_ (.D(net1987),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _5195_ (.D(net1989),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _5196_ (.D(net1991),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _5197_ (.D(net1993),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _5198_ (.D(net1995),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _5199_ (.D(net1997),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _5200_ (.D(net1937),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _5201_ (.D(net1940),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _5202_ (.D(net1941),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _5203_ (.D(net1943),
    .GATE(net1763),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _5204_ (.D(net1946),
    .GATE(net1765),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _5205_ (.D(net1948),
    .GATE(net1765),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _5206_ (.D(net1949),
    .GATE(net1765),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _5207_ (.D(net1955),
    .GATE(net1764),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _5208_ (.D(net1978),
    .GATE(net1767),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _5209_ (.D(net2000),
    .GATE(net1766),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _5210_ (.D(net1951),
    .GATE(net1753),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _5211_ (.D(net1953),
    .GATE(net1756),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _5212_ (.D(net1957),
    .GATE(net1753),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _5213_ (.D(net1959),
    .GATE(net1753),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _5214_ (.D(net1962),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _5215_ (.D(net1963),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _5216_ (.D(net1965),
    .GATE(net1755),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _5217_ (.D(net1967),
    .GATE(net1755),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _5218_ (.D(net1969),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _5219_ (.D(net1971),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _5220_ (.D(net1974),
    .GATE(net1753),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _5221_ (.D(net1976),
    .GATE(net1753),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _5222_ (.D(net1979),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _5223_ (.D(net1981),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _5224_ (.D(net1984),
    .GATE(net1752),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _5225_ (.D(net1986),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _5226_ (.D(net1987),
    .GATE(net1756),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _5227_ (.D(net1989),
    .GATE(net1756),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _5228_ (.D(net1992),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _5229_ (.D(net1994),
    .GATE(net1753),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _5230_ (.D(net1996),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _5231_ (.D(net1998),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _5232_ (.D(net1937),
    .GATE(net1756),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _5233_ (.D(net1939),
    .GATE(net1756),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _5234_ (.D(net1941),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _5235_ (.D(net1943),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _5236_ (.D(net1945),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _5237_ (.D(net1947),
    .GATE(net1751),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _5238_ (.D(net1950),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _5239_ (.D(net1956),
    .GATE(net1754),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _5240_ (.D(net1978),
    .GATE(net1755),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _5241_ (.D(net2000),
    .GATE(net1755),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _5242_ (.D(net1951),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _5243_ (.D(net1953),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _5244_ (.D(net1957),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _5245_ (.D(net1959),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _5246_ (.D(net1962),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _5247_ (.D(net1963),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _5248_ (.D(net1966),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _5249_ (.D(net1968),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _5250_ (.D(net1969),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _5251_ (.D(net1971),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _5252_ (.D(net1974),
    .GATE(net1741),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _5253_ (.D(net1976),
    .GATE(net1741),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _5254_ (.D(net1979),
    .GATE(net1743),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _5255_ (.D(net1981),
    .GATE(net1743),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _5256_ (.D(net1983),
    .GATE(net1744),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _5257_ (.D(net1985),
    .GATE(net1744),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _5258_ (.D(net1987),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _5259_ (.D(net1989),
    .GATE(net1745),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _5260_ (.D(net1992),
    .GATE(net1740),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _5261_ (.D(net1994),
    .GATE(net1740),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _5262_ (.D(net1996),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _5263_ (.D(net1998),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _5264_ (.D(net1937),
    .GATE(net1743),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _5265_ (.D(net1940),
    .GATE(net1743),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _5266_ (.D(net1941),
    .GATE(net1740),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _5267_ (.D(net1943),
    .GATE(net1740),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _5268_ (.D(net1945),
    .GATE(net1740),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _5269_ (.D(net1947),
    .GATE(net1740),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _5270_ (.D(net1949),
    .GATE(net1744),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _5271_ (.D(net1955),
    .GATE(net1744),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _5272_ (.D(net1977),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _5273_ (.D(net2000),
    .GATE(net1742),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _5274_ (.D(net1951),
    .GATE(net1733),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _5275_ (.D(net1953),
    .GATE(net1733),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _5276_ (.D(net1957),
    .GATE(net1733),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _5277_ (.D(net1960),
    .GATE(net1732),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _5278_ (.D(net1961),
    .GATE(net1732),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _5279_ (.D(net1963),
    .GATE(net1732),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _5280_ (.D(net1965),
    .GATE(net1730),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _5281_ (.D(net1967),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _5282_ (.D(net1969),
    .GATE(net1730),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _5283_ (.D(net1971),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _5284_ (.D(net1973),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _5285_ (.D(net1975),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _5286_ (.D(net1979),
    .GATE(net1732),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _5287_ (.D(net1981),
    .GATE(net1732),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _5288_ (.D(net1984),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _5289_ (.D(net1986),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _5290_ (.D(net1988),
    .GATE(net1730),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _5291_ (.D(net1990),
    .GATE(net1730),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _5292_ (.D(net1992),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _5293_ (.D(net1994),
    .GATE(net1732),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _5294_ (.D(net1995),
    .GATE(net1733),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _5295_ (.D(net1997),
    .GATE(net1733),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _5296_ (.D(net1937),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _5297_ (.D(net1939),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _5298_ (.D(net1941),
    .GATE(net1728),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _5299_ (.D(net1943),
    .GATE(net1727),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _5300_ (.D(net1946),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _5301_ (.D(net1948),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _5302_ (.D(net1950),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _5303_ (.D(net1956),
    .GATE(net1731),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _5304_ (.D(net1977),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _5305_ (.D(net1999),
    .GATE(net1729),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _5306_ (.D(net1951),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _5307_ (.D(net1953),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _5308_ (.D(net1957),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _5309_ (.D(net1959),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _5310_ (.D(net1962),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _5311_ (.D(net1963),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _5312_ (.D(net1966),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _5313_ (.D(net1968),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _5314_ (.D(net1970),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _5315_ (.D(net1971),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _5316_ (.D(net1974),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_dlhq_1 _5317_ (.D(net1976),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_dlhq_1 _5318_ (.D(net1980),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19.Q ));
 sg13g2_dlhq_1 _5319_ (.D(net1982),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_dlhq_1 _5320_ (.D(net1983),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17.Q ));
 sg13g2_dlhq_1 _5321_ (.D(net1985),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_dlhq_1 _5322_ (.D(net1988),
    .GATE(net1723),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_dlhq_1 _5323_ (.D(net1989),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_dlhq_1 _5324_ (.D(net1991),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_dlhq_1 _5325_ (.D(net1993),
    .GATE(net1722),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12.Q ));
 sg13g2_dlhq_1 _5326_ (.D(net1996),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_dlhq_1 _5327_ (.D(net1998),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10.Q ));
 sg13g2_dlhq_1 _5328_ (.D(net1938),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9.Q ));
 sg13g2_dlhq_1 _5329_ (.D(net1940),
    .GATE(net1720),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_dlhq_1 _5330_ (.D(net1942),
    .GATE(net1719),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7.Q ));
 sg13g2_dlhq_1 _5331_ (.D(net1944),
    .GATE(net1720),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6.Q ));
 sg13g2_dlhq_1 _5332_ (.D(net1945),
    .GATE(net1720),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5.Q ));
 sg13g2_dlhq_1 _5333_ (.D(net1947),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4.Q ));
 sg13g2_dlhq_1 _5334_ (.D(net1949),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3.Q ));
 sg13g2_dlhq_1 _5335_ (.D(net1955),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_dlhq_1 _5336_ (.D(net1977),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1.Q ));
 sg13g2_dlhq_1 _5337_ (.D(net1999),
    .GATE(net1721),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0.Q ));
 sg13g2_dlhq_1 _5338_ (.D(net1951),
    .GATE(net1840),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31.Q ));
 sg13g2_dlhq_1 _5339_ (.D(net1953),
    .GATE(net1840),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30.Q ));
 sg13g2_dlhq_1 _5340_ (.D(net1957),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29.Q ));
 sg13g2_dlhq_1 _5341_ (.D(net1959),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28.Q ));
 sg13g2_dlhq_1 _5342_ (.D(net1962),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27.Q ));
 sg13g2_dlhq_1 _5343_ (.D(net1963),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26.Q ));
 sg13g2_dlhq_1 _5344_ (.D(net1966),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25.Q ));
 sg13g2_dlhq_1 _5345_ (.D(net1968),
    .GATE(net1840),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24.Q ));
 sg13g2_dlhq_1 _5346_ (.D(net1969),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23.Q ));
 sg13g2_dlhq_1 _5347_ (.D(net1971),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22.Q ));
 sg13g2_dlhq_1 _5348_ (.D(net1974),
    .GATE(net1843),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21.Q ));
 sg13g2_dlhq_1 _5349_ (.D(net1976),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20.Q ));
 sg13g2_dlhq_1 _5350_ (.D(net1979),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19.Q ));
 sg13g2_dlhq_1 _5351_ (.D(net1981),
    .GATE(net1842),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18.Q ));
 sg13g2_dlhq_1 _5352_ (.D(net1984),
    .GATE(net1843),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17.Q ));
 sg13g2_dlhq_1 _5353_ (.D(net1986),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16.Q ));
 sg13g2_dlhq_1 _5354_ (.D(net1987),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15.Q ));
 sg13g2_dlhq_1 _5355_ (.D(net1990),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14.Q ));
 sg13g2_dlhq_1 _5356_ (.D(net1992),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13.Q ));
 sg13g2_dlhq_1 _5357_ (.D(net1994),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12.Q ));
 sg13g2_dlhq_1 _5358_ (.D(net1995),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11.Q ));
 sg13g2_dlhq_1 _5359_ (.D(net1998),
    .GATE(net1839),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10.Q ));
 sg13g2_dlhq_1 _5360_ (.D(net1937),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_dlhq_1 _5361_ (.D(net1939),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8.Q ));
 sg13g2_dlhq_1 _5362_ (.D(net1942),
    .GATE(net1843),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7.Q ));
 sg13g2_dlhq_1 _5363_ (.D(net1943),
    .GATE(net1843),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6.Q ));
 sg13g2_dlhq_1 _5364_ (.D(net1945),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5.Q ));
 sg13g2_dlhq_1 _5365_ (.D(net1947),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4.Q ));
 sg13g2_dlhq_1 _5366_ (.D(net1949),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3.Q ));
 sg13g2_dlhq_1 _5367_ (.D(net1955),
    .GATE(net1841),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2.Q ));
 sg13g2_dlhq_1 _5368_ (.D(net1978),
    .GATE(net1844),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_dlhq_1 _5369_ (.D(net2000),
    .GATE(net1844),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0.Q ));
 sg13g2_dlhq_1 _5370_ (.D(net1952),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31.Q ));
 sg13g2_dlhq_1 _5371_ (.D(net1954),
    .GATE(net1829),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30.Q ));
 sg13g2_dlhq_1 _5372_ (.D(net1958),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29.Q ));
 sg13g2_dlhq_1 _5373_ (.D(net1960),
    .GATE(net1830),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28.Q ));
 sg13g2_dlhq_1 _5374_ (.D(net1961),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27.Q ));
 sg13g2_dlhq_1 _5375_ (.D(net1964),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26.Q ));
 sg13g2_dlhq_1 _5376_ (.D(net1966),
    .GATE(net1829),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25.Q ));
 sg13g2_dlhq_1 _5377_ (.D(net1968),
    .GATE(net1829),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24.Q ));
 sg13g2_dlhq_1 _5378_ (.D(net1969),
    .GATE(net1829),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23.Q ));
 sg13g2_dlhq_1 _5379_ (.D(net1972),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_dlhq_1 _5380_ (.D(net1973),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_dlhq_1 _5381_ (.D(net1975),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20.Q ));
 sg13g2_dlhq_1 _5382_ (.D(net1979),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19.Q ));
 sg13g2_dlhq_1 _5383_ (.D(net1981),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18.Q ));
 sg13g2_dlhq_1 _5384_ (.D(net1983),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17.Q ));
 sg13g2_dlhq_1 _5385_ (.D(net1985),
    .GATE(net1828),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16.Q ));
 sg13g2_dlhq_1 _5386_ (.D(net1988),
    .GATE(net1829),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15.Q ));
 sg13g2_dlhq_1 _5387_ (.D(net1990),
    .GATE(net1829),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14.Q ));
 sg13g2_dlhq_1 _5388_ (.D(net1991),
    .GATE(net1831),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13.Q ));
 sg13g2_dlhq_1 _5389_ (.D(net1993),
    .GATE(net1831),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12.Q ));
 sg13g2_dlhq_1 _5390_ (.D(net1996),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11.Q ));
 sg13g2_dlhq_1 _5391_ (.D(net1998),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10.Q ));
 sg13g2_dlhq_1 _5392_ (.D(net1937),
    .GATE(net1831),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9.Q ));
 sg13g2_dlhq_1 _5393_ (.D(net1939),
    .GATE(net1831),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8.Q ));
 sg13g2_dlhq_1 _5394_ (.D(net1941),
    .GATE(net1831),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7.Q ));
 sg13g2_dlhq_1 _5395_ (.D(net1944),
    .GATE(net1831),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6.Q ));
 sg13g2_dlhq_1 _5396_ (.D(net1945),
    .GATE(net1830),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5.Q ));
 sg13g2_dlhq_1 _5397_ (.D(net1948),
    .GATE(net1830),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4.Q ));
 sg13g2_dlhq_1 _5398_ (.D(net1950),
    .GATE(net1830),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3.Q ));
 sg13g2_dlhq_1 _5399_ (.D(net1956),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2.Q ));
 sg13g2_dlhq_1 _5400_ (.D(net1977),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1.Q ));
 sg13g2_dlhq_1 _5401_ (.D(net1999),
    .GATE(net1827),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0.Q ));
 sg13g2_dlhq_1 _5402_ (.D(net1952),
    .GATE(net1818),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31.Q ));
 sg13g2_dlhq_1 _5403_ (.D(net1954),
    .GATE(net1818),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30.Q ));
 sg13g2_dlhq_1 _5404_ (.D(net1958),
    .GATE(net1818),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29.Q ));
 sg13g2_dlhq_1 _5405_ (.D(net1960),
    .GATE(net1820),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28.Q ));
 sg13g2_dlhq_1 _5406_ (.D(net1961),
    .GATE(net1820),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27.Q ));
 sg13g2_dlhq_1 _5407_ (.D(net1964),
    .GATE(net1818),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26.Q ));
 sg13g2_dlhq_1 _5408_ (.D(net1966),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25.Q ));
 sg13g2_dlhq_1 _5409_ (.D(net1968),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24.Q ));
 sg13g2_dlhq_1 _5410_ (.D(net1970),
    .GATE(net1818),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23.Q ));
 sg13g2_dlhq_1 _5411_ (.D(net1972),
    .GATE(net1818),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22.Q ));
 sg13g2_dlhq_1 _5412_ (.D(net1973),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21.Q ));
 sg13g2_dlhq_1 _5413_ (.D(net1975),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20.Q ));
 sg13g2_dlhq_1 _5414_ (.D(net1980),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19.Q ));
 sg13g2_dlhq_1 _5415_ (.D(net1982),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18.Q ));
 sg13g2_dlhq_1 _5416_ (.D(net1984),
    .GATE(net1819),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17.Q ));
 sg13g2_dlhq_1 _5417_ (.D(net1986),
    .GATE(net1819),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16.Q ));
 sg13g2_dlhq_1 _5418_ (.D(net1988),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15.Q ));
 sg13g2_dlhq_1 _5419_ (.D(net1990),
    .GATE(net1817),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14.Q ));
 sg13g2_dlhq_1 _5420_ (.D(net1991),
    .GATE(net1819),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13.Q ));
 sg13g2_dlhq_1 _5421_ (.D(net1993),
    .GATE(net1819),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12.Q ));
 sg13g2_dlhq_1 _5422_ (.D(net1995),
    .GATE(net1819),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11.Q ));
 sg13g2_dlhq_1 _5423_ (.D(net1997),
    .GATE(net1819),
    .Q(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10.Q ));
 sg13g2_dfrbp_1 _5424_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net574),
    .D(_0038_),
    .Q_N(_0024_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[0] ));
 sg13g2_dfrbp_1 _5425_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net573),
    .D(_0039_),
    .Q_N(_0022_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[1] ));
 sg13g2_dfrbp_1 _5426_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net572),
    .D(_0040_),
    .Q_N(_0020_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[2] ));
 sg13g2_dfrbp_1 _5427_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net571),
    .D(_0041_),
    .Q_N(_0018_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[3] ));
 sg13g2_dfrbp_1 _5428_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net570),
    .D(_0042_),
    .Q_N(_0016_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[4] ));
 sg13g2_dfrbp_1 _5429_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net569),
    .D(_0043_),
    .Q_N(_0014_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[5] ));
 sg13g2_dfrbp_1 _5430_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net568),
    .D(_0044_),
    .Q_N(_0012_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[6] ));
 sg13g2_dfrbp_1 _5431_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net567),
    .D(_0045_),
    .Q_N(_0010_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[7] ));
 sg13g2_dfrbp_1 _5432_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net566),
    .D(_0046_),
    .Q_N(_0008_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[8] ));
 sg13g2_dfrbp_1 _5433_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net565),
    .D(_0047_),
    .Q_N(_0006_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[9] ));
 sg13g2_dfrbp_1 _5434_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net564),
    .D(_0048_),
    .Q_N(_0004_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[10] ));
 sg13g2_dfrbp_1 _5435_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net563),
    .D(_0049_),
    .Q_N(_0002_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[11] ));
 sg13g2_dfrbp_1 _5436_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net562),
    .D(_0050_),
    .Q_N(_0000_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[12] ));
 sg13g2_dfrbp_1 _5437_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net561),
    .D(_0051_),
    .Q_N(_0026_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[13] ));
 sg13g2_dfrbp_1 _5438_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net560),
    .D(_0052_),
    .Q_N(_0028_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[14] ));
 sg13g2_dfrbp_1 _5439_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net559),
    .D(_0053_),
    .Q_N(_0030_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[15] ));
 sg13g2_dfrbp_1 _5440_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net558),
    .D(_0054_),
    .Q_N(_0032_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[16] ));
 sg13g2_dfrbp_1 _5441_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net557),
    .D(_0055_),
    .Q_N(_0034_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[17] ));
 sg13g2_dfrbp_1 _5442_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net556),
    .D(_0056_),
    .Q_N(_0036_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[18] ));
 sg13g2_dfrbp_1 _5443_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net575),
    .D(_0057_),
    .Q_N(_2395_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.ACC[19] ));
 sg13g2_dfrbp_1 _5444_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net576),
    .D(\Tile_X0Y1_DSP_bot.A0 ),
    .Q_N(_2396_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[0] ));
 sg13g2_dfrbp_1 _5445_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net577),
    .D(\Tile_X0Y1_DSP_bot.A1 ),
    .Q_N(_2397_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[1] ));
 sg13g2_dfrbp_1 _5446_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net578),
    .D(\Tile_X0Y1_DSP_bot.A2 ),
    .Q_N(_2398_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[2] ));
 sg13g2_dfrbp_1 _5447_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net579),
    .D(\Tile_X0Y1_DSP_bot.A3 ),
    .Q_N(_2399_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[3] ));
 sg13g2_dfrbp_1 _5448_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net580),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0.X ),
    .Q_N(_2400_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[4] ));
 sg13g2_dfrbp_1 _5449_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net581),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1.X ),
    .Q_N(_2401_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[5] ));
 sg13g2_dfrbp_1 _5450_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net582),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2.X ),
    .Q_N(_2402_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[6] ));
 sg13g2_dfrbp_1 _5451_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net583),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3.X ),
    .Q_N(_2403_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg[7] ));
 sg13g2_dfrbp_1 _5452_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net584),
    .D(\Tile_X0Y1_DSP_bot.B0 ),
    .Q_N(_2404_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[0] ));
 sg13g2_dfrbp_1 _5453_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net585),
    .D(\Tile_X0Y1_DSP_bot.B1 ),
    .Q_N(_2405_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[1] ));
 sg13g2_dfrbp_1 _5454_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net586),
    .D(\Tile_X0Y1_DSP_bot.B2 ),
    .Q_N(_2406_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[2] ));
 sg13g2_dfrbp_1 _5455_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net587),
    .D(\Tile_X0Y1_DSP_bot.B3 ),
    .Q_N(_2407_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[3] ));
 sg13g2_dfrbp_1 _5456_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net588),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4.X ),
    .Q_N(_2408_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[4] ));
 sg13g2_dfrbp_1 _5457_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net589),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5.X ),
    .Q_N(_2409_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[5] ));
 sg13g2_dfrbp_1 _5458_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net590),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6.X ),
    .Q_N(_2410_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[6] ));
 sg13g2_dfrbp_1 _5459_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net591),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7.X ),
    .Q_N(_2411_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg[7] ));
 sg13g2_dfrbp_1 _5460_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net592),
    .D(\Tile_X0Y1_DSP_bot.C0 ),
    .Q_N(_0025_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[0] ));
 sg13g2_dfrbp_1 _5461_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net593),
    .D(\Tile_X0Y1_DSP_bot.C1 ),
    .Q_N(_0023_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[1] ));
 sg13g2_dfrbp_1 _5462_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net594),
    .D(\Tile_X0Y1_DSP_bot.C2 ),
    .Q_N(_0021_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[2] ));
 sg13g2_dfrbp_1 _5463_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net595),
    .D(\Tile_X0Y1_DSP_bot.C3 ),
    .Q_N(_0019_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[3] ));
 sg13g2_dfrbp_1 _5464_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net596),
    .D(\Tile_X0Y1_DSP_bot.C4 ),
    .Q_N(_0017_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[4] ));
 sg13g2_dfrbp_1 _5465_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net597),
    .D(\Tile_X0Y1_DSP_bot.C5 ),
    .Q_N(_0015_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[5] ));
 sg13g2_dfrbp_1 _5466_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net598),
    .D(\Tile_X0Y1_DSP_bot.C6 ),
    .Q_N(_0013_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[6] ));
 sg13g2_dfrbp_1 _5467_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net599),
    .D(\Tile_X0Y1_DSP_bot.C7 ),
    .Q_N(_0011_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[7] ));
 sg13g2_dfrbp_1 _5468_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net600),
    .D(\Tile_X0Y1_DSP_bot.C8 ),
    .Q_N(_0009_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[8] ));
 sg13g2_dfrbp_1 _5469_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net601),
    .D(\Tile_X0Y1_DSP_bot.C9 ),
    .Q_N(_0007_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[9] ));
 sg13g2_dfrbp_1 _5470_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net602),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8.X ),
    .Q_N(_0005_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[10] ));
 sg13g2_dfrbp_1 _5471_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net603),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9.X ),
    .Q_N(_0003_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[11] ));
 sg13g2_dfrbp_1 _5472_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net604),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10.X ),
    .Q_N(_0001_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[12] ));
 sg13g2_dfrbp_1 _5473_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net605),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11.X ),
    .Q_N(_0027_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[13] ));
 sg13g2_dfrbp_1 _5474_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net606),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12.X ),
    .Q_N(_0029_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[14] ));
 sg13g2_dfrbp_1 _5475_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net607),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13.X ),
    .Q_N(_0031_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[15] ));
 sg13g2_dfrbp_1 _5476_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net608),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14.X ),
    .Q_N(_0033_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[16] ));
 sg13g2_dfrbp_1 _5477_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net609),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15.X ),
    .Q_N(_0035_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[17] ));
 sg13g2_dfrbp_1 _5478_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net554),
    .D(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X ),
    .Q_N(_0037_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[18] ));
 sg13g2_dfrbp_1 _5479_ (.CLK(Tile_X0Y1_UserCLK),
    .RESET_B(net555),
    .D(net709),
    .Q_N(_2394_),
    .Q(\Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg[19] ));
 sg13g2_dlhq_1 _5480_ (.D(net1870),
    .GATE(net1846),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dlhq_1 _5481_ (.D(net1872),
    .GATE(net1846),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _5482_ (.D(net1876),
    .GATE(net1847),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _5483_ (.D(net1878),
    .GATE(net1847),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _5484_ (.D(net1881),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _5485_ (.D(net1883),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _5486_ (.D(net1884),
    .GATE(net1849),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _5487_ (.D(net1886),
    .GATE(net1849),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _5488_ (.D(net1888),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _5489_ (.D(net1890),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _5490_ (.D(net1892),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _5491_ (.D(net1894),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _5492_ (.D(net1899),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _5493_ (.D(net1901),
    .GATE(net1846),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _5494_ (.D(net1903),
    .GATE(net1847),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _5495_ (.D(net1905),
    .GATE(net1847),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _5496_ (.D(net1907),
    .GATE(net1850),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _5497_ (.D(net1909),
    .GATE(net1850),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _5498_ (.D(net1911),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _5499_ (.D(net1913),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _5500_ (.D(net1915),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _5501_ (.D(net1917),
    .GATE(net1846),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _5502_ (.D(net1857),
    .GATE(net1849),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _5503_ (.D(net1859),
    .GATE(net1849),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _5504_ (.D(net1860),
    .GATE(net1849),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _5505_ (.D(net1862),
    .GATE(net1849),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _5506_ (.D(net1864),
    .GATE(net1848),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _5507_ (.D(net1866),
    .GATE(net1846),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _5508_ (.D(net1869),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _5509_ (.D(net1874),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _5510_ (.D(net1896),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _5511_ (.D(net1919),
    .GATE(net1845),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _5512_ (.D(net1871),
    .GATE(net1811),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _5513_ (.D(net1873),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _5514_ (.D(net1877),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _5515_ (.D(net1879),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _5516_ (.D(net1881),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _5517_ (.D(net1882),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _5518_ (.D(net1884),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _5519_ (.D(net1886),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _5520_ (.D(net1888),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _5521_ (.D(net1890),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _5522_ (.D(net1893),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _5523_ (.D(net1895),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _5524_ (.D(net1898),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _5525_ (.D(net1900),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _5526_ (.D(net1903),
    .GATE(net1805),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _5527_ (.D(net1904),
    .GATE(net1804),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _5528_ (.D(net1906),
    .GATE(net1802),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _5529_ (.D(net1908),
    .GATE(net1802),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _5530_ (.D(net1910),
    .GATE(net1802),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _5531_ (.D(net1912),
    .GATE(net1802),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _5532_ (.D(net1915),
    .GATE(net1803),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _5533_ (.D(net1917),
    .GATE(net1803),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _5534_ (.D(net1856),
    .GATE(net1803),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _5535_ (.D(net1858),
    .GATE(net1803),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _5536_ (.D(net1860),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _5537_ (.D(net1862),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _5538_ (.D(net1864),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _5539_ (.D(net1866),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _5540_ (.D(net1868),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _5541_ (.D(net1874),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _5542_ (.D(net1896),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _5543_ (.D(net1919),
    .GATE(net1801),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _5544_ (.D(net1870),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _5545_ (.D(net1872),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _5546_ (.D(net1877),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _5547_ (.D(net1878),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _5548_ (.D(net1880),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _5549_ (.D(net1882),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _5550_ (.D(net1884),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _5551_ (.D(net1886),
    .GATE(net1793),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _5552_ (.D(net1888),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _5553_ (.D(net1890),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _5554_ (.D(net1892),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _5555_ (.D(net1894),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _5556_ (.D(net1898),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _5557_ (.D(net1900),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _5558_ (.D(net1902),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _5559_ (.D(net1904),
    .GATE(net1794),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _5560_ (.D(net1906),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _5561_ (.D(net1908),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _5562_ (.D(net1910),
    .GATE(net1791),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _5563_ (.D(net1912),
    .GATE(net1791),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _5564_ (.D(net1915),
    .GATE(net1792),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _5565_ (.D(net1917),
    .GATE(net1792),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _5566_ (.D(net1856),
    .GATE(net1792),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _5567_ (.D(net1858),
    .GATE(net1792),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _5568_ (.D(net1860),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _5569_ (.D(net1862),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _5570_ (.D(net1864),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _5571_ (.D(net1866),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _5572_ (.D(net1868),
    .GATE(net1791),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _5573_ (.D(net1874),
    .GATE(net1791),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _5574_ (.D(net1896),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _5575_ (.D(net1919),
    .GATE(net1790),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _5576_ (.D(net1870),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _5577_ (.D(net1872),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _5578_ (.D(net1876),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _5579_ (.D(net1879),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _5580_ (.D(net1880),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _5581_ (.D(net1882),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _5582_ (.D(net1884),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _5583_ (.D(net1886),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _5584_ (.D(net1888),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _5585_ (.D(net1891),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _5586_ (.D(net1893),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _5587_ (.D(net1895),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _5588_ (.D(net1898),
    .GATE(net1784),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _5589_ (.D(net1901),
    .GATE(net1782),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _5590_ (.D(net1902),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _5591_ (.D(net1904),
    .GATE(net1783),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _5592_ (.D(net1906),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _5593_ (.D(net1908),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _5594_ (.D(net1910),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _5595_ (.D(net1912),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _5596_ (.D(net1915),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _5597_ (.D(net1917),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _5598_ (.D(net1856),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _5599_ (.D(net1858),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _5600_ (.D(net1861),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _5601_ (.D(net1863),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _5602_ (.D(net1865),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _5603_ (.D(net1867),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _5604_ (.D(net1868),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _5605_ (.D(net1874),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _5606_ (.D(net1896),
    .GATE(net1780),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _5607_ (.D(net1919),
    .GATE(net1781),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _5608_ (.D(net1871),
    .GATE(net1774),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _5609_ (.D(net1873),
    .GATE(net1774),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _5610_ (.D(net1877),
    .GATE(net1774),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _5611_ (.D(net1879),
    .GATE(net1774),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _5612_ (.D(net1880),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _5613_ (.D(net1882),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _5614_ (.D(net1884),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _5615_ (.D(net1886),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _5616_ (.D(net1889),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _5617_ (.D(net1890),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _5618_ (.D(net1893),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _5619_ (.D(net1895),
    .GATE(net1772),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _5620_ (.D(net1898),
    .GATE(net1773),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _5621_ (.D(net1900),
    .GATE(net1773),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _5622_ (.D(net1902),
    .GATE(net1773),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _5623_ (.D(net1904),
    .GATE(net1773),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _5624_ (.D(net1906),
    .GATE(net1770),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _5625_ (.D(net1908),
    .GATE(net1770),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _5626_ (.D(net1910),
    .GATE(net1770),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _5627_ (.D(net1912),
    .GATE(net1770),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _5628_ (.D(net1915),
    .GATE(net1771),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _5629_ (.D(net1917),
    .GATE(net1771),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _5630_ (.D(net1856),
    .GATE(net1771),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _5631_ (.D(net1858),
    .GATE(net1771),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _5632_ (.D(net1860),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _5633_ (.D(net1862),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _5634_ (.D(net1864),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _5635_ (.D(net1866),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _5636_ (.D(net1868),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _5637_ (.D(net1874),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _5638_ (.D(net1896),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _5639_ (.D(net1919),
    .GATE(net1769),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _5640_ (.D(net1870),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _5641_ (.D(net1872),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _5642_ (.D(net1876),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _5643_ (.D(net1878),
    .GATE(net1759),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _5644_ (.D(net1881),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _5645_ (.D(net1883),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _5646_ (.D(net1885),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _5647_ (.D(net1887),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _5648_ (.D(net1888),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _5649_ (.D(net1890),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _5650_ (.D(net1892),
    .GATE(net1759),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _5651_ (.D(net1894),
    .GATE(net1759),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _5652_ (.D(net1899),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _5653_ (.D(net1900),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _5654_ (.D(net1903),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _5655_ (.D(net1905),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _5656_ (.D(net1906),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _5657_ (.D(net1908),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _5658_ (.D(net1910),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _5659_ (.D(net1912),
    .GATE(net1758),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _5660_ (.D(net1915),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _5661_ (.D(net1917),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _5662_ (.D(net1857),
    .GATE(net1762),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _5663_ (.D(net1859),
    .GATE(net1762),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _5664_ (.D(net1861),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _5665_ (.D(net1863),
    .GATE(net1761),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _5666_ (.D(net1864),
    .GATE(net1759),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _5667_ (.D(net1866),
    .GATE(net1759),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _5668_ (.D(net1868),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _5669_ (.D(net1875),
    .GATE(net1760),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _5670_ (.D(net1897),
    .GATE(net1762),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _5671_ (.D(net1920),
    .GATE(net1762),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _5672_ (.D(net1871),
    .GATE(net1752),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _5673_ (.D(net1873),
    .GATE(net1752),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _5674_ (.D(net1876),
    .GATE(net1747),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _5675_ (.D(net1878),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _5676_ (.D(net1880),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _5677_ (.D(net1882),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _5678_ (.D(net1885),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _5679_ (.D(net1886),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _5680_ (.D(net1888),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _5681_ (.D(net1890),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _5682_ (.D(net1892),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _5683_ (.D(net1894),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _5684_ (.D(net1898),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _5685_ (.D(net1900),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _5686_ (.D(net1902),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _5687_ (.D(net1904),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _5688_ (.D(net1907),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _5689_ (.D(net1908),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _5690_ (.D(net1910),
    .GATE(net1747),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _5691_ (.D(net1913),
    .GATE(net1747),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _5692_ (.D(net1916),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _5693_ (.D(net1918),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _5694_ (.D(net1857),
    .GATE(net1750),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _5695_ (.D(net1859),
    .GATE(net1750),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _5696_ (.D(net1860),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _5697_ (.D(net1862),
    .GATE(net1749),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _5698_ (.D(net1865),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _5699_ (.D(net1866),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _5700_ (.D(net1868),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _5701_ (.D(net1874),
    .GATE(net1746),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _5702_ (.D(net1897),
    .GATE(net1748),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _5703_ (.D(net1920),
    .GATE(net1750),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _5704_ (.D(net1871),
    .GATE(net1740),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _5705_ (.D(net1873),
    .GATE(net1740),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _5706_ (.D(net1877),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _5707_ (.D(net1879),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _5708_ (.D(net1881),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _5709_ (.D(net1883),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _5710_ (.D(net1884),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _5711_ (.D(net1886),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _5712_ (.D(net1888),
    .GATE(net1736),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _5713_ (.D(net1890),
    .GATE(net1736),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _5714_ (.D(net1892),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _5715_ (.D(net1894),
    .GATE(net1736),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _5716_ (.D(net1899),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _5717_ (.D(net1901),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _5718_ (.D(net1903),
    .GATE(net1738),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _5719_ (.D(net1905),
    .GATE(net1738),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _5720_ (.D(net1906),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _5721_ (.D(net1909),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _5722_ (.D(net1910),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _5723_ (.D(net1912),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _5724_ (.D(net1916),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _5725_ (.D(net1918),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _5726_ (.D(net1857),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _5727_ (.D(net1859),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _5728_ (.D(net1860),
    .GATE(net1736),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _5729_ (.D(net1862),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _5730_ (.D(net1864),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _5731_ (.D(net1866),
    .GATE(net1735),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _5732_ (.D(net1869),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _5733_ (.D(net1875),
    .GATE(net1737),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _5734_ (.D(net1897),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _5735_ (.D(net1920),
    .GATE(net1739),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _5736_ (.D(net1870),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _5737_ (.D(net1872),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _5738_ (.D(net1876),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _5739_ (.D(net1878),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _5740_ (.D(net1880),
    .GATE(net1726),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _5741_ (.D(net1882),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _5742_ (.D(net1884),
    .GATE(net1726),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _5743_ (.D(net1886),
    .GATE(net1726),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _5744_ (.D(net1888),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _5745_ (.D(net1890),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _5746_ (.D(net1892),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _5747_ (.D(net1894),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _5748_ (.D(net1899),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _5749_ (.D(net1901),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _5750_ (.D(net1903),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _5751_ (.D(net1905),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _5752_ (.D(net1907),
    .GATE(net1728),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _5753_ (.D(net1909),
    .GATE(net1728),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _5754_ (.D(net1911),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _5755_ (.D(net1913),
    .GATE(net1727),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _5756_ (.D(net1916),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _5757_ (.D(net1918),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _5758_ (.D(net1856),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _5759_ (.D(net1858),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _5760_ (.D(net1861),
    .GATE(net1726),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _5761_ (.D(net1863),
    .GATE(net1726),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _5762_ (.D(net1865),
    .GATE(net1728),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _5763_ (.D(net1867),
    .GATE(net1728),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _5764_ (.D(net1868),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _5765_ (.D(net1874),
    .GATE(net1724),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _5766_ (.D(net1896),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _5767_ (.D(net1919),
    .GATE(net1725),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _5768_ (.D(net1871),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _5769_ (.D(net1873),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _5770_ (.D(net1877),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _5771_ (.D(net1879),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _5772_ (.D(net1880),
    .GATE(net1718),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _5773_ (.D(net1883),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _5774_ (.D(net1885),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _5775_ (.D(net1887),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _5776_ (.D(net1889),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _5777_ (.D(net1891),
    .GATE(net1718),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _5778_ (.D(net1892),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_dlhq_1 _5779_ (.D(net1894),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_dlhq_1 _5780_ (.D(net1898),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19.Q ));
 sg13g2_dlhq_1 _5781_ (.D(net1900),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_dlhq_1 _5782_ (.D(net1902),
    .GATE(net1715),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17.Q ));
 sg13g2_dlhq_1 _5783_ (.D(net1904),
    .GATE(net1715),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_dlhq_1 _5784_ (.D(net1906),
    .GATE(net1715),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_dlhq_1 _5785_ (.D(net1908),
    .GATE(net1715),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_dlhq_1 _5786_ (.D(net1910),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_dlhq_1 _5787_ (.D(net1912),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12.Q ));
 sg13g2_dlhq_1 _5788_ (.D(net1916),
    .GATE(net1715),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_dlhq_1 _5789_ (.D(net1918),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10.Q ));
 sg13g2_dlhq_1 _5790_ (.D(net1857),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9.Q ));
 sg13g2_dlhq_1 _5791_ (.D(net1859),
    .GATE(net1717),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_dlhq_1 _5792_ (.D(net1860),
    .GATE(net1715),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7.Q ));
 sg13g2_dlhq_1 _5793_ (.D(net1862),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6.Q ));
 sg13g2_dlhq_1 _5794_ (.D(net1864),
    .GATE(net1714),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5.Q ));
 sg13g2_dlhq_1 _5795_ (.D(net1866),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4.Q ));
 sg13g2_dlhq_1 _5796_ (.D(net1868),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3.Q ));
 sg13g2_dlhq_1 _5797_ (.D(net1874),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_dlhq_1 _5798_ (.D(net1896),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1.Q ));
 sg13g2_dlhq_1 _5799_ (.D(net1919),
    .GATE(net1716),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0.Q ));
 sg13g2_dlhq_1 _5800_ (.D(net1870),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31.Q ));
 sg13g2_dlhq_1 _5801_ (.D(net1872),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30.Q ));
 sg13g2_dlhq_1 _5802_ (.D(net1876),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29.Q ));
 sg13g2_dlhq_1 _5803_ (.D(net1878),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28.Q ));
 sg13g2_dlhq_1 _5804_ (.D(net1880),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27.Q ));
 sg13g2_dlhq_1 _5805_ (.D(net1882),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26.Q ));
 sg13g2_dlhq_1 _5806_ (.D(net1885),
    .GATE(net1838),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25.Q ));
 sg13g2_dlhq_1 _5807_ (.D(net1887),
    .GATE(net1835),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24.Q ));
 sg13g2_dlhq_1 _5808_ (.D(net1889),
    .GATE(net1838),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23.Q ));
 sg13g2_dlhq_1 _5809_ (.D(net1891),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22.Q ));
 sg13g2_dlhq_1 _5810_ (.D(net1893),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21.Q ));
 sg13g2_dlhq_1 _5811_ (.D(net1895),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20.Q ));
 sg13g2_dlhq_1 _5812_ (.D(net1898),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19.Q ));
 sg13g2_dlhq_1 _5813_ (.D(net1900),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18.Q ));
 sg13g2_dlhq_1 _5814_ (.D(net1902),
    .GATE(net1833),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17.Q ));
 sg13g2_dlhq_1 _5815_ (.D(net1905),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16.Q ));
 sg13g2_dlhq_1 _5816_ (.D(net1907),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15.Q ));
 sg13g2_dlhq_1 _5817_ (.D(net1909),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14.Q ));
 sg13g2_dlhq_1 _5818_ (.D(net1911),
    .GATE(net1835),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13.Q ));
 sg13g2_dlhq_1 _5819_ (.D(net1912),
    .GATE(net1835),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12.Q ));
 sg13g2_dlhq_1 _5820_ (.D(net1915),
    .GATE(net1834),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11.Q ));
 sg13g2_dlhq_1 _5821_ (.D(net1917),
    .GATE(net1834),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10.Q ));
 sg13g2_dlhq_1 _5822_ (.D(net1856),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_dlhq_1 _5823_ (.D(net1858),
    .GATE(net1834),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8.Q ));
 sg13g2_dlhq_1 _5824_ (.D(net1861),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7.Q ));
 sg13g2_dlhq_1 _5825_ (.D(net1863),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6.Q ));
 sg13g2_dlhq_1 _5826_ (.D(net1864),
    .GATE(net1834),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5.Q ));
 sg13g2_dlhq_1 _5827_ (.D(net1867),
    .GATE(net1836),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4.Q ));
 sg13g2_dlhq_1 _5828_ (.D(net1869),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3.Q ));
 sg13g2_dlhq_1 _5829_ (.D(net1875),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2.Q ));
 sg13g2_dlhq_1 _5830_ (.D(net1896),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_dlhq_1 _5831_ (.D(net1919),
    .GATE(net1837),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0.Q ));
 sg13g2_dlhq_1 _5832_ (.D(net1870),
    .GATE(net1826),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31.Q ));
 sg13g2_dlhq_1 _5833_ (.D(net1872),
    .GATE(net1826),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30.Q ));
 sg13g2_dlhq_1 _5834_ (.D(net1876),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29.Q ));
 sg13g2_dlhq_1 _5835_ (.D(net1878),
    .GATE(net1825),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28.Q ));
 sg13g2_dlhq_1 _5836_ (.D(net1881),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27.Q ));
 sg13g2_dlhq_1 _5837_ (.D(net1883),
    .GATE(net1825),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26.Q ));
 sg13g2_dlhq_1 _5838_ (.D(net1885),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25.Q ));
 sg13g2_dlhq_1 _5839_ (.D(net1887),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24.Q ));
 sg13g2_dlhq_1 _5840_ (.D(net1889),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23.Q ));
 sg13g2_dlhq_1 _5841_ (.D(net1891),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_dlhq_1 _5842_ (.D(net1893),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_dlhq_1 _5843_ (.D(net1895),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20.Q ));
 sg13g2_dlhq_1 _5844_ (.D(net1899),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19.Q ));
 sg13g2_dlhq_1 _5845_ (.D(net1901),
    .GATE(net1832),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18.Q ));
 sg13g2_dlhq_1 _5846_ (.D(net1902),
    .GATE(net1832),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17.Q ));
 sg13g2_dlhq_1 _5847_ (.D(net1904),
    .GATE(net1826),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16.Q ));
 sg13g2_dlhq_1 _5848_ (.D(net1907),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15.Q ));
 sg13g2_dlhq_1 _5849_ (.D(net1909),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14.Q ));
 sg13g2_dlhq_1 _5850_ (.D(net1911),
    .GATE(net1824),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13.Q ));
 sg13g2_dlhq_1 _5851_ (.D(net1914),
    .GATE(net1822),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12.Q ));
 sg13g2_dlhq_1 _5852_ (.D(net1915),
    .GATE(net1822),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11.Q ));
 sg13g2_dlhq_1 _5853_ (.D(net1917),
    .GATE(net1822),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10.Q ));
 sg13g2_dlhq_1 _5854_ (.D(net1856),
    .GATE(net1822),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9.Q ));
 sg13g2_dlhq_1 _5855_ (.D(net1858),
    .GATE(net1823),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8.Q ));
 sg13g2_dlhq_1 _5856_ (.D(net1861),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7.Q ));
 sg13g2_dlhq_1 _5857_ (.D(net1863),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6.Q ));
 sg13g2_dlhq_1 _5858_ (.D(net1865),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5.Q ));
 sg13g2_dlhq_1 _5859_ (.D(net1867),
    .GATE(net1821),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4.Q ));
 sg13g2_dlhq_1 _5860_ (.D(net1869),
    .GATE(net1823),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3.Q ));
 sg13g2_dlhq_1 _5861_ (.D(net1875),
    .GATE(net1823),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2.Q ));
 sg13g2_dlhq_1 _5862_ (.D(net1897),
    .GATE(net1826),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1.Q ));
 sg13g2_dlhq_1 _5863_ (.D(net1920),
    .GATE(net1826),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0.Q ));
 sg13g2_dlhq_1 _5864_ (.D(net1870),
    .GATE(net1815),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31.Q ));
 sg13g2_dlhq_1 _5865_ (.D(net1872),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30.Q ));
 sg13g2_dlhq_1 _5866_ (.D(net1876),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29.Q ));
 sg13g2_dlhq_1 _5867_ (.D(net1878),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28.Q ));
 sg13g2_dlhq_1 _5868_ (.D(net1880),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27.Q ));
 sg13g2_dlhq_1 _5869_ (.D(net1882),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26.Q ));
 sg13g2_dlhq_1 _5870_ (.D(net1884),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25.Q ));
 sg13g2_dlhq_1 _5871_ (.D(net1887),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24.Q ));
 sg13g2_dlhq_1 _5872_ (.D(net1889),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23.Q ));
 sg13g2_dlhq_1 _5873_ (.D(net1891),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22.Q ));
 sg13g2_dlhq_1 _5874_ (.D(net1892),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21.Q ));
 sg13g2_dlhq_1 _5875_ (.D(net1894),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20.Q ));
 sg13g2_dlhq_1 _5876_ (.D(net1898),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19.Q ));
 sg13g2_dlhq_1 _5877_ (.D(net1900),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18.Q ));
 sg13g2_dlhq_1 _5878_ (.D(net1902),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17.Q ));
 sg13g2_dlhq_1 _5879_ (.D(net1904),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16.Q ));
 sg13g2_dlhq_1 _5880_ (.D(net1906),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15.Q ));
 sg13g2_dlhq_1 _5881_ (.D(net1908),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14.Q ));
 sg13g2_dlhq_1 _5882_ (.D(net1911),
    .GATE(net1815),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13.Q ));
 sg13g2_dlhq_1 _5883_ (.D(net1914),
    .GATE(net1816),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12.Q ));
 sg13g2_dlhq_1 _5884_ (.D(net1916),
    .GATE(net1816),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11.Q ));
 sg13g2_dlhq_1 _5885_ (.D(net1918),
    .GATE(net1816),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10.Q ));
 sg13g2_dlhq_1 _5886_ (.D(net1856),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9.Q ));
 sg13g2_dlhq_1 _5887_ (.D(net1859),
    .GATE(net1812),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8.Q ));
 sg13g2_dlhq_1 _5888_ (.D(net1860),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7.Q ));
 sg13g2_dlhq_1 _5889_ (.D(net1862),
    .GATE(net1813),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6.Q ));
 sg13g2_dlhq_1 _5890_ (.D(net1865),
    .GATE(net1816),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ));
 sg13g2_dlhq_1 _5891_ (.D(net1867),
    .GATE(net1819),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4.Q ));
 sg13g2_dlhq_1 _5892_ (.D(net1869),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ));
 sg13g2_dlhq_1 _5893_ (.D(net1875),
    .GATE(net1814),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ));
 sg13g2_dlhq_1 _5894_ (.D(net1897),
    .GATE(net1816),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1.Q ));
 sg13g2_dlhq_1 _5895_ (.D(net1920),
    .GATE(net1816),
    .Q(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ));
 sg13g2_tiehi _5479__555 (.L_HI(net555));
 sg13g2_tiehi _5442__556 (.L_HI(net556));
 sg13g2_tiehi _5441__557 (.L_HI(net557));
 sg13g2_tiehi _5440__558 (.L_HI(net558));
 sg13g2_tiehi _5439__559 (.L_HI(net559));
 sg13g2_tiehi _5438__560 (.L_HI(net560));
 sg13g2_tiehi _5437__561 (.L_HI(net561));
 sg13g2_tiehi _5436__562 (.L_HI(net562));
 sg13g2_tiehi _5435__563 (.L_HI(net563));
 sg13g2_tiehi _5434__564 (.L_HI(net564));
 sg13g2_tiehi _5433__565 (.L_HI(net565));
 sg13g2_tiehi _5432__566 (.L_HI(net566));
 sg13g2_tiehi _5431__567 (.L_HI(net567));
 sg13g2_tiehi _5430__568 (.L_HI(net568));
 sg13g2_tiehi _5429__569 (.L_HI(net569));
 sg13g2_tiehi _5428__570 (.L_HI(net570));
 sg13g2_tiehi _5427__571 (.L_HI(net571));
 sg13g2_tiehi _5426__572 (.L_HI(net572));
 sg13g2_tiehi _5425__573 (.L_HI(net573));
 sg13g2_tiehi _5424__574 (.L_HI(net574));
 sg13g2_tiehi _5443__575 (.L_HI(net575));
 sg13g2_tiehi _5444__576 (.L_HI(net576));
 sg13g2_tiehi _5445__577 (.L_HI(net577));
 sg13g2_tiehi _5446__578 (.L_HI(net578));
 sg13g2_tiehi _5447__579 (.L_HI(net579));
 sg13g2_tiehi _5448__580 (.L_HI(net580));
 sg13g2_tiehi _5449__581 (.L_HI(net581));
 sg13g2_tiehi _5450__582 (.L_HI(net582));
 sg13g2_tiehi _5451__583 (.L_HI(net583));
 sg13g2_tiehi _5452__584 (.L_HI(net584));
 sg13g2_tiehi _5453__585 (.L_HI(net585));
 sg13g2_tiehi _5454__586 (.L_HI(net586));
 sg13g2_tiehi _5455__587 (.L_HI(net587));
 sg13g2_tiehi _5456__588 (.L_HI(net588));
 sg13g2_tiehi _5457__589 (.L_HI(net589));
 sg13g2_tiehi _5458__590 (.L_HI(net590));
 sg13g2_tiehi _5459__591 (.L_HI(net591));
 sg13g2_tiehi _5460__592 (.L_HI(net592));
 sg13g2_tiehi _5461__593 (.L_HI(net593));
 sg13g2_tiehi _5462__594 (.L_HI(net594));
 sg13g2_tiehi _5463__595 (.L_HI(net595));
 sg13g2_tiehi _5464__596 (.L_HI(net596));
 sg13g2_tiehi _5465__597 (.L_HI(net597));
 sg13g2_tiehi _5466__598 (.L_HI(net598));
 sg13g2_tiehi _5467__599 (.L_HI(net599));
 sg13g2_tiehi _5468__600 (.L_HI(net600));
 sg13g2_tiehi _5469__601 (.L_HI(net601));
 sg13g2_tiehi _5470__602 (.L_HI(net602));
 sg13g2_tiehi _5471__603 (.L_HI(net603));
 sg13g2_tiehi _5472__604 (.L_HI(net604));
 sg13g2_tiehi _5473__605 (.L_HI(net605));
 sg13g2_tiehi _5474__606 (.L_HI(net606));
 sg13g2_tiehi _5475__607 (.L_HI(net607));
 sg13g2_tiehi _5476__608 (.L_HI(net608));
 sg13g2_tiehi _5477__609 (.L_HI(net609));
 sg13g2_dlygate4sd1_1 rebuffer1 (.A(_0597_),
    .X(net610));
 sg13g2_dlygate4sd1_1 rebuffer119 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .X(net728));
 sg13g2_buf_2 rebuffer121 (.A(net731),
    .X(net730));
 sg13g2_buf_1 _5954_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG2 ),
    .X(net175));
 sg13g2_buf_8 _5955_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG3 ),
    .X(net176));
 sg13g2_buf_1 _5956_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG0 ),
    .X(net177));
 sg13g2_buf_1 _5957_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG1 ),
    .X(net178));
 sg13g2_buf_1 _5958_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG2 ),
    .X(net179));
 sg13g2_buf_1 _5959_ (.A(net706),
    .X(net180));
 sg13g2_buf_1 _5960_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG4 ),
    .X(net181));
 sg13g2_buf_1 _5961_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG5 ),
    .X(net182));
 sg13g2_buf_1 _5962_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG6 ),
    .X(net183));
 sg13g2_buf_8 _5963_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG7 ),
    .X(net184));
 sg13g2_buf_1 _5964_ (.A(net12),
    .X(net185));
 sg13g2_buf_1 _5965_ (.A(net13),
    .X(net186));
 sg13g2_buf_1 _5966_ (.A(net14),
    .X(net187));
 sg13g2_buf_1 _5967_ (.A(net15),
    .X(net188));
 sg13g2_buf_1 _5968_ (.A(net16),
    .X(net189));
 sg13g2_buf_1 _5969_ (.A(net17),
    .X(net190));
 sg13g2_buf_1 _5970_ (.A(net18),
    .X(net191));
 sg13g2_buf_1 _5971_ (.A(net19),
    .X(net192));
 sg13g2_buf_1 _5972_ (.A(Tile_X0Y0_E6END[2]),
    .X(net193));
 sg13g2_buf_1 _5973_ (.A(Tile_X0Y0_E6END[3]),
    .X(net196));
 sg13g2_buf_1 _5974_ (.A(Tile_X0Y0_E6END[4]),
    .X(net197));
 sg13g2_buf_1 _5975_ (.A(Tile_X0Y0_E6END[5]),
    .X(net198));
 sg13g2_buf_1 _5976_ (.A(Tile_X0Y0_E6END[6]),
    .X(net199));
 sg13g2_buf_1 _5977_ (.A(Tile_X0Y0_E6END[7]),
    .X(net200));
 sg13g2_buf_1 _5978_ (.A(Tile_X0Y0_E6END[8]),
    .X(net201));
 sg13g2_buf_1 _5979_ (.A(Tile_X0Y0_E6END[9]),
    .X(net202));
 sg13g2_buf_1 _5980_ (.A(Tile_X0Y0_E6END[10]),
    .X(net203));
 sg13g2_buf_1 _5981_ (.A(Tile_X0Y0_E6END[11]),
    .X(net204));
 sg13g2_buf_1 _5982_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG0 ),
    .X(net194));
 sg13g2_buf_1 _5983_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E6BEG1 ),
    .X(net195));
 sg13g2_buf_1 _5984_ (.A(Tile_X0Y0_EE4END[4]),
    .X(net205));
 sg13g2_buf_1 _5985_ (.A(Tile_X0Y0_EE4END[5]),
    .X(net212));
 sg13g2_buf_1 _5986_ (.A(Tile_X0Y0_EE4END[6]),
    .X(net213));
 sg13g2_buf_1 _5987_ (.A(Tile_X0Y0_EE4END[7]),
    .X(net214));
 sg13g2_buf_1 _5988_ (.A(Tile_X0Y0_EE4END[8]),
    .X(net215));
 sg13g2_buf_1 _5989_ (.A(Tile_X0Y0_EE4END[9]),
    .X(net216));
 sg13g2_buf_1 _5990_ (.A(Tile_X0Y0_EE4END[10]),
    .X(net217));
 sg13g2_buf_1 _5991_ (.A(Tile_X0Y0_EE4END[11]),
    .X(net218));
 sg13g2_buf_1 _5992_ (.A(Tile_X0Y0_EE4END[12]),
    .X(net219));
 sg13g2_buf_1 _5993_ (.A(Tile_X0Y0_EE4END[13]),
    .X(net220));
 sg13g2_buf_1 _5994_ (.A(Tile_X0Y0_EE4END[14]),
    .X(net206));
 sg13g2_buf_1 _5995_ (.A(Tile_X0Y0_EE4END[15]),
    .X(net207));
 sg13g2_buf_1 _5996_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG0 ),
    .X(net208));
 sg13g2_buf_1 _5997_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG1 ),
    .X(net209));
 sg13g2_buf_2 rebuffer125 (.A(net735),
    .X(net734));
 sg13g2_buf_8 _5999_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG3 ),
    .X(net211));
 sg13g2_buf_1 _6000_ (.A(net2000),
    .X(net221));
 sg13g2_buf_1 _6001_ (.A(net1978),
    .X(net232));
 sg13g2_buf_1 _6002_ (.A(net1956),
    .X(net243));
 sg13g2_buf_1 _6003_ (.A(net1950),
    .X(net246));
 sg13g2_buf_1 _6004_ (.A(net1947),
    .X(net247));
 sg13g2_buf_1 _6005_ (.A(net1946),
    .X(net248));
 sg13g2_buf_1 _6006_ (.A(net1944),
    .X(net249));
 sg13g2_buf_1 _6007_ (.A(net1942),
    .X(net250));
 sg13g2_buf_1 _6008_ (.A(net1940),
    .X(net251));
 sg13g2_buf_1 _6009_ (.A(net1938),
    .X(net252));
 sg13g2_buf_1 _6010_ (.A(net1998),
    .X(net222));
 sg13g2_buf_1 _6011_ (.A(net1996),
    .X(net223));
 sg13g2_buf_1 _6012_ (.A(net1994),
    .X(net224));
 sg13g2_buf_1 _6013_ (.A(net1992),
    .X(net225));
 sg13g2_buf_1 _6014_ (.A(net1990),
    .X(net226));
 sg13g2_buf_1 _6015_ (.A(net1988),
    .X(net227));
 sg13g2_buf_1 _6016_ (.A(net1985),
    .X(net228));
 sg13g2_buf_1 _6017_ (.A(net1983),
    .X(net229));
 sg13g2_buf_1 _6018_ (.A(net1981),
    .X(net230));
 sg13g2_buf_1 _6019_ (.A(net1979),
    .X(net231));
 sg13g2_buf_1 _6020_ (.A(net1975),
    .X(net233));
 sg13g2_buf_1 _6021_ (.A(net1973),
    .X(net234));
 sg13g2_buf_1 _6022_ (.A(net1972),
    .X(net235));
 sg13g2_buf_1 _6023_ (.A(net1969),
    .X(net236));
 sg13g2_buf_1 _6024_ (.A(net1967),
    .X(net237));
 sg13g2_buf_1 _6025_ (.A(net1965),
    .X(net238));
 sg13g2_buf_1 _6026_ (.A(net1963),
    .X(net239));
 sg13g2_buf_1 _6027_ (.A(net1961),
    .X(net240));
 sg13g2_buf_1 _6028_ (.A(net1959),
    .X(net241));
 sg13g2_buf_1 _6029_ (.A(net1958),
    .X(net242));
 sg13g2_buf_1 _6030_ (.A(net1954),
    .X(net244));
 sg13g2_buf_1 _6031_ (.A(net1952),
    .X(net245));
 sg13g2_buf_1 _6032_ (.A(net1854),
    .X(net253));
 sg13g2_buf_1 _6033_ (.A(net1811),
    .X(net264));
 sg13g2_buf_1 _6034_ (.A(net1798),
    .X(net265));
 sg13g2_buf_1 _6035_ (.A(net1787),
    .X(net266));
 sg13g2_buf_1 _6036_ (.A(net1779),
    .X(net267));
 sg13g2_buf_1 _6037_ (.A(net1767),
    .X(net268));
 sg13g2_buf_1 _6038_ (.A(net1755),
    .X(net269));
 sg13g2_buf_1 _6039_ (.A(net1743),
    .X(net270));
 sg13g2_buf_1 _6040_ (.A(net1731),
    .X(net271));
 sg13g2_buf_1 _6041_ (.A(net1722),
    .X(net272));
 sg13g2_buf_1 _6042_ (.A(net1844),
    .X(net254));
 sg13g2_buf_1 _6043_ (.A(net1830),
    .X(net255));
 sg13g2_buf_1 _6044_ (.A(net1818),
    .X(net256));
 sg13g2_buf_1 _6045_ (.A(Tile_X0Y1_FrameStrobe[13]),
    .X(net257));
 sg13g2_buf_1 _6046_ (.A(Tile_X0Y1_FrameStrobe[14]),
    .X(net258));
 sg13g2_buf_1 _6047_ (.A(Tile_X0Y1_FrameStrobe[15]),
    .X(net259));
 sg13g2_buf_1 _6048_ (.A(Tile_X0Y1_FrameStrobe[16]),
    .X(net260));
 sg13g2_buf_1 _6049_ (.A(Tile_X0Y1_FrameStrobe[17]),
    .X(net261));
 sg13g2_buf_1 _6050_ (.A(Tile_X0Y1_FrameStrobe[18]),
    .X(net262));
 sg13g2_buf_1 _6051_ (.A(Tile_X0Y1_FrameStrobe[19]),
    .X(net263));
 sg13g2_buf_1 _6052_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 ),
    .X(net273));
 sg13g2_buf_1 _6053_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 ),
    .X(net274));
 sg13g2_buf_8 rebuffer117 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net726));
 sg13g2_buf_8 _6055_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 ),
    .X(net276));
 sg13g2_buf_1 _6056_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 ),
    .X(net277));
 sg13g2_buf_1 _6057_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 ),
    .X(net278));
 sg13g2_buf_1 _6058_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 ),
    .X(net279));
 sg13g2_buf_1 _6059_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 ),
    .X(net280));
 sg13g2_buf_1 _6060_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 ),
    .X(net281));
 sg13g2_buf_1 _6061_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .X(net282));
 sg13g2_buf_1 _6062_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 ),
    .X(net283));
 sg13g2_buf_2 rebuffer123 (.A(net733),
    .X(net732));
 sg13g2_buf_1 _6064_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 ),
    .X(net285));
 sg13g2_buf_1 _6065_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 ),
    .X(net286));
 sg13g2_buf_8 _6066_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 ),
    .X(net287));
 sg13g2_buf_1 _6067_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 ),
    .X(net288));
 sg13g2_buf_8 _6068_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 ),
    .X(net289));
 sg13g2_buf_1 _6069_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 ),
    .X(net290));
 sg13g2_buf_1 _6070_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 ),
    .X(net291));
 sg13g2_buf_1 _6071_ (.A(net725),
    .X(net292));
 sg13g2_buf_1 _6072_ (.A(Tile_X0Y1_N4END[8]),
    .X(net293));
 sg13g2_buf_1 _6073_ (.A(Tile_X0Y1_N4END[9]),
    .X(net300));
 sg13g2_buf_1 _6074_ (.A(Tile_X0Y1_N4END[10]),
    .X(net301));
 sg13g2_buf_1 _6075_ (.A(Tile_X0Y1_N4END[11]),
    .X(net302));
 sg13g2_buf_1 _6076_ (.A(Tile_X0Y1_N4END[12]),
    .X(net303));
 sg13g2_buf_1 _6077_ (.A(Tile_X0Y1_N4END[13]),
    .X(net304));
 sg13g2_buf_1 _6078_ (.A(Tile_X0Y1_N4END[14]),
    .X(net305));
 sg13g2_buf_1 _6079_ (.A(Tile_X0Y1_N4END[15]),
    .X(net306));
 sg13g2_buf_1 _6080_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_8.A ),
    .X(net307));
 sg13g2_buf_1 _6081_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_9.A ),
    .X(net308));
 sg13g2_buf_1 _6082_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_10.A ),
    .X(net294));
 sg13g2_buf_1 _6083_ (.A(\Tile_X0Y0_DSP_top.N4BEG_outbuf_11.A ),
    .X(net295));
 sg13g2_buf_1 _6084_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 ),
    .X(net296));
 sg13g2_buf_1 _6085_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 ),
    .X(net297));
 sg13g2_buf_1 _6086_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 ),
    .X(net298));
 sg13g2_buf_1 _6087_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 ),
    .X(net299));
 sg13g2_buf_1 _6088_ (.A(Tile_X0Y1_NN4END[8]),
    .X(net309));
 sg13g2_buf_1 _6089_ (.A(Tile_X0Y1_NN4END[9]),
    .X(net316));
 sg13g2_buf_1 _6090_ (.A(Tile_X0Y1_NN4END[10]),
    .X(net317));
 sg13g2_buf_1 _6091_ (.A(Tile_X0Y1_NN4END[11]),
    .X(net318));
 sg13g2_buf_1 _6092_ (.A(Tile_X0Y1_NN4END[12]),
    .X(net319));
 sg13g2_buf_1 _6093_ (.A(Tile_X0Y1_NN4END[13]),
    .X(net320));
 sg13g2_buf_1 _6094_ (.A(Tile_X0Y1_NN4END[14]),
    .X(net321));
 sg13g2_buf_1 _6095_ (.A(Tile_X0Y1_NN4END[15]),
    .X(net322));
 sg13g2_buf_1 _6096_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_8.A ),
    .X(net323));
 sg13g2_buf_8 _6097_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_9.A ),
    .X(net324));
 sg13g2_buf_1 _6098_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_10.A ),
    .X(net310));
 sg13g2_buf_8 _6099_ (.A(\Tile_X0Y0_DSP_top.NN4BEG_outbuf_11.A ),
    .X(net311));
 sg13g2_buf_1 _6100_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 ),
    .X(net312));
 sg13g2_buf_2 _6101_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 ),
    .X(net313));
 sg13g2_buf_2 rebuffer124 (.A(net734),
    .X(net733));
 sg13g2_buf_2 rebuffer127 (.A(net737),
    .X(net736));
 sg13g2_buf_1 _6104_ (.A(Tile_X0Y1_UserCLK),
    .X(net325));
 sg13g2_buf_1 _6105_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 ),
    .X(net326));
 sg13g2_buf_1 _6106_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 ),
    .X(net327));
 sg13g2_buf_1 _6107_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 ),
    .X(net328));
 sg13g2_buf_1 _6108_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 ),
    .X(net329));
 sg13g2_buf_1 _6109_ (.A(net65),
    .X(net330));
 sg13g2_buf_1 _6110_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 ),
    .X(net331));
 sg13g2_buf_1 _6111_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 ),
    .X(net332));
 sg13g2_buf_1 _6112_ (.A(net68),
    .X(net333));
 sg13g2_buf_1 _6113_ (.A(net69),
    .X(net334));
 sg13g2_buf_1 _6114_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 ),
    .X(net335));
 sg13g2_buf_2 _6115_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .X(net336));
 sg13g2_buf_1 _6116_ (.A(net72),
    .X(net337));
 sg13g2_buf_1 _6117_ (.A(net73),
    .X(net338));
 sg13g2_buf_1 _6118_ (.A(net74),
    .X(net339));
 sg13g2_buf_1 _6119_ (.A(net75),
    .X(net340));
 sg13g2_buf_1 _6120_ (.A(net76),
    .X(net341));
 sg13g2_buf_1 _6121_ (.A(net77),
    .X(net342));
 sg13g2_buf_1 _6122_ (.A(net78),
    .X(net343));
 sg13g2_buf_1 _6123_ (.A(net79),
    .X(net344));
 sg13g2_buf_1 _6124_ (.A(net80),
    .X(net345));
 sg13g2_buf_1 _6125_ (.A(Tile_X0Y0_W6END[2]),
    .X(net346));
 sg13g2_buf_1 _6126_ (.A(Tile_X0Y0_W6END[3]),
    .X(net349));
 sg13g2_buf_1 _6127_ (.A(Tile_X0Y0_W6END[4]),
    .X(net350));
 sg13g2_buf_1 _6128_ (.A(Tile_X0Y0_W6END[5]),
    .X(net351));
 sg13g2_buf_1 _6129_ (.A(Tile_X0Y0_W6END[6]),
    .X(net352));
 sg13g2_buf_1 _6130_ (.A(Tile_X0Y0_W6END[7]),
    .X(net353));
 sg13g2_buf_1 _6131_ (.A(Tile_X0Y0_W6END[8]),
    .X(net354));
 sg13g2_buf_1 _6132_ (.A(Tile_X0Y0_W6END[9]),
    .X(net355));
 sg13g2_buf_1 _6133_ (.A(Tile_X0Y0_W6END[10]),
    .X(net356));
 sg13g2_buf_1 _6134_ (.A(Tile_X0Y0_W6END[11]),
    .X(net357));
 sg13g2_buf_1 _6135_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 ),
    .X(net347));
 sg13g2_buf_16 rebuffer39 (.X(net648),
    .A(net1607));
 sg13g2_buf_1 _6137_ (.A(Tile_X0Y0_WW4END[4]),
    .X(net358));
 sg13g2_buf_1 _6138_ (.A(Tile_X0Y0_WW4END[5]),
    .X(net365));
 sg13g2_buf_1 _6139_ (.A(Tile_X0Y0_WW4END[6]),
    .X(net366));
 sg13g2_buf_1 _6140_ (.A(Tile_X0Y0_WW4END[7]),
    .X(net367));
 sg13g2_buf_1 _6141_ (.A(Tile_X0Y0_WW4END[8]),
    .X(net368));
 sg13g2_buf_1 _6142_ (.A(Tile_X0Y0_WW4END[9]),
    .X(net369));
 sg13g2_buf_1 _6143_ (.A(Tile_X0Y0_WW4END[10]),
    .X(net370));
 sg13g2_buf_1 _6144_ (.A(Tile_X0Y0_WW4END[11]),
    .X(net371));
 sg13g2_buf_1 _6145_ (.A(Tile_X0Y0_WW4END[12]),
    .X(net372));
 sg13g2_buf_1 _6146_ (.A(Tile_X0Y0_WW4END[13]),
    .X(net373));
 sg13g2_buf_1 _6147_ (.A(Tile_X0Y0_WW4END[14]),
    .X(net359));
 sg13g2_buf_1 _6148_ (.A(Tile_X0Y0_WW4END[15]),
    .X(net360));
 sg13g2_buf_1 _6149_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 ),
    .X(net361));
 sg13g2_buf_2 _6150_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 ),
    .X(net362));
 sg13g2_buf_2 rebuffer122 (.A(net732),
    .X(net731));
 sg13g2_buf_8 _6152_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 ),
    .X(net364));
 sg13g2_buf_1 _6153_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG0 ),
    .X(net374));
 sg13g2_buf_1 _6154_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG1 ),
    .X(net375));
 sg13g2_buf_1 _6155_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG2 ),
    .X(net376));
 sg13g2_dlygate4sd1_1 rebuffer118 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 ),
    .X(net727));
 sg13g2_buf_1 _6157_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG0 ),
    .X(net378));
 sg13g2_buf_1 _6158_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG1 ),
    .X(net379));
 sg13g2_buf_1 _6159_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .X(net380));
 sg13g2_buf_1 _6160_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG3 ),
    .X(net381));
 sg13g2_buf_1 _6161_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG4 ),
    .X(net382));
 sg13g2_buf_1 _6162_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG5 ),
    .X(net383));
 sg13g2_buf_1 _6163_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG6 ),
    .X(net384));
 sg13g2_buf_8 _6164_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG7 ),
    .X(net385));
 sg13g2_buf_1 _6165_ (.A(net99),
    .X(net386));
 sg13g2_buf_1 _6166_ (.A(net100),
    .X(net387));
 sg13g2_buf_1 _6167_ (.A(net101),
    .X(net388));
 sg13g2_buf_1 _6168_ (.A(net102),
    .X(net389));
 sg13g2_buf_1 _6169_ (.A(net103),
    .X(net390));
 sg13g2_buf_1 _6170_ (.A(net104),
    .X(net391));
 sg13g2_buf_1 _6171_ (.A(net105),
    .X(net392));
 sg13g2_buf_1 _6172_ (.A(net106),
    .X(net393));
 sg13g2_buf_1 _6173_ (.A(Tile_X0Y1_E6END[2]),
    .X(net394));
 sg13g2_buf_1 _6174_ (.A(Tile_X0Y1_E6END[3]),
    .X(net397));
 sg13g2_buf_1 _6175_ (.A(Tile_X0Y1_E6END[4]),
    .X(net398));
 sg13g2_buf_1 _6176_ (.A(Tile_X0Y1_E6END[5]),
    .X(net399));
 sg13g2_buf_1 _6177_ (.A(Tile_X0Y1_E6END[6]),
    .X(net400));
 sg13g2_buf_1 _6178_ (.A(Tile_X0Y1_E6END[7]),
    .X(net401));
 sg13g2_buf_1 _6179_ (.A(Tile_X0Y1_E6END[8]),
    .X(net402));
 sg13g2_buf_1 _6180_ (.A(Tile_X0Y1_E6END[9]),
    .X(net403));
 sg13g2_buf_1 _6181_ (.A(Tile_X0Y1_E6END[10]),
    .X(net404));
 sg13g2_buf_1 _6182_ (.A(Tile_X0Y1_E6END[11]),
    .X(net405));
 sg13g2_buf_8 _6183_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG0 ),
    .X(net395));
 sg13g2_buf_1 _6184_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E6BEG1 ),
    .X(net396));
 sg13g2_buf_1 _6185_ (.A(Tile_X0Y1_EE4END[4]),
    .X(net406));
 sg13g2_buf_1 _6186_ (.A(Tile_X0Y1_EE4END[5]),
    .X(net413));
 sg13g2_buf_1 _6187_ (.A(Tile_X0Y1_EE4END[6]),
    .X(net414));
 sg13g2_buf_1 _6188_ (.A(Tile_X0Y1_EE4END[7]),
    .X(net415));
 sg13g2_buf_1 _6189_ (.A(Tile_X0Y1_EE4END[8]),
    .X(net416));
 sg13g2_buf_1 _6190_ (.A(Tile_X0Y1_EE4END[9]),
    .X(net417));
 sg13g2_buf_1 _6191_ (.A(Tile_X0Y1_EE4END[10]),
    .X(net418));
 sg13g2_buf_1 _6192_ (.A(Tile_X0Y1_EE4END[11]),
    .X(net419));
 sg13g2_buf_1 _6193_ (.A(Tile_X0Y1_EE4END[12]),
    .X(net420));
 sg13g2_buf_1 _6194_ (.A(Tile_X0Y1_EE4END[13]),
    .X(net421));
 sg13g2_buf_1 _6195_ (.A(Tile_X0Y1_EE4END[14]),
    .X(net407));
 sg13g2_buf_1 _6196_ (.A(Tile_X0Y1_EE4END[15]),
    .X(net408));
 sg13g2_buf_1 _6197_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG0 ),
    .X(net409));
 sg13g2_buf_1 _6198_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG1 ),
    .X(net410));
 sg13g2_buf_1 _6199_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG2 ),
    .X(net411));
 sg13g2_buf_1 _6200_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.EE4BEG3 ),
    .X(net412));
 sg13g2_buf_1 _6201_ (.A(net1920),
    .X(net422));
 sg13g2_buf_1 _6202_ (.A(net1897),
    .X(net433));
 sg13g2_buf_1 _6203_ (.A(net1875),
    .X(net444));
 sg13g2_buf_1 _6204_ (.A(net1869),
    .X(net447));
 sg13g2_buf_1 _6205_ (.A(net1867),
    .X(net448));
 sg13g2_buf_1 _6206_ (.A(net1865),
    .X(net449));
 sg13g2_buf_1 _6207_ (.A(net1863),
    .X(net450));
 sg13g2_buf_1 _6208_ (.A(net1861),
    .X(net451));
 sg13g2_buf_1 _6209_ (.A(net1858),
    .X(net452));
 sg13g2_buf_1 _6210_ (.A(net1857),
    .X(net453));
 sg13g2_buf_1 _6211_ (.A(net1918),
    .X(net423));
 sg13g2_buf_1 _6212_ (.A(net1916),
    .X(net424));
 sg13g2_buf_1 _6213_ (.A(net1914),
    .X(net425));
 sg13g2_buf_1 _6214_ (.A(net1911),
    .X(net426));
 sg13g2_buf_1 _6215_ (.A(net1909),
    .X(net427));
 sg13g2_buf_1 _6216_ (.A(net1907),
    .X(net428));
 sg13g2_buf_1 _6217_ (.A(net1905),
    .X(net429));
 sg13g2_buf_1 _6218_ (.A(net1903),
    .X(net430));
 sg13g2_buf_1 _6219_ (.A(net1901),
    .X(net431));
 sg13g2_buf_1 _6220_ (.A(net1899),
    .X(net432));
 sg13g2_buf_1 _6221_ (.A(net1895),
    .X(net434));
 sg13g2_buf_1 _6222_ (.A(net1893),
    .X(net435));
 sg13g2_buf_1 _6223_ (.A(net1891),
    .X(net436));
 sg13g2_buf_1 _6224_ (.A(net1889),
    .X(net437));
 sg13g2_buf_1 _6225_ (.A(net1887),
    .X(net438));
 sg13g2_buf_1 _6226_ (.A(net1885),
    .X(net439));
 sg13g2_buf_1 _6227_ (.A(net1883),
    .X(net440));
 sg13g2_buf_1 _6228_ (.A(net1881),
    .X(net441));
 sg13g2_buf_1 _6229_ (.A(net1879),
    .X(net442));
 sg13g2_buf_1 _6230_ (.A(net1877),
    .X(net443));
 sg13g2_buf_1 _6231_ (.A(net1873),
    .X(net445));
 sg13g2_buf_1 _6232_ (.A(net1871),
    .X(net446));
 sg13g2_buf_8 _6233_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 ),
    .X(net454));
 sg13g2_buf_8 _6234_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 ),
    .X(net455));
 sg13g2_buf_1 _6235_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 ),
    .X(net456));
 sg13g2_dlygate4sd1_1 rebuffer120 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 ),
    .X(net729));
 sg13g2_buf_1 _6237_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 ),
    .X(net458));
 sg13g2_buf_1 _6238_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .X(net459));
 sg13g2_buf_1 _6239_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .X(net460));
 sg13g2_buf_2 _6240_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 ),
    .X(net461));
 sg13g2_buf_2 _6241_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 ),
    .X(net462));
 sg13g2_buf_2 _6242_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 ),
    .X(net463));
 sg13g2_buf_2 _6243_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 ),
    .X(net464));
 sg13g2_buf_8 _6244_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 ),
    .X(net465));
 sg13g2_buf_1 _6245_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .X(net466));
 sg13g2_buf_1 _6246_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 ),
    .X(net467));
 sg13g2_buf_1 _6247_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .X(net468));
 sg13g2_buf_1 _6248_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .X(net469));
 sg13g2_buf_1 _6249_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .X(net470));
 sg13g2_buf_1 _6250_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 ),
    .X(net471));
 sg13g2_buf_1 _6251_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .X(net472));
 sg13g2_buf_1 _6252_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 ),
    .X(net473));
 sg13g2_buf_1 _6253_ (.A(Tile_X0Y0_S4END[8]),
    .X(net474));
 sg13g2_buf_1 _6254_ (.A(Tile_X0Y0_S4END[9]),
    .X(net481));
 sg13g2_buf_1 _6255_ (.A(Tile_X0Y0_S4END[10]),
    .X(net482));
 sg13g2_buf_1 _6256_ (.A(Tile_X0Y0_S4END[11]),
    .X(net483));
 sg13g2_buf_1 _6257_ (.A(Tile_X0Y0_S4END[12]),
    .X(net484));
 sg13g2_buf_1 _6258_ (.A(Tile_X0Y0_S4END[13]),
    .X(net485));
 sg13g2_buf_1 _6259_ (.A(Tile_X0Y0_S4END[14]),
    .X(net486));
 sg13g2_buf_1 _6260_ (.A(Tile_X0Y0_S4END[15]),
    .X(net487));
 sg13g2_buf_1 _6261_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0 ),
    .X(net488));
 sg13g2_buf_1 _6262_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1 ),
    .X(net489));
 sg13g2_buf_1 _6263_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2 ),
    .X(net475));
 sg13g2_buf_1 _6264_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3 ),
    .X(net476));
 sg13g2_buf_1 _6265_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 ),
    .X(net477));
 sg13g2_buf_1 _6266_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 ),
    .X(net478));
 sg13g2_buf_1 _6267_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 ),
    .X(net479));
 sg13g2_buf_1 _6268_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 ),
    .X(net480));
 sg13g2_buf_1 _6269_ (.A(Tile_X0Y0_SS4END[8]),
    .X(net490));
 sg13g2_buf_1 _6270_ (.A(Tile_X0Y0_SS4END[9]),
    .X(net497));
 sg13g2_buf_1 _6271_ (.A(Tile_X0Y0_SS4END[10]),
    .X(net498));
 sg13g2_buf_1 _6272_ (.A(Tile_X0Y0_SS4END[11]),
    .X(net499));
 sg13g2_buf_1 _6273_ (.A(Tile_X0Y0_SS4END[12]),
    .X(net500));
 sg13g2_buf_1 _6274_ (.A(Tile_X0Y0_SS4END[13]),
    .X(net501));
 sg13g2_buf_1 _6275_ (.A(Tile_X0Y0_SS4END[14]),
    .X(net502));
 sg13g2_buf_1 _6276_ (.A(Tile_X0Y0_SS4END[15]),
    .X(net503));
 sg13g2_buf_1 _6277_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 ),
    .X(net504));
 sg13g2_buf_8 _6278_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 ),
    .X(net505));
 sg13g2_buf_8 _6279_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 ),
    .X(net491));
 sg13g2_buf_8 _6280_ (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 ),
    .X(net492));
 sg13g2_buf_1 _6281_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 ),
    .X(net493));
 sg13g2_buf_8 _6282_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 ),
    .X(net494));
 sg13g2_buf_1 _6283_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 ),
    .X(net495));
 sg13g2_buf_1 _6284_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 ),
    .X(net496));
 sg13g2_buf_1 _6285_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 ),
    .X(net506));
 sg13g2_buf_8 _6286_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 ),
    .X(net507));
 sg13g2_buf_1 _6287_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 ),
    .X(net508));
 sg13g2_buf_2 rebuffer126 (.A(net736),
    .X(net735));
 sg13g2_buf_1 _6289_ (.A(net151),
    .X(net510));
 sg13g2_buf_1 _6290_ (.A(net646),
    .X(net511));
 sg13g2_buf_2 _6291_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 ),
    .X(net512));
 sg13g2_buf_1 _6292_ (.A(net154),
    .X(net513));
 sg13g2_buf_1 _6293_ (.A(net155),
    .X(net514));
 sg13g2_buf_8 _6294_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .X(net515));
 sg13g2_buf_2 _6295_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 ),
    .X(net516));
 sg13g2_buf_1 _6296_ (.A(net158),
    .X(net517));
 sg13g2_buf_1 _6297_ (.A(net159),
    .X(net518));
 sg13g2_buf_1 _6298_ (.A(net160),
    .X(net519));
 sg13g2_buf_1 _6299_ (.A(net161),
    .X(net520));
 sg13g2_buf_1 _6300_ (.A(net162),
    .X(net521));
 sg13g2_buf_1 _6301_ (.A(net163),
    .X(net522));
 sg13g2_buf_1 _6302_ (.A(net164),
    .X(net523));
 sg13g2_buf_1 _6303_ (.A(net165),
    .X(net524));
 sg13g2_buf_1 _6304_ (.A(net166),
    .X(net525));
 sg13g2_buf_1 _6305_ (.A(Tile_X0Y1_W6END[2]),
    .X(net526));
 sg13g2_buf_1 _6306_ (.A(Tile_X0Y1_W6END[3]),
    .X(net529));
 sg13g2_buf_1 _6307_ (.A(Tile_X0Y1_W6END[4]),
    .X(net530));
 sg13g2_buf_1 _6308_ (.A(Tile_X0Y1_W6END[5]),
    .X(net531));
 sg13g2_buf_1 _6309_ (.A(Tile_X0Y1_W6END[6]),
    .X(net532));
 sg13g2_buf_1 _6310_ (.A(Tile_X0Y1_W6END[7]),
    .X(net533));
 sg13g2_buf_1 _6311_ (.A(Tile_X0Y1_W6END[8]),
    .X(net534));
 sg13g2_buf_1 _6312_ (.A(Tile_X0Y1_W6END[9]),
    .X(net535));
 sg13g2_buf_1 _6313_ (.A(Tile_X0Y1_W6END[10]),
    .X(net536));
 sg13g2_buf_1 _6314_ (.A(Tile_X0Y1_W6END[11]),
    .X(net537));
 sg13g2_buf_1 _6315_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 ),
    .X(net527));
 sg13g2_buf_1 _6316_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 ),
    .X(net528));
 sg13g2_buf_1 _6317_ (.A(Tile_X0Y1_WW4END[4]),
    .X(net538));
 sg13g2_buf_1 _6318_ (.A(Tile_X0Y1_WW4END[5]),
    .X(net545));
 sg13g2_buf_1 _6319_ (.A(Tile_X0Y1_WW4END[6]),
    .X(net546));
 sg13g2_buf_1 _6320_ (.A(Tile_X0Y1_WW4END[7]),
    .X(net547));
 sg13g2_buf_1 _6321_ (.A(Tile_X0Y1_WW4END[8]),
    .X(net548));
 sg13g2_buf_1 _6322_ (.A(Tile_X0Y1_WW4END[9]),
    .X(net549));
 sg13g2_buf_1 _6323_ (.A(Tile_X0Y1_WW4END[10]),
    .X(net550));
 sg13g2_buf_1 _6324_ (.A(Tile_X0Y1_WW4END[11]),
    .X(net551));
 sg13g2_buf_1 _6325_ (.A(Tile_X0Y1_WW4END[12]),
    .X(net552));
 sg13g2_buf_1 _6326_ (.A(Tile_X0Y1_WW4END[13]),
    .X(net553));
 sg13g2_buf_1 _6327_ (.A(Tile_X0Y1_WW4END[14]),
    .X(net539));
 sg13g2_buf_1 _6328_ (.A(Tile_X0Y1_WW4END[15]),
    .X(net540));
 sg13g2_buf_1 _6329_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 ),
    .X(net541));
 sg13g2_buf_1 _6330_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 ),
    .X(net542));
 sg13g2_buf_1 _6331_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 ),
    .X(net543));
 sg13g2_buf_1 _6332_ (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 ),
    .X(net544));
 sg13g2_buf_8 fanout1511 (.A(_0462_),
    .X(net1511));
 sg13g2_buf_8 fanout1512 (.A(net1514),
    .X(net1512));
 sg13g2_buf_8 fanout1513 (.A(net1514),
    .X(net1513));
 sg13g2_buf_8 fanout1514 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr ),
    .X(net1514));
 sg13g2_buf_8 fanout1515 (.A(_0518_),
    .X(net1515));
 sg13g2_buf_8 fanout1516 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 ),
    .X(net1516));
 sg13g2_buf_1 fanout1517 (.A(_1724_),
    .X(net1517));
 sg13g2_buf_8 fanout1518 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 ),
    .X(net1518));
 sg13g2_buf_2 fanout1519 (.A(net1520),
    .X(net1519));
 sg13g2_buf_16 fanout1520 (.X(net1520),
    .A(net726));
 sg13g2_buf_16 fanout1521 (.X(net1521),
    .A(net1526));
 sg13g2_buf_1 fanout1522 (.A(net1525),
    .X(net1522));
 sg13g2_buf_1 fanout1523 (.A(net1524),
    .X(net1523));
 sg13g2_buf_1 fanout1524 (.A(net1525),
    .X(net1524));
 sg13g2_buf_1 fanout1525 (.A(net1526),
    .X(net1525));
 sg13g2_buf_8 fanout1526 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 ),
    .X(net1526));
 sg13g2_buf_1 fanout1527 (.A(_0376_),
    .X(net1527));
 sg13g2_buf_8 fanout1528 (.A(net1530),
    .X(net1528));
 sg13g2_buf_16 fanout1529 (.X(net1529),
    .A(net1530));
 sg13g2_buf_16 fanout1530 (.X(net1530),
    .A(net1533));
 sg13g2_buf_16 fanout1531 (.X(net1531),
    .A(net1532));
 sg13g2_buf_16 fanout1532 (.X(net1532),
    .A(net1533));
 sg13g2_buf_8 fanout1533 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 ),
    .X(net1533));
 sg13g2_buf_8 fanout1534 (.A(net1535),
    .X(net1534));
 sg13g2_buf_8 fanout1535 (.A(net637),
    .X(net1535));
 sg13g2_buf_8 fanout1536 (.A(net635),
    .X(net1536));
 sg13g2_buf_16 fanout1537 (.X(net1537),
    .A(net635));
 sg13g2_buf_16 rebuffer40 (.X(net649),
    .A(net648));
 sg13g2_buf_16 fanout1539 (.X(net1539),
    .A(net1540));
 sg13g2_buf_16 fanout1540 (.X(net1540),
    .A(net1541));
 sg13g2_buf_8 fanout1541 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 ),
    .X(net1541));
 sg13g2_buf_1 fanout1542 (.A(net1544),
    .X(net1542));
 sg13g2_buf_16 fanout1543 (.X(net1543),
    .A(net1544));
 sg13g2_buf_8 fanout1544 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net1544));
 sg13g2_buf_1 fanout1545 (.A(net1546),
    .X(net1545));
 sg13g2_buf_1 fanout1546 (.A(net1547),
    .X(net1546));
 sg13g2_buf_1 fanout1547 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 ),
    .X(net1547));
 sg13g2_buf_8 fanout1548 (.A(_1282_),
    .X(net1548));
 sg13g2_buf_16 fanout1549 (.X(net1549),
    .A(net1551));
 sg13g2_buf_8 fanout1550 (.A(net1551),
    .X(net1550));
 sg13g2_buf_16 fanout1551 (.X(net1551),
    .A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ));
 sg13g2_buf_1 fanout1552 (.A(net1553),
    .X(net1552));
 sg13g2_buf_1 fanout1553 (.A(net1554),
    .X(net1553));
 sg13g2_buf_1 fanout1554 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 ),
    .X(net1554));
 sg13g2_buf_8 fanout1555 (.A(_0171_),
    .X(net1555));
 sg13g2_buf_16 fanout1556 (.X(net1556),
    .A(net1557));
 sg13g2_buf_16 fanout1557 (.X(net1557),
    .A(net1558));
 sg13g2_buf_16 fanout1558 (.X(net1558),
    .A(net721));
 sg13g2_buf_8 fanout1559 (.A(net1560),
    .X(net1559));
 sg13g2_buf_1 fanout1560 (.A(net719),
    .X(net1560));
 sg13g2_buf_16 fanout1561 (.X(net1561),
    .A(_0172_));
 sg13g2_buf_1 fanout1562 (.A(_0172_),
    .X(net1562));
 sg13g2_buf_16 fanout1563 (.X(net1563),
    .A(net1564));
 sg13g2_buf_16 fanout1564 (.X(net1564),
    .A(net1567));
 sg13g2_buf_1 fanout1565 (.A(net1567),
    .X(net1565));
 sg13g2_buf_1 fanout1566 (.A(net1567),
    .X(net1566));
 sg13g2_buf_8 fanout1567 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 ),
    .X(net1567));
 sg13g2_buf_8 fanout1568 (.A(_1331_),
    .X(net1568));
 sg13g2_buf_1 fanout1569 (.A(net1571),
    .X(net1569));
 sg13g2_buf_1 fanout1570 (.A(net1571),
    .X(net1570));
 sg13g2_buf_1 fanout1571 (.A(_0173_),
    .X(net1571));
 sg13g2_buf_1 fanout1572 (.A(net1573),
    .X(net1572));
 sg13g2_buf_16 fanout1573 (.X(net1573),
    .A(net1574));
 sg13g2_buf_8 fanout1574 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 ),
    .X(net1574));
 sg13g2_buf_1 fanout1575 (.A(_0973_),
    .X(net1575));
 sg13g2_buf_8 fanout1576 (.A(_0681_),
    .X(net1576));
 sg13g2_buf_16 fanout1577 (.X(net1577),
    .A(net1578));
 sg13g2_buf_16 fanout1578 (.X(net1578),
    .A(net1580));
 sg13g2_buf_1 fanout1579 (.A(net1580),
    .X(net1579));
 sg13g2_buf_8 fanout1580 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .X(net1580));
 sg13g2_buf_1 fanout1581 (.A(net1582),
    .X(net1581));
 sg13g2_buf_1 fanout1582 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 ),
    .X(net1582));
 sg13g2_buf_16 fanout1583 (.X(net1583),
    .A(net1584));
 sg13g2_buf_16 fanout1584 (.X(net1584),
    .A(net1589));
 sg13g2_buf_1 fanout1585 (.A(net1587),
    .X(net1585));
 sg13g2_buf_1 fanout1586 (.A(net1587),
    .X(net1586));
 sg13g2_buf_1 fanout1587 (.A(net1589),
    .X(net1587));
 sg13g2_buf_1 fanout1588 (.A(net1589),
    .X(net1588));
 sg13g2_buf_8 fanout1589 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 ),
    .X(net1589));
 sg13g2_buf_1 fanout1590 (.A(_0174_),
    .X(net1590));
 sg13g2_buf_16 fanout1591 (.X(net1591),
    .A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ));
 sg13g2_buf_8 fanout1592 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net1592));
 sg13g2_buf_1 fanout1593 (.A(net1594),
    .X(net1593));
 sg13g2_buf_1 fanout1594 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net1594));
 sg13g2_buf_2 rebuffer8 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 ),
    .X(net617));
 sg13g2_buf_16 fanout1596 (.X(net1596),
    .A(net1601));
 sg13g2_buf_1 fanout1597 (.A(net1598),
    .X(net1597));
 sg13g2_buf_1 fanout1598 (.A(net1601),
    .X(net1598));
 sg13g2_buf_1 fanout1599 (.A(net1600),
    .X(net1599));
 sg13g2_buf_1 fanout1600 (.A(net1601),
    .X(net1600));
 sg13g2_buf_8 fanout1601 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 ),
    .X(net1601));
 sg13g2_buf_8 fanout1602 (.A(net1607),
    .X(net1602));
 sg13g2_buf_1 fanout1603 (.A(net648),
    .X(net1603));
 sg13g2_buf_8 rebuffer78 (.A(_0328_),
    .X(net687));
 sg13g2_buf_1 fanout1605 (.A(net1606),
    .X(net1605));
 sg13g2_buf_1 fanout1606 (.A(net1607),
    .X(net1606));
 sg13g2_buf_8 fanout1607 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 ),
    .X(net1607));
 sg13g2_buf_8 fanout1608 (.A(_0768_),
    .X(net1608));
 sg13g2_buf_16 fanout1609 (.X(net1609),
    .A(net1614));
 sg13g2_buf_1 fanout1610 (.A(net1611),
    .X(net1610));
 sg13g2_buf_1 fanout1611 (.A(net1614),
    .X(net1611));
 sg13g2_buf_1 fanout1612 (.A(net1613),
    .X(net1612));
 sg13g2_buf_1 fanout1613 (.A(net1614),
    .X(net1613));
 sg13g2_buf_8 fanout1614 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 ),
    .X(net1614));
 sg13g2_buf_16 fanout1615 (.X(net1615),
    .A(net1616));
 sg13g2_buf_8 fanout1616 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 ),
    .X(net1616));
 sg13g2_buf_16 fanout1617 (.X(net1617),
    .A(net1618));
 sg13g2_buf_16 fanout1618 (.X(net1618),
    .A(net1620));
 sg13g2_buf_1 fanout1619 (.A(net1620),
    .X(net1619));
 sg13g2_buf_8 fanout1620 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 ),
    .X(net1620));
 sg13g2_buf_16 fanout1621 (.X(net1621),
    .A(net1622));
 sg13g2_buf_16 fanout1622 (.X(net1622),
    .A(net1627));
 sg13g2_buf_1 fanout1623 (.A(net1627),
    .X(net1623));
 sg13g2_buf_1 fanout1624 (.A(net1627),
    .X(net1624));
 sg13g2_buf_1 fanout1625 (.A(net1626),
    .X(net1625));
 sg13g2_buf_1 fanout1626 (.A(net1627),
    .X(net1626));
 sg13g2_buf_8 fanout1627 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 ),
    .X(net1627));
 sg13g2_buf_8 fanout1628 (.A(_1148_),
    .X(net1628));
 sg13g2_buf_1 fanout1629 (.A(net1631),
    .X(net1629));
 sg13g2_buf_16 fanout1630 (.X(net1630),
    .A(net1631));
 sg13g2_buf_8 fanout1631 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .X(net1631));
 sg13g2_buf_1 fanout1632 (.A(net1635),
    .X(net1632));
 sg13g2_buf_1 fanout1633 (.A(net1635),
    .X(net1633));
 sg13g2_buf_1 fanout1634 (.A(net1635),
    .X(net1634));
 sg13g2_buf_1 fanout1635 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 ),
    .X(net1635));
 sg13g2_buf_1 fanout1636 (.A(_0135_),
    .X(net1636));
 sg13g2_buf_1 fanout1637 (.A(net1639),
    .X(net1637));
 sg13g2_buf_1 fanout1638 (.A(net1639),
    .X(net1638));
 sg13g2_buf_1 fanout1639 (.A(_0134_),
    .X(net1639));
 sg13g2_buf_1 fanout1640 (.A(_0123_),
    .X(net1640));
 sg13g2_buf_1 fanout1641 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .X(net1641));
 sg13g2_buf_1 fanout1642 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0.Q ),
    .X(net1642));
 sg13g2_buf_1 fanout1643 (.A(net1646),
    .X(net1643));
 sg13g2_buf_1 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_1 fanout1645 (.A(net1646),
    .X(net1645));
 sg13g2_buf_1 fanout1646 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2.Q ),
    .X(net1646));
 sg13g2_buf_1 fanout1647 (.A(net1648),
    .X(net1647));
 sg13g2_buf_1 fanout1648 (.A(net1651),
    .X(net1648));
 sg13g2_buf_1 fanout1649 (.A(net1650),
    .X(net1649));
 sg13g2_buf_1 fanout1650 (.A(net1651),
    .X(net1650));
 sg13g2_buf_1 fanout1651 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3.Q ),
    .X(net1651));
 sg13g2_buf_1 fanout1652 (.A(net1653),
    .X(net1652));
 sg13g2_buf_1 fanout1653 (.A(net1654),
    .X(net1653));
 sg13g2_buf_1 fanout1654 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .X(net1654));
 sg13g2_buf_1 fanout1655 (.A(net1656),
    .X(net1655));
 sg13g2_buf_1 fanout1656 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5.Q ),
    .X(net1656));
 sg13g2_buf_1 fanout1657 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4.Q ),
    .X(net1657));
 sg13g2_buf_1 fanout1658 (.A(net1659),
    .X(net1658));
 sg13g2_buf_1 fanout1659 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12.Q ),
    .X(net1659));
 sg13g2_buf_1 fanout1660 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16.Q ),
    .X(net1660));
 sg13g2_buf_1 fanout1661 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24.Q ),
    .X(net1661));
 sg13g2_buf_1 fanout1662 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28.Q ),
    .X(net1662));
 sg13g2_buf_1 fanout1663 (.A(net1664),
    .X(net1663));
 sg13g2_buf_1 fanout1664 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0.Q ),
    .X(net1664));
 sg13g2_buf_1 fanout1665 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4.Q ),
    .X(net1665));
 sg13g2_buf_1 fanout1666 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8.Q ),
    .X(net1666));
 sg13g2_buf_1 fanout1667 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4.Q ),
    .X(net1667));
 sg13g2_buf_1 fanout1668 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16.Q ),
    .X(net1668));
 sg13g2_buf_1 fanout1669 (.A(net1670),
    .X(net1669));
 sg13g2_buf_1 fanout1670 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20.Q ),
    .X(net1670));
 sg13g2_buf_1 fanout1671 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28.Q ),
    .X(net1671));
 sg13g2_buf_1 fanout1672 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .X(net1672));
 sg13g2_buf_1 fanout1673 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0.Q ),
    .X(net1673));
 sg13g2_buf_1 fanout1674 (.A(net1675),
    .X(net1674));
 sg13g2_buf_1 fanout1675 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4.Q ),
    .X(net1675));
 sg13g2_buf_1 fanout1676 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8.Q ),
    .X(net1676));
 sg13g2_buf_1 fanout1677 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16.Q ),
    .X(net1677));
 sg13g2_buf_1 fanout1678 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24.Q ),
    .X(net1678));
 sg13g2_buf_1 fanout1679 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28.Q ),
    .X(net1679));
 sg13g2_buf_1 fanout1680 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(net1680));
 sg13g2_buf_1 fanout1681 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0.Q ),
    .X(net1681));
 sg13g2_buf_1 fanout1682 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4.Q ),
    .X(net1682));
 sg13g2_buf_1 fanout1683 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8.Q ),
    .X(net1683));
 sg13g2_buf_1 fanout1684 (.A(net1685),
    .X(net1684));
 sg13g2_buf_1 fanout1685 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12.Q ),
    .X(net1685));
 sg13g2_buf_1 fanout1686 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16.Q ),
    .X(net1686));
 sg13g2_buf_1 fanout1687 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20.Q ),
    .X(net1687));
 sg13g2_buf_1 fanout1688 (.A(net1689),
    .X(net1688));
 sg13g2_buf_1 fanout1689 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8.Q ),
    .X(net1689));
 sg13g2_buf_1 fanout1690 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16.Q ),
    .X(net1690));
 sg13g2_buf_1 fanout1691 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24.Q ),
    .X(net1691));
 sg13g2_buf_1 fanout1692 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28.Q ),
    .X(net1692));
 sg13g2_buf_1 fanout1693 (.A(net1694),
    .X(net1693));
 sg13g2_buf_1 fanout1694 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0.Q ),
    .X(net1694));
 sg13g2_buf_1 fanout1695 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(net1695));
 sg13g2_buf_1 fanout1696 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4.Q ),
    .X(net1696));
 sg13g2_buf_1 fanout1697 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(net1697));
 sg13g2_buf_1 fanout1698 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8.Q ),
    .X(net1698));
 sg13g2_buf_1 fanout1699 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20.Q ),
    .X(net1699));
 sg13g2_buf_1 fanout1700 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24.Q ),
    .X(net1700));
 sg13g2_buf_1 fanout1701 (.A(net1702),
    .X(net1701));
 sg13g2_buf_1 fanout1702 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28.Q ),
    .X(net1702));
 sg13g2_buf_1 fanout1703 (.A(net168),
    .X(net1703));
 sg13g2_buf_1 fanout1704 (.A(net150),
    .X(net1704));
 sg13g2_buf_1 fanout1705 (.A(net149),
    .X(net1705));
 sg13g2_buf_1 fanout1706 (.A(net130),
    .X(net1706));
 sg13g2_buf_1 fanout1707 (.A(net129),
    .X(net1707));
 sg13g2_buf_1 fanout1708 (.A(net127),
    .X(net1708));
 sg13g2_buf_1 fanout1709 (.A(net123),
    .X(net1709));
 sg13g2_buf_1 fanout1710 (.A(net114),
    .X(net1710));
 sg13g2_buf_1 fanout1711 (.A(net113),
    .X(net1711));
 sg13g2_buf_1 fanout1712 (.A(net112),
    .X(net1712));
 sg13g2_buf_1 fanout1713 (.A(net111),
    .X(net1713));
 sg13g2_buf_1 fanout1714 (.A(net1715),
    .X(net1714));
 sg13g2_buf_1 fanout1715 (.A(net1718),
    .X(net1715));
 sg13g2_buf_1 fanout1716 (.A(net1718),
    .X(net1716));
 sg13g2_buf_1 fanout1717 (.A(net1718),
    .X(net1717));
 sg13g2_buf_1 fanout1718 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1718));
 sg13g2_buf_1 fanout1719 (.A(net1720),
    .X(net1719));
 sg13g2_buf_1 fanout1720 (.A(net1721),
    .X(net1720));
 sg13g2_buf_1 fanout1721 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1721));
 sg13g2_buf_1 fanout1722 (.A(net1723),
    .X(net1722));
 sg13g2_buf_1 fanout1723 (.A(Tile_X0Y1_FrameStrobe[9]),
    .X(net1723));
 sg13g2_buf_1 fanout1724 (.A(net1726),
    .X(net1724));
 sg13g2_buf_1 fanout1725 (.A(net1726),
    .X(net1725));
 sg13g2_buf_1 fanout1726 (.A(net1734),
    .X(net1726));
 sg13g2_buf_1 fanout1727 (.A(net1728),
    .X(net1727));
 sg13g2_buf_1 fanout1728 (.A(net1734),
    .X(net1728));
 sg13g2_buf_1 fanout1729 (.A(net1734),
    .X(net1729));
 sg13g2_buf_1 fanout1730 (.A(net1734),
    .X(net1730));
 sg13g2_buf_1 fanout1731 (.A(net1733),
    .X(net1731));
 sg13g2_buf_1 fanout1732 (.A(net1733),
    .X(net1732));
 sg13g2_buf_1 fanout1733 (.A(net1734),
    .X(net1733));
 sg13g2_buf_1 fanout1734 (.A(Tile_X0Y1_FrameStrobe[8]),
    .X(net1734));
 sg13g2_buf_1 fanout1735 (.A(net1738),
    .X(net1735));
 sg13g2_buf_1 fanout1736 (.A(net1738),
    .X(net1736));
 sg13g2_buf_1 fanout1737 (.A(net1738),
    .X(net1737));
 sg13g2_buf_1 fanout1738 (.A(net1741),
    .X(net1738));
 sg13g2_buf_1 fanout1739 (.A(net1741),
    .X(net1739));
 sg13g2_buf_1 fanout1740 (.A(net1741),
    .X(net1740));
 sg13g2_buf_1 fanout1741 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1741));
 sg13g2_buf_1 fanout1742 (.A(net1744),
    .X(net1742));
 sg13g2_buf_1 fanout1743 (.A(net1744),
    .X(net1743));
 sg13g2_buf_1 fanout1744 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1744));
 sg13g2_buf_1 fanout1745 (.A(Tile_X0Y1_FrameStrobe[7]),
    .X(net1745));
 sg13g2_buf_1 fanout1746 (.A(net1747),
    .X(net1746));
 sg13g2_buf_1 fanout1747 (.A(net1757),
    .X(net1747));
 sg13g2_buf_1 fanout1748 (.A(net1750),
    .X(net1748));
 sg13g2_buf_1 fanout1749 (.A(net1757),
    .X(net1749));
 sg13g2_buf_1 fanout1750 (.A(net1757),
    .X(net1750));
 sg13g2_buf_1 fanout1751 (.A(net1752),
    .X(net1751));
 sg13g2_buf_1 fanout1752 (.A(net1753),
    .X(net1752));
 sg13g2_buf_1 fanout1753 (.A(net1757),
    .X(net1753));
 sg13g2_buf_1 fanout1754 (.A(net1755),
    .X(net1754));
 sg13g2_buf_1 fanout1755 (.A(net1756),
    .X(net1755));
 sg13g2_buf_1 fanout1756 (.A(net1757),
    .X(net1756));
 sg13g2_buf_1 fanout1757 (.A(Tile_X0Y1_FrameStrobe[6]),
    .X(net1757));
 sg13g2_buf_1 fanout1758 (.A(net1762),
    .X(net1758));
 sg13g2_buf_1 fanout1759 (.A(net1762),
    .X(net1759));
 sg13g2_buf_1 fanout1760 (.A(net1761),
    .X(net1760));
 sg13g2_buf_1 fanout1761 (.A(net1762),
    .X(net1761));
 sg13g2_buf_1 fanout1762 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1762));
 sg13g2_buf_1 fanout1763 (.A(net1768),
    .X(net1763));
 sg13g2_buf_1 fanout1764 (.A(net1765),
    .X(net1764));
 sg13g2_buf_1 fanout1765 (.A(net1768),
    .X(net1765));
 sg13g2_buf_1 fanout1766 (.A(net1767),
    .X(net1766));
 sg13g2_buf_1 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_1 fanout1768 (.A(Tile_X0Y1_FrameStrobe[5]),
    .X(net1768));
 sg13g2_buf_1 fanout1769 (.A(net1771),
    .X(net1769));
 sg13g2_buf_1 fanout1770 (.A(net1771),
    .X(net1770));
 sg13g2_buf_1 fanout1771 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1771));
 sg13g2_buf_1 fanout1772 (.A(net1774),
    .X(net1772));
 sg13g2_buf_1 fanout1773 (.A(net1774),
    .X(net1773));
 sg13g2_buf_1 fanout1774 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1774));
 sg13g2_buf_1 fanout1775 (.A(net1776),
    .X(net1775));
 sg13g2_buf_1 fanout1776 (.A(net1779),
    .X(net1776));
 sg13g2_buf_1 fanout1777 (.A(net1779),
    .X(net1777));
 sg13g2_buf_1 fanout1778 (.A(net1779),
    .X(net1778));
 sg13g2_buf_1 fanout1779 (.A(Tile_X0Y1_FrameStrobe[4]),
    .X(net1779));
 sg13g2_buf_1 fanout1780 (.A(net1784),
    .X(net1780));
 sg13g2_buf_1 fanout1781 (.A(net1784),
    .X(net1781));
 sg13g2_buf_1 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_1 fanout1783 (.A(net1784),
    .X(net1783));
 sg13g2_buf_1 fanout1784 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net1784));
 sg13g2_buf_1 fanout1785 (.A(net1786),
    .X(net1785));
 sg13g2_buf_1 fanout1786 (.A(net1788),
    .X(net1786));
 sg13g2_buf_1 fanout1787 (.A(net1788),
    .X(net1787));
 sg13g2_buf_1 fanout1788 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net1788));
 sg13g2_buf_1 fanout1789 (.A(Tile_X0Y1_FrameStrobe[3]),
    .X(net1789));
 sg13g2_buf_1 fanout1790 (.A(net1791),
    .X(net1790));
 sg13g2_buf_1 fanout1791 (.A(net1792),
    .X(net1791));
 sg13g2_buf_1 fanout1792 (.A(net1800),
    .X(net1792));
 sg13g2_buf_1 fanout1793 (.A(net1800),
    .X(net1793));
 sg13g2_buf_1 fanout1794 (.A(net1800),
    .X(net1794));
 sg13g2_buf_1 fanout1795 (.A(net1796),
    .X(net1795));
 sg13g2_buf_1 fanout1796 (.A(net1797),
    .X(net1796));
 sg13g2_buf_1 fanout1797 (.A(net1800),
    .X(net1797));
 sg13g2_buf_1 fanout1798 (.A(net1799),
    .X(net1798));
 sg13g2_buf_1 fanout1799 (.A(net1800),
    .X(net1799));
 sg13g2_buf_1 fanout1800 (.A(Tile_X0Y1_FrameStrobe[2]),
    .X(net1800));
 sg13g2_buf_1 fanout1801 (.A(net1803),
    .X(net1801));
 sg13g2_buf_1 fanout1802 (.A(net1803),
    .X(net1802));
 sg13g2_buf_1 fanout1803 (.A(net1811),
    .X(net1803));
 sg13g2_buf_1 fanout1804 (.A(net1805),
    .X(net1804));
 sg13g2_buf_1 fanout1805 (.A(net1811),
    .X(net1805));
 sg13g2_buf_1 fanout1806 (.A(net1808),
    .X(net1806));
 sg13g2_buf_1 fanout1807 (.A(net1808),
    .X(net1807));
 sg13g2_buf_1 fanout1808 (.A(net1811),
    .X(net1808));
 sg13g2_buf_1 fanout1809 (.A(net1811),
    .X(net1809));
 sg13g2_buf_1 fanout1810 (.A(net1811),
    .X(net1810));
 sg13g2_buf_1 fanout1811 (.A(Tile_X0Y1_FrameStrobe[1]),
    .X(net1811));
 sg13g2_buf_1 fanout1812 (.A(net1813),
    .X(net1812));
 sg13g2_buf_1 fanout1813 (.A(net1815),
    .X(net1813));
 sg13g2_buf_1 fanout1814 (.A(net1815),
    .X(net1814));
 sg13g2_buf_1 fanout1815 (.A(net1816),
    .X(net1815));
 sg13g2_buf_1 fanout1816 (.A(net1820),
    .X(net1816));
 sg13g2_buf_1 fanout1817 (.A(net1818),
    .X(net1817));
 sg13g2_buf_1 fanout1818 (.A(net1819),
    .X(net1818));
 sg13g2_buf_1 fanout1819 (.A(net1820),
    .X(net1819));
 sg13g2_buf_1 fanout1820 (.A(Tile_X0Y1_FrameStrobe[12]),
    .X(net1820));
 sg13g2_buf_1 fanout1821 (.A(net1823),
    .X(net1821));
 sg13g2_buf_1 fanout1822 (.A(net1823),
    .X(net1822));
 sg13g2_buf_1 fanout1823 (.A(net1825),
    .X(net1823));
 sg13g2_buf_1 fanout1824 (.A(net1825),
    .X(net1824));
 sg13g2_buf_1 fanout1825 (.A(net1826),
    .X(net1825));
 sg13g2_buf_1 fanout1826 (.A(net1832),
    .X(net1826));
 sg13g2_buf_1 fanout1827 (.A(net1830),
    .X(net1827));
 sg13g2_buf_1 fanout1828 (.A(net1829),
    .X(net1828));
 sg13g2_buf_1 fanout1829 (.A(net1830),
    .X(net1829));
 sg13g2_buf_1 fanout1830 (.A(net1831),
    .X(net1830));
 sg13g2_buf_1 fanout1831 (.A(net1832),
    .X(net1831));
 sg13g2_buf_1 fanout1832 (.A(Tile_X0Y1_FrameStrobe[11]),
    .X(net1832));
 sg13g2_buf_1 fanout1833 (.A(net1835),
    .X(net1833));
 sg13g2_buf_1 fanout1834 (.A(net1835),
    .X(net1834));
 sg13g2_buf_1 fanout1835 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1835));
 sg13g2_buf_1 fanout1836 (.A(net1838),
    .X(net1836));
 sg13g2_buf_1 fanout1837 (.A(net1838),
    .X(net1837));
 sg13g2_buf_1 fanout1838 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1838));
 sg13g2_buf_1 fanout1839 (.A(net1840),
    .X(net1839));
 sg13g2_buf_1 fanout1840 (.A(net1841),
    .X(net1840));
 sg13g2_buf_1 fanout1841 (.A(net1844),
    .X(net1841));
 sg13g2_buf_1 fanout1842 (.A(net1843),
    .X(net1842));
 sg13g2_buf_1 fanout1843 (.A(net1844),
    .X(net1843));
 sg13g2_buf_1 fanout1844 (.A(Tile_X0Y1_FrameStrobe[10]),
    .X(net1844));
 sg13g2_buf_1 fanout1845 (.A(net1846),
    .X(net1845));
 sg13g2_buf_1 fanout1846 (.A(net1847),
    .X(net1846));
 sg13g2_buf_1 fanout1847 (.A(net1848),
    .X(net1847));
 sg13g2_buf_1 fanout1848 (.A(net1850),
    .X(net1848));
 sg13g2_buf_1 fanout1849 (.A(net1850),
    .X(net1849));
 sg13g2_buf_1 fanout1850 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net1850));
 sg13g2_buf_1 fanout1851 (.A(net1853),
    .X(net1851));
 sg13g2_buf_1 fanout1852 (.A(net1853),
    .X(net1852));
 sg13g2_buf_1 fanout1853 (.A(net1855),
    .X(net1853));
 sg13g2_buf_1 fanout1854 (.A(net1855),
    .X(net1854));
 sg13g2_buf_1 fanout1855 (.A(Tile_X0Y1_FrameStrobe[0]),
    .X(net1855));
 sg13g2_buf_1 fanout1856 (.A(Tile_X0Y1_FrameData[9]),
    .X(net1856));
 sg13g2_buf_1 fanout1857 (.A(Tile_X0Y1_FrameData[9]),
    .X(net1857));
 sg13g2_buf_1 fanout1858 (.A(net1859),
    .X(net1858));
 sg13g2_buf_1 fanout1859 (.A(Tile_X0Y1_FrameData[8]),
    .X(net1859));
 sg13g2_buf_1 fanout1860 (.A(Tile_X0Y1_FrameData[7]),
    .X(net1860));
 sg13g2_buf_1 fanout1861 (.A(Tile_X0Y1_FrameData[7]),
    .X(net1861));
 sg13g2_buf_1 fanout1862 (.A(Tile_X0Y1_FrameData[6]),
    .X(net1862));
 sg13g2_buf_1 fanout1863 (.A(Tile_X0Y1_FrameData[6]),
    .X(net1863));
 sg13g2_buf_1 fanout1864 (.A(Tile_X0Y1_FrameData[5]),
    .X(net1864));
 sg13g2_buf_1 fanout1865 (.A(Tile_X0Y1_FrameData[5]),
    .X(net1865));
 sg13g2_buf_1 fanout1866 (.A(net1867),
    .X(net1866));
 sg13g2_buf_1 fanout1867 (.A(Tile_X0Y1_FrameData[4]),
    .X(net1867));
 sg13g2_buf_1 fanout1868 (.A(Tile_X0Y1_FrameData[3]),
    .X(net1868));
 sg13g2_buf_1 fanout1869 (.A(Tile_X0Y1_FrameData[3]),
    .X(net1869));
 sg13g2_buf_1 fanout1870 (.A(Tile_X0Y1_FrameData[31]),
    .X(net1870));
 sg13g2_buf_1 fanout1871 (.A(Tile_X0Y1_FrameData[31]),
    .X(net1871));
 sg13g2_buf_1 fanout1872 (.A(Tile_X0Y1_FrameData[30]),
    .X(net1872));
 sg13g2_buf_1 fanout1873 (.A(Tile_X0Y1_FrameData[30]),
    .X(net1873));
 sg13g2_buf_1 fanout1874 (.A(Tile_X0Y1_FrameData[2]),
    .X(net1874));
 sg13g2_buf_1 fanout1875 (.A(Tile_X0Y1_FrameData[2]),
    .X(net1875));
 sg13g2_buf_1 fanout1876 (.A(Tile_X0Y1_FrameData[29]),
    .X(net1876));
 sg13g2_buf_1 fanout1877 (.A(Tile_X0Y1_FrameData[29]),
    .X(net1877));
 sg13g2_buf_1 fanout1878 (.A(Tile_X0Y1_FrameData[28]),
    .X(net1878));
 sg13g2_buf_1 fanout1879 (.A(Tile_X0Y1_FrameData[28]),
    .X(net1879));
 sg13g2_buf_1 fanout1880 (.A(net1881),
    .X(net1880));
 sg13g2_buf_1 fanout1881 (.A(Tile_X0Y1_FrameData[27]),
    .X(net1881));
 sg13g2_buf_1 fanout1882 (.A(Tile_X0Y1_FrameData[26]),
    .X(net1882));
 sg13g2_buf_1 fanout1883 (.A(Tile_X0Y1_FrameData[26]),
    .X(net1883));
 sg13g2_buf_1 fanout1884 (.A(Tile_X0Y1_FrameData[25]),
    .X(net1884));
 sg13g2_buf_1 fanout1885 (.A(Tile_X0Y1_FrameData[25]),
    .X(net1885));
 sg13g2_buf_1 fanout1886 (.A(Tile_X0Y1_FrameData[24]),
    .X(net1886));
 sg13g2_buf_1 fanout1887 (.A(Tile_X0Y1_FrameData[24]),
    .X(net1887));
 sg13g2_buf_1 fanout1888 (.A(net1889),
    .X(net1888));
 sg13g2_buf_1 fanout1889 (.A(Tile_X0Y1_FrameData[23]),
    .X(net1889));
 sg13g2_buf_1 fanout1890 (.A(net1891),
    .X(net1890));
 sg13g2_buf_1 fanout1891 (.A(Tile_X0Y1_FrameData[22]),
    .X(net1891));
 sg13g2_buf_1 fanout1892 (.A(net1893),
    .X(net1892));
 sg13g2_buf_1 fanout1893 (.A(Tile_X0Y1_FrameData[21]),
    .X(net1893));
 sg13g2_buf_1 fanout1894 (.A(net1895),
    .X(net1894));
 sg13g2_buf_1 fanout1895 (.A(Tile_X0Y1_FrameData[20]),
    .X(net1895));
 sg13g2_buf_1 fanout1896 (.A(Tile_X0Y1_FrameData[1]),
    .X(net1896));
 sg13g2_buf_1 fanout1897 (.A(Tile_X0Y1_FrameData[1]),
    .X(net1897));
 sg13g2_buf_1 fanout1898 (.A(Tile_X0Y1_FrameData[19]),
    .X(net1898));
 sg13g2_buf_1 fanout1899 (.A(Tile_X0Y1_FrameData[19]),
    .X(net1899));
 sg13g2_buf_1 fanout1900 (.A(Tile_X0Y1_FrameData[18]),
    .X(net1900));
 sg13g2_buf_1 fanout1901 (.A(Tile_X0Y1_FrameData[18]),
    .X(net1901));
 sg13g2_buf_1 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_1 fanout1903 (.A(Tile_X0Y1_FrameData[17]),
    .X(net1903));
 sg13g2_buf_1 fanout1904 (.A(Tile_X0Y1_FrameData[16]),
    .X(net1904));
 sg13g2_buf_1 fanout1905 (.A(Tile_X0Y1_FrameData[16]),
    .X(net1905));
 sg13g2_buf_1 fanout1906 (.A(net1907),
    .X(net1906));
 sg13g2_buf_1 fanout1907 (.A(Tile_X0Y1_FrameData[15]),
    .X(net1907));
 sg13g2_buf_1 fanout1908 (.A(net1909),
    .X(net1908));
 sg13g2_buf_1 fanout1909 (.A(Tile_X0Y1_FrameData[14]),
    .X(net1909));
 sg13g2_buf_1 fanout1910 (.A(net1911),
    .X(net1910));
 sg13g2_buf_1 fanout1911 (.A(Tile_X0Y1_FrameData[13]),
    .X(net1911));
 sg13g2_buf_1 fanout1912 (.A(net1913),
    .X(net1912));
 sg13g2_buf_1 fanout1913 (.A(net1914),
    .X(net1913));
 sg13g2_buf_1 fanout1914 (.A(Tile_X0Y1_FrameData[12]),
    .X(net1914));
 sg13g2_buf_1 fanout1915 (.A(net1916),
    .X(net1915));
 sg13g2_buf_1 fanout1916 (.A(Tile_X0Y1_FrameData[11]),
    .X(net1916));
 sg13g2_buf_1 fanout1917 (.A(net1918),
    .X(net1917));
 sg13g2_buf_1 fanout1918 (.A(Tile_X0Y1_FrameData[10]),
    .X(net1918));
 sg13g2_buf_1 fanout1919 (.A(Tile_X0Y1_FrameData[0]),
    .X(net1919));
 sg13g2_buf_1 fanout1920 (.A(Tile_X0Y1_FrameData[0]),
    .X(net1920));
 sg13g2_buf_1 fanout1921 (.A(Tile_X0Y1_E6END[1]),
    .X(net1921));
 sg13g2_buf_1 fanout1922 (.A(Tile_X0Y1_E6END[1]),
    .X(net1922));
 sg13g2_buf_1 fanout1923 (.A(net1924),
    .X(net1923));
 sg13g2_buf_1 fanout1924 (.A(Tile_X0Y1_E6END[0]),
    .X(net1924));
 sg13g2_buf_1 fanout1925 (.A(net90),
    .X(net1925));
 sg13g2_buf_1 fanout1926 (.A(net89),
    .X(net1926));
 sg13g2_buf_1 fanout1927 (.A(net88),
    .X(net1927));
 sg13g2_buf_1 fanout1928 (.A(net87),
    .X(net1928));
 sg13g2_buf_1 fanout1929 (.A(net81),
    .X(net1929));
 sg13g2_buf_1 fanout1930 (.A(net1931),
    .X(net1930));
 sg13g2_buf_1 fanout1931 (.A(Tile_X0Y0_W1END[3]),
    .X(net1931));
 sg13g2_buf_1 fanout1932 (.A(net64),
    .X(net1932));
 sg13g2_buf_1 fanout1933 (.A(net63),
    .X(net1933));
 sg13g2_buf_1 fanout1934 (.A(net45),
    .X(net1934));
 sg13g2_buf_1 fanout1935 (.A(net40),
    .X(net1935));
 sg13g2_buf_1 fanout1936 (.A(net39),
    .X(net1936));
 sg13g2_buf_1 fanout1937 (.A(net1938),
    .X(net1937));
 sg13g2_buf_1 fanout1938 (.A(Tile_X0Y0_FrameData[9]),
    .X(net1938));
 sg13g2_buf_1 fanout1939 (.A(net1940),
    .X(net1939));
 sg13g2_buf_1 fanout1940 (.A(Tile_X0Y0_FrameData[8]),
    .X(net1940));
 sg13g2_buf_1 fanout1941 (.A(net1942),
    .X(net1941));
 sg13g2_buf_1 fanout1942 (.A(Tile_X0Y0_FrameData[7]),
    .X(net1942));
 sg13g2_buf_1 fanout1943 (.A(net1944),
    .X(net1943));
 sg13g2_buf_1 fanout1944 (.A(Tile_X0Y0_FrameData[6]),
    .X(net1944));
 sg13g2_buf_1 fanout1945 (.A(Tile_X0Y0_FrameData[5]),
    .X(net1945));
 sg13g2_buf_1 fanout1946 (.A(Tile_X0Y0_FrameData[5]),
    .X(net1946));
 sg13g2_buf_1 fanout1947 (.A(Tile_X0Y0_FrameData[4]),
    .X(net1947));
 sg13g2_buf_1 fanout1948 (.A(Tile_X0Y0_FrameData[4]),
    .X(net1948));
 sg13g2_buf_1 fanout1949 (.A(net1950),
    .X(net1949));
 sg13g2_buf_1 fanout1950 (.A(Tile_X0Y0_FrameData[3]),
    .X(net1950));
 sg13g2_buf_1 fanout1951 (.A(Tile_X0Y0_FrameData[31]),
    .X(net1951));
 sg13g2_buf_1 fanout1952 (.A(Tile_X0Y0_FrameData[31]),
    .X(net1952));
 sg13g2_buf_1 fanout1953 (.A(Tile_X0Y0_FrameData[30]),
    .X(net1953));
 sg13g2_buf_1 fanout1954 (.A(Tile_X0Y0_FrameData[30]),
    .X(net1954));
 sg13g2_buf_1 fanout1955 (.A(net1956),
    .X(net1955));
 sg13g2_buf_1 fanout1956 (.A(Tile_X0Y0_FrameData[2]),
    .X(net1956));
 sg13g2_buf_1 fanout1957 (.A(Tile_X0Y0_FrameData[29]),
    .X(net1957));
 sg13g2_buf_1 fanout1958 (.A(Tile_X0Y0_FrameData[29]),
    .X(net1958));
 sg13g2_buf_1 fanout1959 (.A(Tile_X0Y0_FrameData[28]),
    .X(net1959));
 sg13g2_buf_1 fanout1960 (.A(Tile_X0Y0_FrameData[28]),
    .X(net1960));
 sg13g2_buf_1 fanout1961 (.A(net1962),
    .X(net1961));
 sg13g2_buf_1 fanout1962 (.A(Tile_X0Y0_FrameData[27]),
    .X(net1962));
 sg13g2_buf_1 fanout1963 (.A(Tile_X0Y0_FrameData[26]),
    .X(net1963));
 sg13g2_buf_1 fanout1964 (.A(Tile_X0Y0_FrameData[26]),
    .X(net1964));
 sg13g2_buf_1 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_1 fanout1966 (.A(Tile_X0Y0_FrameData[25]),
    .X(net1966));
 sg13g2_buf_1 fanout1967 (.A(net1968),
    .X(net1967));
 sg13g2_buf_1 fanout1968 (.A(Tile_X0Y0_FrameData[24]),
    .X(net1968));
 sg13g2_buf_1 fanout1969 (.A(Tile_X0Y0_FrameData[23]),
    .X(net1969));
 sg13g2_buf_1 fanout1970 (.A(Tile_X0Y0_FrameData[23]),
    .X(net1970));
 sg13g2_buf_1 fanout1971 (.A(Tile_X0Y0_FrameData[22]),
    .X(net1971));
 sg13g2_buf_1 fanout1972 (.A(Tile_X0Y0_FrameData[22]),
    .X(net1972));
 sg13g2_buf_1 fanout1973 (.A(net1974),
    .X(net1973));
 sg13g2_buf_1 fanout1974 (.A(Tile_X0Y0_FrameData[21]),
    .X(net1974));
 sg13g2_buf_1 fanout1975 (.A(net1976),
    .X(net1975));
 sg13g2_buf_1 fanout1976 (.A(Tile_X0Y0_FrameData[20]),
    .X(net1976));
 sg13g2_buf_1 fanout1977 (.A(net1978),
    .X(net1977));
 sg13g2_buf_1 fanout1978 (.A(Tile_X0Y0_FrameData[1]),
    .X(net1978));
 sg13g2_buf_1 fanout1979 (.A(net1980),
    .X(net1979));
 sg13g2_buf_1 fanout1980 (.A(Tile_X0Y0_FrameData[19]),
    .X(net1980));
 sg13g2_buf_1 fanout1981 (.A(net1982),
    .X(net1981));
 sg13g2_buf_1 fanout1982 (.A(Tile_X0Y0_FrameData[18]),
    .X(net1982));
 sg13g2_buf_1 fanout1983 (.A(net1984),
    .X(net1983));
 sg13g2_buf_1 fanout1984 (.A(Tile_X0Y0_FrameData[17]),
    .X(net1984));
 sg13g2_buf_1 fanout1985 (.A(net1986),
    .X(net1985));
 sg13g2_buf_1 fanout1986 (.A(Tile_X0Y0_FrameData[16]),
    .X(net1986));
 sg13g2_buf_1 fanout1987 (.A(net1988),
    .X(net1987));
 sg13g2_buf_1 fanout1988 (.A(Tile_X0Y0_FrameData[15]),
    .X(net1988));
 sg13g2_buf_1 fanout1989 (.A(net1990),
    .X(net1989));
 sg13g2_buf_1 fanout1990 (.A(Tile_X0Y0_FrameData[14]),
    .X(net1990));
 sg13g2_buf_1 fanout1991 (.A(net1992),
    .X(net1991));
 sg13g2_buf_1 fanout1992 (.A(Tile_X0Y0_FrameData[13]),
    .X(net1992));
 sg13g2_buf_1 fanout1993 (.A(net1994),
    .X(net1993));
 sg13g2_buf_1 fanout1994 (.A(Tile_X0Y0_FrameData[12]),
    .X(net1994));
 sg13g2_buf_1 fanout1995 (.A(net1996),
    .X(net1995));
 sg13g2_buf_1 fanout1996 (.A(Tile_X0Y0_FrameData[11]),
    .X(net1996));
 sg13g2_buf_1 fanout1997 (.A(Tile_X0Y0_FrameData[10]),
    .X(net1997));
 sg13g2_buf_1 fanout1998 (.A(Tile_X0Y0_FrameData[10]),
    .X(net1998));
 sg13g2_buf_1 fanout1999 (.A(Tile_X0Y0_FrameData[0]),
    .X(net1999));
 sg13g2_buf_1 fanout2000 (.A(Tile_X0Y0_FrameData[0]),
    .X(net2000));
 sg13g2_buf_1 fanout2001 (.A(net2002),
    .X(net2001));
 sg13g2_buf_1 fanout2002 (.A(Tile_X0Y0_E1END[3]),
    .X(net2002));
 sg13g2_buf_1 fanout2003 (.A(net3),
    .X(net2003));
 sg13g2_buf_1 fanout2004 (.A(net2),
    .X(net2004));
 sg13g2_buf_1 fanout2005 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24.Q ),
    .X(net2005));
 sg13g2_buf_2 input1 (.A(Tile_X0Y0_E1END[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(Tile_X0Y0_E1END[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(Tile_X0Y0_E1END[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(Tile_X0Y0_E2END[0]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(Tile_X0Y0_E2END[1]),
    .X(net5));
 sg13g2_buf_8 input6 (.A(Tile_X0Y0_E2END[2]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(Tile_X0Y0_E2END[3]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(Tile_X0Y0_E2END[4]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(Tile_X0Y0_E2END[5]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(Tile_X0Y0_E2END[6]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(Tile_X0Y0_E2END[7]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(Tile_X0Y0_E2MID[0]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(Tile_X0Y0_E2MID[1]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(Tile_X0Y0_E2MID[2]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(Tile_X0Y0_E2MID[3]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(Tile_X0Y0_E2MID[4]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(Tile_X0Y0_E2MID[5]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(Tile_X0Y0_E2MID[6]),
    .X(net18));
 sg13g2_buf_1 input19 (.A(Tile_X0Y0_E2MID[7]),
    .X(net19));
 sg13g2_buf_2 input20 (.A(Tile_X0Y0_E6END[0]),
    .X(net20));
 sg13g2_buf_1 input21 (.A(Tile_X0Y0_E6END[1]),
    .X(net21));
 sg13g2_buf_1 input22 (.A(Tile_X0Y0_EE4END[0]),
    .X(net22));
 sg13g2_buf_1 input23 (.A(Tile_X0Y0_EE4END[1]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(Tile_X0Y0_EE4END[2]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(Tile_X0Y0_EE4END[3]),
    .X(net25));
 sg13g2_buf_1 input26 (.A(Tile_X0Y0_S1END[0]),
    .X(net26));
 sg13g2_buf_1 input27 (.A(Tile_X0Y0_S1END[1]),
    .X(net27));
 sg13g2_buf_1 input28 (.A(Tile_X0Y0_S1END[2]),
    .X(net28));
 sg13g2_buf_1 input29 (.A(Tile_X0Y0_S1END[3]),
    .X(net29));
 sg13g2_buf_1 input30 (.A(Tile_X0Y0_S2END[0]),
    .X(net30));
 sg13g2_buf_1 input31 (.A(Tile_X0Y0_S2END[1]),
    .X(net31));
 sg13g2_buf_16 input32 (.X(net32),
    .A(Tile_X0Y0_S2END[2]));
 sg13g2_buf_1 input33 (.A(Tile_X0Y0_S2END[3]),
    .X(net33));
 sg13g2_buf_1 input34 (.A(Tile_X0Y0_S2END[4]),
    .X(net34));
 sg13g2_buf_1 input35 (.A(Tile_X0Y0_S2END[5]),
    .X(net35));
 sg13g2_buf_1 input36 (.A(Tile_X0Y0_S2END[6]),
    .X(net36));
 sg13g2_buf_1 input37 (.A(Tile_X0Y0_S2END[7]),
    .X(net37));
 sg13g2_buf_1 input38 (.A(Tile_X0Y0_S2MID[0]),
    .X(net38));
 sg13g2_buf_1 input39 (.A(Tile_X0Y0_S2MID[1]),
    .X(net39));
 sg13g2_buf_1 input40 (.A(Tile_X0Y0_S2MID[2]),
    .X(net40));
 sg13g2_buf_1 input41 (.A(Tile_X0Y0_S2MID[3]),
    .X(net41));
 sg13g2_buf_1 input42 (.A(Tile_X0Y0_S2MID[4]),
    .X(net42));
 sg13g2_buf_1 input43 (.A(Tile_X0Y0_S2MID[5]),
    .X(net43));
 sg13g2_buf_1 input44 (.A(Tile_X0Y0_S2MID[6]),
    .X(net44));
 sg13g2_buf_1 input45 (.A(Tile_X0Y0_S2MID[7]),
    .X(net45));
 sg13g2_buf_1 input46 (.A(Tile_X0Y0_S4END[0]),
    .X(net46));
 sg13g2_buf_1 input47 (.A(Tile_X0Y0_S4END[1]),
    .X(net47));
 sg13g2_buf_1 input48 (.A(Tile_X0Y0_S4END[2]),
    .X(net48));
 sg13g2_buf_1 input49 (.A(Tile_X0Y0_S4END[3]),
    .X(net49));
 sg13g2_buf_1 input50 (.A(Tile_X0Y0_S4END[4]),
    .X(net50));
 sg13g2_buf_1 input51 (.A(Tile_X0Y0_S4END[5]),
    .X(net51));
 sg13g2_buf_1 input52 (.A(Tile_X0Y0_S4END[6]),
    .X(net52));
 sg13g2_buf_1 input53 (.A(Tile_X0Y0_S4END[7]),
    .X(net53));
 sg13g2_buf_1 input54 (.A(Tile_X0Y0_SS4END[0]),
    .X(net54));
 sg13g2_buf_1 input55 (.A(Tile_X0Y0_SS4END[1]),
    .X(net55));
 sg13g2_buf_1 input56 (.A(Tile_X0Y0_SS4END[2]),
    .X(net56));
 sg13g2_buf_1 input57 (.A(Tile_X0Y0_SS4END[3]),
    .X(net57));
 sg13g2_buf_1 input58 (.A(Tile_X0Y0_SS4END[4]),
    .X(net58));
 sg13g2_buf_1 input59 (.A(Tile_X0Y0_SS4END[5]),
    .X(net59));
 sg13g2_buf_1 input60 (.A(Tile_X0Y0_SS4END[6]),
    .X(net60));
 sg13g2_buf_1 input61 (.A(Tile_X0Y0_SS4END[7]),
    .X(net61));
 sg13g2_buf_1 input62 (.A(Tile_X0Y0_W1END[0]),
    .X(net62));
 sg13g2_buf_1 input63 (.A(Tile_X0Y0_W1END[1]),
    .X(net63));
 sg13g2_buf_1 input64 (.A(Tile_X0Y0_W1END[2]),
    .X(net64));
 sg13g2_buf_1 input65 (.A(Tile_X0Y0_W2END[0]),
    .X(net65));
 sg13g2_buf_1 input66 (.A(Tile_X0Y0_W2END[1]),
    .X(net66));
 sg13g2_buf_8 input67 (.A(Tile_X0Y0_W2END[2]),
    .X(net67));
 sg13g2_buf_1 input68 (.A(Tile_X0Y0_W2END[3]),
    .X(net68));
 sg13g2_buf_1 input69 (.A(Tile_X0Y0_W2END[4]),
    .X(net69));
 sg13g2_buf_1 input70 (.A(Tile_X0Y0_W2END[5]),
    .X(net70));
 sg13g2_buf_1 input71 (.A(Tile_X0Y0_W2END[6]),
    .X(net71));
 sg13g2_buf_1 input72 (.A(Tile_X0Y0_W2END[7]),
    .X(net72));
 sg13g2_buf_1 input73 (.A(Tile_X0Y0_W2MID[0]),
    .X(net73));
 sg13g2_buf_1 input74 (.A(Tile_X0Y0_W2MID[1]),
    .X(net74));
 sg13g2_buf_1 input75 (.A(Tile_X0Y0_W2MID[2]),
    .X(net75));
 sg13g2_buf_1 input76 (.A(Tile_X0Y0_W2MID[3]),
    .X(net76));
 sg13g2_buf_1 input77 (.A(Tile_X0Y0_W2MID[4]),
    .X(net77));
 sg13g2_buf_1 input78 (.A(Tile_X0Y0_W2MID[5]),
    .X(net78));
 sg13g2_buf_1 input79 (.A(Tile_X0Y0_W2MID[6]),
    .X(net79));
 sg13g2_buf_1 input80 (.A(Tile_X0Y0_W2MID[7]),
    .X(net80));
 sg13g2_buf_8 input81 (.A(Tile_X0Y0_W6END[0]),
    .X(net81));
 sg13g2_buf_1 input82 (.A(Tile_X0Y0_W6END[1]),
    .X(net82));
 sg13g2_buf_1 input83 (.A(Tile_X0Y0_WW4END[0]),
    .X(net83));
 sg13g2_buf_1 input84 (.A(Tile_X0Y0_WW4END[1]),
    .X(net84));
 sg13g2_buf_1 input85 (.A(Tile_X0Y0_WW4END[2]),
    .X(net85));
 sg13g2_buf_1 input86 (.A(Tile_X0Y0_WW4END[3]),
    .X(net86));
 sg13g2_buf_1 input87 (.A(Tile_X0Y1_E1END[0]),
    .X(net87));
 sg13g2_buf_1 input88 (.A(Tile_X0Y1_E1END[1]),
    .X(net88));
 sg13g2_buf_1 input89 (.A(Tile_X0Y1_E1END[2]),
    .X(net89));
 sg13g2_buf_1 input90 (.A(Tile_X0Y1_E1END[3]),
    .X(net90));
 sg13g2_buf_1 input91 (.A(Tile_X0Y1_E2END[0]),
    .X(net91));
 sg13g2_buf_1 input92 (.A(Tile_X0Y1_E2END[1]),
    .X(net92));
 sg13g2_buf_1 input93 (.A(Tile_X0Y1_E2END[2]),
    .X(net93));
 sg13g2_buf_1 input94 (.A(Tile_X0Y1_E2END[3]),
    .X(net94));
 sg13g2_buf_1 input95 (.A(Tile_X0Y1_E2END[4]),
    .X(net95));
 sg13g2_buf_1 input96 (.A(Tile_X0Y1_E2END[5]),
    .X(net96));
 sg13g2_buf_1 input97 (.A(Tile_X0Y1_E2END[6]),
    .X(net97));
 sg13g2_buf_1 input98 (.A(Tile_X0Y1_E2END[7]),
    .X(net98));
 sg13g2_buf_1 input99 (.A(Tile_X0Y1_E2MID[0]),
    .X(net99));
 sg13g2_buf_1 input100 (.A(Tile_X0Y1_E2MID[1]),
    .X(net100));
 sg13g2_buf_1 input101 (.A(Tile_X0Y1_E2MID[2]),
    .X(net101));
 sg13g2_buf_1 input102 (.A(Tile_X0Y1_E2MID[3]),
    .X(net102));
 sg13g2_buf_1 input103 (.A(Tile_X0Y1_E2MID[4]),
    .X(net103));
 sg13g2_buf_1 input104 (.A(Tile_X0Y1_E2MID[5]),
    .X(net104));
 sg13g2_buf_1 input105 (.A(Tile_X0Y1_E2MID[6]),
    .X(net105));
 sg13g2_buf_1 input106 (.A(Tile_X0Y1_E2MID[7]),
    .X(net106));
 sg13g2_buf_1 input107 (.A(Tile_X0Y1_EE4END[0]),
    .X(net107));
 sg13g2_buf_1 input108 (.A(Tile_X0Y1_EE4END[1]),
    .X(net108));
 sg13g2_buf_1 input109 (.A(Tile_X0Y1_EE4END[2]),
    .X(net109));
 sg13g2_buf_1 input110 (.A(Tile_X0Y1_EE4END[3]),
    .X(net110));
 sg13g2_buf_1 input111 (.A(Tile_X0Y1_N1END[0]),
    .X(net111));
 sg13g2_buf_1 input112 (.A(Tile_X0Y1_N1END[1]),
    .X(net112));
 sg13g2_buf_1 input113 (.A(Tile_X0Y1_N1END[2]),
    .X(net113));
 sg13g2_buf_1 input114 (.A(Tile_X0Y1_N1END[3]),
    .X(net114));
 sg13g2_buf_1 input115 (.A(Tile_X0Y1_N2END[0]),
    .X(net115));
 sg13g2_buf_1 input116 (.A(Tile_X0Y1_N2END[1]),
    .X(net116));
 sg13g2_buf_1 input117 (.A(Tile_X0Y1_N2END[2]),
    .X(net117));
 sg13g2_buf_1 input118 (.A(Tile_X0Y1_N2END[3]),
    .X(net118));
 sg13g2_buf_1 input119 (.A(Tile_X0Y1_N2END[4]),
    .X(net119));
 sg13g2_buf_1 input120 (.A(Tile_X0Y1_N2END[5]),
    .X(net120));
 sg13g2_buf_1 input121 (.A(Tile_X0Y1_N2END[6]),
    .X(net121));
 sg13g2_buf_1 input122 (.A(Tile_X0Y1_N2END[7]),
    .X(net122));
 sg13g2_buf_1 input123 (.A(Tile_X0Y1_N2MID[0]),
    .X(net123));
 sg13g2_buf_1 input124 (.A(Tile_X0Y1_N2MID[1]),
    .X(net124));
 sg13g2_buf_8 input125 (.A(Tile_X0Y1_N2MID[2]),
    .X(net125));
 sg13g2_buf_1 input126 (.A(Tile_X0Y1_N2MID[3]),
    .X(net126));
 sg13g2_buf_1 input127 (.A(Tile_X0Y1_N2MID[4]),
    .X(net127));
 sg13g2_buf_1 input128 (.A(Tile_X0Y1_N2MID[5]),
    .X(net128));
 sg13g2_buf_1 input129 (.A(Tile_X0Y1_N2MID[6]),
    .X(net129));
 sg13g2_buf_1 input130 (.A(Tile_X0Y1_N2MID[7]),
    .X(net130));
 sg13g2_buf_1 input131 (.A(Tile_X0Y1_N4END[0]),
    .X(net131));
 sg13g2_buf_1 input132 (.A(Tile_X0Y1_N4END[1]),
    .X(net132));
 sg13g2_buf_1 input133 (.A(Tile_X0Y1_N4END[2]),
    .X(net133));
 sg13g2_buf_1 input134 (.A(Tile_X0Y1_N4END[3]),
    .X(net134));
 sg13g2_buf_1 input135 (.A(Tile_X0Y1_N4END[4]),
    .X(net135));
 sg13g2_buf_1 input136 (.A(Tile_X0Y1_N4END[5]),
    .X(net136));
 sg13g2_buf_16 input137 (.X(net137),
    .A(Tile_X0Y1_N4END[6]));
 sg13g2_buf_1 input138 (.A(Tile_X0Y1_N4END[7]),
    .X(net138));
 sg13g2_buf_1 input139 (.A(Tile_X0Y1_NN4END[0]),
    .X(net139));
 sg13g2_buf_1 input140 (.A(Tile_X0Y1_NN4END[1]),
    .X(net140));
 sg13g2_buf_1 input141 (.A(Tile_X0Y1_NN4END[2]),
    .X(net141));
 sg13g2_buf_1 input142 (.A(Tile_X0Y1_NN4END[3]),
    .X(net142));
 sg13g2_buf_1 input143 (.A(Tile_X0Y1_NN4END[4]),
    .X(net143));
 sg13g2_buf_1 input144 (.A(Tile_X0Y1_NN4END[5]),
    .X(net144));
 sg13g2_buf_1 input145 (.A(Tile_X0Y1_NN4END[6]),
    .X(net145));
 sg13g2_buf_1 input146 (.A(Tile_X0Y1_NN4END[7]),
    .X(net146));
 sg13g2_buf_1 input147 (.A(Tile_X0Y1_W1END[0]),
    .X(net147));
 sg13g2_buf_1 input148 (.A(Tile_X0Y1_W1END[1]),
    .X(net148));
 sg13g2_buf_1 input149 (.A(Tile_X0Y1_W1END[2]),
    .X(net149));
 sg13g2_buf_1 input150 (.A(Tile_X0Y1_W1END[3]),
    .X(net150));
 sg13g2_buf_1 input151 (.A(Tile_X0Y1_W2END[0]),
    .X(net151));
 sg13g2_buf_1 input152 (.A(Tile_X0Y1_W2END[1]),
    .X(net152));
 sg13g2_buf_1 input153 (.A(Tile_X0Y1_W2END[2]),
    .X(net153));
 sg13g2_buf_1 input154 (.A(Tile_X0Y1_W2END[3]),
    .X(net154));
 sg13g2_buf_1 input155 (.A(Tile_X0Y1_W2END[4]),
    .X(net155));
 sg13g2_buf_1 input156 (.A(Tile_X0Y1_W2END[5]),
    .X(net156));
 sg13g2_buf_1 input157 (.A(Tile_X0Y1_W2END[6]),
    .X(net157));
 sg13g2_buf_1 input158 (.A(Tile_X0Y1_W2END[7]),
    .X(net158));
 sg13g2_buf_1 input159 (.A(Tile_X0Y1_W2MID[0]),
    .X(net159));
 sg13g2_buf_1 input160 (.A(Tile_X0Y1_W2MID[1]),
    .X(net160));
 sg13g2_buf_1 input161 (.A(Tile_X0Y1_W2MID[2]),
    .X(net161));
 sg13g2_buf_1 input162 (.A(Tile_X0Y1_W2MID[3]),
    .X(net162));
 sg13g2_buf_1 input163 (.A(Tile_X0Y1_W2MID[4]),
    .X(net163));
 sg13g2_buf_1 input164 (.A(Tile_X0Y1_W2MID[5]),
    .X(net164));
 sg13g2_buf_1 input165 (.A(Tile_X0Y1_W2MID[6]),
    .X(net165));
 sg13g2_buf_1 input166 (.A(Tile_X0Y1_W2MID[7]),
    .X(net166));
 sg13g2_buf_1 input167 (.A(Tile_X0Y1_W6END[0]),
    .X(net167));
 sg13g2_buf_1 input168 (.A(Tile_X0Y1_W6END[1]),
    .X(net168));
 sg13g2_buf_1 input169 (.A(Tile_X0Y1_WW4END[0]),
    .X(net169));
 sg13g2_buf_1 input170 (.A(Tile_X0Y1_WW4END[1]),
    .X(net170));
 sg13g2_buf_1 input171 (.A(Tile_X0Y1_WW4END[2]),
    .X(net171));
 sg13g2_buf_1 input172 (.A(Tile_X0Y1_WW4END[3]),
    .X(net172));
 sg13g2_buf_1 output173 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG0 ),
    .X(Tile_X0Y0_E1BEG[0]));
 sg13g2_buf_1 output174 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E1BEG1 ),
    .X(Tile_X0Y0_E1BEG[1]));
 sg13g2_buf_1 output175 (.A(net175),
    .X(Tile_X0Y0_E1BEG[2]));
 sg13g2_buf_1 output176 (.A(net176),
    .X(Tile_X0Y0_E1BEG[3]));
 sg13g2_buf_1 output177 (.A(net177),
    .X(Tile_X0Y0_E2BEG[0]));
 sg13g2_buf_1 output178 (.A(net178),
    .X(Tile_X0Y0_E2BEG[1]));
 sg13g2_buf_1 output179 (.A(net179),
    .X(Tile_X0Y0_E2BEG[2]));
 sg13g2_buf_1 output180 (.A(net180),
    .X(Tile_X0Y0_E2BEG[3]));
 sg13g2_buf_1 output181 (.A(net181),
    .X(Tile_X0Y0_E2BEG[4]));
 sg13g2_buf_1 output182 (.A(net182),
    .X(Tile_X0Y0_E2BEG[5]));
 sg13g2_buf_1 output183 (.A(net183),
    .X(Tile_X0Y0_E2BEG[6]));
 sg13g2_buf_1 output184 (.A(net184),
    .X(Tile_X0Y0_E2BEG[7]));
 sg13g2_buf_1 output185 (.A(net185),
    .X(Tile_X0Y0_E2BEGb[0]));
 sg13g2_buf_1 output186 (.A(net186),
    .X(Tile_X0Y0_E2BEGb[1]));
 sg13g2_buf_1 output187 (.A(net187),
    .X(Tile_X0Y0_E2BEGb[2]));
 sg13g2_buf_1 output188 (.A(net188),
    .X(Tile_X0Y0_E2BEGb[3]));
 sg13g2_buf_1 output189 (.A(net189),
    .X(Tile_X0Y0_E2BEGb[4]));
 sg13g2_buf_1 output190 (.A(net190),
    .X(Tile_X0Y0_E2BEGb[5]));
 sg13g2_buf_1 output191 (.A(net191),
    .X(Tile_X0Y0_E2BEGb[6]));
 sg13g2_buf_1 output192 (.A(net192),
    .X(Tile_X0Y0_E2BEGb[7]));
 sg13g2_buf_1 output193 (.A(net193),
    .X(Tile_X0Y0_E6BEG[0]));
 sg13g2_buf_1 output194 (.A(net194),
    .X(Tile_X0Y0_E6BEG[10]));
 sg13g2_buf_1 output195 (.A(net195),
    .X(Tile_X0Y0_E6BEG[11]));
 sg13g2_buf_1 output196 (.A(net196),
    .X(Tile_X0Y0_E6BEG[1]));
 sg13g2_buf_1 output197 (.A(net197),
    .X(Tile_X0Y0_E6BEG[2]));
 sg13g2_buf_1 output198 (.A(net198),
    .X(Tile_X0Y0_E6BEG[3]));
 sg13g2_buf_1 output199 (.A(net199),
    .X(Tile_X0Y0_E6BEG[4]));
 sg13g2_buf_1 output200 (.A(net200),
    .X(Tile_X0Y0_E6BEG[5]));
 sg13g2_buf_1 output201 (.A(net201),
    .X(Tile_X0Y0_E6BEG[6]));
 sg13g2_buf_1 output202 (.A(net202),
    .X(Tile_X0Y0_E6BEG[7]));
 sg13g2_buf_1 output203 (.A(net203),
    .X(Tile_X0Y0_E6BEG[8]));
 sg13g2_buf_1 output204 (.A(net204),
    .X(Tile_X0Y0_E6BEG[9]));
 sg13g2_buf_1 output205 (.A(net205),
    .X(Tile_X0Y0_EE4BEG[0]));
 sg13g2_buf_1 output206 (.A(net206),
    .X(Tile_X0Y0_EE4BEG[10]));
 sg13g2_buf_1 output207 (.A(net207),
    .X(Tile_X0Y0_EE4BEG[11]));
 sg13g2_buf_1 output208 (.A(net208),
    .X(Tile_X0Y0_EE4BEG[12]));
 sg13g2_buf_1 output209 (.A(net209),
    .X(Tile_X0Y0_EE4BEG[13]));
 sg13g2_buf_1 output210 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.EE4BEG2 ),
    .X(Tile_X0Y0_EE4BEG[14]));
 sg13g2_buf_1 output211 (.A(net211),
    .X(Tile_X0Y0_EE4BEG[15]));
 sg13g2_buf_1 output212 (.A(net212),
    .X(Tile_X0Y0_EE4BEG[1]));
 sg13g2_buf_1 output213 (.A(net213),
    .X(Tile_X0Y0_EE4BEG[2]));
 sg13g2_buf_1 output214 (.A(net214),
    .X(Tile_X0Y0_EE4BEG[3]));
 sg13g2_buf_1 output215 (.A(net215),
    .X(Tile_X0Y0_EE4BEG[4]));
 sg13g2_buf_1 output216 (.A(net216),
    .X(Tile_X0Y0_EE4BEG[5]));
 sg13g2_buf_1 output217 (.A(net217),
    .X(Tile_X0Y0_EE4BEG[6]));
 sg13g2_buf_1 output218 (.A(net218),
    .X(Tile_X0Y0_EE4BEG[7]));
 sg13g2_buf_1 output219 (.A(net219),
    .X(Tile_X0Y0_EE4BEG[8]));
 sg13g2_buf_1 output220 (.A(net220),
    .X(Tile_X0Y0_EE4BEG[9]));
 sg13g2_buf_1 output221 (.A(net221),
    .X(Tile_X0Y0_FrameData_O[0]));
 sg13g2_buf_1 output222 (.A(net222),
    .X(Tile_X0Y0_FrameData_O[10]));
 sg13g2_buf_1 output223 (.A(net223),
    .X(Tile_X0Y0_FrameData_O[11]));
 sg13g2_buf_1 output224 (.A(net224),
    .X(Tile_X0Y0_FrameData_O[12]));
 sg13g2_buf_1 output225 (.A(net225),
    .X(Tile_X0Y0_FrameData_O[13]));
 sg13g2_buf_1 output226 (.A(net226),
    .X(Tile_X0Y0_FrameData_O[14]));
 sg13g2_buf_1 output227 (.A(net227),
    .X(Tile_X0Y0_FrameData_O[15]));
 sg13g2_buf_1 output228 (.A(net228),
    .X(Tile_X0Y0_FrameData_O[16]));
 sg13g2_buf_1 output229 (.A(net229),
    .X(Tile_X0Y0_FrameData_O[17]));
 sg13g2_buf_1 output230 (.A(net230),
    .X(Tile_X0Y0_FrameData_O[18]));
 sg13g2_buf_1 output231 (.A(net231),
    .X(Tile_X0Y0_FrameData_O[19]));
 sg13g2_buf_1 output232 (.A(net232),
    .X(Tile_X0Y0_FrameData_O[1]));
 sg13g2_buf_1 output233 (.A(net233),
    .X(Tile_X0Y0_FrameData_O[20]));
 sg13g2_buf_1 output234 (.A(net234),
    .X(Tile_X0Y0_FrameData_O[21]));
 sg13g2_buf_1 output235 (.A(net235),
    .X(Tile_X0Y0_FrameData_O[22]));
 sg13g2_buf_1 output236 (.A(net236),
    .X(Tile_X0Y0_FrameData_O[23]));
 sg13g2_buf_1 output237 (.A(net237),
    .X(Tile_X0Y0_FrameData_O[24]));
 sg13g2_buf_1 output238 (.A(net238),
    .X(Tile_X0Y0_FrameData_O[25]));
 sg13g2_buf_1 output239 (.A(net239),
    .X(Tile_X0Y0_FrameData_O[26]));
 sg13g2_buf_1 output240 (.A(net240),
    .X(Tile_X0Y0_FrameData_O[27]));
 sg13g2_buf_1 output241 (.A(net241),
    .X(Tile_X0Y0_FrameData_O[28]));
 sg13g2_buf_1 output242 (.A(net242),
    .X(Tile_X0Y0_FrameData_O[29]));
 sg13g2_buf_1 output243 (.A(net243),
    .X(Tile_X0Y0_FrameData_O[2]));
 sg13g2_buf_1 output244 (.A(net244),
    .X(Tile_X0Y0_FrameData_O[30]));
 sg13g2_buf_1 output245 (.A(net245),
    .X(Tile_X0Y0_FrameData_O[31]));
 sg13g2_buf_1 output246 (.A(net246),
    .X(Tile_X0Y0_FrameData_O[3]));
 sg13g2_buf_1 output247 (.A(net247),
    .X(Tile_X0Y0_FrameData_O[4]));
 sg13g2_buf_1 output248 (.A(net248),
    .X(Tile_X0Y0_FrameData_O[5]));
 sg13g2_buf_1 output249 (.A(net249),
    .X(Tile_X0Y0_FrameData_O[6]));
 sg13g2_buf_1 output250 (.A(net250),
    .X(Tile_X0Y0_FrameData_O[7]));
 sg13g2_buf_1 output251 (.A(net251),
    .X(Tile_X0Y0_FrameData_O[8]));
 sg13g2_buf_1 output252 (.A(net252),
    .X(Tile_X0Y0_FrameData_O[9]));
 sg13g2_buf_1 output253 (.A(net253),
    .X(Tile_X0Y0_FrameStrobe_O[0]));
 sg13g2_buf_1 output254 (.A(net254),
    .X(Tile_X0Y0_FrameStrobe_O[10]));
 sg13g2_buf_1 output255 (.A(net255),
    .X(Tile_X0Y0_FrameStrobe_O[11]));
 sg13g2_buf_1 output256 (.A(net256),
    .X(Tile_X0Y0_FrameStrobe_O[12]));
 sg13g2_buf_1 output257 (.A(net257),
    .X(Tile_X0Y0_FrameStrobe_O[13]));
 sg13g2_buf_1 output258 (.A(net258),
    .X(Tile_X0Y0_FrameStrobe_O[14]));
 sg13g2_buf_1 output259 (.A(net259),
    .X(Tile_X0Y0_FrameStrobe_O[15]));
 sg13g2_buf_1 output260 (.A(net260),
    .X(Tile_X0Y0_FrameStrobe_O[16]));
 sg13g2_buf_1 output261 (.A(net261),
    .X(Tile_X0Y0_FrameStrobe_O[17]));
 sg13g2_buf_1 output262 (.A(net262),
    .X(Tile_X0Y0_FrameStrobe_O[18]));
 sg13g2_buf_1 output263 (.A(net263),
    .X(Tile_X0Y0_FrameStrobe_O[19]));
 sg13g2_buf_1 output264 (.A(net264),
    .X(Tile_X0Y0_FrameStrobe_O[1]));
 sg13g2_buf_1 output265 (.A(net265),
    .X(Tile_X0Y0_FrameStrobe_O[2]));
 sg13g2_buf_1 output266 (.A(net266),
    .X(Tile_X0Y0_FrameStrobe_O[3]));
 sg13g2_buf_1 output267 (.A(net267),
    .X(Tile_X0Y0_FrameStrobe_O[4]));
 sg13g2_buf_1 output268 (.A(net268),
    .X(Tile_X0Y0_FrameStrobe_O[5]));
 sg13g2_buf_1 output269 (.A(net269),
    .X(Tile_X0Y0_FrameStrobe_O[6]));
 sg13g2_buf_1 output270 (.A(net270),
    .X(Tile_X0Y0_FrameStrobe_O[7]));
 sg13g2_buf_1 output271 (.A(net271),
    .X(Tile_X0Y0_FrameStrobe_O[8]));
 sg13g2_buf_1 output272 (.A(net272),
    .X(Tile_X0Y0_FrameStrobe_O[9]));
 sg13g2_buf_1 output273 (.A(net273),
    .X(Tile_X0Y0_N1BEG[0]));
 sg13g2_buf_1 output274 (.A(net274),
    .X(Tile_X0Y0_N1BEG[1]));
 sg13g2_buf_1 output275 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 ),
    .X(Tile_X0Y0_N1BEG[2]));
 sg13g2_buf_8 output276 (.A(net276),
    .X(Tile_X0Y0_N1BEG[3]));
 sg13g2_buf_1 output277 (.A(net277),
    .X(Tile_X0Y0_N2BEG[0]));
 sg13g2_buf_1 output278 (.A(net278),
    .X(Tile_X0Y0_N2BEG[1]));
 sg13g2_buf_1 output279 (.A(net279),
    .X(Tile_X0Y0_N2BEG[2]));
 sg13g2_buf_1 output280 (.A(net280),
    .X(Tile_X0Y0_N2BEG[3]));
 sg13g2_buf_1 output281 (.A(net281),
    .X(Tile_X0Y0_N2BEG[4]));
 sg13g2_buf_1 output282 (.A(net282),
    .X(Tile_X0Y0_N2BEG[5]));
 sg13g2_buf_1 output283 (.A(net283),
    .X(Tile_X0Y0_N2BEG[6]));
 sg13g2_buf_1 output284 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 ),
    .X(Tile_X0Y0_N2BEG[7]));
 sg13g2_buf_1 output285 (.A(net285),
    .X(Tile_X0Y0_N2BEGb[0]));
 sg13g2_buf_1 output286 (.A(net286),
    .X(Tile_X0Y0_N2BEGb[1]));
 sg13g2_buf_1 output287 (.A(net287),
    .X(Tile_X0Y0_N2BEGb[2]));
 sg13g2_buf_1 output288 (.A(net288),
    .X(Tile_X0Y0_N2BEGb[3]));
 sg13g2_buf_8 output289 (.A(net289),
    .X(Tile_X0Y0_N2BEGb[4]));
 sg13g2_buf_1 output290 (.A(net290),
    .X(Tile_X0Y0_N2BEGb[5]));
 sg13g2_buf_1 output291 (.A(net291),
    .X(Tile_X0Y0_N2BEGb[6]));
 sg13g2_buf_1 output292 (.A(net292),
    .X(Tile_X0Y0_N2BEGb[7]));
 sg13g2_buf_1 output293 (.A(net293),
    .X(Tile_X0Y0_N4BEG[0]));
 sg13g2_buf_1 output294 (.A(net294),
    .X(Tile_X0Y0_N4BEG[10]));
 sg13g2_buf_1 output295 (.A(net295),
    .X(Tile_X0Y0_N4BEG[11]));
 sg13g2_buf_1 output296 (.A(net296),
    .X(Tile_X0Y0_N4BEG[12]));
 sg13g2_buf_1 output297 (.A(net297),
    .X(Tile_X0Y0_N4BEG[13]));
 sg13g2_buf_1 output298 (.A(net298),
    .X(Tile_X0Y0_N4BEG[14]));
 sg13g2_buf_1 output299 (.A(net299),
    .X(Tile_X0Y0_N4BEG[15]));
 sg13g2_buf_1 output300 (.A(net300),
    .X(Tile_X0Y0_N4BEG[1]));
 sg13g2_buf_1 output301 (.A(net301),
    .X(Tile_X0Y0_N4BEG[2]));
 sg13g2_buf_1 output302 (.A(net302),
    .X(Tile_X0Y0_N4BEG[3]));
 sg13g2_buf_1 output303 (.A(net303),
    .X(Tile_X0Y0_N4BEG[4]));
 sg13g2_buf_1 output304 (.A(net304),
    .X(Tile_X0Y0_N4BEG[5]));
 sg13g2_buf_1 output305 (.A(net305),
    .X(Tile_X0Y0_N4BEG[6]));
 sg13g2_buf_1 output306 (.A(net306),
    .X(Tile_X0Y0_N4BEG[7]));
 sg13g2_buf_1 output307 (.A(net307),
    .X(Tile_X0Y0_N4BEG[8]));
 sg13g2_buf_1 output308 (.A(net308),
    .X(Tile_X0Y0_N4BEG[9]));
 sg13g2_buf_1 output309 (.A(net309),
    .X(Tile_X0Y0_NN4BEG[0]));
 sg13g2_buf_1 output310 (.A(net310),
    .X(Tile_X0Y0_NN4BEG[10]));
 sg13g2_buf_1 output311 (.A(net311),
    .X(Tile_X0Y0_NN4BEG[11]));
 sg13g2_buf_1 output312 (.A(net312),
    .X(Tile_X0Y0_NN4BEG[12]));
 sg13g2_buf_1 output313 (.A(net313),
    .X(Tile_X0Y0_NN4BEG[13]));
 sg13g2_buf_1 output314 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 ),
    .X(Tile_X0Y0_NN4BEG[14]));
 sg13g2_buf_1 output315 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 ),
    .X(Tile_X0Y0_NN4BEG[15]));
 sg13g2_buf_1 output316 (.A(net316),
    .X(Tile_X0Y0_NN4BEG[1]));
 sg13g2_buf_1 output317 (.A(net317),
    .X(Tile_X0Y0_NN4BEG[2]));
 sg13g2_buf_1 output318 (.A(net318),
    .X(Tile_X0Y0_NN4BEG[3]));
 sg13g2_buf_1 output319 (.A(net319),
    .X(Tile_X0Y0_NN4BEG[4]));
 sg13g2_buf_1 output320 (.A(net320),
    .X(Tile_X0Y0_NN4BEG[5]));
 sg13g2_buf_1 output321 (.A(net321),
    .X(Tile_X0Y0_NN4BEG[6]));
 sg13g2_buf_1 output322 (.A(net322),
    .X(Tile_X0Y0_NN4BEG[7]));
 sg13g2_buf_1 output323 (.A(net323),
    .X(Tile_X0Y0_NN4BEG[8]));
 sg13g2_buf_1 output324 (.A(net324),
    .X(Tile_X0Y0_NN4BEG[9]));
 sg13g2_buf_1 output325 (.A(net325),
    .X(Tile_X0Y0_UserCLKo));
 sg13g2_buf_1 output326 (.A(net326),
    .X(Tile_X0Y0_W1BEG[0]));
 sg13g2_buf_1 output327 (.A(net327),
    .X(Tile_X0Y0_W1BEG[1]));
 sg13g2_buf_1 output328 (.A(net328),
    .X(Tile_X0Y0_W1BEG[2]));
 sg13g2_buf_1 output329 (.A(net329),
    .X(Tile_X0Y0_W1BEG[3]));
 sg13g2_buf_1 output330 (.A(net330),
    .X(Tile_X0Y0_W2BEG[0]));
 sg13g2_buf_1 output331 (.A(net331),
    .X(Tile_X0Y0_W2BEG[1]));
 sg13g2_buf_1 output332 (.A(net332),
    .X(Tile_X0Y0_W2BEG[2]));
 sg13g2_buf_1 output333 (.A(net333),
    .X(Tile_X0Y0_W2BEG[3]));
 sg13g2_buf_1 output334 (.A(net334),
    .X(Tile_X0Y0_W2BEG[4]));
 sg13g2_buf_1 output335 (.A(net335),
    .X(Tile_X0Y0_W2BEG[5]));
 sg13g2_buf_1 output336 (.A(net336),
    .X(Tile_X0Y0_W2BEG[6]));
 sg13g2_buf_1 output337 (.A(net337),
    .X(Tile_X0Y0_W2BEG[7]));
 sg13g2_buf_1 output338 (.A(net338),
    .X(Tile_X0Y0_W2BEGb[0]));
 sg13g2_buf_1 output339 (.A(net339),
    .X(Tile_X0Y0_W2BEGb[1]));
 sg13g2_buf_1 output340 (.A(net340),
    .X(Tile_X0Y0_W2BEGb[2]));
 sg13g2_buf_1 output341 (.A(net341),
    .X(Tile_X0Y0_W2BEGb[3]));
 sg13g2_buf_1 output342 (.A(net342),
    .X(Tile_X0Y0_W2BEGb[4]));
 sg13g2_buf_1 output343 (.A(net343),
    .X(Tile_X0Y0_W2BEGb[5]));
 sg13g2_buf_1 output344 (.A(net344),
    .X(Tile_X0Y0_W2BEGb[6]));
 sg13g2_buf_1 output345 (.A(net345),
    .X(Tile_X0Y0_W2BEGb[7]));
 sg13g2_buf_1 output346 (.A(net346),
    .X(Tile_X0Y0_W6BEG[0]));
 sg13g2_buf_1 output347 (.A(net347),
    .X(Tile_X0Y0_W6BEG[10]));
 sg13g2_buf_1 output348 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 ),
    .X(Tile_X0Y0_W6BEG[11]));
 sg13g2_buf_1 output349 (.A(net349),
    .X(Tile_X0Y0_W6BEG[1]));
 sg13g2_buf_1 output350 (.A(net350),
    .X(Tile_X0Y0_W6BEG[2]));
 sg13g2_buf_1 output351 (.A(net351),
    .X(Tile_X0Y0_W6BEG[3]));
 sg13g2_buf_1 output352 (.A(net352),
    .X(Tile_X0Y0_W6BEG[4]));
 sg13g2_buf_1 output353 (.A(net353),
    .X(Tile_X0Y0_W6BEG[5]));
 sg13g2_buf_1 output354 (.A(net354),
    .X(Tile_X0Y0_W6BEG[6]));
 sg13g2_buf_1 output355 (.A(net355),
    .X(Tile_X0Y0_W6BEG[7]));
 sg13g2_buf_1 output356 (.A(net356),
    .X(Tile_X0Y0_W6BEG[8]));
 sg13g2_buf_1 output357 (.A(net357),
    .X(Tile_X0Y0_W6BEG[9]));
 sg13g2_buf_1 output358 (.A(net358),
    .X(Tile_X0Y0_WW4BEG[0]));
 sg13g2_buf_1 output359 (.A(net359),
    .X(Tile_X0Y0_WW4BEG[10]));
 sg13g2_buf_1 output360 (.A(net360),
    .X(Tile_X0Y0_WW4BEG[11]));
 sg13g2_buf_1 output361 (.A(net361),
    .X(Tile_X0Y0_WW4BEG[12]));
 sg13g2_buf_1 output362 (.A(net362),
    .X(Tile_X0Y0_WW4BEG[13]));
 sg13g2_buf_1 output363 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 ),
    .X(Tile_X0Y0_WW4BEG[14]));
 sg13g2_buf_8 output364 (.A(net364),
    .X(Tile_X0Y0_WW4BEG[15]));
 sg13g2_buf_1 output365 (.A(net365),
    .X(Tile_X0Y0_WW4BEG[1]));
 sg13g2_buf_1 output366 (.A(net366),
    .X(Tile_X0Y0_WW4BEG[2]));
 sg13g2_buf_1 output367 (.A(net367),
    .X(Tile_X0Y0_WW4BEG[3]));
 sg13g2_buf_1 output368 (.A(net368),
    .X(Tile_X0Y0_WW4BEG[4]));
 sg13g2_buf_1 output369 (.A(net369),
    .X(Tile_X0Y0_WW4BEG[5]));
 sg13g2_buf_1 output370 (.A(net370),
    .X(Tile_X0Y0_WW4BEG[6]));
 sg13g2_buf_1 output371 (.A(net371),
    .X(Tile_X0Y0_WW4BEG[7]));
 sg13g2_buf_1 output372 (.A(net372),
    .X(Tile_X0Y0_WW4BEG[8]));
 sg13g2_buf_1 output373 (.A(net373),
    .X(Tile_X0Y0_WW4BEG[9]));
 sg13g2_buf_1 output374 (.A(net374),
    .X(Tile_X0Y1_E1BEG[0]));
 sg13g2_buf_1 output375 (.A(net375),
    .X(Tile_X0Y1_E1BEG[1]));
 sg13g2_buf_1 output376 (.A(net376),
    .X(Tile_X0Y1_E1BEG[2]));
 sg13g2_buf_1 output377 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E1BEG3 ),
    .X(Tile_X0Y1_E1BEG[3]));
 sg13g2_buf_1 output378 (.A(net378),
    .X(Tile_X0Y1_E2BEG[0]));
 sg13g2_buf_1 output379 (.A(net379),
    .X(Tile_X0Y1_E2BEG[1]));
 sg13g2_buf_1 output380 (.A(net380),
    .X(Tile_X0Y1_E2BEG[2]));
 sg13g2_buf_1 output381 (.A(net381),
    .X(Tile_X0Y1_E2BEG[3]));
 sg13g2_buf_1 output382 (.A(net382),
    .X(Tile_X0Y1_E2BEG[4]));
 sg13g2_buf_1 output383 (.A(net383),
    .X(Tile_X0Y1_E2BEG[5]));
 sg13g2_buf_1 output384 (.A(net384),
    .X(Tile_X0Y1_E2BEG[6]));
 sg13g2_buf_8 output385 (.A(net385),
    .X(Tile_X0Y1_E2BEG[7]));
 sg13g2_buf_1 output386 (.A(net386),
    .X(Tile_X0Y1_E2BEGb[0]));
 sg13g2_buf_1 output387 (.A(net387),
    .X(Tile_X0Y1_E2BEGb[1]));
 sg13g2_buf_1 output388 (.A(net388),
    .X(Tile_X0Y1_E2BEGb[2]));
 sg13g2_buf_1 output389 (.A(net389),
    .X(Tile_X0Y1_E2BEGb[3]));
 sg13g2_buf_1 output390 (.A(net390),
    .X(Tile_X0Y1_E2BEGb[4]));
 sg13g2_buf_1 output391 (.A(net391),
    .X(Tile_X0Y1_E2BEGb[5]));
 sg13g2_buf_1 output392 (.A(net392),
    .X(Tile_X0Y1_E2BEGb[6]));
 sg13g2_buf_1 output393 (.A(net393),
    .X(Tile_X0Y1_E2BEGb[7]));
 sg13g2_buf_1 output394 (.A(net394),
    .X(Tile_X0Y1_E6BEG[0]));
 sg13g2_buf_8 output395 (.A(net395),
    .X(Tile_X0Y1_E6BEG[10]));
 sg13g2_buf_1 output396 (.A(net396),
    .X(Tile_X0Y1_E6BEG[11]));
 sg13g2_buf_1 output397 (.A(net397),
    .X(Tile_X0Y1_E6BEG[1]));
 sg13g2_buf_1 output398 (.A(net398),
    .X(Tile_X0Y1_E6BEG[2]));
 sg13g2_buf_1 output399 (.A(net399),
    .X(Tile_X0Y1_E6BEG[3]));
 sg13g2_buf_1 output400 (.A(net400),
    .X(Tile_X0Y1_E6BEG[4]));
 sg13g2_buf_1 output401 (.A(net401),
    .X(Tile_X0Y1_E6BEG[5]));
 sg13g2_buf_1 output402 (.A(net402),
    .X(Tile_X0Y1_E6BEG[6]));
 sg13g2_buf_1 output403 (.A(net403),
    .X(Tile_X0Y1_E6BEG[7]));
 sg13g2_buf_1 output404 (.A(net404),
    .X(Tile_X0Y1_E6BEG[8]));
 sg13g2_buf_1 output405 (.A(net405),
    .X(Tile_X0Y1_E6BEG[9]));
 sg13g2_buf_1 output406 (.A(net406),
    .X(Tile_X0Y1_EE4BEG[0]));
 sg13g2_buf_1 output407 (.A(net407),
    .X(Tile_X0Y1_EE4BEG[10]));
 sg13g2_buf_1 output408 (.A(net408),
    .X(Tile_X0Y1_EE4BEG[11]));
 sg13g2_buf_1 output409 (.A(net409),
    .X(Tile_X0Y1_EE4BEG[12]));
 sg13g2_buf_1 output410 (.A(net410),
    .X(Tile_X0Y1_EE4BEG[13]));
 sg13g2_buf_1 output411 (.A(net411),
    .X(Tile_X0Y1_EE4BEG[14]));
 sg13g2_buf_1 output412 (.A(net412),
    .X(Tile_X0Y1_EE4BEG[15]));
 sg13g2_buf_1 output413 (.A(net413),
    .X(Tile_X0Y1_EE4BEG[1]));
 sg13g2_buf_1 output414 (.A(net414),
    .X(Tile_X0Y1_EE4BEG[2]));
 sg13g2_buf_1 output415 (.A(net415),
    .X(Tile_X0Y1_EE4BEG[3]));
 sg13g2_buf_1 output416 (.A(net416),
    .X(Tile_X0Y1_EE4BEG[4]));
 sg13g2_buf_1 output417 (.A(net417),
    .X(Tile_X0Y1_EE4BEG[5]));
 sg13g2_buf_1 output418 (.A(net418),
    .X(Tile_X0Y1_EE4BEG[6]));
 sg13g2_buf_1 output419 (.A(net419),
    .X(Tile_X0Y1_EE4BEG[7]));
 sg13g2_buf_1 output420 (.A(net420),
    .X(Tile_X0Y1_EE4BEG[8]));
 sg13g2_buf_1 output421 (.A(net421),
    .X(Tile_X0Y1_EE4BEG[9]));
 sg13g2_buf_1 output422 (.A(net422),
    .X(Tile_X0Y1_FrameData_O[0]));
 sg13g2_buf_1 output423 (.A(net423),
    .X(Tile_X0Y1_FrameData_O[10]));
 sg13g2_buf_1 output424 (.A(net424),
    .X(Tile_X0Y1_FrameData_O[11]));
 sg13g2_buf_1 output425 (.A(net425),
    .X(Tile_X0Y1_FrameData_O[12]));
 sg13g2_buf_1 output426 (.A(net426),
    .X(Tile_X0Y1_FrameData_O[13]));
 sg13g2_buf_1 output427 (.A(net427),
    .X(Tile_X0Y1_FrameData_O[14]));
 sg13g2_buf_1 output428 (.A(net428),
    .X(Tile_X0Y1_FrameData_O[15]));
 sg13g2_buf_1 output429 (.A(net429),
    .X(Tile_X0Y1_FrameData_O[16]));
 sg13g2_buf_1 output430 (.A(net430),
    .X(Tile_X0Y1_FrameData_O[17]));
 sg13g2_buf_1 output431 (.A(net431),
    .X(Tile_X0Y1_FrameData_O[18]));
 sg13g2_buf_1 output432 (.A(net432),
    .X(Tile_X0Y1_FrameData_O[19]));
 sg13g2_buf_1 output433 (.A(net433),
    .X(Tile_X0Y1_FrameData_O[1]));
 sg13g2_buf_1 output434 (.A(net434),
    .X(Tile_X0Y1_FrameData_O[20]));
 sg13g2_buf_1 output435 (.A(net435),
    .X(Tile_X0Y1_FrameData_O[21]));
 sg13g2_buf_1 output436 (.A(net436),
    .X(Tile_X0Y1_FrameData_O[22]));
 sg13g2_buf_1 output437 (.A(net437),
    .X(Tile_X0Y1_FrameData_O[23]));
 sg13g2_buf_1 output438 (.A(net438),
    .X(Tile_X0Y1_FrameData_O[24]));
 sg13g2_buf_1 output439 (.A(net439),
    .X(Tile_X0Y1_FrameData_O[25]));
 sg13g2_buf_1 output440 (.A(net440),
    .X(Tile_X0Y1_FrameData_O[26]));
 sg13g2_buf_1 output441 (.A(net441),
    .X(Tile_X0Y1_FrameData_O[27]));
 sg13g2_buf_1 output442 (.A(net442),
    .X(Tile_X0Y1_FrameData_O[28]));
 sg13g2_buf_1 output443 (.A(net443),
    .X(Tile_X0Y1_FrameData_O[29]));
 sg13g2_buf_1 output444 (.A(net444),
    .X(Tile_X0Y1_FrameData_O[2]));
 sg13g2_buf_1 output445 (.A(net445),
    .X(Tile_X0Y1_FrameData_O[30]));
 sg13g2_buf_1 output446 (.A(net446),
    .X(Tile_X0Y1_FrameData_O[31]));
 sg13g2_buf_1 output447 (.A(net447),
    .X(Tile_X0Y1_FrameData_O[3]));
 sg13g2_buf_1 output448 (.A(net448),
    .X(Tile_X0Y1_FrameData_O[4]));
 sg13g2_buf_1 output449 (.A(net449),
    .X(Tile_X0Y1_FrameData_O[5]));
 sg13g2_buf_1 output450 (.A(net450),
    .X(Tile_X0Y1_FrameData_O[6]));
 sg13g2_buf_1 output451 (.A(net451),
    .X(Tile_X0Y1_FrameData_O[7]));
 sg13g2_buf_1 output452 (.A(net452),
    .X(Tile_X0Y1_FrameData_O[8]));
 sg13g2_buf_1 output453 (.A(net453),
    .X(Tile_X0Y1_FrameData_O[9]));
 sg13g2_buf_8 output454 (.A(net454),
    .X(Tile_X0Y1_S1BEG[0]));
 sg13g2_buf_8 output455 (.A(net455),
    .X(Tile_X0Y1_S1BEG[1]));
 sg13g2_buf_1 output456 (.A(net456),
    .X(Tile_X0Y1_S1BEG[2]));
 sg13g2_buf_1 output457 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 ),
    .X(Tile_X0Y1_S1BEG[3]));
 sg13g2_buf_1 output458 (.A(net458),
    .X(Tile_X0Y1_S2BEG[0]));
 sg13g2_buf_1 output459 (.A(net459),
    .X(Tile_X0Y1_S2BEG[1]));
 sg13g2_buf_1 output460 (.A(net460),
    .X(Tile_X0Y1_S2BEG[2]));
 sg13g2_buf_1 output461 (.A(net461),
    .X(Tile_X0Y1_S2BEG[3]));
 sg13g2_buf_1 output462 (.A(net462),
    .X(Tile_X0Y1_S2BEG[4]));
 sg13g2_buf_1 output463 (.A(net463),
    .X(Tile_X0Y1_S2BEG[5]));
 sg13g2_buf_1 output464 (.A(net464),
    .X(Tile_X0Y1_S2BEG[6]));
 sg13g2_buf_1 output465 (.A(net465),
    .X(Tile_X0Y1_S2BEG[7]));
 sg13g2_buf_1 output466 (.A(net466),
    .X(Tile_X0Y1_S2BEGb[0]));
 sg13g2_buf_1 output467 (.A(net467),
    .X(Tile_X0Y1_S2BEGb[1]));
 sg13g2_buf_1 output468 (.A(net468),
    .X(Tile_X0Y1_S2BEGb[2]));
 sg13g2_buf_1 output469 (.A(net469),
    .X(Tile_X0Y1_S2BEGb[3]));
 sg13g2_buf_1 output470 (.A(net470),
    .X(Tile_X0Y1_S2BEGb[4]));
 sg13g2_buf_1 output471 (.A(net471),
    .X(Tile_X0Y1_S2BEGb[5]));
 sg13g2_buf_1 output472 (.A(net472),
    .X(Tile_X0Y1_S2BEGb[6]));
 sg13g2_buf_1 output473 (.A(net473),
    .X(Tile_X0Y1_S2BEGb[7]));
 sg13g2_buf_1 output474 (.A(net474),
    .X(Tile_X0Y1_S4BEG[0]));
 sg13g2_buf_1 output475 (.A(net475),
    .X(Tile_X0Y1_S4BEG[10]));
 sg13g2_buf_1 output476 (.A(net476),
    .X(Tile_X0Y1_S4BEG[11]));
 sg13g2_buf_1 output477 (.A(net477),
    .X(Tile_X0Y1_S4BEG[12]));
 sg13g2_buf_1 output478 (.A(net478),
    .X(Tile_X0Y1_S4BEG[13]));
 sg13g2_buf_1 output479 (.A(net479),
    .X(Tile_X0Y1_S4BEG[14]));
 sg13g2_buf_1 output480 (.A(net480),
    .X(Tile_X0Y1_S4BEG[15]));
 sg13g2_buf_1 output481 (.A(net481),
    .X(Tile_X0Y1_S4BEG[1]));
 sg13g2_buf_1 output482 (.A(net482),
    .X(Tile_X0Y1_S4BEG[2]));
 sg13g2_buf_1 output483 (.A(net483),
    .X(Tile_X0Y1_S4BEG[3]));
 sg13g2_buf_1 output484 (.A(net484),
    .X(Tile_X0Y1_S4BEG[4]));
 sg13g2_buf_1 output485 (.A(net485),
    .X(Tile_X0Y1_S4BEG[5]));
 sg13g2_buf_1 output486 (.A(net486),
    .X(Tile_X0Y1_S4BEG[6]));
 sg13g2_buf_1 output487 (.A(net487),
    .X(Tile_X0Y1_S4BEG[7]));
 sg13g2_buf_1 output488 (.A(net488),
    .X(Tile_X0Y1_S4BEG[8]));
 sg13g2_buf_1 output489 (.A(net489),
    .X(Tile_X0Y1_S4BEG[9]));
 sg13g2_buf_1 output490 (.A(net490),
    .X(Tile_X0Y1_SS4BEG[0]));
 sg13g2_buf_8 output491 (.A(net491),
    .X(Tile_X0Y1_SS4BEG[10]));
 sg13g2_buf_8 output492 (.A(net492),
    .X(Tile_X0Y1_SS4BEG[11]));
 sg13g2_buf_1 output493 (.A(net493),
    .X(Tile_X0Y1_SS4BEG[12]));
 sg13g2_buf_8 output494 (.A(net494),
    .X(Tile_X0Y1_SS4BEG[13]));
 sg13g2_buf_1 output495 (.A(net495),
    .X(Tile_X0Y1_SS4BEG[14]));
 sg13g2_buf_1 output496 (.A(net496),
    .X(Tile_X0Y1_SS4BEG[15]));
 sg13g2_buf_1 output497 (.A(net497),
    .X(Tile_X0Y1_SS4BEG[1]));
 sg13g2_buf_1 output498 (.A(net498),
    .X(Tile_X0Y1_SS4BEG[2]));
 sg13g2_buf_1 output499 (.A(net499),
    .X(Tile_X0Y1_SS4BEG[3]));
 sg13g2_buf_1 output500 (.A(net500),
    .X(Tile_X0Y1_SS4BEG[4]));
 sg13g2_buf_1 output501 (.A(net501),
    .X(Tile_X0Y1_SS4BEG[5]));
 sg13g2_buf_1 output502 (.A(net502),
    .X(Tile_X0Y1_SS4BEG[6]));
 sg13g2_buf_1 output503 (.A(net503),
    .X(Tile_X0Y1_SS4BEG[7]));
 sg13g2_buf_1 output504 (.A(net504),
    .X(Tile_X0Y1_SS4BEG[8]));
 sg13g2_buf_8 output505 (.A(net505),
    .X(Tile_X0Y1_SS4BEG[9]));
 sg13g2_buf_1 output506 (.A(net506),
    .X(Tile_X0Y1_W1BEG[0]));
 sg13g2_buf_1 output507 (.A(net507),
    .X(Tile_X0Y1_W1BEG[1]));
 sg13g2_buf_1 output508 (.A(net508),
    .X(Tile_X0Y1_W1BEG[2]));
 sg13g2_buf_1 output509 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 ),
    .X(Tile_X0Y1_W1BEG[3]));
 sg13g2_buf_1 output510 (.A(net510),
    .X(Tile_X0Y1_W2BEG[0]));
 sg13g2_buf_1 output511 (.A(net511),
    .X(Tile_X0Y1_W2BEG[1]));
 sg13g2_buf_1 output512 (.A(net512),
    .X(Tile_X0Y1_W2BEG[2]));
 sg13g2_buf_1 output513 (.A(net513),
    .X(Tile_X0Y1_W2BEG[3]));
 sg13g2_buf_1 output514 (.A(net514),
    .X(Tile_X0Y1_W2BEG[4]));
 sg13g2_buf_1 output515 (.A(net515),
    .X(Tile_X0Y1_W2BEG[5]));
 sg13g2_buf_1 output516 (.A(net516),
    .X(Tile_X0Y1_W2BEG[6]));
 sg13g2_buf_1 output517 (.A(net517),
    .X(Tile_X0Y1_W2BEG[7]));
 sg13g2_buf_1 output518 (.A(net518),
    .X(Tile_X0Y1_W2BEGb[0]));
 sg13g2_buf_1 output519 (.A(net519),
    .X(Tile_X0Y1_W2BEGb[1]));
 sg13g2_buf_1 output520 (.A(net520),
    .X(Tile_X0Y1_W2BEGb[2]));
 sg13g2_buf_1 output521 (.A(net521),
    .X(Tile_X0Y1_W2BEGb[3]));
 sg13g2_buf_1 output522 (.A(net522),
    .X(Tile_X0Y1_W2BEGb[4]));
 sg13g2_buf_1 output523 (.A(net523),
    .X(Tile_X0Y1_W2BEGb[5]));
 sg13g2_buf_1 output524 (.A(net524),
    .X(Tile_X0Y1_W2BEGb[6]));
 sg13g2_buf_1 output525 (.A(net525),
    .X(Tile_X0Y1_W2BEGb[7]));
 sg13g2_buf_1 output526 (.A(net526),
    .X(Tile_X0Y1_W6BEG[0]));
 sg13g2_buf_1 output527 (.A(net527),
    .X(Tile_X0Y1_W6BEG[10]));
 sg13g2_buf_1 output528 (.A(net528),
    .X(Tile_X0Y1_W6BEG[11]));
 sg13g2_buf_1 output529 (.A(net529),
    .X(Tile_X0Y1_W6BEG[1]));
 sg13g2_buf_1 output530 (.A(net530),
    .X(Tile_X0Y1_W6BEG[2]));
 sg13g2_buf_1 output531 (.A(net531),
    .X(Tile_X0Y1_W6BEG[3]));
 sg13g2_buf_1 output532 (.A(net532),
    .X(Tile_X0Y1_W6BEG[4]));
 sg13g2_buf_1 output533 (.A(net533),
    .X(Tile_X0Y1_W6BEG[5]));
 sg13g2_buf_1 output534 (.A(net534),
    .X(Tile_X0Y1_W6BEG[6]));
 sg13g2_buf_1 output535 (.A(net535),
    .X(Tile_X0Y1_W6BEG[7]));
 sg13g2_buf_1 output536 (.A(net536),
    .X(Tile_X0Y1_W6BEG[8]));
 sg13g2_buf_1 output537 (.A(net537),
    .X(Tile_X0Y1_W6BEG[9]));
 sg13g2_buf_1 output538 (.A(net538),
    .X(Tile_X0Y1_WW4BEG[0]));
 sg13g2_buf_1 output539 (.A(net539),
    .X(Tile_X0Y1_WW4BEG[10]));
 sg13g2_buf_1 output540 (.A(net540),
    .X(Tile_X0Y1_WW4BEG[11]));
 sg13g2_buf_1 output541 (.A(net541),
    .X(Tile_X0Y1_WW4BEG[12]));
 sg13g2_buf_1 output542 (.A(net542),
    .X(Tile_X0Y1_WW4BEG[13]));
 sg13g2_buf_1 output543 (.A(net543),
    .X(Tile_X0Y1_WW4BEG[14]));
 sg13g2_buf_1 output544 (.A(net544),
    .X(Tile_X0Y1_WW4BEG[15]));
 sg13g2_buf_1 output545 (.A(net545),
    .X(Tile_X0Y1_WW4BEG[1]));
 sg13g2_buf_1 output546 (.A(net546),
    .X(Tile_X0Y1_WW4BEG[2]));
 sg13g2_buf_1 output547 (.A(net547),
    .X(Tile_X0Y1_WW4BEG[3]));
 sg13g2_buf_1 output548 (.A(net548),
    .X(Tile_X0Y1_WW4BEG[4]));
 sg13g2_buf_1 output549 (.A(net549),
    .X(Tile_X0Y1_WW4BEG[5]));
 sg13g2_buf_1 output550 (.A(net550),
    .X(Tile_X0Y1_WW4BEG[6]));
 sg13g2_buf_1 output551 (.A(net551),
    .X(Tile_X0Y1_WW4BEG[7]));
 sg13g2_buf_1 output552 (.A(net552),
    .X(Tile_X0Y1_WW4BEG[8]));
 sg13g2_buf_1 output553 (.A(net553),
    .X(Tile_X0Y1_WW4BEG[9]));
 sg13g2_tiehi _5478__554 (.L_HI(net554));
 sg13g2_buf_16 rebuffer2 (.X(net611),
    .A(net667));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(net611),
    .X(net612));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(net611),
    .X(net613));
 sg13g2_dlygate4sd1_1 rebuffer5 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.E2BEG2 ),
    .X(net614));
 sg13g2_buf_8 rebuffer6 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 ),
    .X(net615));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(net634),
    .X(net616));
 sg13g2_buf_2 rebuffer9 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .X(net618));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(net624),
    .X(net619));
 sg13g2_dlygate4sd1_1 rebuffer11 (.A(_0597_),
    .X(net620));
 sg13g2_dlygate4sd1_1 rebuffer12 (.A(_0597_),
    .X(net621));
 sg13g2_buf_8 rebuffer13 (.A(_0597_),
    .X(net622));
 sg13g2_buf_8 rebuffer14 (.A(_1943_),
    .X(net623));
 sg13g2_buf_8 rebuffer15 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 ),
    .X(net624));
 sg13g2_buf_2 rebuffer16 (.A(_0928_),
    .X(net625));
 sg13g2_buf_8 rebuffer24 (.A(_0680_),
    .X(net633));
 sg13g2_dlygate4sd1_1 rebuffer25 (.A(net633),
    .X(net634));
 sg13g2_buf_16 rebuffer26 (.X(net635),
    .A(net698));
 sg13g2_buf_2 rebuffer27 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .X(net636));
 sg13g2_buf_2 rebuffer28 (.A(net636),
    .X(net637));
 sg13g2_buf_2 rebuffer29 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 ),
    .X(net638));
 sg13g2_buf_1 rebuffer30 (.A(net638),
    .X(net639));
 sg13g2_buf_8 rebuffer33 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 ),
    .X(net642));
 sg13g2_dlygate4sd1_1 rebuffer34 (.A(_0595_),
    .X(net643));
 sg13g2_buf_2 rebuffer35 (.A(_1804_),
    .X(net644));
 sg13g2_buf_2 rebuffer36 (.A(_0615_),
    .X(net645));
 sg13g2_dlygate4sd1_1 rebuffer37 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 ),
    .X(net646));
 sg13g2_buf_8 rebuffer38 (.A(net716),
    .X(net647));
 sg13g2_buf_8 rebuffer58 (.A(net728),
    .X(net667));
 sg13g2_dlygate4sd1_1 rebuffer59 (.A(_0565_),
    .X(net668));
 sg13g2_dlygate4sd1_1 rebuffer60 (.A(_0565_),
    .X(net669));
 sg13g2_buf_8 rebuffer72 (.A(_0327_),
    .X(net681));
 sg13g2_dlygate4sd1_1 rebuffer73 (.A(_1433_),
    .X(net682));
 sg13g2_dlygate4sd1_1 rebuffer74 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 ),
    .X(net683));
 sg13g2_dlygate4sd1_1 rebuffer75 (.A(_0565_),
    .X(net684));
 sg13g2_dlygate4sd1_1 rebuffer76 (.A(_1433_),
    .X(net685));
 sg13g2_buf_2 rebuffer77 (.A(_1804_),
    .X(net686));
 sg13g2_buf_8 rebuffer79 (.A(net687),
    .X(net688));
 sg13g2_dlygate4sd1_1 rebuffer80 (.A(_0348_),
    .X(net689));
 sg13g2_dlygate4sd1_1 rebuffer81 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net690));
 sg13g2_dlygate4sd1_1 rebuffer82 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 ),
    .X(net691));
 sg13g2_dlygate4sd1_1 rebuffer83 (.A(_0289_),
    .X(net692));
 sg13g2_dlygate4sd1_1 rebuffer84 (.A(_0289_),
    .X(net693));
 sg13g2_dlygate4sd1_1 rebuffer85 (.A(_0681_),
    .X(net694));
 sg13g2_dlygate4sd1_1 rebuffer86 (.A(_0288_),
    .X(net695));
 sg13g2_dlygate4sd1_1 rebuffer87 (.A(_0288_),
    .X(net696));
 sg13g2_buf_1 rebuffer88 (.A(_1462_),
    .X(net697));
 sg13g2_buf_2 rebuffer89 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 ),
    .X(net698));
 sg13g2_dlygate4sd1_1 rebuffer90 (.A(net1541),
    .X(net699));
 sg13g2_buf_8 rebuffer91 (.A(_1931_),
    .X(net700));
 sg13g2_buf_8 rebuffer92 (.A(_0411_),
    .X(net701));
 sg13g2_dlygate4sd1_1 rebuffer94 (.A(_0417_),
    .X(net703));
 sg13g2_dlygate4sd1_1 rebuffer95 (.A(_1801_),
    .X(net704));
 sg13g2_dlygate4sd1_1 rebuffer96 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .X(net705));
 sg13g2_dlygate4sd1_1 rebuffer97 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .X(net706));
 sg13g2_dlygate4sd1_1 rebuffer98 (.A(_0460_),
    .X(net707));
 sg13g2_dlygate4sd1_1 rebuffer99 (.A(_0417_),
    .X(net708));
 sg13g2_dlygate4sd1_1 rebuffer100 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X ),
    .X(net709));
 sg13g2_dlygate4sd1_1 rebuffer101 (.A(_0323_),
    .X(net710));
 sg13g2_dlygate4sd1_1 rebuffer102 (.A(_2053_),
    .X(net711));
 sg13g2_buf_8 rebuffer103 (.A(_0324_),
    .X(net712));
 sg13g2_buf_2 rebuffer104 (.A(_0323_),
    .X(net713));
 sg13g2_buf_8 rebuffer105 (.A(_0929_),
    .X(net714));
 sg13g2_buf_8 rebuffer106 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 ),
    .X(net715));
 sg13g2_buf_2 rebuffer107 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.E2BEG3 ),
    .X(net716));
 sg13g2_dlygate4sd1_1 rebuffer108 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 ),
    .X(net717));
 sg13g2_dlygate4sd1_1 rebuffer109 (.A(_0416_),
    .X(net718));
 sg13g2_dlygate4sd1_1 rebuffer110 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net719));
 sg13g2_buf_2 rebuffer111 (.A(_0682_),
    .X(net720));
 sg13g2_buf_2 rebuffer112 (.A(\Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 ),
    .X(net721));
 sg13g2_dlygate4sd1_1 rebuffer113 (.A(_0230_),
    .X(net722));
 sg13g2_buf_2 rebuffer114 (.A(net730),
    .X(net723));
 sg13g2_dlygate4sd1_1 rebuffer115 (.A(net723),
    .X(net724));
 sg13g2_dlygate4sd1_1 rebuffer116 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .X(net725));
 sg13g2_buf_2 rebuffer128 (.A(net738),
    .X(net737));
 sg13g2_buf_2 rebuffer129 (.A(net739),
    .X(net738));
 sg13g2_buf_2 rebuffer130 (.A(net740),
    .X(net739));
 sg13g2_buf_2 rebuffer131 (.A(net741),
    .X(net740));
 sg13g2_buf_2 rebuffer132 (.A(net742),
    .X(net741));
 sg13g2_buf_2 rebuffer133 (.A(net743),
    .X(net742));
 sg13g2_buf_2 rebuffer134 (.A(net744),
    .X(net743));
 sg13g2_buf_2 rebuffer135 (.A(\Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0024_),
    .X(net745));
 sg13g2_fill_1 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_26 ();
 sg13g2_fill_2 FILLER_0_95 ();
 sg13g2_fill_1 FILLER_0_97 ();
 sg13g2_fill_2 FILLER_0_119 ();
 sg13g2_fill_1 FILLER_0_164 ();
 sg13g2_fill_1 FILLER_0_182 ();
 sg13g2_fill_1 FILLER_0_220 ();
 sg13g2_fill_2 FILLER_0_258 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_307 ();
 sg13g2_fill_1 FILLER_0_330 ();
 sg13g2_fill_1 FILLER_1_80 ();
 sg13g2_fill_2 FILLER_1_115 ();
 sg13g2_fill_1 FILLER_1_168 ();
 sg13g2_fill_2 FILLER_1_186 ();
 sg13g2_fill_2 FILLER_1_221 ();
 sg13g2_fill_2 FILLER_1_257 ();
 sg13g2_fill_1 FILLER_1_259 ();
 sg13g2_fill_2 FILLER_1_306 ();
 sg13g2_fill_1 FILLER_1_308 ();
 sg13g2_fill_2 FILLER_1_326 ();
 sg13g2_fill_2 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_376 ();
 sg13g2_fill_2 FILLER_2_12 ();
 sg13g2_fill_2 FILLER_2_71 ();
 sg13g2_fill_1 FILLER_2_93 ();
 sg13g2_fill_2 FILLER_2_162 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_fill_1 FILLER_2_213 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_fill_2 FILLER_2_308 ();
 sg13g2_fill_2 FILLER_2_358 ();
 sg13g2_fill_1 FILLER_2_360 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_95 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_3_236 ();
 sg13g2_fill_2 FILLER_3_250 ();
 sg13g2_fill_2 FILLER_3_262 ();
 sg13g2_fill_1 FILLER_3_264 ();
 sg13g2_fill_2 FILLER_3_303 ();
 sg13g2_fill_1 FILLER_3_305 ();
 sg13g2_fill_2 FILLER_3_345 ();
 sg13g2_fill_1 FILLER_3_347 ();
 sg13g2_fill_2 FILLER_4_4 ();
 sg13g2_fill_1 FILLER_4_6 ();
 sg13g2_fill_1 FILLER_4_104 ();
 sg13g2_fill_1 FILLER_4_136 ();
 sg13g2_fill_2 FILLER_4_197 ();
 sg13g2_fill_2 FILLER_4_214 ();
 sg13g2_fill_2 FILLER_4_257 ();
 sg13g2_fill_2 FILLER_4_325 ();
 sg13g2_fill_2 FILLER_4_371 ();
 sg13g2_fill_2 FILLER_5_8 ();
 sg13g2_fill_1 FILLER_5_10 ();
 sg13g2_fill_1 FILLER_5_118 ();
 sg13g2_fill_1 FILLER_5_123 ();
 sg13g2_fill_1 FILLER_5_128 ();
 sg13g2_fill_1 FILLER_5_188 ();
 sg13g2_fill_1 FILLER_5_207 ();
 sg13g2_fill_2 FILLER_5_255 ();
 sg13g2_fill_1 FILLER_5_269 ();
 sg13g2_fill_2 FILLER_5_346 ();
 sg13g2_fill_1 FILLER_5_348 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_fill_1 FILLER_6_45 ();
 sg13g2_fill_2 FILLER_6_76 ();
 sg13g2_fill_1 FILLER_6_122 ();
 sg13g2_fill_1 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_149 ();
 sg13g2_fill_1 FILLER_6_151 ();
 sg13g2_fill_2 FILLER_6_186 ();
 sg13g2_fill_2 FILLER_6_192 ();
 sg13g2_fill_1 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_225 ();
 sg13g2_fill_2 FILLER_6_246 ();
 sg13g2_fill_2 FILLER_6_279 ();
 sg13g2_fill_2 FILLER_6_344 ();
 sg13g2_fill_1 FILLER_6_365 ();
 sg13g2_fill_2 FILLER_6_378 ();
 sg13g2_fill_1 FILLER_6_380 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_31 ();
 sg13g2_fill_2 FILLER_7_48 ();
 sg13g2_fill_2 FILLER_7_90 ();
 sg13g2_fill_1 FILLER_7_189 ();
 sg13g2_fill_1 FILLER_7_310 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_fill_2 FILLER_7_344 ();
 sg13g2_fill_1 FILLER_7_361 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_1 FILLER_7_380 ();
 sg13g2_fill_2 FILLER_8_25 ();
 sg13g2_fill_2 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_75 ();
 sg13g2_fill_2 FILLER_8_114 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_fill_2 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_fill_2 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_375 ();
 sg13g2_fill_2 FILLER_9_4 ();
 sg13g2_fill_2 FILLER_9_44 ();
 sg13g2_fill_1 FILLER_9_46 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_fill_1 FILLER_9_107 ();
 sg13g2_fill_2 FILLER_9_134 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_fill_2 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_343 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_fill_1 FILLER_10_43 ();
 sg13g2_fill_2 FILLER_10_53 ();
 sg13g2_fill_1 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_fill_2 FILLER_10_105 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_213 ();
 sg13g2_fill_1 FILLER_10_231 ();
 sg13g2_fill_1 FILLER_10_303 ();
 sg13g2_fill_2 FILLER_10_325 ();
 sg13g2_fill_2 FILLER_10_354 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_375 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_19 ();
 sg13g2_fill_1 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_43 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_fill_2 FILLER_11_69 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_fill_2 FILLER_11_139 ();
 sg13g2_fill_2 FILLER_11_145 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_222 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_326 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_40 ();
 sg13g2_fill_1 FILLER_12_42 ();
 sg13g2_fill_1 FILLER_12_60 ();
 sg13g2_fill_1 FILLER_12_82 ();
 sg13g2_fill_2 FILLER_12_184 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_1 FILLER_12_338 ();
 sg13g2_fill_2 FILLER_12_360 ();
 sg13g2_fill_2 FILLER_12_383 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_18 ();
 sg13g2_fill_2 FILLER_13_48 ();
 sg13g2_fill_1 FILLER_13_50 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_2 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_244 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_315 ();
 sg13g2_fill_1 FILLER_13_380 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_fill_1 FILLER_14_41 ();
 sg13g2_fill_2 FILLER_14_150 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_fill_1 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_335 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_1 FILLER_15_24 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_fill_2 FILLER_15_104 ();
 sg13g2_fill_2 FILLER_15_127 ();
 sg13g2_fill_2 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_181 ();
 sg13g2_fill_1 FILLER_15_216 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_240 ();
 sg13g2_fill_1 FILLER_15_249 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_383 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_2 FILLER_16_68 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_fill_2 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_108 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_255 ();
 sg13g2_fill_2 FILLER_16_287 ();
 sg13g2_fill_1 FILLER_16_289 ();
 sg13g2_fill_2 FILLER_16_298 ();
 sg13g2_fill_1 FILLER_16_300 ();
 sg13g2_fill_1 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_339 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_1 FILLER_16_384 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_157 ();
 sg13g2_fill_2 FILLER_17_196 ();
 sg13g2_fill_1 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_fill_2 FILLER_17_250 ();
 sg13g2_fill_1 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_270 ();
 sg13g2_fill_1 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_379 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_18 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_1 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_117 ();
 sg13g2_fill_2 FILLER_18_139 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_167 ();
 sg13g2_fill_1 FILLER_18_169 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_297 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_352 ();
 sg13g2_fill_2 FILLER_18_374 ();
 sg13g2_fill_1 FILLER_18_376 ();
 sg13g2_fill_1 FILLER_19_8 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_120 ();
 sg13g2_fill_2 FILLER_19_138 ();
 sg13g2_fill_2 FILLER_19_161 ();
 sg13g2_fill_1 FILLER_19_163 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_205 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_fill_2 FILLER_19_382 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_20_117 ();
 sg13g2_fill_2 FILLER_20_135 ();
 sg13g2_fill_1 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_246 ();
 sg13g2_fill_2 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_320 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_21_64 ();
 sg13g2_fill_1 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_133 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_fill_1 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_179 ();
 sg13g2_fill_1 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_203 ();
 sg13g2_fill_2 FILLER_21_213 ();
 sg13g2_decap_4 FILLER_21_243 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_27 ();
 sg13g2_fill_2 FILLER_22_54 ();
 sg13g2_fill_1 FILLER_22_56 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_decap_8 FILLER_22_225 ();
 sg13g2_fill_2 FILLER_22_232 ();
 sg13g2_fill_2 FILLER_22_339 ();
 sg13g2_fill_2 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_175 ();
 sg13g2_fill_1 FILLER_23_177 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_fill_2 FILLER_23_298 ();
 sg13g2_fill_1 FILLER_24_8 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_1 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_fill_1 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_341 ();
 sg13g2_fill_1 FILLER_24_372 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_1 FILLER_25_90 ();
 sg13g2_fill_2 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_fill_2 FILLER_25_174 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_2 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_26_4 ();
 sg13g2_fill_1 FILLER_26_22 ();
 sg13g2_fill_1 FILLER_26_44 ();
 sg13g2_fill_2 FILLER_26_95 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_fill_2 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_220 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_4 FILLER_26_242 ();
 sg13g2_fill_2 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_fill_2 FILLER_26_383 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_22 ();
 sg13g2_fill_1 FILLER_27_24 ();
 sg13g2_fill_2 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_45 ();
 sg13g2_fill_2 FILLER_27_94 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_171 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_4 FILLER_27_203 ();
 sg13g2_fill_1 FILLER_27_207 ();
 sg13g2_decap_4 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_292 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_fill_1 FILLER_27_384 ();
 sg13g2_fill_2 FILLER_28_25 ();
 sg13g2_fill_1 FILLER_28_27 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_fill_2 FILLER_28_80 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_100 ();
 sg13g2_decap_8 FILLER_28_107 ();
 sg13g2_decap_8 FILLER_28_114 ();
 sg13g2_decap_8 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_128 ();
 sg13g2_fill_2 FILLER_28_133 ();
 sg13g2_fill_1 FILLER_28_135 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_40 ();
 sg13g2_fill_1 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_47 ();
 sg13g2_decap_4 FILLER_29_54 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_79 ();
 sg13g2_decap_4 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_88 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_162 ();
 sg13g2_fill_1 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_181 ();
 sg13g2_fill_2 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_decap_4 FILLER_30_60 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_fill_1 FILLER_30_149 ();
 sg13g2_decap_4 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_230 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_fill_2 FILLER_30_275 ();
 sg13g2_fill_2 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_341 ();
 sg13g2_fill_1 FILLER_30_343 ();
 sg13g2_fill_2 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_20 ();
 sg13g2_fill_2 FILLER_31_31 ();
 sg13g2_fill_1 FILLER_31_33 ();
 sg13g2_fill_1 FILLER_31_51 ();
 sg13g2_decap_4 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_decap_4 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_200 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_1 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_fill_2 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_354 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_6 ();
 sg13g2_fill_2 FILLER_32_19 ();
 sg13g2_fill_1 FILLER_32_26 ();
 sg13g2_fill_2 FILLER_32_36 ();
 sg13g2_fill_1 FILLER_32_38 ();
 sg13g2_fill_1 FILLER_32_53 ();
 sg13g2_decap_4 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_88 ();
 sg13g2_decap_4 FILLER_32_104 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_fill_2 FILLER_32_126 ();
 sg13g2_fill_1 FILLER_32_128 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_162 ();
 sg13g2_decap_8 FILLER_32_174 ();
 sg13g2_decap_8 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_188 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_246 ();
 sg13g2_fill_2 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_1 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_67 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_76 ();
 sg13g2_fill_2 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_130 ();
 sg13g2_decap_8 FILLER_33_148 ();
 sg13g2_decap_4 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_181 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_4 FILLER_33_209 ();
 sg13g2_fill_2 FILLER_33_247 ();
 sg13g2_fill_1 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_289 ();
 sg13g2_fill_2 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_1 FILLER_33_335 ();
 sg13g2_fill_2 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_384 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_38 ();
 sg13g2_fill_2 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_107 ();
 sg13g2_fill_2 FILLER_34_142 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_fill_2 FILLER_34_222 ();
 sg13g2_fill_1 FILLER_34_224 ();
 sg13g2_fill_2 FILLER_34_242 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_2 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_fill_1 FILLER_35_20 ();
 sg13g2_decap_4 FILLER_35_45 ();
 sg13g2_fill_2 FILLER_35_53 ();
 sg13g2_fill_2 FILLER_35_59 ();
 sg13g2_fill_2 FILLER_35_78 ();
 sg13g2_fill_1 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_101 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_136 ();
 sg13g2_fill_1 FILLER_35_138 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_11 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_decap_4 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_236 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_318 ();
 sg13g2_fill_1 FILLER_36_376 ();
 sg13g2_fill_1 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_18 ();
 sg13g2_fill_1 FILLER_37_20 ();
 sg13g2_decap_8 FILLER_37_24 ();
 sg13g2_decap_4 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_159 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_4 FILLER_37_224 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_fill_2 FILLER_37_359 ();
 sg13g2_fill_1 FILLER_37_361 ();
 sg13g2_fill_2 FILLER_37_383 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_24 ();
 sg13g2_decap_4 FILLER_38_33 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_2 FILLER_38_251 ();
 sg13g2_fill_1 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_fill_2 FILLER_38_357 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_2 ();
 sg13g2_fill_2 FILLER_39_61 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_fill_2 FILLER_39_85 ();
 sg13g2_fill_2 FILLER_39_129 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_fill_1 FILLER_39_166 ();
 sg13g2_fill_2 FILLER_39_184 ();
 sg13g2_decap_4 FILLER_39_199 ();
 sg13g2_decap_8 FILLER_39_220 ();
 sg13g2_fill_1 FILLER_39_246 ();
 sg13g2_fill_2 FILLER_39_298 ();
 sg13g2_fill_1 FILLER_39_300 ();
 sg13g2_fill_1 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_fill_1 FILLER_39_365 ();
 sg13g2_fill_2 FILLER_39_375 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_fill_2 FILLER_39_383 ();
 sg13g2_fill_2 FILLER_40_17 ();
 sg13g2_fill_1 FILLER_40_19 ();
 sg13g2_fill_1 FILLER_40_41 ();
 sg13g2_decap_8 FILLER_40_75 ();
 sg13g2_decap_8 FILLER_40_82 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_186 ();
 sg13g2_fill_1 FILLER_40_188 ();
 sg13g2_fill_1 FILLER_40_233 ();
 sg13g2_fill_1 FILLER_40_291 ();
 sg13g2_fill_2 FILLER_40_359 ();
 sg13g2_fill_1 FILLER_40_361 ();
 sg13g2_fill_2 FILLER_40_375 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_4 ();
 sg13g2_fill_2 FILLER_41_45 ();
 sg13g2_fill_1 FILLER_41_47 ();
 sg13g2_fill_1 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_74 ();
 sg13g2_fill_2 FILLER_41_81 ();
 sg13g2_fill_1 FILLER_41_87 ();
 sg13g2_fill_2 FILLER_41_113 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_fill_2 FILLER_41_177 ();
 sg13g2_fill_2 FILLER_41_203 ();
 sg13g2_fill_2 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_fill_2 FILLER_41_224 ();
 sg13g2_fill_1 FILLER_41_226 ();
 sg13g2_fill_2 FILLER_41_269 ();
 sg13g2_fill_1 FILLER_41_304 ();
 sg13g2_fill_2 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_319 ();
 sg13g2_fill_2 FILLER_41_357 ();
 sg13g2_fill_2 FILLER_42_17 ();
 sg13g2_fill_1 FILLER_42_19 ();
 sg13g2_fill_2 FILLER_42_41 ();
 sg13g2_fill_2 FILLER_42_90 ();
 sg13g2_decap_8 FILLER_42_104 ();
 sg13g2_decap_8 FILLER_42_111 ();
 sg13g2_fill_2 FILLER_42_118 ();
 sg13g2_fill_1 FILLER_42_216 ();
 sg13g2_decap_8 FILLER_42_234 ();
 sg13g2_decap_8 FILLER_42_241 ();
 sg13g2_fill_2 FILLER_42_248 ();
 sg13g2_fill_1 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_fill_1 FILLER_43_117 ();
 sg13g2_fill_2 FILLER_43_139 ();
 sg13g2_fill_1 FILLER_43_141 ();
 sg13g2_decap_8 FILLER_43_157 ();
 sg13g2_decap_8 FILLER_43_164 ();
 sg13g2_decap_8 FILLER_43_171 ();
 sg13g2_decap_4 FILLER_43_178 ();
 sg13g2_fill_2 FILLER_43_216 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_fill_2 FILLER_43_274 ();
 sg13g2_fill_2 FILLER_43_291 ();
 sg13g2_fill_2 FILLER_43_328 ();
 sg13g2_fill_1 FILLER_43_363 ();
 sg13g2_fill_1 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_33 ();
 sg13g2_fill_1 FILLER_44_35 ();
 sg13g2_fill_2 FILLER_44_44 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_fill_2 FILLER_44_64 ();
 sg13g2_fill_1 FILLER_44_73 ();
 sg13g2_fill_1 FILLER_44_79 ();
 sg13g2_fill_2 FILLER_44_111 ();
 sg13g2_decap_4 FILLER_44_121 ();
 sg13g2_fill_1 FILLER_44_141 ();
 sg13g2_decap_4 FILLER_44_151 ();
 sg13g2_fill_1 FILLER_44_165 ();
 sg13g2_fill_1 FILLER_44_218 ();
 sg13g2_decap_8 FILLER_44_223 ();
 sg13g2_fill_2 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_232 ();
 sg13g2_decap_4 FILLER_44_250 ();
 sg13g2_fill_1 FILLER_44_254 ();
 sg13g2_fill_2 FILLER_44_294 ();
 sg13g2_fill_2 FILLER_44_335 ();
 sg13g2_fill_1 FILLER_44_337 ();
 sg13g2_fill_1 FILLER_44_384 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_27 ();
 sg13g2_decap_4 FILLER_45_56 ();
 sg13g2_fill_1 FILLER_45_60 ();
 sg13g2_fill_2 FILLER_45_96 ();
 sg13g2_fill_1 FILLER_45_107 ();
 sg13g2_decap_8 FILLER_45_129 ();
 sg13g2_fill_2 FILLER_45_136 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_fill_2 FILLER_45_180 ();
 sg13g2_fill_2 FILLER_45_206 ();
 sg13g2_fill_1 FILLER_45_208 ();
 sg13g2_decap_4 FILLER_45_213 ();
 sg13g2_decap_4 FILLER_45_260 ();
 sg13g2_fill_1 FILLER_45_264 ();
 sg13g2_fill_2 FILLER_45_299 ();
 sg13g2_fill_1 FILLER_45_313 ();
 sg13g2_fill_1 FILLER_45_362 ();
 sg13g2_fill_1 FILLER_45_367 ();
 sg13g2_fill_2 FILLER_45_383 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_36 ();
 sg13g2_fill_1 FILLER_46_38 ();
 sg13g2_fill_2 FILLER_46_90 ();
 sg13g2_fill_1 FILLER_46_92 ();
 sg13g2_fill_1 FILLER_46_119 ();
 sg13g2_fill_1 FILLER_46_130 ();
 sg13g2_fill_2 FILLER_46_171 ();
 sg13g2_fill_2 FILLER_46_179 ();
 sg13g2_fill_2 FILLER_46_187 ();
 sg13g2_decap_4 FILLER_46_194 ();
 sg13g2_fill_2 FILLER_46_249 ();
 sg13g2_fill_1 FILLER_46_264 ();
 sg13g2_fill_1 FILLER_46_269 ();
 sg13g2_fill_2 FILLER_46_329 ();
 sg13g2_fill_1 FILLER_46_331 ();
 sg13g2_fill_2 FILLER_46_339 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_18 ();
 sg13g2_fill_2 FILLER_47_52 ();
 sg13g2_fill_1 FILLER_47_54 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_fill_1 FILLER_47_116 ();
 sg13g2_fill_2 FILLER_47_152 ();
 sg13g2_fill_1 FILLER_47_159 ();
 sg13g2_decap_4 FILLER_47_164 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_fill_2 FILLER_47_195 ();
 sg13g2_fill_2 FILLER_47_238 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_1 FILLER_47_288 ();
 sg13g2_fill_1 FILLER_47_317 ();
 sg13g2_fill_2 FILLER_47_344 ();
 sg13g2_fill_2 FILLER_47_365 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_379 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_23 ();
 sg13g2_fill_1 FILLER_48_25 ();
 sg13g2_fill_2 FILLER_48_31 ();
 sg13g2_fill_2 FILLER_48_105 ();
 sg13g2_fill_2 FILLER_48_127 ();
 sg13g2_decap_8 FILLER_48_146 ();
 sg13g2_decap_8 FILLER_48_153 ();
 sg13g2_decap_8 FILLER_48_160 ();
 sg13g2_decap_8 FILLER_48_198 ();
 sg13g2_decap_4 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_209 ();
 sg13g2_fill_2 FILLER_48_215 ();
 sg13g2_fill_1 FILLER_48_217 ();
 sg13g2_fill_2 FILLER_48_235 ();
 sg13g2_fill_1 FILLER_48_237 ();
 sg13g2_decap_4 FILLER_48_265 ();
 sg13g2_fill_1 FILLER_48_269 ();
 sg13g2_fill_2 FILLER_48_336 ();
 sg13g2_fill_1 FILLER_48_362 ();
 sg13g2_fill_1 FILLER_48_384 ();
 sg13g2_fill_2 FILLER_49_68 ();
 sg13g2_fill_1 FILLER_49_70 ();
 sg13g2_fill_2 FILLER_49_75 ();
 sg13g2_fill_2 FILLER_49_86 ();
 sg13g2_fill_1 FILLER_49_88 ();
 sg13g2_fill_1 FILLER_49_138 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_decap_4 FILLER_49_192 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_fill_2 FILLER_49_223 ();
 sg13g2_fill_1 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_fill_2 FILLER_49_358 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_172 ();
 sg13g2_decap_8 FILLER_50_179 ();
 sg13g2_fill_1 FILLER_50_203 ();
 sg13g2_fill_2 FILLER_50_250 ();
 sg13g2_decap_8 FILLER_50_269 ();
 sg13g2_decap_8 FILLER_50_276 ();
 sg13g2_fill_1 FILLER_50_283 ();
 sg13g2_fill_2 FILLER_50_310 ();
 sg13g2_fill_2 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_349 ();
 sg13g2_fill_1 FILLER_50_366 ();
 sg13g2_fill_2 FILLER_50_383 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_72 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_fill_2 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_174 ();
 sg13g2_decap_4 FILLER_51_181 ();
 sg13g2_fill_2 FILLER_51_185 ();
 sg13g2_fill_2 FILLER_51_212 ();
 sg13g2_decap_4 FILLER_51_219 ();
 sg13g2_fill_2 FILLER_51_223 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_fill_2 FILLER_51_254 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_2 FILLER_51_314 ();
 sg13g2_fill_2 FILLER_51_336 ();
 sg13g2_fill_1 FILLER_51_366 ();
 sg13g2_fill_2 FILLER_51_375 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_2 ();
 sg13g2_decap_8 FILLER_52_20 ();
 sg13g2_fill_1 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_68 ();
 sg13g2_fill_2 FILLER_52_74 ();
 sg13g2_fill_1 FILLER_52_76 ();
 sg13g2_fill_2 FILLER_52_96 ();
 sg13g2_fill_1 FILLER_52_98 ();
 sg13g2_fill_1 FILLER_52_116 ();
 sg13g2_decap_4 FILLER_52_194 ();
 sg13g2_fill_1 FILLER_52_206 ();
 sg13g2_fill_1 FILLER_52_259 ();
 sg13g2_fill_2 FILLER_52_305 ();
 sg13g2_fill_1 FILLER_52_307 ();
 sg13g2_fill_2 FILLER_52_322 ();
 sg13g2_fill_1 FILLER_52_324 ();
 sg13g2_fill_1 FILLER_52_370 ();
 sg13g2_fill_1 FILLER_52_384 ();
 sg13g2_decap_4 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_4 ();
 sg13g2_decap_4 FILLER_53_22 ();
 sg13g2_fill_2 FILLER_53_80 ();
 sg13g2_decap_8 FILLER_53_92 ();
 sg13g2_decap_8 FILLER_53_99 ();
 sg13g2_decap_8 FILLER_53_106 ();
 sg13g2_fill_2 FILLER_53_120 ();
 sg13g2_fill_1 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_221 ();
 sg13g2_decap_8 FILLER_53_228 ();
 sg13g2_fill_1 FILLER_53_235 ();
 sg13g2_fill_2 FILLER_53_364 ();
 sg13g2_fill_1 FILLER_53_366 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_29 ();
 sg13g2_decap_4 FILLER_54_36 ();
 sg13g2_fill_1 FILLER_54_40 ();
 sg13g2_fill_2 FILLER_54_86 ();
 sg13g2_fill_1 FILLER_54_88 ();
 sg13g2_decap_8 FILLER_54_110 ();
 sg13g2_fill_2 FILLER_54_117 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_180 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_238 ();
 sg13g2_fill_1 FILLER_54_240 ();
 sg13g2_decap_8 FILLER_54_255 ();
 sg13g2_fill_2 FILLER_54_262 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_4 FILLER_54_287 ();
 sg13g2_fill_1 FILLER_54_299 ();
 sg13g2_fill_1 FILLER_54_308 ();
 sg13g2_fill_2 FILLER_54_354 ();
 sg13g2_fill_1 FILLER_54_356 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_40 ();
 sg13g2_fill_1 FILLER_55_44 ();
 sg13g2_decap_8 FILLER_55_132 ();
 sg13g2_fill_2 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_175 ();
 sg13g2_fill_2 FILLER_55_191 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_328 ();
 sg13g2_fill_1 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_19 ();
 sg13g2_decap_8 FILLER_56_34 ();
 sg13g2_decap_4 FILLER_56_41 ();
 sg13g2_fill_2 FILLER_56_45 ();
 sg13g2_fill_2 FILLER_56_97 ();
 sg13g2_fill_2 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_129 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_146 ();
 sg13g2_fill_2 FILLER_56_176 ();
 sg13g2_decap_8 FILLER_56_202 ();
 sg13g2_fill_2 FILLER_56_209 ();
 sg13g2_fill_1 FILLER_56_211 ();
 sg13g2_fill_2 FILLER_56_222 ();
 sg13g2_fill_1 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_242 ();
 sg13g2_fill_2 FILLER_56_310 ();
 sg13g2_fill_1 FILLER_56_320 ();
 sg13g2_fill_1 FILLER_56_337 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_fill_2 FILLER_56_382 ();
 sg13g2_fill_1 FILLER_56_384 ();
 sg13g2_fill_2 FILLER_57_48 ();
 sg13g2_fill_1 FILLER_57_50 ();
 sg13g2_fill_1 FILLER_57_103 ();
 sg13g2_fill_1 FILLER_57_109 ();
 sg13g2_decap_4 FILLER_57_161 ();
 sg13g2_fill_2 FILLER_57_168 ();
 sg13g2_fill_1 FILLER_57_170 ();
 sg13g2_fill_1 FILLER_57_196 ();
 sg13g2_fill_2 FILLER_57_208 ();
 sg13g2_fill_1 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_283 ();
 sg13g2_decap_4 FILLER_57_290 ();
 sg13g2_fill_1 FILLER_57_294 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_1 FILLER_57_344 ();
 sg13g2_fill_2 FILLER_57_369 ();
 sg13g2_fill_1 FILLER_57_371 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_4 ();
 sg13g2_fill_1 FILLER_58_31 ();
 sg13g2_fill_2 FILLER_58_44 ();
 sg13g2_fill_2 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_70 ();
 sg13g2_fill_2 FILLER_58_77 ();
 sg13g2_fill_2 FILLER_58_113 ();
 sg13g2_fill_1 FILLER_58_131 ();
 sg13g2_decap_4 FILLER_58_158 ();
 sg13g2_fill_2 FILLER_58_162 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_fill_2 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_250 ();
 sg13g2_decap_8 FILLER_58_276 ();
 sg13g2_fill_1 FILLER_58_352 ();
 sg13g2_fill_1 FILLER_58_366 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_decap_4 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_67 ();
 sg13g2_decap_8 FILLER_59_79 ();
 sg13g2_decap_4 FILLER_59_86 ();
 sg13g2_decap_4 FILLER_59_94 ();
 sg13g2_fill_1 FILLER_59_98 ();
 sg13g2_fill_2 FILLER_59_124 ();
 sg13g2_decap_8 FILLER_59_136 ();
 sg13g2_decap_8 FILLER_59_143 ();
 sg13g2_fill_1 FILLER_59_150 ();
 sg13g2_fill_2 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_156 ();
 sg13g2_decap_8 FILLER_59_181 ();
 sg13g2_decap_4 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_192 ();
 sg13g2_fill_2 FILLER_59_238 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_fill_2 FILLER_59_290 ();
 sg13g2_fill_1 FILLER_59_292 ();
 sg13g2_fill_1 FILLER_59_305 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_2 ();
 sg13g2_fill_1 FILLER_60_45 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_94 ();
 sg13g2_decap_8 FILLER_60_101 ();
 sg13g2_decap_8 FILLER_60_108 ();
 sg13g2_decap_4 FILLER_60_115 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_fill_1 FILLER_60_151 ();
 sg13g2_fill_2 FILLER_60_169 ();
 sg13g2_fill_2 FILLER_60_198 ();
 sg13g2_fill_1 FILLER_60_200 ();
 sg13g2_fill_2 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_384 ();
 sg13g2_decap_4 FILLER_61_17 ();
 sg13g2_fill_2 FILLER_61_21 ();
 sg13g2_fill_2 FILLER_61_26 ();
 sg13g2_decap_8 FILLER_61_45 ();
 sg13g2_decap_8 FILLER_61_52 ();
 sg13g2_fill_2 FILLER_61_59 ();
 sg13g2_fill_1 FILLER_61_61 ();
 sg13g2_decap_4 FILLER_61_100 ();
 sg13g2_fill_1 FILLER_61_104 ();
 sg13g2_decap_4 FILLER_61_109 ();
 sg13g2_decap_4 FILLER_61_172 ();
 sg13g2_fill_1 FILLER_61_180 ();
 sg13g2_fill_2 FILLER_61_202 ();
 sg13g2_fill_1 FILLER_61_204 ();
 sg13g2_decap_4 FILLER_61_211 ();
 sg13g2_fill_1 FILLER_61_215 ();
 sg13g2_fill_2 FILLER_61_237 ();
 sg13g2_fill_1 FILLER_61_264 ();
 sg13g2_decap_4 FILLER_61_284 ();
 sg13g2_fill_1 FILLER_61_293 ();
 sg13g2_fill_2 FILLER_61_312 ();
 sg13g2_fill_1 FILLER_61_314 ();
 sg13g2_fill_1 FILLER_61_327 ();
 sg13g2_fill_1 FILLER_61_333 ();
 sg13g2_fill_1 FILLER_61_339 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_53 ();
 sg13g2_decap_4 FILLER_62_64 ();
 sg13g2_fill_1 FILLER_62_85 ();
 sg13g2_decap_4 FILLER_62_147 ();
 sg13g2_fill_1 FILLER_62_151 ();
 sg13g2_decap_8 FILLER_62_156 ();
 sg13g2_fill_2 FILLER_62_189 ();
 sg13g2_decap_4 FILLER_62_195 ();
 sg13g2_decap_8 FILLER_62_207 ();
 sg13g2_decap_4 FILLER_62_214 ();
 sg13g2_decap_8 FILLER_62_222 ();
 sg13g2_decap_4 FILLER_62_229 ();
 sg13g2_fill_2 FILLER_62_233 ();
 sg13g2_decap_4 FILLER_62_239 ();
 sg13g2_fill_2 FILLER_62_247 ();
 sg13g2_fill_2 FILLER_62_269 ();
 sg13g2_decap_4 FILLER_62_274 ();
 sg13g2_fill_1 FILLER_62_278 ();
 sg13g2_fill_2 FILLER_62_305 ();
 sg13g2_fill_1 FILLER_62_307 ();
 sg13g2_fill_1 FILLER_62_315 ();
 sg13g2_fill_1 FILLER_62_339 ();
 sg13g2_fill_2 FILLER_62_356 ();
 sg13g2_fill_1 FILLER_62_358 ();
 sg13g2_fill_2 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_2 ();
 sg13g2_fill_1 FILLER_63_24 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_fill_2 FILLER_63_86 ();
 sg13g2_fill_1 FILLER_63_88 ();
 sg13g2_fill_1 FILLER_63_127 ();
 sg13g2_fill_2 FILLER_63_132 ();
 sg13g2_fill_1 FILLER_63_134 ();
 sg13g2_decap_4 FILLER_63_139 ();
 sg13g2_decap_4 FILLER_63_146 ();
 sg13g2_fill_2 FILLER_63_150 ();
 sg13g2_decap_4 FILLER_63_187 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_fill_2 FILLER_63_196 ();
 sg13g2_fill_1 FILLER_63_198 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_4 FILLER_63_238 ();
 sg13g2_fill_2 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_259 ();
 sg13g2_fill_1 FILLER_63_289 ();
 sg13g2_fill_2 FILLER_63_294 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_fill_2 FILLER_63_352 ();
 sg13g2_fill_1 FILLER_63_354 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_374 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_1 FILLER_64_24 ();
 sg13g2_fill_1 FILLER_64_38 ();
 sg13g2_fill_2 FILLER_64_48 ();
 sg13g2_decap_4 FILLER_64_127 ();
 sg13g2_decap_8 FILLER_64_148 ();
 sg13g2_fill_1 FILLER_64_242 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_2 FILLER_64_330 ();
 sg13g2_fill_1 FILLER_64_332 ();
 sg13g2_decap_4 FILLER_64_355 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_36 ();
 sg13g2_fill_1 FILLER_65_52 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_decap_8 FILLER_65_81 ();
 sg13g2_decap_8 FILLER_65_88 ();
 sg13g2_decap_8 FILLER_65_95 ();
 sg13g2_decap_8 FILLER_65_102 ();
 sg13g2_fill_2 FILLER_65_109 ();
 sg13g2_fill_2 FILLER_65_135 ();
 sg13g2_decap_8 FILLER_65_162 ();
 sg13g2_decap_8 FILLER_65_169 ();
 sg13g2_decap_8 FILLER_65_176 ();
 sg13g2_decap_8 FILLER_65_183 ();
 sg13g2_fill_2 FILLER_65_190 ();
 sg13g2_fill_2 FILLER_65_264 ();
 sg13g2_fill_1 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_306 ();
 sg13g2_fill_2 FILLER_65_338 ();
 sg13g2_fill_2 FILLER_65_355 ();
 sg13g2_fill_1 FILLER_65_357 ();
 sg13g2_fill_1 FILLER_65_371 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_19 ();
 sg13g2_fill_2 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_51 ();
 sg13g2_fill_2 FILLER_66_60 ();
 sg13g2_fill_1 FILLER_66_62 ();
 sg13g2_decap_4 FILLER_66_80 ();
 sg13g2_fill_2 FILLER_66_111 ();
 sg13g2_fill_1 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_159 ();
 sg13g2_fill_1 FILLER_66_166 ();
 sg13g2_fill_2 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_fill_1 FILLER_66_192 ();
 sg13g2_fill_2 FILLER_66_210 ();
 sg13g2_fill_1 FILLER_66_216 ();
 sg13g2_fill_1 FILLER_66_221 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_fill_2 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_329 ();
 sg13g2_fill_1 FILLER_66_371 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_19 ();
 sg13g2_fill_1 FILLER_67_21 ();
 sg13g2_fill_1 FILLER_67_60 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_fill_2 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_121 ();
 sg13g2_fill_2 FILLER_67_148 ();
 sg13g2_fill_1 FILLER_67_150 ();
 sg13g2_decap_4 FILLER_67_168 ();
 sg13g2_fill_1 FILLER_67_189 ();
 sg13g2_fill_2 FILLER_67_194 ();
 sg13g2_fill_1 FILLER_67_241 ();
 sg13g2_fill_2 FILLER_67_293 ();
 sg13g2_fill_2 FILLER_67_317 ();
 sg13g2_fill_1 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_328 ();
 sg13g2_fill_1 FILLER_67_339 ();
 sg13g2_fill_2 FILLER_67_351 ();
 sg13g2_fill_2 FILLER_67_383 ();
 sg13g2_decap_4 FILLER_68_50 ();
 sg13g2_fill_2 FILLER_68_95 ();
 sg13g2_fill_2 FILLER_68_102 ();
 sg13g2_fill_1 FILLER_68_104 ();
 sg13g2_fill_2 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_131 ();
 sg13g2_fill_2 FILLER_68_158 ();
 sg13g2_fill_1 FILLER_68_160 ();
 sg13g2_fill_1 FILLER_68_192 ();
 sg13g2_decap_4 FILLER_68_214 ();
 sg13g2_fill_1 FILLER_68_267 ();
 sg13g2_fill_2 FILLER_68_318 ();
 sg13g2_fill_1 FILLER_68_320 ();
 sg13g2_fill_1 FILLER_68_337 ();
 sg13g2_fill_2 FILLER_68_362 ();
 sg13g2_fill_1 FILLER_68_364 ();
 sg13g2_fill_2 FILLER_68_372 ();
 sg13g2_fill_2 FILLER_68_382 ();
 sg13g2_fill_1 FILLER_68_384 ();
 sg13g2_fill_2 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_2 ();
 sg13g2_decap_8 FILLER_69_66 ();
 sg13g2_decap_8 FILLER_69_73 ();
 sg13g2_decap_8 FILLER_69_80 ();
 sg13g2_decap_4 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_91 ();
 sg13g2_fill_1 FILLER_69_147 ();
 sg13g2_fill_2 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_224 ();
 sg13g2_fill_2 FILLER_69_230 ();
 sg13g2_fill_1 FILLER_69_269 ();
 sg13g2_fill_2 FILLER_69_296 ();
 sg13g2_fill_2 FILLER_69_319 ();
 sg13g2_fill_1 FILLER_69_329 ();
 sg13g2_fill_2 FILLER_69_343 ();
 sg13g2_fill_1 FILLER_69_345 ();
 sg13g2_fill_2 FILLER_69_366 ();
 sg13g2_fill_1 FILLER_69_368 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_18 ();
 sg13g2_fill_2 FILLER_70_24 ();
 sg13g2_fill_1 FILLER_70_34 ();
 sg13g2_fill_2 FILLER_70_58 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_fill_2 FILLER_70_78 ();
 sg13g2_fill_1 FILLER_70_80 ();
 sg13g2_decap_4 FILLER_70_102 ();
 sg13g2_decap_8 FILLER_70_127 ();
 sg13g2_fill_1 FILLER_70_134 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_197 ();
 sg13g2_decap_8 FILLER_70_204 ();
 sg13g2_decap_8 FILLER_70_211 ();
 sg13g2_decap_8 FILLER_70_218 ();
 sg13g2_fill_2 FILLER_70_225 ();
 sg13g2_fill_1 FILLER_70_227 ();
 sg13g2_fill_1 FILLER_70_295 ();
 sg13g2_fill_1 FILLER_70_309 ();
 sg13g2_fill_2 FILLER_70_327 ();
 sg13g2_fill_1 FILLER_70_384 ();
 sg13g2_fill_1 FILLER_71_17 ();
 sg13g2_fill_2 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_39 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_131 ();
 sg13g2_fill_1 FILLER_71_165 ();
 sg13g2_fill_1 FILLER_71_174 ();
 sg13g2_decap_8 FILLER_71_213 ();
 sg13g2_decap_4 FILLER_71_220 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_fill_1 FILLER_71_243 ();
 sg13g2_fill_2 FILLER_71_296 ();
 sg13g2_fill_1 FILLER_71_298 ();
 sg13g2_fill_2 FILLER_71_326 ();
 sg13g2_fill_1 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_369 ();
 sg13g2_fill_1 FILLER_71_378 ();
 sg13g2_fill_1 FILLER_71_384 ();
 sg13g2_fill_1 FILLER_72_34 ();
 sg13g2_decap_4 FILLER_72_61 ();
 sg13g2_fill_2 FILLER_72_82 ();
 sg13g2_fill_1 FILLER_72_84 ();
 sg13g2_fill_1 FILLER_72_139 ();
 sg13g2_decap_4 FILLER_72_161 ();
 sg13g2_decap_4 FILLER_72_186 ();
 sg13g2_fill_1 FILLER_72_190 ();
 sg13g2_fill_2 FILLER_72_237 ();
 sg13g2_fill_1 FILLER_72_239 ();
 sg13g2_fill_2 FILLER_72_288 ();
 sg13g2_fill_2 FILLER_72_295 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_fill_1 FILLER_72_318 ();
 sg13g2_fill_2 FILLER_72_331 ();
 sg13g2_fill_2 FILLER_72_354 ();
 sg13g2_decap_4 FILLER_73_55 ();
 sg13g2_fill_1 FILLER_73_59 ();
 sg13g2_fill_2 FILLER_73_77 ();
 sg13g2_fill_2 FILLER_73_88 ();
 sg13g2_fill_1 FILLER_73_90 ();
 sg13g2_fill_2 FILLER_73_97 ();
 sg13g2_decap_8 FILLER_73_116 ();
 sg13g2_fill_2 FILLER_73_123 ();
 sg13g2_fill_1 FILLER_73_125 ();
 sg13g2_fill_2 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_215 ();
 sg13g2_decap_8 FILLER_73_222 ();
 sg13g2_decap_4 FILLER_73_229 ();
 sg13g2_fill_1 FILLER_73_233 ();
 sg13g2_fill_2 FILLER_73_282 ();
 sg13g2_fill_2 FILLER_73_338 ();
 sg13g2_fill_1 FILLER_73_340 ();
 sg13g2_fill_2 FILLER_73_382 ();
 sg13g2_fill_1 FILLER_73_384 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_decap_4 FILLER_74_54 ();
 sg13g2_fill_2 FILLER_74_100 ();
 sg13g2_fill_1 FILLER_74_102 ();
 sg13g2_fill_2 FILLER_74_106 ();
 sg13g2_fill_1 FILLER_74_108 ();
 sg13g2_fill_2 FILLER_74_143 ();
 sg13g2_fill_1 FILLER_74_162 ();
 sg13g2_fill_2 FILLER_74_171 ();
 sg13g2_fill_1 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_fill_2 FILLER_74_326 ();
 sg13g2_fill_2 FILLER_74_340 ();
 sg13g2_fill_2 FILLER_74_383 ();
 sg13g2_fill_2 FILLER_75_17 ();
 sg13g2_fill_2 FILLER_75_59 ();
 sg13g2_fill_2 FILLER_75_104 ();
 sg13g2_fill_2 FILLER_75_123 ();
 sg13g2_fill_1 FILLER_75_125 ();
 sg13g2_fill_2 FILLER_75_145 ();
 sg13g2_fill_2 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_166 ();
 sg13g2_fill_1 FILLER_75_195 ();
 sg13g2_fill_2 FILLER_75_234 ();
 sg13g2_fill_2 FILLER_75_348 ();
 sg13g2_fill_1 FILLER_75_350 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_2 ();
 sg13g2_fill_2 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_83 ();
 sg13g2_fill_2 FILLER_76_112 ();
 sg13g2_fill_2 FILLER_76_159 ();
 sg13g2_fill_1 FILLER_76_161 ();
 sg13g2_fill_2 FILLER_76_179 ();
 sg13g2_decap_8 FILLER_76_198 ();
 sg13g2_decap_8 FILLER_76_205 ();
 sg13g2_decap_4 FILLER_76_212 ();
 sg13g2_fill_2 FILLER_76_272 ();
 sg13g2_fill_2 FILLER_76_311 ();
 sg13g2_fill_1 FILLER_76_313 ();
 sg13g2_fill_2 FILLER_76_327 ();
 sg13g2_fill_2 FILLER_76_350 ();
 sg13g2_fill_1 FILLER_76_364 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_2 ();
 sg13g2_fill_1 FILLER_77_41 ();
 sg13g2_fill_2 FILLER_77_52 ();
 sg13g2_fill_2 FILLER_77_123 ();
 sg13g2_fill_2 FILLER_77_150 ();
 sg13g2_fill_2 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_222 ();
 sg13g2_fill_1 FILLER_77_229 ();
 sg13g2_fill_1 FILLER_77_272 ();
 sg13g2_fill_1 FILLER_77_289 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_2 FILLER_77_351 ();
 sg13g2_fill_2 FILLER_77_361 ();
 sg13g2_fill_1 FILLER_77_380 ();
 sg13g2_fill_2 FILLER_78_42 ();
 sg13g2_fill_2 FILLER_78_63 ();
 sg13g2_fill_1 FILLER_78_65 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_fill_1 FILLER_78_77 ();
 sg13g2_decap_4 FILLER_78_81 ();
 sg13g2_fill_1 FILLER_78_85 ();
 sg13g2_decap_4 FILLER_78_122 ();
 sg13g2_fill_2 FILLER_78_139 ();
 sg13g2_fill_1 FILLER_78_141 ();
 sg13g2_fill_2 FILLER_78_159 ();
 sg13g2_fill_1 FILLER_78_182 ();
 sg13g2_decap_4 FILLER_78_225 ();
 sg13g2_fill_1 FILLER_78_229 ();
 sg13g2_fill_1 FILLER_78_240 ();
 sg13g2_fill_1 FILLER_78_261 ();
 sg13g2_fill_2 FILLER_78_309 ();
 sg13g2_fill_1 FILLER_78_329 ();
 sg13g2_fill_1 FILLER_78_358 ();
 sg13g2_fill_2 FILLER_79_25 ();
 sg13g2_fill_1 FILLER_79_27 ();
 sg13g2_fill_2 FILLER_79_102 ();
 sg13g2_fill_1 FILLER_79_104 ();
 sg13g2_decap_4 FILLER_79_126 ();
 sg13g2_fill_2 FILLER_79_202 ();
 sg13g2_fill_1 FILLER_79_204 ();
 sg13g2_decap_8 FILLER_79_226 ();
 sg13g2_fill_2 FILLER_79_271 ();
 sg13g2_fill_1 FILLER_79_347 ();
 sg13g2_fill_2 FILLER_79_383 ();
 sg13g2_fill_1 FILLER_80_12 ();
 sg13g2_fill_1 FILLER_80_57 ();
 sg13g2_decap_8 FILLER_80_75 ();
 sg13g2_decap_4 FILLER_80_82 ();
 sg13g2_fill_2 FILLER_80_86 ();
 sg13g2_fill_2 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_158 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_fill_2 FILLER_80_254 ();
 sg13g2_fill_2 FILLER_81_0 ();
 sg13g2_fill_2 FILLER_81_43 ();
 sg13g2_fill_1 FILLER_81_45 ();
 sg13g2_fill_2 FILLER_81_63 ();
 sg13g2_fill_1 FILLER_81_65 ();
 sg13g2_decap_4 FILLER_81_87 ();
 sg13g2_fill_2 FILLER_81_91 ();
 sg13g2_decap_4 FILLER_81_114 ();
 sg13g2_fill_2 FILLER_81_118 ();
 sg13g2_decap_4 FILLER_81_124 ();
 sg13g2_fill_1 FILLER_81_128 ();
 sg13g2_fill_1 FILLER_81_170 ();
 sg13g2_decap_4 FILLER_81_203 ();
 sg13g2_fill_2 FILLER_81_207 ();
 sg13g2_fill_1 FILLER_81_239 ();
 sg13g2_fill_2 FILLER_81_244 ();
 sg13g2_fill_1 FILLER_81_246 ();
 sg13g2_fill_1 FILLER_81_264 ();
 sg13g2_fill_2 FILLER_81_361 ();
 sg13g2_fill_1 FILLER_81_384 ();
 sg13g2_fill_2 FILLER_82_0 ();
 sg13g2_fill_1 FILLER_82_2 ();
 sg13g2_fill_2 FILLER_82_20 ();
 sg13g2_decap_4 FILLER_82_162 ();
 sg13g2_fill_1 FILLER_82_166 ();
 sg13g2_fill_1 FILLER_82_196 ();
 sg13g2_decap_4 FILLER_82_249 ();
 sg13g2_fill_1 FILLER_82_253 ();
 sg13g2_fill_1 FILLER_82_271 ();
 sg13g2_fill_1 FILLER_82_306 ();
 sg13g2_fill_2 FILLER_82_336 ();
 sg13g2_fill_2 FILLER_83_4 ();
 sg13g2_fill_1 FILLER_83_6 ();
 sg13g2_fill_1 FILLER_83_116 ();
 sg13g2_fill_1 FILLER_83_151 ();
 sg13g2_fill_1 FILLER_83_177 ();
 sg13g2_decap_8 FILLER_83_235 ();
 sg13g2_fill_1 FILLER_83_246 ();
 sg13g2_fill_2 FILLER_83_290 ();
 sg13g2_fill_2 FILLER_84_0 ();
 sg13g2_fill_2 FILLER_84_19 ();
 sg13g2_fill_1 FILLER_84_21 ();
 sg13g2_fill_2 FILLER_84_36 ();
 sg13g2_fill_1 FILLER_84_84 ();
 sg13g2_decap_4 FILLER_84_95 ();
 sg13g2_fill_2 FILLER_84_99 ();
 sg13g2_fill_1 FILLER_84_131 ();
 sg13g2_fill_2 FILLER_84_149 ();
 sg13g2_fill_1 FILLER_84_151 ();
 sg13g2_decap_8 FILLER_84_219 ();
 sg13g2_decap_4 FILLER_84_226 ();
 sg13g2_fill_1 FILLER_84_230 ();
 sg13g2_fill_2 FILLER_84_248 ();
 sg13g2_fill_1 FILLER_84_250 ();
 sg13g2_fill_2 FILLER_84_268 ();
 sg13g2_fill_2 FILLER_84_287 ();
 sg13g2_fill_2 FILLER_84_304 ();
 sg13g2_fill_2 FILLER_84_328 ();
 sg13g2_fill_1 FILLER_84_356 ();
 sg13g2_fill_2 FILLER_85_95 ();
 sg13g2_fill_1 FILLER_85_139 ();
 sg13g2_fill_2 FILLER_85_186 ();
 sg13g2_decap_8 FILLER_85_222 ();
 sg13g2_fill_2 FILLER_85_229 ();
 sg13g2_fill_1 FILLER_85_231 ();
 sg13g2_fill_1 FILLER_85_354 ();
 sg13g2_fill_1 FILLER_85_384 ();
 sg13g2_fill_2 FILLER_86_21 ();
 sg13g2_fill_2 FILLER_86_37 ();
 sg13g2_fill_1 FILLER_86_39 ();
 sg13g2_fill_2 FILLER_86_99 ();
 sg13g2_fill_1 FILLER_86_101 ();
 sg13g2_fill_2 FILLER_86_124 ();
 sg13g2_fill_2 FILLER_86_134 ();
 sg13g2_fill_2 FILLER_86_180 ();
 sg13g2_fill_1 FILLER_86_200 ();
 sg13g2_fill_2 FILLER_86_223 ();
 sg13g2_fill_1 FILLER_86_225 ();
 sg13g2_decap_8 FILLER_86_243 ();
 sg13g2_decap_8 FILLER_86_250 ();
 sg13g2_fill_1 FILLER_86_269 ();
 sg13g2_fill_2 FILLER_86_295 ();
 sg13g2_fill_1 FILLER_86_319 ();
 sg13g2_fill_1 FILLER_86_330 ();
 sg13g2_fill_1 FILLER_86_344 ();
 sg13g2_fill_1 FILLER_86_358 ();
 sg13g2_fill_1 FILLER_87_13 ();
 sg13g2_fill_2 FILLER_87_35 ();
 sg13g2_fill_2 FILLER_87_53 ();
 sg13g2_fill_1 FILLER_87_55 ();
 sg13g2_fill_2 FILLER_87_111 ();
 sg13g2_fill_2 FILLER_87_173 ();
 sg13g2_fill_2 FILLER_87_212 ();
 sg13g2_fill_1 FILLER_87_214 ();
 sg13g2_fill_1 FILLER_87_327 ();
 sg13g2_fill_1 FILLER_87_368 ();
 sg13g2_fill_2 FILLER_88_0 ();
 sg13g2_fill_2 FILLER_88_38 ();
 sg13g2_fill_1 FILLER_88_40 ();
 sg13g2_fill_2 FILLER_88_46 ();
 sg13g2_fill_2 FILLER_88_164 ();
 sg13g2_fill_2 FILLER_88_214 ();
 sg13g2_decap_8 FILLER_88_254 ();
 sg13g2_decap_4 FILLER_88_261 ();
 sg13g2_fill_1 FILLER_88_265 ();
 sg13g2_fill_2 FILLER_88_283 ();
 sg13g2_fill_1 FILLER_88_311 ();
 sg13g2_fill_1 FILLER_88_338 ();
 sg13g2_fill_1 FILLER_89_4 ();
 sg13g2_fill_2 FILLER_89_57 ();
 sg13g2_fill_1 FILLER_89_59 ();
 sg13g2_fill_2 FILLER_89_73 ();
 sg13g2_fill_1 FILLER_89_75 ();
 sg13g2_fill_2 FILLER_89_103 ();
 sg13g2_fill_1 FILLER_89_169 ();
 sg13g2_fill_1 FILLER_89_310 ();
 sg13g2_fill_2 FILLER_89_341 ();
 sg13g2_fill_2 FILLER_90_40 ();
 sg13g2_fill_1 FILLER_90_63 ();
 sg13g2_fill_1 FILLER_90_111 ();
 sg13g2_fill_1 FILLER_90_171 ();
 sg13g2_decap_4 FILLER_90_218 ();
 sg13g2_decap_8 FILLER_90_260 ();
 sg13g2_decap_4 FILLER_90_267 ();
 sg13g2_fill_2 FILLER_90_271 ();
 sg13g2_fill_1 FILLER_90_318 ();
 sg13g2_fill_1 FILLER_91_0 ();
 sg13g2_fill_2 FILLER_91_29 ();
 sg13g2_fill_1 FILLER_91_31 ();
 sg13g2_fill_2 FILLER_91_42 ();
 sg13g2_fill_1 FILLER_91_125 ();
 sg13g2_fill_1 FILLER_91_187 ();
 sg13g2_fill_1 FILLER_91_231 ();
 sg13g2_decap_8 FILLER_91_270 ();
 sg13g2_fill_1 FILLER_91_277 ();
 sg13g2_fill_2 FILLER_91_307 ();
 sg13g2_fill_1 FILLER_91_309 ();
 sg13g2_fill_2 FILLER_91_372 ();
 sg13g2_fill_2 FILLER_91_379 ();
 sg13g2_fill_2 FILLER_92_0 ();
 sg13g2_fill_1 FILLER_92_2 ();
 sg13g2_fill_2 FILLER_92_141 ();
 sg13g2_fill_1 FILLER_92_143 ();
 sg13g2_fill_2 FILLER_92_161 ();
 sg13g2_fill_1 FILLER_92_163 ();
 sg13g2_decap_4 FILLER_92_195 ();
 sg13g2_fill_2 FILLER_92_204 ();
 sg13g2_fill_1 FILLER_92_206 ();
 sg13g2_fill_2 FILLER_92_228 ();
 sg13g2_fill_1 FILLER_92_251 ();
 sg13g2_decap_4 FILLER_92_269 ();
 sg13g2_fill_1 FILLER_92_273 ();
 sg13g2_fill_1 FILLER_92_299 ();
 sg13g2_fill_1 FILLER_92_339 ();
 sg13g2_fill_1 FILLER_92_358 ();
 sg13g2_fill_2 FILLER_93_0 ();
 sg13g2_fill_1 FILLER_93_2 ();
 sg13g2_fill_1 FILLER_93_28 ();
 sg13g2_fill_1 FILLER_93_44 ();
 sg13g2_decap_4 FILLER_93_95 ();
 sg13g2_fill_2 FILLER_93_99 ();
 sg13g2_fill_1 FILLER_93_105 ();
 sg13g2_fill_2 FILLER_93_182 ();
 sg13g2_fill_1 FILLER_93_184 ();
 sg13g2_fill_2 FILLER_93_202 ();
 sg13g2_fill_1 FILLER_93_226 ();
 sg13g2_fill_2 FILLER_93_257 ();
 sg13g2_fill_1 FILLER_93_259 ();
 sg13g2_fill_2 FILLER_93_319 ();
 sg13g2_fill_1 FILLER_93_376 ();
 sg13g2_fill_2 FILLER_94_0 ();
 sg13g2_fill_1 FILLER_94_2 ();
 sg13g2_fill_2 FILLER_94_20 ();
 sg13g2_fill_1 FILLER_94_22 ();
 sg13g2_fill_1 FILLER_94_49 ();
 sg13g2_decap_4 FILLER_94_95 ();
 sg13g2_fill_2 FILLER_94_99 ();
 sg13g2_decap_8 FILLER_94_118 ();
 sg13g2_decap_8 FILLER_94_125 ();
 sg13g2_fill_2 FILLER_94_166 ();
 sg13g2_fill_1 FILLER_94_168 ();
 sg13g2_fill_2 FILLER_94_186 ();
 sg13g2_fill_1 FILLER_94_188 ();
 sg13g2_fill_2 FILLER_94_203 ();
 sg13g2_fill_2 FILLER_94_215 ();
 sg13g2_fill_2 FILLER_94_255 ();
 sg13g2_fill_2 FILLER_94_310 ();
 sg13g2_fill_1 FILLER_94_312 ();
 sg13g2_fill_2 FILLER_94_346 ();
 sg13g2_fill_1 FILLER_94_380 ();
 sg13g2_fill_1 FILLER_95_21 ();
 sg13g2_fill_2 FILLER_95_80 ();
 sg13g2_fill_1 FILLER_95_99 ();
 sg13g2_fill_2 FILLER_95_121 ();
 sg13g2_decap_4 FILLER_95_148 ();
 sg13g2_fill_2 FILLER_95_152 ();
 sg13g2_fill_2 FILLER_95_210 ();
 sg13g2_decap_8 FILLER_95_229 ();
 sg13g2_fill_2 FILLER_95_265 ();
 sg13g2_fill_1 FILLER_95_267 ();
 sg13g2_fill_2 FILLER_95_285 ();
 sg13g2_fill_1 FILLER_95_321 ();
 sg13g2_fill_1 FILLER_95_347 ();
 sg13g2_fill_2 FILLER_95_366 ();
 sg13g2_fill_1 FILLER_95_368 ();
 sg13g2_fill_1 FILLER_95_384 ();
 sg13g2_fill_2 FILLER_96_42 ();
 sg13g2_fill_1 FILLER_96_81 ();
 sg13g2_decap_8 FILLER_96_97 ();
 sg13g2_decap_4 FILLER_96_104 ();
 sg13g2_fill_2 FILLER_96_108 ();
 sg13g2_fill_2 FILLER_96_115 ();
 sg13g2_fill_1 FILLER_96_117 ();
 sg13g2_fill_2 FILLER_96_132 ();
 sg13g2_decap_8 FILLER_96_176 ();
 sg13g2_decap_4 FILLER_96_183 ();
 sg13g2_fill_1 FILLER_96_191 ();
 sg13g2_fill_2 FILLER_96_205 ();
 sg13g2_fill_1 FILLER_96_207 ();
 sg13g2_decap_4 FILLER_96_212 ();
 sg13g2_fill_1 FILLER_96_216 ();
 sg13g2_decap_8 FILLER_96_221 ();
 sg13g2_decap_4 FILLER_96_228 ();
 sg13g2_fill_2 FILLER_96_232 ();
 sg13g2_decap_4 FILLER_96_244 ();
 sg13g2_fill_1 FILLER_96_248 ();
 sg13g2_fill_1 FILLER_96_292 ();
 sg13g2_fill_2 FILLER_96_300 ();
 sg13g2_decap_8 FILLER_96_306 ();
 sg13g2_fill_2 FILLER_97_0 ();
 sg13g2_fill_2 FILLER_97_23 ();
 sg13g2_fill_1 FILLER_97_25 ();
 sg13g2_fill_2 FILLER_97_46 ();
 sg13g2_fill_2 FILLER_97_56 ();
 sg13g2_fill_2 FILLER_97_127 ();
 sg13g2_fill_1 FILLER_97_129 ();
 sg13g2_decap_4 FILLER_97_147 ();
 sg13g2_fill_2 FILLER_97_151 ();
 sg13g2_decap_8 FILLER_97_170 ();
 sg13g2_fill_2 FILLER_97_177 ();
 sg13g2_decap_8 FILLER_97_217 ();
 sg13g2_fill_2 FILLER_97_224 ();
 sg13g2_fill_1 FILLER_97_226 ();
 sg13g2_fill_1 FILLER_97_231 ();
 sg13g2_decap_8 FILLER_97_248 ();
 sg13g2_decap_8 FILLER_97_255 ();
 sg13g2_decap_4 FILLER_97_278 ();
 sg13g2_fill_2 FILLER_97_282 ();
 sg13g2_fill_2 FILLER_97_288 ();
 sg13g2_fill_2 FILLER_97_299 ();
 sg13g2_fill_2 FILLER_97_322 ();
 sg13g2_fill_2 FILLER_97_383 ();
 sg13g2_fill_2 FILLER_98_21 ();
 sg13g2_fill_1 FILLER_98_23 ();
 sg13g2_fill_2 FILLER_98_45 ();
 sg13g2_fill_1 FILLER_98_47 ();
 sg13g2_fill_2 FILLER_98_73 ();
 sg13g2_fill_2 FILLER_98_86 ();
 sg13g2_fill_2 FILLER_98_130 ();
 sg13g2_fill_1 FILLER_98_132 ();
 sg13g2_decap_4 FILLER_98_158 ();
 sg13g2_fill_1 FILLER_98_162 ();
 sg13g2_fill_2 FILLER_98_184 ();
 sg13g2_fill_1 FILLER_98_186 ();
 sg13g2_fill_2 FILLER_98_256 ();
 sg13g2_fill_1 FILLER_98_258 ();
 sg13g2_fill_2 FILLER_98_264 ();
 sg13g2_fill_1 FILLER_98_266 ();
 sg13g2_fill_2 FILLER_98_272 ();
 sg13g2_fill_1 FILLER_98_317 ();
 sg13g2_fill_1 FILLER_98_376 ();
 sg13g2_fill_1 FILLER_99_4 ();
 sg13g2_fill_1 FILLER_99_26 ();
 sg13g2_fill_1 FILLER_99_46 ();
 sg13g2_fill_1 FILLER_99_68 ();
 sg13g2_fill_1 FILLER_99_78 ();
 sg13g2_fill_2 FILLER_99_84 ();
 sg13g2_fill_1 FILLER_99_113 ();
 sg13g2_decap_8 FILLER_99_133 ();
 sg13g2_decap_8 FILLER_99_140 ();
 sg13g2_decap_8 FILLER_99_147 ();
 sg13g2_decap_4 FILLER_99_154 ();
 sg13g2_fill_2 FILLER_99_158 ();
 sg13g2_fill_2 FILLER_99_164 ();
 sg13g2_fill_1 FILLER_99_166 ();
 sg13g2_fill_2 FILLER_99_184 ();
 sg13g2_fill_1 FILLER_99_186 ();
 sg13g2_decap_8 FILLER_99_204 ();
 sg13g2_decap_8 FILLER_99_211 ();
 sg13g2_fill_1 FILLER_99_218 ();
 sg13g2_fill_2 FILLER_99_241 ();
 sg13g2_fill_2 FILLER_99_265 ();
 sg13g2_fill_1 FILLER_99_267 ();
 sg13g2_decap_4 FILLER_99_285 ();
 sg13g2_fill_1 FILLER_99_289 ();
 sg13g2_fill_1 FILLER_99_294 ();
 sg13g2_decap_4 FILLER_99_323 ();
 sg13g2_fill_2 FILLER_99_331 ();
 sg13g2_fill_1 FILLER_99_333 ();
 sg13g2_fill_1 FILLER_99_354 ();
 sg13g2_fill_2 FILLER_99_375 ();
 sg13g2_fill_2 FILLER_100_0 ();
 sg13g2_fill_1 FILLER_100_2 ();
 sg13g2_fill_1 FILLER_100_52 ();
 sg13g2_fill_1 FILLER_100_73 ();
 sg13g2_decap_8 FILLER_100_95 ();
 sg13g2_decap_4 FILLER_100_102 ();
 sg13g2_fill_2 FILLER_100_106 ();
 sg13g2_decap_4 FILLER_100_161 ();
 sg13g2_fill_2 FILLER_100_165 ();
 sg13g2_decap_4 FILLER_100_192 ();
 sg13g2_decap_8 FILLER_100_213 ();
 sg13g2_decap_8 FILLER_100_220 ();
 sg13g2_fill_2 FILLER_100_230 ();
 sg13g2_fill_1 FILLER_100_232 ();
 sg13g2_decap_4 FILLER_100_242 ();
 sg13g2_decap_8 FILLER_100_277 ();
 sg13g2_fill_1 FILLER_100_284 ();
 sg13g2_decap_8 FILLER_100_294 ();
 sg13g2_decap_4 FILLER_100_301 ();
 sg13g2_fill_2 FILLER_100_305 ();
 sg13g2_fill_1 FILLER_100_324 ();
 sg13g2_fill_2 FILLER_100_342 ();
 sg13g2_fill_1 FILLER_100_352 ();
 sg13g2_fill_2 FILLER_101_4 ();
 sg13g2_fill_1 FILLER_101_53 ();
 sg13g2_decap_8 FILLER_101_80 ();
 sg13g2_decap_4 FILLER_101_87 ();
 sg13g2_fill_1 FILLER_101_91 ();
 sg13g2_fill_1 FILLER_101_96 ();
 sg13g2_fill_1 FILLER_101_118 ();
 sg13g2_fill_1 FILLER_101_157 ();
 sg13g2_fill_2 FILLER_101_175 ();
 sg13g2_fill_1 FILLER_101_177 ();
 sg13g2_decap_8 FILLER_101_198 ();
 sg13g2_decap_8 FILLER_101_205 ();
 sg13g2_fill_2 FILLER_101_212 ();
 sg13g2_decap_4 FILLER_101_266 ();
 sg13g2_fill_1 FILLER_101_270 ();
 sg13g2_fill_2 FILLER_101_321 ();
 sg13g2_fill_1 FILLER_101_323 ();
 sg13g2_fill_2 FILLER_101_338 ();
 sg13g2_fill_2 FILLER_101_356 ();
 sg13g2_fill_2 FILLER_101_368 ();
 sg13g2_fill_1 FILLER_101_370 ();
 sg13g2_fill_2 FILLER_101_379 ();
 sg13g2_fill_1 FILLER_102_8 ();
 sg13g2_fill_2 FILLER_102_46 ();
 sg13g2_decap_8 FILLER_102_64 ();
 sg13g2_fill_1 FILLER_102_71 ();
 sg13g2_decap_4 FILLER_102_77 ();
 sg13g2_fill_2 FILLER_102_81 ();
 sg13g2_fill_1 FILLER_102_104 ();
 sg13g2_decap_8 FILLER_102_110 ();
 sg13g2_fill_2 FILLER_102_117 ();
 sg13g2_fill_2 FILLER_102_140 ();
 sg13g2_decap_4 FILLER_102_159 ();
 sg13g2_fill_1 FILLER_102_163 ();
 sg13g2_decap_8 FILLER_102_251 ();
 sg13g2_decap_8 FILLER_102_258 ();
 sg13g2_fill_2 FILLER_102_265 ();
 sg13g2_fill_1 FILLER_102_309 ();
 sg13g2_fill_2 FILLER_102_383 ();
 sg13g2_fill_2 FILLER_103_0 ();
 sg13g2_fill_1 FILLER_103_2 ();
 sg13g2_fill_2 FILLER_103_20 ();
 sg13g2_fill_1 FILLER_103_22 ();
 sg13g2_fill_1 FILLER_103_27 ();
 sg13g2_fill_1 FILLER_103_41 ();
 sg13g2_fill_2 FILLER_103_50 ();
 sg13g2_decap_4 FILLER_103_77 ();
 sg13g2_fill_2 FILLER_103_144 ();
 sg13g2_decap_8 FILLER_103_163 ();
 sg13g2_fill_2 FILLER_103_170 ();
 sg13g2_fill_1 FILLER_103_172 ();
 sg13g2_decap_8 FILLER_103_198 ();
 sg13g2_decap_4 FILLER_103_222 ();
 sg13g2_fill_1 FILLER_103_226 ();
 sg13g2_decap_8 FILLER_103_244 ();
 sg13g2_decap_4 FILLER_103_251 ();
 sg13g2_fill_1 FILLER_103_255 ();
 sg13g2_decap_4 FILLER_103_287 ();
 sg13g2_fill_2 FILLER_103_299 ();
 sg13g2_fill_1 FILLER_103_301 ();
 sg13g2_fill_1 FILLER_103_319 ();
 sg13g2_fill_1 FILLER_103_376 ();
 sg13g2_fill_1 FILLER_104_58 ();
 sg13g2_fill_2 FILLER_104_69 ();
 sg13g2_fill_1 FILLER_104_71 ();
 sg13g2_decap_8 FILLER_104_96 ();
 sg13g2_decap_8 FILLER_104_103 ();
 sg13g2_fill_2 FILLER_104_110 ();
 sg13g2_fill_1 FILLER_104_112 ();
 sg13g2_fill_2 FILLER_104_129 ();
 sg13g2_decap_8 FILLER_104_137 ();
 sg13g2_fill_1 FILLER_104_144 ();
 sg13g2_decap_4 FILLER_104_166 ();
 sg13g2_fill_1 FILLER_104_170 ();
 sg13g2_decap_8 FILLER_104_175 ();
 sg13g2_decap_8 FILLER_104_187 ();
 sg13g2_decap_8 FILLER_104_194 ();
 sg13g2_decap_8 FILLER_104_201 ();
 sg13g2_decap_4 FILLER_104_225 ();
 sg13g2_fill_1 FILLER_104_229 ();
 sg13g2_fill_2 FILLER_104_238 ();
 sg13g2_decap_8 FILLER_104_278 ();
 sg13g2_fill_1 FILLER_104_285 ();
 sg13g2_fill_2 FILLER_104_300 ();
 sg13g2_fill_1 FILLER_104_319 ();
 sg13g2_fill_1 FILLER_104_348 ();
 sg13g2_fill_2 FILLER_104_362 ();
 sg13g2_fill_2 FILLER_105_5 ();
 sg13g2_decap_4 FILLER_105_75 ();
 sg13g2_fill_1 FILLER_105_121 ();
 sg13g2_fill_1 FILLER_105_155 ();
 sg13g2_decap_4 FILLER_105_177 ();
 sg13g2_fill_1 FILLER_105_181 ();
 sg13g2_fill_1 FILLER_105_254 ();
 sg13g2_fill_1 FILLER_105_318 ();
 sg13g2_fill_1 FILLER_105_344 ();
 sg13g2_fill_2 FILLER_105_370 ();
 sg13g2_fill_1 FILLER_105_372 ();
 sg13g2_fill_1 FILLER_106_0 ();
 sg13g2_fill_2 FILLER_106_18 ();
 sg13g2_fill_1 FILLER_106_20 ();
 sg13g2_fill_1 FILLER_106_89 ();
 sg13g2_fill_2 FILLER_106_115 ();
 sg13g2_fill_1 FILLER_106_141 ();
 sg13g2_fill_1 FILLER_106_159 ();
 sg13g2_decap_8 FILLER_106_168 ();
 sg13g2_fill_2 FILLER_106_175 ();
 sg13g2_decap_8 FILLER_106_219 ();
 sg13g2_decap_8 FILLER_106_226 ();
 sg13g2_decap_4 FILLER_106_233 ();
 sg13g2_fill_1 FILLER_106_237 ();
 sg13g2_decap_4 FILLER_106_255 ();
 sg13g2_fill_2 FILLER_106_259 ();
 sg13g2_fill_2 FILLER_106_278 ();
 sg13g2_fill_1 FILLER_106_283 ();
 sg13g2_fill_2 FILLER_107_12 ();
 sg13g2_fill_1 FILLER_107_14 ();
 sg13g2_fill_2 FILLER_107_23 ();
 sg13g2_fill_1 FILLER_107_25 ();
 sg13g2_fill_2 FILLER_107_64 ();
 sg13g2_decap_8 FILLER_107_83 ();
 sg13g2_fill_2 FILLER_107_161 ();
 sg13g2_decap_8 FILLER_107_214 ();
 sg13g2_fill_2 FILLER_107_221 ();
 sg13g2_fill_2 FILLER_107_240 ();
 sg13g2_fill_1 FILLER_107_267 ();
 sg13g2_fill_1 FILLER_107_285 ();
 sg13g2_decap_4 FILLER_107_290 ();
 sg13g2_fill_1 FILLER_107_310 ();
 sg13g2_fill_2 FILLER_107_330 ();
 sg13g2_fill_2 FILLER_107_353 ();
 sg13g2_fill_2 FILLER_108_0 ();
 sg13g2_fill_1 FILLER_108_40 ();
 sg13g2_fill_2 FILLER_108_50 ();
 sg13g2_fill_1 FILLER_108_52 ();
 sg13g2_fill_2 FILLER_108_95 ();
 sg13g2_fill_1 FILLER_108_115 ();
 sg13g2_fill_2 FILLER_108_153 ();
 sg13g2_decap_4 FILLER_108_159 ();
 sg13g2_fill_1 FILLER_108_163 ();
 sg13g2_fill_1 FILLER_108_181 ();
 sg13g2_fill_2 FILLER_108_209 ();
 sg13g2_fill_1 FILLER_108_211 ();
 sg13g2_fill_1 FILLER_108_237 ();
 sg13g2_fill_1 FILLER_108_269 ();
 sg13g2_fill_2 FILLER_108_283 ();
 sg13g2_fill_1 FILLER_108_285 ();
 sg13g2_fill_2 FILLER_108_360 ();
 sg13g2_fill_2 FILLER_108_378 ();
 sg13g2_fill_2 FILLER_109_0 ();
 sg13g2_fill_2 FILLER_109_23 ();
 sg13g2_fill_1 FILLER_109_25 ();
 sg13g2_fill_2 FILLER_109_44 ();
 sg13g2_fill_2 FILLER_109_57 ();
 sg13g2_decap_4 FILLER_109_63 ();
 sg13g2_fill_2 FILLER_109_67 ();
 sg13g2_decap_4 FILLER_109_72 ();
 sg13g2_fill_1 FILLER_109_76 ();
 sg13g2_fill_2 FILLER_109_94 ();
 sg13g2_fill_1 FILLER_109_101 ();
 sg13g2_decap_4 FILLER_109_138 ();
 sg13g2_fill_1 FILLER_109_149 ();
 sg13g2_fill_2 FILLER_109_165 ();
 sg13g2_fill_1 FILLER_109_167 ();
 sg13g2_decap_8 FILLER_109_211 ();
 sg13g2_fill_1 FILLER_109_218 ();
 sg13g2_fill_2 FILLER_109_240 ();
 sg13g2_decap_8 FILLER_109_246 ();
 sg13g2_decap_8 FILLER_109_253 ();
 sg13g2_fill_1 FILLER_109_297 ();
 sg13g2_fill_1 FILLER_109_307 ();
 sg13g2_fill_1 FILLER_109_384 ();
 sg13g2_fill_2 FILLER_110_4 ();
 sg13g2_fill_1 FILLER_110_6 ();
 sg13g2_fill_2 FILLER_110_24 ();
 sg13g2_fill_2 FILLER_110_36 ();
 sg13g2_fill_1 FILLER_110_38 ();
 sg13g2_fill_2 FILLER_110_68 ();
 sg13g2_fill_1 FILLER_110_104 ();
 sg13g2_fill_1 FILLER_110_159 ();
 sg13g2_fill_1 FILLER_110_178 ();
 sg13g2_fill_2 FILLER_110_184 ();
 sg13g2_decap_8 FILLER_110_190 ();
 sg13g2_fill_2 FILLER_110_197 ();
 sg13g2_fill_2 FILLER_110_203 ();
 sg13g2_fill_2 FILLER_110_226 ();
 sg13g2_fill_1 FILLER_110_228 ();
 sg13g2_decap_4 FILLER_110_237 ();
 sg13g2_fill_2 FILLER_110_325 ();
 sg13g2_fill_2 FILLER_110_365 ();
 sg13g2_fill_2 FILLER_111_117 ();
 sg13g2_decap_8 FILLER_111_134 ();
 sg13g2_fill_1 FILLER_111_187 ();
 sg13g2_decap_4 FILLER_111_227 ();
 sg13g2_fill_2 FILLER_111_235 ();
 sg13g2_fill_1 FILLER_111_237 ();
 sg13g2_fill_2 FILLER_111_296 ();
 sg13g2_fill_2 FILLER_111_365 ();
 sg13g2_fill_1 FILLER_112_0 ();
 sg13g2_fill_1 FILLER_112_18 ();
 sg13g2_decap_4 FILLER_112_23 ();
 sg13g2_fill_1 FILLER_112_27 ();
 sg13g2_fill_1 FILLER_112_32 ();
 sg13g2_decap_4 FILLER_112_47 ();
 sg13g2_decap_8 FILLER_112_56 ();
 sg13g2_decap_8 FILLER_112_63 ();
 sg13g2_fill_1 FILLER_112_70 ();
 sg13g2_decap_8 FILLER_112_75 ();
 sg13g2_decap_8 FILLER_112_82 ();
 sg13g2_fill_2 FILLER_112_93 ();
 sg13g2_fill_1 FILLER_112_95 ();
 sg13g2_fill_2 FILLER_112_110 ();
 sg13g2_decap_8 FILLER_112_129 ();
 sg13g2_decap_4 FILLER_112_136 ();
 sg13g2_fill_2 FILLER_112_140 ();
 sg13g2_fill_1 FILLER_112_188 ();
 sg13g2_fill_1 FILLER_112_267 ();
 sg13g2_fill_1 FILLER_112_278 ();
 sg13g2_fill_2 FILLER_112_324 ();
 sg13g2_fill_2 FILLER_112_382 ();
 sg13g2_fill_1 FILLER_112_384 ();
 sg13g2_fill_2 FILLER_113_0 ();
 sg13g2_decap_4 FILLER_113_27 ();
 sg13g2_fill_2 FILLER_113_40 ();
 sg13g2_decap_4 FILLER_113_84 ();
 sg13g2_decap_8 FILLER_113_92 ();
 sg13g2_decap_4 FILLER_113_99 ();
 sg13g2_decap_4 FILLER_113_108 ();
 sg13g2_fill_1 FILLER_113_182 ();
 sg13g2_fill_2 FILLER_113_208 ();
 sg13g2_fill_2 FILLER_113_252 ();
 sg13g2_fill_1 FILLER_113_279 ();
 sg13g2_fill_1 FILLER_113_320 ();
 sg13g2_fill_2 FILLER_113_353 ();
 sg13g2_fill_2 FILLER_113_373 ();
 sg13g2_fill_1 FILLER_113_384 ();
 sg13g2_fill_2 FILLER_114_0 ();
 sg13g2_fill_1 FILLER_114_2 ();
 sg13g2_fill_2 FILLER_114_61 ();
 sg13g2_fill_1 FILLER_114_67 ();
 sg13g2_fill_1 FILLER_114_102 ();
 sg13g2_fill_1 FILLER_114_150 ();
 sg13g2_fill_1 FILLER_114_204 ();
 sg13g2_fill_2 FILLER_114_213 ();
 sg13g2_fill_1 FILLER_114_215 ();
 sg13g2_fill_2 FILLER_114_233 ();
 sg13g2_fill_1 FILLER_114_273 ();
 sg13g2_fill_2 FILLER_114_282 ();
 sg13g2_fill_2 FILLER_114_349 ();
 sg13g2_fill_1 FILLER_115_0 ();
 sg13g2_decap_8 FILLER_115_56 ();
 sg13g2_fill_2 FILLER_115_63 ();
 sg13g2_fill_2 FILLER_115_82 ();
 sg13g2_fill_1 FILLER_115_84 ();
 sg13g2_fill_1 FILLER_115_131 ();
 sg13g2_fill_2 FILLER_115_149 ();
 sg13g2_decap_8 FILLER_115_156 ();
 sg13g2_fill_2 FILLER_115_163 ();
 sg13g2_fill_1 FILLER_115_165 ();
 sg13g2_fill_2 FILLER_115_169 ();
 sg13g2_fill_1 FILLER_115_188 ();
 sg13g2_fill_2 FILLER_115_194 ();
 sg13g2_fill_2 FILLER_115_234 ();
 sg13g2_fill_2 FILLER_115_253 ();
 sg13g2_fill_2 FILLER_115_290 ();
 sg13g2_fill_1 FILLER_115_313 ();
 sg13g2_fill_2 FILLER_115_359 ();
 sg13g2_fill_2 FILLER_115_371 ();
 sg13g2_fill_1 FILLER_116_0 ();
 sg13g2_fill_1 FILLER_116_18 ();
 sg13g2_fill_2 FILLER_116_48 ();
 sg13g2_fill_1 FILLER_116_134 ();
 sg13g2_fill_1 FILLER_116_139 ();
 sg13g2_fill_1 FILLER_116_188 ();
 sg13g2_fill_1 FILLER_116_193 ();
 sg13g2_fill_1 FILLER_116_219 ();
 sg13g2_fill_1 FILLER_116_283 ();
 sg13g2_fill_2 FILLER_116_324 ();
 sg13g2_fill_2 FILLER_117_0 ();
 sg13g2_fill_1 FILLER_117_2 ();
 sg13g2_fill_1 FILLER_117_11 ();
 sg13g2_fill_2 FILLER_117_16 ();
 sg13g2_fill_1 FILLER_117_18 ();
 sg13g2_fill_1 FILLER_117_48 ();
 sg13g2_fill_1 FILLER_117_76 ();
 sg13g2_fill_1 FILLER_117_85 ();
 sg13g2_fill_2 FILLER_117_148 ();
 sg13g2_fill_2 FILLER_117_218 ();
 sg13g2_fill_1 FILLER_117_220 ();
 sg13g2_fill_2 FILLER_117_246 ();
 sg13g2_fill_2 FILLER_117_252 ();
 sg13g2_fill_1 FILLER_117_254 ();
 sg13g2_fill_2 FILLER_117_259 ();
 sg13g2_fill_1 FILLER_117_261 ();
 sg13g2_fill_1 FILLER_117_278 ();
 sg13g2_fill_1 FILLER_117_312 ();
 sg13g2_fill_1 FILLER_117_321 ();
 sg13g2_fill_1 FILLER_117_326 ();
 sg13g2_fill_2 FILLER_117_353 ();
 sg13g2_fill_2 FILLER_118_0 ();
 sg13g2_fill_1 FILLER_118_2 ();
 sg13g2_fill_2 FILLER_118_11 ();
 sg13g2_fill_1 FILLER_118_51 ();
 sg13g2_fill_2 FILLER_118_57 ();
 sg13g2_fill_1 FILLER_118_59 ();
 sg13g2_fill_1 FILLER_118_86 ();
 sg13g2_fill_1 FILLER_118_105 ();
 sg13g2_fill_2 FILLER_118_141 ();
 sg13g2_fill_1 FILLER_118_143 ();
 sg13g2_fill_2 FILLER_118_220 ();
 sg13g2_fill_1 FILLER_118_222 ();
 sg13g2_fill_2 FILLER_118_273 ();
 sg13g2_fill_1 FILLER_118_275 ();
 sg13g2_fill_2 FILLER_118_344 ();
 sg13g2_fill_1 FILLER_118_373 ();
 sg13g2_fill_1 FILLER_119_0 ();
 sg13g2_fill_2 FILLER_119_75 ();
 sg13g2_fill_2 FILLER_119_94 ();
 sg13g2_fill_1 FILLER_119_96 ();
 sg13g2_fill_1 FILLER_119_110 ();
 sg13g2_fill_2 FILLER_119_194 ();
 sg13g2_fill_1 FILLER_119_196 ();
 sg13g2_fill_1 FILLER_119_214 ();
 sg13g2_fill_2 FILLER_119_219 ();
 sg13g2_fill_1 FILLER_119_221 ();
 sg13g2_fill_2 FILLER_119_288 ();
 sg13g2_fill_2 FILLER_120_0 ();
 sg13g2_fill_1 FILLER_120_2 ();
 sg13g2_fill_1 FILLER_120_61 ();
 sg13g2_fill_2 FILLER_120_92 ();
 sg13g2_fill_2 FILLER_120_119 ();
 sg13g2_fill_1 FILLER_120_136 ();
 sg13g2_fill_2 FILLER_120_314 ();
 sg13g2_fill_1 FILLER_120_316 ();
 sg13g2_fill_1 FILLER_120_357 ();
 sg13g2_fill_2 FILLER_121_0 ();
 sg13g2_fill_2 FILLER_121_105 ();
 sg13g2_fill_2 FILLER_121_128 ();
 sg13g2_fill_1 FILLER_121_135 ();
 sg13g2_fill_2 FILLER_121_239 ();
 sg13g2_fill_1 FILLER_121_258 ();
 sg13g2_fill_1 FILLER_121_301 ();
 sg13g2_fill_2 FILLER_122_0 ();
 sg13g2_fill_1 FILLER_122_2 ();
 sg13g2_fill_2 FILLER_122_67 ();
 sg13g2_fill_1 FILLER_122_69 ();
 sg13g2_fill_1 FILLER_122_119 ();
 sg13g2_fill_1 FILLER_122_166 ();
 sg13g2_fill_2 FILLER_122_189 ();
 sg13g2_fill_1 FILLER_122_191 ();
 sg13g2_fill_1 FILLER_122_213 ();
 sg13g2_fill_1 FILLER_122_218 ();
 sg13g2_fill_1 FILLER_122_235 ();
 sg13g2_fill_2 FILLER_122_303 ();
 sg13g2_fill_2 FILLER_122_359 ();
 sg13g2_fill_1 FILLER_122_361 ();
 sg13g2_fill_2 FILLER_123_0 ();
 sg13g2_fill_1 FILLER_123_2 ();
 sg13g2_fill_2 FILLER_123_44 ();
 sg13g2_fill_1 FILLER_123_46 ();
 sg13g2_fill_2 FILLER_123_70 ();
 sg13g2_fill_1 FILLER_123_72 ();
 sg13g2_fill_2 FILLER_123_81 ();
 sg13g2_fill_1 FILLER_123_83 ();
 sg13g2_fill_2 FILLER_123_113 ();
 sg13g2_fill_2 FILLER_123_166 ();
 sg13g2_fill_2 FILLER_123_227 ();
 sg13g2_fill_2 FILLER_123_281 ();
 sg13g2_fill_1 FILLER_123_283 ();
 sg13g2_fill_2 FILLER_123_374 ();
 sg13g2_fill_1 FILLER_123_376 ();
endmodule
