module S_CPU_IF (Co,
    I_top0,
    I_top1,
    I_top10,
    I_top11,
    I_top12,
    I_top13,
    I_top14,
    I_top15,
    I_top2,
    I_top3,
    I_top4,
    I_top5,
    I_top6,
    I_top7,
    I_top8,
    I_top9,
    O_top0,
    O_top1,
    O_top10,
    O_top11,
    O_top12,
    O_top13,
    O_top14,
    O_top15,
    O_top2,
    O_top3,
    O_top4,
    O_top5,
    O_top6,
    O_top7,
    O_top8,
    O_top9,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output Co;
 output I_top0;
 output I_top1;
 output I_top10;
 output I_top11;
 output I_top12;
 output I_top13;
 output I_top14;
 output I_top15;
 output I_top2;
 output I_top3;
 output I_top4;
 output I_top5;
 output I_top6;
 output I_top7;
 output I_top8;
 output I_top9;
 input O_top0;
 input O_top1;
 input O_top10;
 input O_top11;
 input O_top12;
 input O_top13;
 input O_top14;
 input O_top15;
 input O_top2;
 input O_top3;
 input O_top4;
 input O_top5;
 input O_top6;
 input O_top7;
 input O_top8;
 input O_top9;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG4 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG5 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG6 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG7 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb4 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb5 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb6 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb7 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG10 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG11 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG12 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG13 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG14 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG15 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG4 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG5 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG6 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG7 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG8 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG9 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG10 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG11 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG12 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG13 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG14 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG15 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG4 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG5 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG6 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG7 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG8 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG9 ;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net233;

 sky130_fd_sc_hd__mux4_1 _000_ (.A0(net63),
    .A1(net79),
    .A2(net86),
    .A3(net102),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .X(net171));
 sky130_fd_sc_hd__mux4_1 _001_ (.A0(net62),
    .A1(net78),
    .A2(net85),
    .A3(net101),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .X(net170));
 sky130_fd_sc_hd__mux4_1 _002_ (.A0(net61),
    .A1(net77),
    .A2(net84),
    .A3(net100),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 _003_ (.A0(net60),
    .A1(net76),
    .A2(net83),
    .A3(net99),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .X(net168));
 sky130_fd_sc_hd__mux4_1 _004_ (.A0(net63),
    .A1(net71),
    .A2(net82),
    .A3(net98),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q ),
    .X(net167));
 sky130_fd_sc_hd__mux4_1 _005_ (.A0(net62),
    .A1(net70),
    .A2(net81),
    .A3(net97),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q ),
    .X(net166));
 sky130_fd_sc_hd__mux4_1 _006_ (.A0(net61),
    .A1(net69),
    .A2(net95),
    .A3(net111),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q ),
    .X(net179));
 sky130_fd_sc_hd__mux4_1 _007_ (.A0(net60),
    .A1(net68),
    .A2(net94),
    .A3(net110),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q ),
    .X(net178));
 sky130_fd_sc_hd__mux4_1 _008_ (.A0(net63),
    .A1(net67),
    .A2(net93),
    .A3(net109),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q ),
    .X(net177));
 sky130_fd_sc_hd__mux4_1 _009_ (.A0(net62),
    .A1(net66),
    .A2(net92),
    .A3(net108),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q ),
    .X(net176));
 sky130_fd_sc_hd__mux4_1 _010_ (.A0(net61),
    .A1(net65),
    .A2(net91),
    .A3(net107),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q ),
    .X(net175));
 sky130_fd_sc_hd__mux4_1 _011_ (.A0(net60),
    .A1(net64),
    .A2(net90),
    .A3(net106),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q ),
    .X(net174));
 sky130_fd_sc_hd__mux4_1 _012_ (.A0(net63),
    .A1(net75),
    .A2(net89),
    .A3(net105),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q ),
    .X(net173));
 sky130_fd_sc_hd__mux4_1 _013_ (.A0(net62),
    .A1(net74),
    .A2(net88),
    .A3(net104),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q ),
    .X(net172));
 sky130_fd_sc_hd__mux4_1 _014_ (.A0(net61),
    .A1(net73),
    .A2(net87),
    .A3(net103),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q ),
    .X(net165));
 sky130_fd_sc_hd__mux4_1 _015_ (.A0(net60),
    .A1(net72),
    .A2(net80),
    .A3(net96),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q ),
    .X(net164));
 sky130_fd_sc_hd__mux2_1 _016_ (.A0(net96),
    .A1(net33),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG15 ));
 sky130_fd_sc_hd__mux2_1 _017_ (.A0(net103),
    .A1(net34),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG14 ));
 sky130_fd_sc_hd__mux2_1 _018_ (.A0(net104),
    .A1(net52),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG13 ));
 sky130_fd_sc_hd__mux2_1 _019_ (.A0(net105),
    .A1(net53),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG12 ));
 sky130_fd_sc_hd__mux2_1 _020_ (.A0(net106),
    .A1(net54),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG11 ));
 sky130_fd_sc_hd__mux2_1 _021_ (.A0(net107),
    .A1(net55),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG10 ));
 sky130_fd_sc_hd__mux2_1 _022_ (.A0(net108),
    .A1(net56),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG9 ));
 sky130_fd_sc_hd__mux2_1 _023_ (.A0(net109),
    .A1(net57),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG8 ));
 sky130_fd_sc_hd__mux2_1 _024_ (.A0(net110),
    .A1(net58),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG7 ));
 sky130_fd_sc_hd__mux2_1 _025_ (.A0(net111),
    .A1(net59),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG6 ));
 sky130_fd_sc_hd__mux2_1 _026_ (.A0(net97),
    .A1(net46),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG5 ));
 sky130_fd_sc_hd__mux2_1 _027_ (.A0(net98),
    .A1(net47),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG4 ));
 sky130_fd_sc_hd__mux2_1 _028_ (.A0(net99),
    .A1(net48),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _029_ (.A0(net100),
    .A1(net49),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__mux2_1 _030_ (.A0(net101),
    .A1(net50),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _031_ (.A0(net102),
    .A1(net51),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__mux2_1 _032_ (.A0(net80),
    .A1(net33),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG15 ));
 sky130_fd_sc_hd__mux2_1 _033_ (.A0(net87),
    .A1(net34),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG14 ));
 sky130_fd_sc_hd__mux2_1 _034_ (.A0(net88),
    .A1(net52),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG13 ));
 sky130_fd_sc_hd__mux2_1 _035_ (.A0(net89),
    .A1(net53),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG12 ));
 sky130_fd_sc_hd__mux2_1 _036_ (.A0(net90),
    .A1(net54),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG11 ));
 sky130_fd_sc_hd__mux2_1 _037_ (.A0(net91),
    .A1(net55),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG10 ));
 sky130_fd_sc_hd__mux2_1 _038_ (.A0(net92),
    .A1(net56),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG9 ));
 sky130_fd_sc_hd__mux2_1 _039_ (.A0(net93),
    .A1(net57),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG8 ));
 sky130_fd_sc_hd__mux2_1 _040_ (.A0(net94),
    .A1(net58),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG7 ));
 sky130_fd_sc_hd__mux2_1 _041_ (.A0(net95),
    .A1(net59),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG6 ));
 sky130_fd_sc_hd__mux2_1 _042_ (.A0(net81),
    .A1(net46),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG5 ));
 sky130_fd_sc_hd__mux2_1 _043_ (.A0(net82),
    .A1(net47),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG4 ));
 sky130_fd_sc_hd__mux2_1 _044_ (.A0(net83),
    .A1(net48),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux2_1 _045_ (.A0(net84),
    .A1(net49),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux2_1 _046_ (.A0(net85),
    .A1(net50),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux2_1 _047_ (.A0(net86),
    .A1(net51),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux2_1 _048_ (.A0(net64),
    .A1(net58),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__mux2_1 _049_ (.A0(net65),
    .A1(net59),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__mux2_1 _050_ (.A0(net66),
    .A1(net46),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__mux2_1 _051_ (.A0(net67),
    .A1(net47),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__mux2_1 _052_ (.A0(net68),
    .A1(net48),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__mux2_1 _053_ (.A0(net69),
    .A1(net49),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__mux2_1 _054_ (.A0(net70),
    .A1(net50),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__mux2_1 _055_ (.A0(net71),
    .A1(net51),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__mux2_1 _056_ (.A0(net72),
    .A1(net33),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG7 ));
 sky130_fd_sc_hd__mux2_1 _057_ (.A0(net73),
    .A1(net34),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG6 ));
 sky130_fd_sc_hd__mux2_1 _058_ (.A0(net74),
    .A1(net52),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG5 ));
 sky130_fd_sc_hd__mux2_1 _059_ (.A0(net75),
    .A1(net53),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG4 ));
 sky130_fd_sc_hd__mux2_1 _060_ (.A0(net76),
    .A1(net54),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG3 ));
 sky130_fd_sc_hd__mux2_1 _061_ (.A0(net77),
    .A1(net55),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG2 ));
 sky130_fd_sc_hd__mux2_1 _062_ (.A0(net78),
    .A1(net56),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG1 ));
 sky130_fd_sc_hd__mux2_1 _063_ (.A0(net79),
    .A1(net57),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG0 ));
 sky130_fd_sc_hd__mux4_1 _064_ (.A0(net60),
    .A1(net33),
    .A2(net54),
    .A3(net48),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_1 _065_ (.A0(net61),
    .A1(net34),
    .A2(net55),
    .A3(net49),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_1 _066_ (.A0(net62),
    .A1(net52),
    .A2(net56),
    .A3(net50),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_1 _067_ (.A0(net63),
    .A1(net53),
    .A2(net57),
    .A3(net51),
    .S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__dlxtp_1 _068_ (.D(net31),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _069_ (.D(net32),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _070_ (.D(net2),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _071_ (.D(net3),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _072_ (.D(net4),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _073_ (.D(net5),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _074_ (.D(net6),
    .GATE(net37),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _075_ (.D(net7),
    .GATE(net37),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _076_ (.D(net8),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _077_ (.D(net9),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _078_ (.D(net10),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _079_ (.D(net11),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _080_ (.D(net13),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _081_ (.D(net14),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _082_ (.D(net15),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _083_ (.D(net16),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _084_ (.D(net17),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _085_ (.D(net18),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _086_ (.D(net19),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _087_ (.D(net20),
    .GATE(net36),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _088_ (.D(net21),
    .GATE(net37),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _089_ (.D(net22),
    .GATE(net37),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _090_ (.D(net24),
    .GATE(net37),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _091_ (.D(net25),
    .GATE(net35),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _092_ (.D(net1),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _093_ (.D(net12),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _094_ (.D(net23),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _095_ (.D(net26),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _096_ (.D(net27),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _097_ (.D(net28),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _098_ (.D(net29),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _099_ (.D(net30),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _100_ (.D(net31),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _101_ (.D(net32),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _102_ (.D(net2),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _103_ (.D(net3),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _104_ (.D(net4),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _105_ (.D(net5),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _106_ (.D(net6),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _107_ (.D(net7),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _108_ (.D(net8),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _109_ (.D(net9),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _110_ (.D(net10),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _111_ (.D(net11),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _112_ (.D(net13),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _113_ (.D(net14),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _114_ (.D(net15),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _115_ (.D(net16),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _116_ (.D(net17),
    .GATE(net38),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _117_ (.D(net18),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _118_ (.D(net19),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _119_ (.D(net20),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _120_ (.D(net21),
    .GATE(net39),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _121_ (.D(net22),
    .GATE(net41),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _122_ (.D(net24),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _123_ (.D(net25),
    .GATE(net40),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q ));
 sky130_fd_sc_hd__dlxtp_1 _124_ (.D(net1),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q ));
 sky130_fd_sc_hd__dlxtp_1 _125_ (.D(net12),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q ));
 sky130_fd_sc_hd__dlxtp_1 _126_ (.D(net23),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q ));
 sky130_fd_sc_hd__dlxtp_1 _127_ (.D(net26),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q ));
 sky130_fd_sc_hd__dlxtp_1 _128_ (.D(net27),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q ));
 sky130_fd_sc_hd__dlxtp_1 _129_ (.D(net28),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q ));
 sky130_fd_sc_hd__dlxtp_1 _130_ (.D(net29),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q ));
 sky130_fd_sc_hd__dlxtp_1 _131_ (.D(net30),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q ));
 sky130_fd_sc_hd__dlxtp_1 _132_ (.D(net31),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q ));
 sky130_fd_sc_hd__dlxtp_1 _133_ (.D(net32),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q ));
 sky130_fd_sc_hd__dlxtp_1 _134_ (.D(net2),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q ));
 sky130_fd_sc_hd__dlxtp_1 _135_ (.D(net3),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q ));
 sky130_fd_sc_hd__dlxtp_1 _136_ (.D(net4),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q ));
 sky130_fd_sc_hd__dlxtp_1 _137_ (.D(net5),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q ));
 sky130_fd_sc_hd__dlxtp_1 _138_ (.D(net6),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q ));
 sky130_fd_sc_hd__dlxtp_1 _139_ (.D(net7),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q ));
 sky130_fd_sc_hd__dlxtp_1 _140_ (.D(net8),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q ));
 sky130_fd_sc_hd__dlxtp_1 _141_ (.D(net9),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q ));
 sky130_fd_sc_hd__dlxtp_1 _142_ (.D(net10),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q ));
 sky130_fd_sc_hd__dlxtp_1 _143_ (.D(net11),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q ));
 sky130_fd_sc_hd__dlxtp_1 _144_ (.D(net13),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q ));
 sky130_fd_sc_hd__dlxtp_1 _145_ (.D(net14),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q ));
 sky130_fd_sc_hd__dlxtp_1 _146_ (.D(net15),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q ));
 sky130_fd_sc_hd__dlxtp_1 _147_ (.D(net16),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q ));
 sky130_fd_sc_hd__dlxtp_1 _148_ (.D(net17),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q ));
 sky130_fd_sc_hd__dlxtp_1 _149_ (.D(net18),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sky130_fd_sc_hd__dlxtp_1 _150_ (.D(net19),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q ));
 sky130_fd_sc_hd__dlxtp_1 _151_ (.D(net20),
    .GATE(net43),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sky130_fd_sc_hd__dlxtp_1 _152_ (.D(net21),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q ));
 sky130_fd_sc_hd__dlxtp_1 _153_ (.D(net22),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sky130_fd_sc_hd__dlxtp_1 _154_ (.D(net24),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q ));
 sky130_fd_sc_hd__dlxtp_1 _155_ (.D(net25),
    .GATE(net42),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net128));
 sky130_fd_sc_hd__buf_1 _157_ (.A(net1),
    .X(net112));
 sky130_fd_sc_hd__buf_1 _158_ (.A(net12),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 _159_ (.A(net23),
    .X(net134));
 sky130_fd_sc_hd__buf_1 _160_ (.A(net26),
    .X(net137));
 sky130_fd_sc_hd__buf_1 _161_ (.A(net27),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _162_ (.A(net28),
    .X(net139));
 sky130_fd_sc_hd__buf_1 _163_ (.A(net29),
    .X(net140));
 sky130_fd_sc_hd__buf_1 _164_ (.A(net30),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 _165_ (.A(net31),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 _166_ (.A(net32),
    .X(net143));
 sky130_fd_sc_hd__buf_1 _167_ (.A(net2),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 _168_ (.A(net3),
    .X(net114));
 sky130_fd_sc_hd__buf_1 _169_ (.A(net4),
    .X(net115));
 sky130_fd_sc_hd__buf_1 _170_ (.A(net5),
    .X(net116));
 sky130_fd_sc_hd__buf_1 _171_ (.A(net6),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 _172_ (.A(net7),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 _173_ (.A(net8),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 _174_ (.A(net9),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 _175_ (.A(net10),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 _176_ (.A(net11),
    .X(net122));
 sky130_fd_sc_hd__buf_1 _177_ (.A(net13),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _178_ (.A(net14),
    .X(net125));
 sky130_fd_sc_hd__buf_1 _179_ (.A(net15),
    .X(net126));
 sky130_fd_sc_hd__buf_1 _180_ (.A(net16),
    .X(net127));
 sky130_fd_sc_hd__buf_1 _181_ (.A(net17),
    .X(net128));
 sky130_fd_sc_hd__buf_1 _182_ (.A(net18),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 _183_ (.A(net19),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 _184_ (.A(net20),
    .X(net131));
 sky130_fd_sc_hd__buf_1 _185_ (.A(net21),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _186_ (.A(net22),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 _187_ (.A(net24),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 _188_ (.A(net25),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _189_ (.A(net44),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(net41),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _191_ (.A(net37),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(FrameStrobe[3]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _193_ (.A(FrameStrobe[4]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(FrameStrobe[5]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _195_ (.A(FrameStrobe[6]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(FrameStrobe[7]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _197_ (.A(FrameStrobe[8]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _198_ (.A(FrameStrobe[9]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _199_ (.A(FrameStrobe[10]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(FrameStrobe[11]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _201_ (.A(FrameStrobe[12]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _202_ (.A(FrameStrobe[13]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _203_ (.A(FrameStrobe[14]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(FrameStrobe[15]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _205_ (.A(FrameStrobe[16]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _206_ (.A(FrameStrobe[17]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _207_ (.A(FrameStrobe[18]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _208_ (.A(FrameStrobe[19]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _209_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG0 ),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 _210_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG1 ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG2 ),
    .X(net182));
 sky130_fd_sc_hd__buf_1 _212_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG3 ),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _213_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG0 ),
    .X(net184));
 sky130_fd_sc_hd__buf_1 _214_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG1 ),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _215_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG2 ),
    .X(net186));
 sky130_fd_sc_hd__buf_1 _216_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG3 ),
    .X(net187));
 sky130_fd_sc_hd__buf_1 _217_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG4 ),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 _218_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG5 ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 _219_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG6 ),
    .X(net190));
 sky130_fd_sc_hd__buf_1 _220_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG7 ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 _221_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb0 ),
    .X(net192));
 sky130_fd_sc_hd__buf_1 _222_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb1 ),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 _223_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb2 ),
    .X(net194));
 sky130_fd_sc_hd__buf_1 _224_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb3 ),
    .X(net195));
 sky130_fd_sc_hd__buf_1 _225_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb4 ),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 _226_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb5 ),
    .X(net197));
 sky130_fd_sc_hd__buf_1 _227_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb6 ),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _228_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb7 ),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 _229_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG0 ),
    .X(net200));
 sky130_fd_sc_hd__buf_1 _230_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG1 ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 _231_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG2 ),
    .X(net208));
 sky130_fd_sc_hd__buf_1 _232_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG3 ),
    .X(net209));
 sky130_fd_sc_hd__buf_1 _233_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG4 ),
    .X(net210));
 sky130_fd_sc_hd__buf_1 _234_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG5 ),
    .X(net211));
 sky130_fd_sc_hd__buf_1 _235_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG6 ),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 _236_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG7 ),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 _237_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG8 ),
    .X(net214));
 sky130_fd_sc_hd__buf_1 _238_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG9 ),
    .X(net215));
 sky130_fd_sc_hd__buf_1 _239_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG10 ),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 _240_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG11 ),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 _241_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG12 ),
    .X(net203));
 sky130_fd_sc_hd__buf_1 _242_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG13 ),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 _243_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG14 ),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 _244_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG15 ),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG0 ),
    .X(net216));
 sky130_fd_sc_hd__buf_1 _246_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG1 ),
    .X(net223));
 sky130_fd_sc_hd__buf_1 _247_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG2 ),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 _248_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG3 ),
    .X(net225));
 sky130_fd_sc_hd__buf_1 _249_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG4 ),
    .X(net226));
 sky130_fd_sc_hd__buf_1 _250_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG5 ),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 _251_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG6 ),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 _252_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG7 ),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 _253_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG8 ),
    .X(net230));
 sky130_fd_sc_hd__buf_1 _254_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG9 ),
    .X(net231));
 sky130_fd_sc_hd__buf_1 _255_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG10 ),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 _256_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG11 ),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 _257_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG12 ),
    .X(net219));
 sky130_fd_sc_hd__buf_1 _258_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG13 ),
    .X(net220));
 sky130_fd_sc_hd__buf_1 _259_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG14 ),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 _260_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG15 ),
    .X(net222));
 sky130_fd_sc_hd__buf_2 _261_ (.A(UserCLK),
    .X(net232));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_121 ();
 sky130_fd_sc_hd__clkbuf_2 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__buf_2 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(FrameStrobe[2]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(FrameStrobe[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(FrameStrobe[0]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input1 (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(FrameData[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(FrameData[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(FrameData[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(FrameData[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(FrameData[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(FrameData[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(FrameData[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(FrameData[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(FrameData[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(FrameData[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(FrameData[2]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(FrameData[30]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(FrameData[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(FrameData[3]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(FrameData[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(FrameData[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(FrameData[6]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(FrameData[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(FrameData[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(FrameData[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(O_top0),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(O_top1),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(O_top10),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input36 (.A(O_top11),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input37 (.A(O_top12),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input38 (.A(O_top13),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(O_top14),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input40 (.A(O_top15),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(O_top2),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(O_top3),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(O_top4),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input44 (.A(O_top5),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(O_top6),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input46 (.A(O_top7),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(O_top8),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input48 (.A(O_top9),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input49 (.A(S1END[0]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(S1END[1]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(S1END[2]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(S1END[3]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input53 (.A(S2END[0]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input54 (.A(S2END[1]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input55 (.A(S2END[2]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input56 (.A(S2END[3]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(S2END[4]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input58 (.A(S2END[5]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input59 (.A(S2END[6]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input60 (.A(S2END[7]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(S2MID[0]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input62 (.A(S2MID[1]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input63 (.A(S2MID[2]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(S2MID[3]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(S2MID[4]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input66 (.A(S2MID[5]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input67 (.A(S2MID[6]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input68 (.A(S2MID[7]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(S4END[0]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input70 (.A(S4END[10]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(S4END[11]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input72 (.A(S4END[12]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input73 (.A(S4END[13]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(S4END[14]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input75 (.A(S4END[15]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input76 (.A(S4END[1]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input77 (.A(S4END[2]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(S4END[3]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input79 (.A(S4END[4]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input80 (.A(S4END[5]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(S4END[6]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input82 (.A(S4END[7]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input83 (.A(S4END[8]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input84 (.A(S4END[9]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input85 (.A(SS4END[0]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(SS4END[10]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input87 (.A(SS4END[11]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input88 (.A(SS4END[12]),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(SS4END[13]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(SS4END[14]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input91 (.A(SS4END[15]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input92 (.A(SS4END[1]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(SS4END[2]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input94 (.A(SS4END[3]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input95 (.A(SS4END[4]),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 input96 (.A(SS4END[5]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(SS4END[6]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input98 (.A(SS4END[7]),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input99 (.A(SS4END[8]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input100 (.A(SS4END[9]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 output101 (.A(net112),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net113),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net114),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net115),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net116),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net117),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net118),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net119),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net120),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net121),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net122),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net123),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net124),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net125),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net126),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net127),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net128),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net129),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net130),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net131),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net132),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net133),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net134),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net135),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net136),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net137),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net138),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net139),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net140),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net141),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net142),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net143),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net144),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net145),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net146),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net147),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net148),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net149),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net150),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net151),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net152),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net153),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net154),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net155),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net156),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net157),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net158),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net159),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net160),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net161),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net162),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net163),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net164),
    .X(I_top0));
 sky130_fd_sc_hd__buf_2 output154 (.A(net165),
    .X(I_top1));
 sky130_fd_sc_hd__buf_2 output155 (.A(net166),
    .X(I_top10));
 sky130_fd_sc_hd__buf_2 output156 (.A(net167),
    .X(I_top11));
 sky130_fd_sc_hd__buf_2 output157 (.A(net168),
    .X(I_top12));
 sky130_fd_sc_hd__buf_2 output158 (.A(net169),
    .X(I_top13));
 sky130_fd_sc_hd__buf_2 output159 (.A(net170),
    .X(I_top14));
 sky130_fd_sc_hd__buf_2 output160 (.A(net171),
    .X(I_top15));
 sky130_fd_sc_hd__buf_2 output161 (.A(net172),
    .X(I_top2));
 sky130_fd_sc_hd__buf_2 output162 (.A(net173),
    .X(I_top3));
 sky130_fd_sc_hd__buf_2 output163 (.A(net174),
    .X(I_top4));
 sky130_fd_sc_hd__buf_2 output164 (.A(net175),
    .X(I_top5));
 sky130_fd_sc_hd__buf_2 output165 (.A(net176),
    .X(I_top6));
 sky130_fd_sc_hd__buf_2 output166 (.A(net177),
    .X(I_top7));
 sky130_fd_sc_hd__buf_2 output167 (.A(net178),
    .X(I_top8));
 sky130_fd_sc_hd__buf_2 output168 (.A(net179),
    .X(I_top9));
 sky130_fd_sc_hd__buf_2 output169 (.A(net180),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net181),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net182),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net183),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net184),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net185),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net186),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net187),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net188),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net189),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net190),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net191),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net192),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net193),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net194),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net195),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net196),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net197),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net198),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net199),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net200),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net201),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net202),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net203),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net204),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net205),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net206),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net207),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net208),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net209),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net210),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net211),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net212),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net213),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net214),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net215),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net216),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net217),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net218),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net219),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net220),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net221),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net222),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net223),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net224),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net225),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net226),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net227),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net228),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net229),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net230),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net231),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__buf_1 output221 (.A(net232),
    .X(UserCLKo));
 sky130_fd_sc_hd__conb_1 S_CPU_IF_222 (.LO(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameStrobe[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net195));
 sky130_fd_sc_hd__fill_1 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_409 ();
 assign Co = net233;
endmodule
