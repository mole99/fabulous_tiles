magic
tech sky130A
magscale 1 2
timestamp 1739717529
<< viali >>
rect 3065 8585 3099 8619
rect 3433 8585 3467 8619
rect 6745 8585 6779 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15301 8585 15335 8619
rect 16037 8585 16071 8619
rect 16313 8585 16347 8619
rect 17693 8585 17727 8619
rect 17969 8585 18003 8619
rect 42165 8585 42199 8619
rect 43453 8585 43487 8619
rect 10885 8517 10919 8551
rect 22293 8517 22327 8551
rect 26525 8517 26559 8551
rect 29009 8517 29043 8551
rect 29193 8517 29227 8551
rect 32229 8517 32263 8551
rect 34345 8517 34379 8551
rect 1409 8449 1443 8483
rect 2881 8449 2915 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 5825 8449 5859 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8033 8449 8067 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9321 8449 9355 8483
rect 9413 8449 9447 8483
rect 9781 8449 9815 8483
rect 10425 8449 10459 8483
rect 11805 8449 11839 8483
rect 13185 8449 13219 8483
rect 14105 8449 14139 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15117 8449 15151 8483
rect 15761 8449 15795 8483
rect 15853 8449 15887 8483
rect 16497 8449 16531 8483
rect 17141 8449 17175 8483
rect 17509 8449 17543 8483
rect 18153 8449 18187 8483
rect 18797 8449 18831 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 21649 8449 21683 8483
rect 22017 8449 22051 8483
rect 22477 8449 22511 8483
rect 23397 8449 23431 8483
rect 23673 8449 23707 8483
rect 24685 8449 24719 8483
rect 25513 8449 25547 8483
rect 26985 8449 27019 8483
rect 27261 8449 27295 8483
rect 28181 8449 28215 8483
rect 30021 8449 30055 8483
rect 30849 8449 30883 8483
rect 31953 8449 31987 8483
rect 33425 8449 33459 8483
rect 33885 8449 33919 8483
rect 34161 8449 34195 8483
rect 34713 8449 34747 8483
rect 35633 8449 35667 8483
rect 35909 8449 35943 8483
rect 36829 8449 36863 8483
rect 36921 8449 36955 8483
rect 37289 8449 37323 8483
rect 38485 8449 38519 8483
rect 38853 8449 38887 8483
rect 38945 8449 38979 8483
rect 39589 8449 39623 8483
rect 40141 8449 40175 8483
rect 40509 8449 40543 8483
rect 40877 8449 40911 8483
rect 41245 8449 41279 8483
rect 41613 8449 41647 8483
rect 41981 8449 42015 8483
rect 42809 8449 42843 8483
rect 42901 8449 42935 8483
rect 43269 8449 43303 8483
rect 1685 8381 1719 8415
rect 10701 8381 10735 8415
rect 10793 8381 10827 8415
rect 11529 8381 11563 8415
rect 12909 8381 12943 8415
rect 16957 8381 16991 8415
rect 19073 8381 19107 8415
rect 20177 8381 20211 8415
rect 21373 8381 21407 8415
rect 22753 8381 22787 8415
rect 24409 8381 24443 8415
rect 25789 8381 25823 8415
rect 26709 8381 26743 8415
rect 27905 8381 27939 8415
rect 29745 8381 29779 8415
rect 33701 8381 33735 8415
rect 34989 8381 35023 8415
rect 37565 8381 37599 8415
rect 2697 8313 2731 8347
rect 4537 8313 4571 8347
rect 6009 8313 6043 8347
rect 7113 8313 7147 8347
rect 7481 8313 7515 8347
rect 8217 8313 8251 8347
rect 8585 8313 8619 8347
rect 9597 8313 9631 8347
rect 9965 8313 9999 8347
rect 10241 8313 10275 8347
rect 12541 8313 12575 8347
rect 14289 8313 14323 8347
rect 15577 8313 15611 8347
rect 17325 8313 17359 8347
rect 19441 8313 19475 8347
rect 21833 8313 21867 8347
rect 28917 8313 28951 8347
rect 32689 8313 32723 8347
rect 34069 8313 34103 8347
rect 36645 8313 36679 8347
rect 38301 8313 38335 8347
rect 38669 8313 38703 8347
rect 39129 8313 39163 8347
rect 39405 8313 39439 8347
rect 39957 8313 39991 8347
rect 41429 8313 41463 8347
rect 43085 8313 43119 8347
rect 4169 8245 4203 8279
rect 4905 8245 4939 8279
rect 5273 8245 5307 8279
rect 5641 8245 5675 8279
rect 7849 8245 7883 8279
rect 11253 8245 11287 8279
rect 13921 8245 13955 8279
rect 22201 8245 22235 8279
rect 25421 8245 25455 8279
rect 30757 8245 30791 8279
rect 31079 8245 31113 8279
rect 31769 8245 31803 8279
rect 32321 8245 32355 8279
rect 37105 8245 37139 8279
rect 40325 8245 40359 8279
rect 40693 8245 40727 8279
rect 41061 8245 41095 8279
rect 3065 8041 3099 8075
rect 3893 8041 3927 8075
rect 6101 8041 6135 8075
rect 6469 8041 6503 8075
rect 8217 8041 8251 8075
rect 8585 8041 8619 8075
rect 15301 8041 15335 8075
rect 18889 8041 18923 8075
rect 19441 8041 19475 8075
rect 19625 8041 19659 8075
rect 22109 8041 22143 8075
rect 34345 8041 34379 8075
rect 34805 8041 34839 8075
rect 37565 8041 37599 8075
rect 37933 8041 37967 8075
rect 38669 8041 38703 8075
rect 39405 8041 39439 8075
rect 41061 8041 41095 8075
rect 41521 8041 41555 8075
rect 42717 8041 42751 8075
rect 3617 7973 3651 8007
rect 5181 7973 5215 8007
rect 10609 7973 10643 8007
rect 13369 7973 13403 8007
rect 16589 7973 16623 8007
rect 17877 7973 17911 8007
rect 22201 7973 22235 8007
rect 25697 7973 25731 8007
rect 30665 7973 30699 8007
rect 31953 7973 31987 8007
rect 35173 7973 35207 8007
rect 38209 7973 38243 8007
rect 39129 7973 39163 8007
rect 41981 7973 42015 8007
rect 42349 7973 42383 8007
rect 1685 7905 1719 7939
rect 5549 7905 5583 7939
rect 6745 7905 6779 7939
rect 8953 7905 8987 7939
rect 11989 7905 12023 7939
rect 15577 7905 15611 7939
rect 21005 7905 21039 7939
rect 23305 7905 23339 7939
rect 26090 7905 26124 7939
rect 26985 7905 27019 7939
rect 30021 7905 30055 7939
rect 30941 7905 30975 7939
rect 31217 7905 31251 7939
rect 32965 7905 32999 7939
rect 35541 7905 35575 7939
rect 36185 7905 36219 7939
rect 1501 7837 1535 7871
rect 2053 7837 2087 7871
rect 2605 7837 2639 7871
rect 2973 7837 3007 7871
rect 4077 7837 4111 7871
rect 4169 7837 4203 7871
rect 4445 7837 4479 7871
rect 6285 7837 6319 7871
rect 6653 7837 6687 7871
rect 7008 7837 7042 7871
rect 8401 7837 8435 7871
rect 8769 7837 8803 7871
rect 9229 7837 9263 7871
rect 11897 7837 11931 7871
rect 12256 7837 12290 7871
rect 13921 7837 13955 7871
rect 14841 7837 14875 7871
rect 15117 7837 15151 7871
rect 15485 7837 15519 7871
rect 15840 7837 15874 7871
rect 17325 7837 17359 7871
rect 17463 7837 17497 7871
rect 17601 7837 17635 7871
rect 18337 7837 18371 7871
rect 18521 7837 18555 7871
rect 19073 7837 19107 7871
rect 19257 7837 19291 7871
rect 19809 7837 19843 7871
rect 20637 7837 20671 7871
rect 20913 7837 20947 7871
rect 21281 7837 21315 7871
rect 21925 7837 21959 7871
rect 22937 7837 22971 7871
rect 23213 7837 23247 7871
rect 23581 7837 23615 7871
rect 24777 7837 24811 7871
rect 25053 7837 25087 7871
rect 25237 7837 25271 7871
rect 25973 7837 26007 7871
rect 26249 7837 26283 7871
rect 27261 7837 27295 7871
rect 27905 7837 27939 7871
rect 28181 7837 28215 7871
rect 29745 7837 29779 7871
rect 30205 7837 30239 7871
rect 31058 7837 31092 7871
rect 32689 7837 32723 7871
rect 33057 7837 33091 7871
rect 33333 7837 33367 7871
rect 34529 7837 34563 7871
rect 34989 7837 35023 7871
rect 35357 7837 35391 7871
rect 35725 7837 35759 7871
rect 36461 7837 36495 7871
rect 36578 7837 36612 7871
rect 36737 7837 36771 7871
rect 37749 7837 37783 7871
rect 38117 7837 38151 7871
rect 38853 7837 38887 7871
rect 38945 7837 38979 7871
rect 39589 7837 39623 7871
rect 39865 7837 39899 7871
rect 40141 7837 40175 7871
rect 41245 7837 41279 7871
rect 41705 7837 41739 7871
rect 41797 7837 41831 7871
rect 42165 7837 42199 7871
rect 42533 7837 42567 7871
rect 42901 7837 42935 7871
rect 43269 7837 43303 7871
rect 2237 7769 2271 7803
rect 2421 7769 2455 7803
rect 2789 7769 2823 7803
rect 3433 7769 3467 7803
rect 5365 7769 5399 7803
rect 5733 7769 5767 7803
rect 24501 7769 24535 7803
rect 24685 7769 24719 7803
rect 26893 7769 26927 7803
rect 29193 7769 29227 7803
rect 37381 7769 37415 7803
rect 38393 7769 38427 7803
rect 1869 7701 1903 7735
rect 5825 7701 5859 7735
rect 7757 7701 7791 7735
rect 9965 7701 9999 7735
rect 13737 7701 13771 7735
rect 14105 7701 14139 7735
rect 16681 7701 16715 7735
rect 19901 7701 19935 7735
rect 24961 7701 24995 7735
rect 28917 7701 28951 7735
rect 29101 7701 29135 7735
rect 29561 7701 29595 7735
rect 31861 7701 31895 7735
rect 34069 7701 34103 7735
rect 40877 7701 40911 7735
rect 43085 7701 43119 7735
rect 43453 7701 43487 7735
rect 6745 7497 6779 7531
rect 7113 7497 7147 7531
rect 7941 7497 7975 7531
rect 8309 7497 8343 7531
rect 9781 7497 9815 7531
rect 11069 7497 11103 7531
rect 11161 7497 11195 7531
rect 16313 7497 16347 7531
rect 17693 7497 17727 7531
rect 19165 7497 19199 7531
rect 19717 7497 19751 7531
rect 23857 7497 23891 7531
rect 25145 7497 25179 7531
rect 31769 7497 31803 7531
rect 35357 7497 35391 7531
rect 36461 7497 36495 7531
rect 36921 7497 36955 7531
rect 40417 7497 40451 7531
rect 40693 7497 40727 7531
rect 42073 7497 42107 7531
rect 42717 7497 42751 7531
rect 43085 7497 43119 7531
rect 2789 7429 2823 7463
rect 3157 7429 3191 7463
rect 3341 7429 3375 7463
rect 26617 7429 26651 7463
rect 26801 7429 26835 7463
rect 28089 7429 28123 7463
rect 35081 7429 35115 7463
rect 40233 7429 40267 7463
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 4537 7361 4571 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 6193 7361 6227 7395
rect 6929 7361 6963 7395
rect 7297 7361 7331 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 8125 7361 8159 7395
rect 8769 7361 8803 7395
rect 9965 7361 9999 7395
rect 10057 7361 10091 7395
rect 10333 7361 10367 7395
rect 11345 7361 11379 7395
rect 13277 7361 13311 7395
rect 13645 7361 13679 7395
rect 13737 7361 13771 7395
rect 14013 7361 14047 7395
rect 15393 7361 15427 7395
rect 16497 7361 16531 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 18061 7361 18095 7395
rect 19257 7361 19291 7395
rect 20499 7361 20533 7395
rect 22293 7361 22327 7395
rect 22385 7361 22419 7395
rect 23297 7361 23331 7395
rect 23581 7361 23615 7395
rect 24032 7361 24066 7395
rect 24133 7361 24167 7395
rect 24409 7361 24443 7395
rect 25513 7361 25547 7395
rect 26985 7361 27019 7395
rect 29561 7361 29595 7395
rect 30389 7361 30423 7395
rect 31493 7361 31527 7395
rect 31585 7361 31619 7395
rect 32137 7361 32171 7395
rect 32413 7361 32447 7395
rect 35173 7361 35207 7395
rect 35725 7361 35759 7395
rect 36829 7361 36863 7395
rect 37105 7361 37139 7395
rect 37565 7361 37599 7395
rect 39313 7361 39347 7395
rect 39451 7361 39485 7395
rect 40601 7361 40635 7395
rect 40877 7361 40911 7395
rect 42257 7361 42291 7395
rect 42533 7361 42567 7395
rect 42901 7361 42935 7395
rect 43269 7361 43303 7395
rect 1409 7293 1443 7327
rect 1685 7293 1719 7327
rect 4261 7293 4295 7327
rect 8493 7293 8527 7327
rect 11529 7293 11563 7327
rect 15117 7293 15151 7327
rect 17785 7293 17819 7327
rect 19073 7293 19107 7327
rect 20361 7293 20395 7327
rect 20637 7293 20671 7327
rect 21373 7293 21407 7327
rect 21557 7293 21591 7327
rect 22661 7293 22695 7327
rect 25237 7293 25271 7327
rect 28365 7293 28399 7327
rect 28549 7293 28583 7327
rect 29009 7293 29043 7327
rect 29285 7293 29319 7327
rect 29423 7293 29457 7327
rect 30665 7293 30699 7327
rect 33241 7293 33275 7327
rect 33425 7293 33459 7327
rect 33885 7293 33919 7327
rect 34161 7293 34195 7327
rect 34278 7293 34312 7327
rect 34437 7293 34471 7327
rect 35449 7293 35483 7327
rect 37289 7293 37323 7327
rect 38393 7293 38427 7327
rect 38577 7293 38611 7327
rect 39589 7293 39623 7327
rect 7481 7225 7515 7259
rect 20913 7225 20947 7259
rect 22109 7225 22143 7259
rect 23489 7225 23523 7259
rect 31309 7225 31343 7259
rect 36645 7225 36679 7259
rect 39037 7225 39071 7259
rect 2881 7157 2915 7191
rect 5273 7157 5307 7191
rect 9505 7157 9539 7191
rect 13461 7157 13495 7191
rect 14749 7157 14783 7191
rect 16129 7157 16163 7191
rect 18797 7157 18831 7191
rect 19625 7157 19659 7191
rect 23765 7157 23799 7191
rect 26249 7157 26283 7191
rect 27215 7157 27249 7191
rect 27997 7157 28031 7191
rect 30205 7157 30239 7191
rect 33149 7157 33183 7191
rect 38301 7157 38335 7191
rect 43453 7157 43487 7191
rect 13461 6953 13495 6987
rect 38853 6953 38887 6987
rect 42349 6953 42383 6987
rect 3985 6885 4019 6919
rect 5089 6885 5123 6919
rect 25421 6885 25455 6919
rect 28549 6885 28583 6919
rect 28641 6885 28675 6919
rect 37749 6885 37783 6919
rect 39405 6885 39439 6919
rect 39681 6885 39715 6919
rect 1409 6817 1443 6851
rect 2973 6817 3007 6851
rect 4445 6817 4479 6851
rect 5365 6817 5399 6851
rect 5503 6817 5537 6851
rect 5641 6817 5675 6851
rect 7757 6817 7791 6851
rect 9848 6817 9882 6851
rect 10241 6817 10275 6851
rect 10977 6817 11011 6851
rect 17693 6817 17727 6851
rect 20453 6817 20487 6851
rect 20913 6817 20947 6851
rect 22477 6817 22511 6851
rect 24409 6817 24443 6851
rect 26157 6817 26191 6851
rect 27537 6817 27571 6851
rect 32597 6817 32631 6851
rect 33701 6817 33735 6851
rect 34713 6817 34747 6851
rect 35909 6817 35943 6851
rect 36093 6817 36127 6851
rect 36553 6817 36587 6851
rect 36829 6817 36863 6851
rect 36967 6817 37001 6851
rect 37841 6817 37875 6851
rect 1685 6749 1719 6783
rect 2329 6749 2363 6783
rect 2789 6749 2823 6783
rect 3801 6749 3835 6783
rect 4629 6749 4663 6783
rect 6469 6749 6503 6783
rect 6745 6749 6779 6783
rect 8033 6749 8067 6783
rect 9689 6749 9723 6783
rect 9965 6749 9999 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 11253 6749 11287 6783
rect 12173 6749 12207 6783
rect 13921 6749 13955 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 14933 6749 14967 6783
rect 16497 6749 16531 6783
rect 16773 6749 16807 6783
rect 17417 6749 17451 6783
rect 17785 6749 17819 6783
rect 18061 6749 18095 6783
rect 19073 6749 19107 6783
rect 19901 6749 19935 6783
rect 20039 6749 20073 6783
rect 20177 6749 20211 6783
rect 21097 6749 21131 6783
rect 21925 6749 21959 6783
rect 22201 6749 22235 6783
rect 22753 6749 22787 6783
rect 24685 6749 24719 6783
rect 25513 6749 25547 6783
rect 25697 6749 25731 6783
rect 26433 6749 26467 6783
rect 26550 6749 26584 6783
rect 26709 6749 26743 6783
rect 27813 6749 27847 6783
rect 28825 6749 28859 6783
rect 28917 6749 28951 6783
rect 29193 6749 29227 6783
rect 29745 6749 29779 6783
rect 30021 6749 30055 6783
rect 30113 6749 30147 6783
rect 30573 6749 30607 6783
rect 30665 6749 30699 6783
rect 30941 6749 30975 6783
rect 31953 6749 31987 6783
rect 32229 6749 32263 6783
rect 32505 6749 32539 6783
rect 32873 6749 32907 6783
rect 33977 6749 34011 6783
rect 34989 6749 35023 6783
rect 35817 6765 35851 6799
rect 37105 6749 37139 6783
rect 38117 6749 38151 6783
rect 39129 6749 39163 6783
rect 39221 6749 39255 6783
rect 39497 6749 39531 6783
rect 42533 6749 42567 6783
rect 42717 6749 42751 6783
rect 43177 6749 43211 6783
rect 43269 6749 43303 6783
rect 3157 6681 3191 6715
rect 3341 6681 3375 6715
rect 27353 6681 27387 6715
rect 43085 6681 43119 6715
rect 2513 6613 2547 6647
rect 6285 6613 6319 6647
rect 7481 6613 7515 6647
rect 8769 6613 8803 6647
rect 9045 6613 9079 6647
rect 11989 6613 12023 6647
rect 14381 6613 14415 6647
rect 15669 6613 15703 6647
rect 15761 6613 15795 6647
rect 17233 6613 17267 6647
rect 18797 6613 18831 6647
rect 18889 6613 18923 6647
rect 19257 6613 19291 6647
rect 21189 6613 21223 6647
rect 23489 6613 23523 6647
rect 29101 6613 29135 6647
rect 29377 6613 29411 6647
rect 29561 6613 29595 6647
rect 29837 6613 29871 6647
rect 30297 6613 30331 6647
rect 30389 6613 30423 6647
rect 31677 6613 31711 6647
rect 31769 6613 31803 6647
rect 32045 6613 32079 6647
rect 32321 6613 32355 6647
rect 33609 6613 33643 6647
rect 35633 6613 35667 6647
rect 38945 6613 38979 6647
rect 42901 6613 42935 6647
rect 43453 6613 43487 6647
rect 6561 6409 6595 6443
rect 6745 6409 6779 6443
rect 9321 6409 9355 6443
rect 11989 6409 12023 6443
rect 13461 6409 13495 6443
rect 13829 6409 13863 6443
rect 19257 6409 19291 6443
rect 23765 6409 23799 6443
rect 31677 6409 31711 6443
rect 36921 6409 36955 6443
rect 40509 6409 40543 6443
rect 42625 6409 42659 6443
rect 43453 6409 43487 6443
rect 14289 6341 14323 6375
rect 18797 6341 18831 6375
rect 24041 6341 24075 6375
rect 24409 6341 24443 6375
rect 24593 6341 24627 6375
rect 32413 6341 32447 6375
rect 1501 6273 1535 6307
rect 1777 6273 1811 6307
rect 3642 6273 3676 6307
rect 3801 6273 3835 6307
rect 4445 6273 4479 6307
rect 4537 6273 4571 6307
rect 5181 6273 5215 6307
rect 5457 6273 5491 6307
rect 6377 6273 6411 6307
rect 6929 6273 6963 6307
rect 7665 6273 7699 6307
rect 7941 6273 7975 6307
rect 8677 6273 8711 6307
rect 9045 6273 9079 6307
rect 9137 6273 9171 6307
rect 9781 6273 9815 6307
rect 11089 6273 11123 6307
rect 13277 6273 13311 6307
rect 13645 6273 13679 6307
rect 14013 6273 14047 6307
rect 17601 6273 17635 6307
rect 17877 6273 17911 6307
rect 19441 6273 19475 6307
rect 19717 6273 19751 6307
rect 19809 6273 19843 6307
rect 20729 6273 20763 6307
rect 21833 6273 21867 6307
rect 22109 6273 22143 6307
rect 23489 6273 23523 6307
rect 23949 6273 23983 6307
rect 24133 6273 24167 6307
rect 24317 6273 24351 6307
rect 24777 6273 24811 6307
rect 25421 6273 25455 6307
rect 26249 6273 26283 6307
rect 26617 6273 26651 6307
rect 27721 6273 27755 6307
rect 27997 6273 28031 6307
rect 28181 6273 28215 6307
rect 28365 6273 28399 6307
rect 29377 6273 29411 6307
rect 30389 6273 30423 6307
rect 31217 6273 31251 6307
rect 31493 6273 31527 6307
rect 31769 6273 31803 6307
rect 32229 6273 32263 6307
rect 32689 6273 32723 6307
rect 32873 6273 32907 6307
rect 35541 6273 35575 6307
rect 35817 6273 35851 6307
rect 36185 6273 36219 6307
rect 37749 6273 37783 6307
rect 38577 6273 38611 6307
rect 38761 6273 38795 6307
rect 39614 6273 39648 6307
rect 40417 6273 40451 6307
rect 40693 6273 40727 6307
rect 42809 6273 42843 6307
rect 42901 6273 42935 6307
rect 43269 6273 43303 6307
rect 2605 6205 2639 6239
rect 2789 6205 2823 6239
rect 3525 6205 3559 6239
rect 7803 6205 7837 6239
rect 8217 6205 8251 6239
rect 8861 6205 8895 6239
rect 11345 6205 11379 6239
rect 19993 6205 20027 6239
rect 20867 6205 20901 6239
rect 21005 6205 21039 6239
rect 23581 6205 23615 6239
rect 25145 6205 25179 6239
rect 29101 6205 29135 6239
rect 29239 6205 29273 6239
rect 30113 6205 30147 6239
rect 33057 6205 33091 6239
rect 33517 6205 33551 6239
rect 33793 6205 33827 6239
rect 33910 6205 33944 6239
rect 34069 6205 34103 6239
rect 35909 6205 35943 6239
rect 37473 6205 37507 6239
rect 39497 6205 39531 6239
rect 39773 6205 39807 6239
rect 3249 6137 3283 6171
rect 4721 6137 4755 6171
rect 15577 6137 15611 6171
rect 18981 6137 19015 6171
rect 20453 6137 20487 6171
rect 26157 6137 26191 6171
rect 26433 6137 26467 6171
rect 28825 6137 28859 6171
rect 31953 6137 31987 6171
rect 32505 6137 32539 6171
rect 39221 6137 39255 6171
rect 2513 6069 2547 6103
rect 6193 6069 6227 6103
rect 7021 6069 7055 6103
rect 9045 6069 9079 6103
rect 9597 6069 9631 6103
rect 9965 6069 9999 6103
rect 18613 6069 18647 6103
rect 19533 6069 19567 6103
rect 21649 6069 21683 6103
rect 22017 6069 22051 6103
rect 22293 6069 22327 6103
rect 26709 6069 26743 6103
rect 26985 6069 27019 6103
rect 30021 6069 30055 6103
rect 31125 6069 31159 6103
rect 31401 6069 31435 6103
rect 32321 6069 32355 6103
rect 34713 6069 34747 6103
rect 34805 6069 34839 6103
rect 38485 6069 38519 6103
rect 43085 6069 43119 6103
rect 3065 5865 3099 5899
rect 4445 5865 4479 5899
rect 7941 5865 7975 5899
rect 12909 5865 12943 5899
rect 13369 5865 13403 5899
rect 13645 5865 13679 5899
rect 15117 5865 15151 5899
rect 18889 5865 18923 5899
rect 19257 5865 19291 5899
rect 23581 5865 23615 5899
rect 23949 5865 23983 5899
rect 24409 5865 24443 5899
rect 33701 5865 33735 5899
rect 34345 5865 34379 5899
rect 34713 5865 34747 5899
rect 36829 5865 36863 5899
rect 37381 5865 37415 5899
rect 38117 5865 38151 5899
rect 39221 5865 39255 5899
rect 3433 5797 3467 5831
rect 6377 5797 6411 5831
rect 7849 5797 7883 5831
rect 10149 5797 10183 5831
rect 12081 5797 12115 5831
rect 14841 5797 14875 5831
rect 16313 5797 16347 5831
rect 18429 5797 18463 5831
rect 20453 5797 20487 5831
rect 31401 5797 31435 5831
rect 33977 5797 34011 5831
rect 43453 5797 43487 5831
rect 2053 5729 2087 5763
rect 4629 5729 4663 5763
rect 5733 5729 5767 5763
rect 5917 5729 5951 5763
rect 6791 5729 6825 5763
rect 9597 5729 9631 5763
rect 9873 5729 9907 5763
rect 10793 5729 10827 5763
rect 11688 5729 11722 5763
rect 12541 5729 12575 5763
rect 12725 5729 12759 5763
rect 13553 5729 13587 5763
rect 14289 5729 14323 5763
rect 16037 5729 16071 5763
rect 16957 5729 16991 5763
rect 18521 5729 18555 5763
rect 19993 5729 20027 5763
rect 21649 5729 21683 5763
rect 22109 5729 22143 5763
rect 23489 5729 23523 5763
rect 24961 5729 24995 5763
rect 25329 5729 25363 5763
rect 26065 5729 26099 5763
rect 26249 5729 26283 5763
rect 26709 5729 26743 5763
rect 27123 5729 27157 5763
rect 27997 5729 28031 5763
rect 30757 5729 30791 5763
rect 31953 5729 31987 5763
rect 32689 5729 32723 5763
rect 38209 5729 38243 5763
rect 1501 5661 1535 5695
rect 2329 5661 2363 5695
rect 4353 5661 4387 5695
rect 4905 5661 4939 5695
rect 6653 5661 6687 5695
rect 6929 5661 6963 5695
rect 7573 5661 7607 5695
rect 7665 5661 7699 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 8953 5661 8987 5695
rect 9756 5661 9790 5695
rect 10609 5661 10643 5695
rect 11529 5661 11563 5695
rect 11805 5661 11839 5695
rect 13093 5661 13127 5695
rect 13185 5661 13219 5695
rect 14473 5661 14507 5695
rect 15761 5661 15795 5695
rect 15920 5661 15954 5695
rect 16773 5661 16807 5695
rect 17417 5661 17451 5695
rect 17693 5661 17727 5695
rect 19441 5661 19475 5695
rect 19717 5661 19751 5695
rect 19809 5661 19843 5695
rect 20729 5661 20763 5695
rect 20867 5661 20901 5695
rect 21005 5661 21039 5695
rect 21925 5661 21959 5695
rect 22201 5661 22235 5695
rect 23765 5661 23799 5695
rect 24869 5661 24903 5695
rect 25237 5661 25271 5695
rect 27003 5661 27037 5695
rect 27261 5661 27295 5695
rect 28273 5661 28307 5695
rect 29745 5661 29779 5695
rect 30941 5661 30975 5695
rect 31677 5661 31711 5695
rect 31794 5661 31828 5695
rect 32965 5661 32999 5695
rect 33793 5661 33827 5695
rect 34529 5661 34563 5695
rect 35449 5661 35483 5695
rect 35725 5661 35759 5695
rect 35817 5661 35851 5695
rect 36093 5661 36127 5695
rect 37565 5661 37599 5695
rect 37933 5661 37967 5695
rect 38485 5661 38519 5695
rect 39313 5661 39347 5695
rect 42901 5661 42935 5695
rect 43269 5661 43303 5695
rect 3249 5593 3283 5627
rect 3893 5593 3927 5627
rect 4077 5593 4111 5627
rect 8585 5593 8619 5627
rect 13737 5593 13771 5627
rect 14381 5593 14415 5627
rect 18889 5593 18923 5627
rect 1593 5525 1627 5559
rect 5641 5525 5675 5559
rect 8217 5525 8251 5559
rect 8677 5525 8711 5559
rect 10885 5525 10919 5559
rect 18429 5525 18463 5559
rect 19073 5525 19107 5559
rect 19533 5525 19567 5559
rect 21741 5525 21775 5559
rect 24777 5525 24811 5559
rect 27905 5525 27939 5559
rect 29561 5525 29595 5559
rect 32597 5525 32631 5559
rect 39497 5525 39531 5559
rect 43085 5525 43119 5559
rect 1593 5321 1627 5355
rect 7389 5321 7423 5355
rect 10057 5321 10091 5355
rect 11345 5321 11379 5355
rect 13829 5321 13863 5355
rect 18245 5321 18279 5355
rect 19625 5321 19659 5355
rect 21649 5321 21683 5355
rect 22523 5321 22557 5355
rect 24777 5321 24811 5355
rect 30757 5321 30791 5355
rect 31769 5321 31803 5355
rect 43453 5321 43487 5355
rect 14197 5253 14231 5287
rect 18337 5253 18371 5287
rect 19073 5253 19107 5287
rect 25605 5253 25639 5287
rect 25973 5253 26007 5287
rect 1409 5185 1443 5219
rect 2421 5185 2455 5219
rect 2789 5185 2823 5219
rect 3709 5185 3743 5219
rect 3847 5185 3881 5219
rect 4813 5185 4847 5219
rect 5089 5185 5123 5219
rect 6377 5185 6411 5219
rect 6653 5185 6687 5219
rect 7481 5185 7515 5219
rect 8125 5185 8159 5219
rect 9137 5185 9171 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 10609 5185 10643 5219
rect 11529 5185 11563 5219
rect 12725 5185 12759 5219
rect 14013 5185 14047 5219
rect 14381 5185 14415 5219
rect 15853 5185 15887 5219
rect 16681 5185 16715 5219
rect 16957 5185 16991 5219
rect 18061 5185 18095 5219
rect 18429 5185 18463 5219
rect 18521 5185 18555 5219
rect 18613 5185 18647 5219
rect 18797 5185 18831 5219
rect 19349 5185 19383 5219
rect 19533 5185 19567 5219
rect 22017 5185 22051 5219
rect 22109 5185 22143 5219
rect 22201 5185 22235 5219
rect 22385 5185 22419 5219
rect 22594 5185 22628 5219
rect 22937 5185 22971 5219
rect 23974 5185 24008 5219
rect 24133 5185 24167 5219
rect 25697 5185 25731 5219
rect 27721 5185 27755 5219
rect 28273 5185 28307 5219
rect 29745 5185 29779 5219
rect 30021 5185 30055 5219
rect 30665 5185 30699 5219
rect 30941 5185 30975 5219
rect 31953 5185 31987 5219
rect 32413 5185 32447 5219
rect 33425 5185 33459 5219
rect 33701 5185 33735 5219
rect 34621 5185 34655 5219
rect 34897 5185 34931 5219
rect 35541 5185 35575 5219
rect 35817 5185 35851 5219
rect 36093 5185 36127 5219
rect 36369 5185 36403 5219
rect 37565 5185 37599 5219
rect 39221 5185 39255 5219
rect 42901 5185 42935 5219
rect 43269 5185 43303 5219
rect 2697 5117 2731 5151
rect 2973 5117 3007 5151
rect 3985 5117 4019 5151
rect 7941 5117 7975 5151
rect 8861 5117 8895 5151
rect 8999 5117 9033 5151
rect 11713 5117 11747 5151
rect 12449 5117 12483 5151
rect 12587 5117 12621 5151
rect 14657 5117 14691 5151
rect 14841 5117 14875 5151
rect 15577 5117 15611 5151
rect 15715 5117 15749 5151
rect 17969 5117 18003 5151
rect 18889 5117 18923 5151
rect 19073 5117 19107 5151
rect 19809 5117 19843 5151
rect 19993 5117 20027 5151
rect 20453 5117 20487 5151
rect 20729 5117 20763 5151
rect 20867 5117 20901 5151
rect 21005 5117 21039 5151
rect 23121 5117 23155 5151
rect 23857 5117 23891 5151
rect 25329 5117 25363 5151
rect 27997 5117 28031 5151
rect 28825 5117 28859 5151
rect 29009 5117 29043 5151
rect 29862 5117 29896 5151
rect 32137 5117 32171 5151
rect 33885 5117 33919 5151
rect 34345 5117 34379 5151
rect 34759 5117 34793 5151
rect 37289 5117 37323 5151
rect 39497 5117 39531 5151
rect 3433 5049 3467 5083
rect 7665 5049 7699 5083
rect 8585 5049 8619 5083
rect 12173 5049 12207 5083
rect 13645 5049 13679 5083
rect 15301 5049 15335 5083
rect 17693 5049 17727 5083
rect 18981 5049 19015 5083
rect 23581 5049 23615 5083
rect 26341 5049 26375 5083
rect 29469 5049 29503 5083
rect 38485 5049 38519 5083
rect 1685 4981 1719 5015
rect 4629 4981 4663 5015
rect 5825 4981 5859 5015
rect 9781 4981 9815 5015
rect 13369 4981 13403 5015
rect 14289 4981 14323 5015
rect 16497 4981 16531 5015
rect 17785 4981 17819 5015
rect 19257 4981 19291 5015
rect 21833 4981 21867 5015
rect 25329 4981 25363 5015
rect 25421 4981 25455 5015
rect 25789 4981 25823 5015
rect 25973 4981 26007 5015
rect 26985 4981 27019 5015
rect 28089 4981 28123 5015
rect 33149 4981 33183 5015
rect 33241 4981 33275 5015
rect 35633 4981 35667 5015
rect 37105 4981 37139 5015
rect 38301 4981 38335 5015
rect 43085 4981 43119 5015
rect 3433 4777 3467 4811
rect 7113 4777 7147 4811
rect 8769 4777 8803 4811
rect 8953 4777 8987 4811
rect 11437 4777 11471 4811
rect 14105 4777 14139 4811
rect 15945 4777 15979 4811
rect 17509 4777 17543 4811
rect 19625 4777 19659 4811
rect 22201 4777 22235 4811
rect 25053 4777 25087 4811
rect 25329 4777 25363 4811
rect 26617 4777 26651 4811
rect 29285 4777 29319 4811
rect 33333 4777 33367 4811
rect 39497 4777 39531 4811
rect 5917 4709 5951 4743
rect 13921 4709 13955 4743
rect 15209 4709 15243 4743
rect 15485 4709 15519 4743
rect 17785 4709 17819 4743
rect 18245 4709 18279 4743
rect 19257 4709 19291 4743
rect 23581 4709 23615 4743
rect 30205 4709 30239 4743
rect 35081 4709 35115 4743
rect 36829 4709 36863 4743
rect 43453 4709 43487 4743
rect 3801 4641 3835 4675
rect 5457 4641 5491 4675
rect 6193 4641 6227 4675
rect 6469 4641 6503 4675
rect 7757 4641 7791 4675
rect 9965 4641 9999 4675
rect 12909 4641 12943 4675
rect 16497 4641 16531 4675
rect 18107 4641 18141 4675
rect 18705 4641 18739 4675
rect 18797 4641 18831 4675
rect 19533 4641 19567 4675
rect 20085 4641 20119 4675
rect 20545 4641 20579 4675
rect 20821 4641 20855 4675
rect 23029 4641 23063 4675
rect 23188 4641 23222 4675
rect 23305 4641 23339 4675
rect 26433 4630 26467 4664
rect 27813 4641 27847 4675
rect 28273 4641 28307 4675
rect 30481 4641 30515 4675
rect 30619 4641 30653 4675
rect 31677 4641 31711 4675
rect 32137 4641 32171 4675
rect 32413 4641 32447 4675
rect 37222 4641 37256 4675
rect 37381 4641 37415 4675
rect 38485 4641 38519 4675
rect 1501 4573 1535 4607
rect 1869 4573 1903 4607
rect 2421 4573 2455 4607
rect 2697 4573 2731 4607
rect 4077 4573 4111 4607
rect 5273 4573 5307 4607
rect 6310 4573 6344 4607
rect 8033 4573 8067 4607
rect 9686 4573 9720 4607
rect 10425 4573 10459 4607
rect 10701 4573 10735 4607
rect 11805 4573 11839 4607
rect 12081 4573 12115 4607
rect 13185 4573 13219 4607
rect 14841 4573 14875 4607
rect 15117 4573 15151 4607
rect 15393 4573 15427 4607
rect 15669 4573 15703 4607
rect 16129 4573 16163 4607
rect 16773 4573 16807 4607
rect 17693 4573 17727 4607
rect 17877 4573 17911 4607
rect 18020 4573 18054 4607
rect 19809 4573 19843 4607
rect 19901 4573 19935 4607
rect 20938 4573 20972 4607
rect 21097 4573 21131 4607
rect 22017 4573 22051 4607
rect 24041 4573 24075 4607
rect 24225 4573 24259 4607
rect 24685 4573 24719 4607
rect 25053 4573 25087 4607
rect 26065 4573 26099 4607
rect 26341 4573 26375 4607
rect 26709 4573 26743 4607
rect 27537 4573 27571 4607
rect 28549 4573 28583 4607
rect 29561 4573 29595 4607
rect 29745 4573 29779 4607
rect 30757 4573 30791 4607
rect 31493 4573 31527 4607
rect 32551 4573 32585 4607
rect 32689 4573 32723 4607
rect 34069 4573 34103 4607
rect 35265 4573 35299 4607
rect 36185 4573 36219 4607
rect 36369 4573 36403 4607
rect 37105 4573 37139 4607
rect 38761 4573 38795 4607
rect 42901 4573 42935 4607
rect 43269 4573 43303 4607
rect 2053 4505 2087 4539
rect 7481 4505 7515 4539
rect 10149 4505 10183 4539
rect 21833 4505 21867 4539
rect 34253 4505 34287 4539
rect 38025 4505 38059 4539
rect 38301 4505 38335 4539
rect 1593 4437 1627 4471
rect 4813 4437 4847 4471
rect 5089 4437 5123 4471
rect 7573 4437 7607 4471
rect 10241 4437 10275 4471
rect 12817 4437 12851 4471
rect 18613 4437 18647 4471
rect 21741 4437 21775 4471
rect 22385 4437 22419 4471
rect 25237 4437 25271 4471
rect 26433 4437 26467 4471
rect 26801 4437 26835 4471
rect 31401 4437 31435 4471
rect 38209 4437 38243 4471
rect 43085 4437 43119 4471
rect 2697 4233 2731 4267
rect 5825 4233 5859 4267
rect 18613 4233 18647 4267
rect 21649 4233 21683 4267
rect 22201 4233 22235 4267
rect 22569 4233 22603 4267
rect 25973 4233 26007 4267
rect 26157 4233 26191 4267
rect 27445 4233 27479 4267
rect 29285 4233 29319 4267
rect 30481 4233 30515 4267
rect 34253 4233 34287 4267
rect 1501 4165 1535 4199
rect 1869 4165 1903 4199
rect 2237 4165 2271 4199
rect 2881 4165 2915 4199
rect 8585 4165 8619 4199
rect 2513 4097 2547 4131
rect 3157 4097 3191 4131
rect 3433 4097 3467 4131
rect 4261 4097 4295 4131
rect 5089 4097 5123 4131
rect 9735 4097 9769 4131
rect 9873 4097 9907 4131
rect 10793 4097 10827 4131
rect 11069 4097 11103 4131
rect 12265 4097 12299 4131
rect 12725 4097 12759 4131
rect 13645 4097 13679 4131
rect 14565 4097 14599 4131
rect 16865 4097 16899 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 18797 4097 18831 4131
rect 22109 4097 22143 4131
rect 22937 4097 22971 4131
rect 24133 4097 24167 4131
rect 25237 4097 25271 4131
rect 25421 4097 25455 4131
rect 25793 4097 25827 4131
rect 26642 4097 26676 4131
rect 27353 4097 27387 4131
rect 28273 4097 28307 4131
rect 28549 4097 28583 4131
rect 30665 4097 30699 4131
rect 32413 4097 32447 4131
rect 32597 4097 32631 4131
rect 33450 4097 33484 4131
rect 35382 4097 35416 4131
rect 36921 4097 36955 4131
rect 38393 4097 38427 4131
rect 38485 4097 38519 4131
rect 39037 4097 39071 4131
rect 42257 4097 42291 4131
rect 42625 4097 42659 4131
rect 42901 4097 42935 4131
rect 43269 4097 43303 4131
rect 4813 4029 4847 4063
rect 8677 4029 8711 4063
rect 8861 4029 8895 4063
rect 9597 4029 9631 4063
rect 10517 4029 10551 4063
rect 12909 4029 12943 4063
rect 13369 4029 13403 4063
rect 13762 4029 13796 4063
rect 13921 4029 13955 4063
rect 16681 4029 16715 4063
rect 17325 4029 17359 4063
rect 17601 4029 17635 4063
rect 17718 4029 17752 4063
rect 19809 4029 19843 4063
rect 19993 4029 20027 4063
rect 20729 4029 20763 4063
rect 20867 4029 20901 4063
rect 21005 4029 21039 4063
rect 22017 4029 22051 4063
rect 23121 4029 23155 4063
rect 23581 4029 23615 4063
rect 23857 4029 23891 4063
rect 23995 4029 24029 4063
rect 24777 4029 24811 4063
rect 25329 4029 25363 4063
rect 25881 4029 25915 4063
rect 26249 4029 26283 4063
rect 27629 4029 27663 4063
rect 33057 4029 33091 4063
rect 33333 4029 33367 4063
rect 33609 4029 33643 4063
rect 34345 4029 34379 4063
rect 34529 4029 34563 4063
rect 35265 4029 35299 4063
rect 35541 4029 35575 4063
rect 36185 4029 36219 4063
rect 2053 3961 2087 3995
rect 4169 3961 4203 3995
rect 4445 3961 4479 3995
rect 9321 3961 9355 3995
rect 20453 3961 20487 3995
rect 25605 3961 25639 3995
rect 34989 3961 35023 3995
rect 36737 3961 36771 3995
rect 38853 3961 38887 3995
rect 42073 3961 42107 3995
rect 43453 3961 43487 3995
rect 1593 3893 1627 3927
rect 2329 3893 2363 3927
rect 2697 3893 2731 3927
rect 2973 3893 3007 3927
rect 7297 3893 7331 3927
rect 10609 3893 10643 3927
rect 10885 3893 10919 3927
rect 12081 3893 12115 3927
rect 26571 3893 26605 3927
rect 26985 3893 27019 3927
rect 38301 3893 38335 3927
rect 38669 3893 38703 3927
rect 42441 3893 42475 3927
rect 43085 3893 43119 3927
rect 7849 3689 7883 3723
rect 9965 3689 9999 3723
rect 11529 3689 11563 3723
rect 13369 3689 13403 3723
rect 14105 3689 14139 3723
rect 16497 3689 16531 3723
rect 29285 3689 29319 3723
rect 30573 3689 30607 3723
rect 32597 3689 32631 3723
rect 35265 3689 35299 3723
rect 38301 3689 38335 3723
rect 42073 3689 42107 3723
rect 2789 3621 2823 3655
rect 5825 3621 5859 3655
rect 19349 3621 19383 3655
rect 20637 3621 20671 3655
rect 42625 3621 42659 3655
rect 43453 3621 43487 3655
rect 2421 3553 2455 3587
rect 4813 3553 4847 3587
rect 6561 3553 6595 3587
rect 6720 3553 6754 3587
rect 7113 3553 7147 3587
rect 7573 3553 7607 3587
rect 8953 3553 8987 3587
rect 10517 3553 10551 3587
rect 11621 3553 11655 3587
rect 15485 3553 15519 3587
rect 19625 3553 19659 3587
rect 22661 3553 22695 3587
rect 25697 3553 25731 3587
rect 25881 3553 25915 3587
rect 26341 3553 26375 3587
rect 26617 3553 26651 3587
rect 26755 3553 26789 3587
rect 26893 3553 26927 3587
rect 28273 3553 28307 3587
rect 29561 3553 29595 3587
rect 31585 3553 31619 3587
rect 32689 3553 32723 3587
rect 36277 3553 36311 3587
rect 37289 3553 37323 3587
rect 1501 3485 1535 3519
rect 3249 3485 3283 3519
rect 5089 3485 5123 3519
rect 6837 3485 6871 3519
rect 7757 3485 7791 3519
rect 8033 3485 8067 3519
rect 9229 3485 9263 3519
rect 10333 3485 10367 3519
rect 10793 3485 10827 3519
rect 11897 3485 11931 3519
rect 13185 3485 13219 3519
rect 13737 3485 13771 3519
rect 14289 3485 14323 3519
rect 14657 3485 14691 3519
rect 15761 3485 15795 3519
rect 17509 3485 17543 3519
rect 17785 3485 17819 3519
rect 19533 3485 19567 3519
rect 19901 3485 19935 3519
rect 21833 3485 21867 3519
rect 22937 3485 22971 3519
rect 24961 3485 24995 3519
rect 28549 3485 28583 3519
rect 29837 3485 29871 3519
rect 31861 3485 31895 3519
rect 32965 3485 32999 3519
rect 34897 3485 34931 3519
rect 36001 3485 36035 3519
rect 37565 3485 37599 3519
rect 38393 3485 38427 3519
rect 39129 3485 39163 3519
rect 42257 3485 42291 3519
rect 42533 3485 42567 3519
rect 42809 3485 42843 3519
rect 42901 3485 42935 3519
rect 43269 3485 43303 3519
rect 1869 3417 1903 3451
rect 2237 3417 2271 3451
rect 2605 3417 2639 3451
rect 3433 3417 3467 3451
rect 8585 3417 8619 3451
rect 8769 3417 8803 3451
rect 12817 3417 12851 3451
rect 14841 3417 14875 3451
rect 38761 3417 38795 3451
rect 1593 3349 1627 3383
rect 1961 3349 1995 3383
rect 5917 3349 5951 3383
rect 10149 3349 10183 3383
rect 12633 3349 12667 3383
rect 12909 3349 12943 3383
rect 13369 3349 13403 3383
rect 13553 3349 13587 3383
rect 18521 3349 18555 3383
rect 22017 3349 22051 3383
rect 23673 3349 23707 3383
rect 25145 3349 25179 3383
rect 27537 3349 27571 3383
rect 33701 3349 33735 3383
rect 34713 3349 34747 3383
rect 38945 3349 38979 3383
rect 42349 3349 42383 3383
rect 43085 3349 43119 3383
rect 2881 3145 2915 3179
rect 7389 3145 7423 3179
rect 13369 3145 13403 3179
rect 14933 3145 14967 3179
rect 16497 3145 16531 3179
rect 16865 3145 16899 3179
rect 17233 3145 17267 3179
rect 17509 3145 17543 3179
rect 25973 3145 26007 3179
rect 30297 3145 30331 3179
rect 31493 3145 31527 3179
rect 36185 3145 36219 3179
rect 38577 3145 38611 3179
rect 38945 3145 38979 3179
rect 40417 3145 40451 3179
rect 41153 3145 41187 3179
rect 41613 3145 41647 3179
rect 41797 3145 41831 3179
rect 43453 3145 43487 3179
rect 2789 3077 2823 3111
rect 22109 3077 22143 3111
rect 2329 3009 2363 3043
rect 6653 3009 6687 3043
rect 7757 3009 7791 3043
rect 8125 3009 8159 3043
rect 10241 3009 10275 3043
rect 10609 3009 10643 3043
rect 11713 3009 11747 3043
rect 12587 3009 12621 3043
rect 13461 3009 13495 3043
rect 13737 3009 13771 3043
rect 14933 3009 14967 3043
rect 15025 3009 15059 3043
rect 15485 3009 15519 3043
rect 15761 3009 15795 3043
rect 16773 3009 16807 3043
rect 17141 3009 17175 3043
rect 18153 3009 18187 3043
rect 18312 3009 18346 3043
rect 19165 3009 19199 3043
rect 19625 3009 19659 3043
rect 20478 3009 20512 3043
rect 21281 3009 21315 3043
rect 21557 3009 21591 3043
rect 21925 3009 21959 3043
rect 22937 3009 22971 3043
rect 23213 3009 23247 3043
rect 23305 3009 23339 3043
rect 23857 3009 23891 3043
rect 24133 3009 24167 3043
rect 24961 3009 24995 3043
rect 25237 3009 25271 3043
rect 26065 3009 26099 3043
rect 27353 3009 27387 3043
rect 27537 3009 27571 3043
rect 27721 3009 27755 3043
rect 28574 3009 28608 3043
rect 29377 3009 29411 3043
rect 29653 3009 29687 3043
rect 30113 3009 30147 3043
rect 30481 3009 30515 3043
rect 30757 3009 30791 3043
rect 32413 3009 32447 3043
rect 32597 3009 32631 3043
rect 33333 3009 33367 3043
rect 33609 3009 33643 3043
rect 34345 3009 34379 3043
rect 34529 3009 34563 3043
rect 35265 3009 35299 3043
rect 38393 3009 38427 3043
rect 38761 3009 38795 3043
rect 40601 3009 40635 3043
rect 41337 3009 41371 3043
rect 41429 3009 41463 3043
rect 41981 3009 42015 3043
rect 42257 3009 42291 3043
rect 42533 3009 42567 3043
rect 42901 3009 42935 3043
rect 43269 3009 43303 3043
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 6377 2941 6411 2975
rect 7941 2941 7975 2975
rect 8861 2941 8895 2975
rect 8978 2941 9012 2975
rect 9137 2941 9171 2975
rect 9781 2941 9815 2975
rect 10333 2941 10367 2975
rect 11529 2941 11563 2975
rect 12449 2941 12483 2975
rect 12725 2941 12759 2975
rect 15117 2941 15151 2975
rect 18429 2941 18463 2975
rect 19349 2941 19383 2975
rect 19441 2941 19475 2975
rect 20361 2941 20395 2975
rect 20637 2941 20671 2975
rect 28457 2941 28491 2975
rect 28733 2941 28767 2975
rect 33057 2941 33091 2975
rect 33450 2941 33484 2975
rect 35382 2941 35416 2975
rect 35541 2941 35575 2975
rect 2513 2873 2547 2907
rect 8585 2873 8619 2907
rect 11345 2873 11379 2907
rect 12173 2873 12207 2907
rect 14473 2873 14507 2907
rect 18705 2873 18739 2907
rect 20085 2873 20119 2907
rect 22201 2873 22235 2907
rect 24869 2873 24903 2907
rect 26249 2873 26283 2907
rect 27169 2873 27203 2907
rect 28181 2873 28215 2907
rect 34989 2873 35023 2907
rect 42717 2873 42751 2907
rect 7573 2805 7607 2839
rect 10057 2805 10091 2839
rect 14565 2805 14599 2839
rect 21373 2805 21407 2839
rect 23489 2805 23523 2839
rect 29469 2805 29503 2839
rect 34253 2805 34287 2839
rect 42073 2805 42107 2839
rect 43085 2805 43119 2839
rect 3433 2601 3467 2635
rect 7389 2601 7423 2635
rect 8493 2601 8527 2635
rect 8953 2601 8987 2635
rect 10241 2601 10275 2635
rect 11345 2601 11379 2635
rect 12541 2601 12575 2635
rect 18613 2601 18647 2635
rect 20269 2601 20303 2635
rect 21373 2601 21407 2635
rect 23397 2601 23431 2635
rect 25973 2601 26007 2635
rect 28181 2601 28215 2635
rect 31401 2601 31435 2635
rect 33149 2601 33183 2635
rect 34713 2601 34747 2635
rect 35817 2601 35851 2635
rect 5549 2533 5583 2567
rect 14565 2533 14599 2567
rect 28089 2533 28123 2567
rect 42165 2533 42199 2567
rect 43453 2533 43487 2567
rect 1685 2465 1719 2499
rect 2605 2465 2639 2499
rect 6377 2465 6411 2499
rect 7481 2465 7515 2499
rect 11529 2465 11563 2499
rect 20361 2465 20395 2499
rect 22385 2465 22419 2499
rect 24961 2465 24995 2499
rect 27077 2465 27111 2499
rect 29193 2465 29227 2499
rect 30389 2465 30423 2499
rect 32137 2465 32171 2499
rect 1409 2397 1443 2431
rect 2329 2397 2363 2431
rect 4077 2397 4111 2431
rect 4905 2397 4939 2431
rect 6193 2397 6227 2431
rect 6653 2397 6687 2431
rect 7757 2397 7791 2431
rect 9689 2397 9723 2431
rect 9965 2397 9999 2431
rect 10057 2397 10091 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 11805 2397 11839 2431
rect 12633 2397 12667 2431
rect 13001 2397 13035 2431
rect 13737 2397 13771 2431
rect 14749 2397 14783 2431
rect 15669 2397 15703 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 17601 2397 17635 2431
rect 17877 2397 17911 2431
rect 19257 2397 19291 2431
rect 19533 2397 19567 2431
rect 20637 2397 20671 2431
rect 22293 2397 22327 2431
rect 22661 2397 22695 2431
rect 25237 2397 25271 2431
rect 27353 2397 27387 2431
rect 28917 2397 28951 2431
rect 30665 2397 30699 2431
rect 32413 2397 32447 2431
rect 34161 2397 34195 2431
rect 35449 2397 35483 2431
rect 35725 2397 35759 2431
rect 36553 2397 36587 2431
rect 36829 2397 36863 2431
rect 41981 2397 42015 2431
rect 42533 2397 42567 2431
rect 42901 2397 42935 2431
rect 43269 2397 43303 2431
rect 3341 2329 3375 2363
rect 5733 2329 5767 2363
rect 14197 2329 14231 2363
rect 14381 2329 14415 2363
rect 3893 2261 3927 2295
rect 4721 2261 4755 2295
rect 6009 2261 6043 2295
rect 12817 2261 12851 2295
rect 13185 2261 13219 2295
rect 13553 2261 13587 2295
rect 15485 2261 15519 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 22109 2261 22143 2295
rect 33977 2261 34011 2295
rect 42717 2261 42751 2295
rect 43085 2261 43119 2295
<< metal1 >>
rect 14090 10888 14096 10940
rect 14148 10928 14154 10940
rect 30098 10928 30104 10940
rect 14148 10900 30104 10928
rect 14148 10888 14154 10900
rect 30098 10888 30104 10900
rect 30156 10888 30162 10940
rect 11146 10820 11152 10872
rect 11204 10860 11210 10872
rect 36998 10860 37004 10872
rect 11204 10832 37004 10860
rect 11204 10820 11210 10832
rect 36998 10820 37004 10832
rect 37056 10820 37062 10872
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 26878 10792 26884 10804
rect 4488 10764 26884 10792
rect 4488 10752 4494 10764
rect 26878 10752 26884 10764
rect 26936 10752 26942 10804
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 34054 10724 34060 10736
rect 5132 10696 34060 10724
rect 5132 10684 5138 10696
rect 34054 10684 34060 10696
rect 34112 10684 34118 10736
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 37090 10656 37096 10668
rect 6420 10628 37096 10656
rect 6420 10616 6426 10628
rect 37090 10616 37096 10628
rect 37148 10616 37154 10668
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 19150 10588 19156 10600
rect 8720 10560 19156 10588
rect 8720 10548 8726 10560
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 30742 10520 30748 10532
rect 26712 10492 30748 10520
rect 26712 10464 26740 10492
rect 30742 10480 30748 10492
rect 30800 10480 30806 10532
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 11514 10452 11520 10464
rect 9272 10424 11520 10452
rect 9272 10412 9278 10424
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 16850 10412 16856 10464
rect 16908 10452 16914 10464
rect 21910 10452 21916 10464
rect 16908 10424 21916 10452
rect 16908 10412 16914 10424
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 26694 10412 26700 10464
rect 26752 10412 26758 10464
rect 33226 10452 33232 10464
rect 26804 10424 33232 10452
rect 8110 10344 8116 10396
rect 8168 10384 8174 10396
rect 12158 10384 12164 10396
rect 8168 10356 12164 10384
rect 8168 10344 8174 10356
rect 12158 10344 12164 10356
rect 12216 10344 12222 10396
rect 14366 10344 14372 10396
rect 14424 10384 14430 10396
rect 19610 10384 19616 10396
rect 14424 10356 19616 10384
rect 14424 10344 14430 10356
rect 19610 10344 19616 10356
rect 19668 10344 19674 10396
rect 25130 10344 25136 10396
rect 25188 10384 25194 10396
rect 26804 10384 26832 10424
rect 33226 10412 33232 10424
rect 33284 10412 33290 10464
rect 33870 10412 33876 10464
rect 33928 10452 33934 10464
rect 37274 10452 37280 10464
rect 33928 10424 37280 10452
rect 33928 10412 33934 10424
rect 37274 10412 37280 10424
rect 37332 10412 37338 10464
rect 37734 10412 37740 10464
rect 37792 10452 37798 10464
rect 39758 10452 39764 10464
rect 37792 10424 39764 10452
rect 37792 10412 37798 10424
rect 39758 10412 39764 10424
rect 39816 10412 39822 10464
rect 25188 10356 26832 10384
rect 25188 10344 25194 10356
rect 30006 10344 30012 10396
rect 30064 10384 30070 10396
rect 32582 10384 32588 10396
rect 30064 10356 32588 10384
rect 30064 10344 30070 10356
rect 32582 10344 32588 10356
rect 32640 10344 32646 10396
rect 36906 10344 36912 10396
rect 36964 10384 36970 10396
rect 39206 10384 39212 10396
rect 36964 10356 39212 10384
rect 36964 10344 36970 10356
rect 39206 10344 39212 10356
rect 39264 10344 39270 10396
rect 42518 10384 42524 10396
rect 41386 10356 42524 10384
rect 7834 10276 7840 10328
rect 7892 10316 7898 10328
rect 11790 10316 11796 10328
rect 7892 10288 11796 10316
rect 7892 10276 7898 10288
rect 11790 10276 11796 10288
rect 11848 10276 11854 10328
rect 29178 10276 29184 10328
rect 29236 10316 29242 10328
rect 31846 10316 31852 10328
rect 29236 10288 31852 10316
rect 29236 10276 29242 10288
rect 31846 10276 31852 10288
rect 31904 10276 31910 10328
rect 36630 10276 36636 10328
rect 36688 10316 36694 10328
rect 39022 10316 39028 10328
rect 36688 10288 39028 10316
rect 36688 10276 36694 10288
rect 39022 10276 39028 10288
rect 39080 10276 39086 10328
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 10962 10248 10968 10260
rect 7340 10220 10968 10248
rect 7340 10208 7346 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11054 10208 11060 10260
rect 11112 10248 11118 10260
rect 12618 10248 12624 10260
rect 11112 10220 12624 10248
rect 11112 10208 11118 10220
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 16206 10248 16212 10260
rect 13320 10220 16212 10248
rect 13320 10208 13326 10220
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 29730 10208 29736 10260
rect 29788 10248 29794 10260
rect 31570 10248 31576 10260
rect 29788 10220 31576 10248
rect 29788 10208 29794 10220
rect 31570 10208 31576 10220
rect 31628 10208 31634 10260
rect 32766 10208 32772 10260
rect 32824 10248 32830 10260
rect 36906 10248 36912 10260
rect 32824 10220 36912 10248
rect 32824 10208 32830 10220
rect 36906 10208 36912 10220
rect 36964 10208 36970 10260
rect 37458 10208 37464 10260
rect 37516 10248 37522 10260
rect 39482 10248 39488 10260
rect 37516 10220 39488 10248
rect 37516 10208 37522 10220
rect 39482 10208 39488 10220
rect 39540 10208 39546 10260
rect 7190 10140 7196 10192
rect 7248 10180 7254 10192
rect 10410 10180 10416 10192
rect 7248 10152 10416 10180
rect 7248 10140 7254 10152
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 22186 10140 22192 10192
rect 22244 10180 22250 10192
rect 35342 10180 35348 10192
rect 22244 10152 35348 10180
rect 22244 10140 22250 10152
rect 35342 10140 35348 10152
rect 35400 10140 35406 10192
rect 36078 10140 36084 10192
rect 36136 10180 36142 10192
rect 37826 10180 37832 10192
rect 36136 10152 37832 10180
rect 36136 10140 36142 10152
rect 37826 10140 37832 10152
rect 37884 10140 37890 10192
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 10686 10112 10692 10124
rect 7800 10084 10692 10112
rect 7800 10072 7806 10084
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 15102 10112 15108 10124
rect 13596 10084 15108 10112
rect 13596 10072 13602 10084
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19484 10084 21496 10112
rect 19484 10072 19490 10084
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 10134 10044 10140 10056
rect 6696 10016 10140 10044
rect 6696 10004 6702 10016
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 10226 10004 10232 10056
rect 10284 10044 10290 10056
rect 13998 10044 14004 10056
rect 10284 10016 14004 10044
rect 10284 10004 10290 10016
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 14108 10016 17172 10044
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 9858 9976 9864 9988
rect 8352 9948 9864 9976
rect 8352 9936 8358 9948
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 9950 9936 9956 9988
rect 10008 9976 10014 9988
rect 13722 9976 13728 9988
rect 10008 9948 13728 9976
rect 10008 9936 10014 9948
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 6454 9868 6460 9920
rect 6512 9908 6518 9920
rect 8754 9908 8760 9920
rect 6512 9880 8760 9908
rect 6512 9868 6518 9880
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 11054 9908 11060 9920
rect 9180 9880 11060 9908
rect 9180 9868 9186 9880
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11330 9868 11336 9920
rect 11388 9908 11394 9920
rect 14108 9908 14136 10016
rect 15470 9936 15476 9988
rect 15528 9976 15534 9988
rect 17144 9976 17172 10016
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 21358 10044 21364 10056
rect 19392 10016 21364 10044
rect 19392 10004 19398 10016
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 21468 10044 21496 10084
rect 24670 10072 24676 10124
rect 24728 10112 24734 10124
rect 30466 10112 30472 10124
rect 24728 10084 30472 10112
rect 24728 10072 24734 10084
rect 30466 10072 30472 10084
rect 30524 10072 30530 10124
rect 31386 10072 31392 10124
rect 31444 10112 31450 10124
rect 34882 10112 34888 10124
rect 31444 10084 34888 10112
rect 31444 10072 31450 10084
rect 34882 10072 34888 10084
rect 34940 10072 34946 10124
rect 35526 10072 35532 10124
rect 35584 10112 35590 10124
rect 38194 10112 38200 10124
rect 35584 10084 38200 10112
rect 35584 10072 35590 10084
rect 38194 10072 38200 10084
rect 38252 10072 38258 10124
rect 38286 10072 38292 10124
rect 38344 10112 38350 10124
rect 40034 10112 40040 10124
rect 38344 10084 40040 10112
rect 38344 10072 38350 10084
rect 40034 10072 40040 10084
rect 40092 10072 40098 10124
rect 23198 10044 23204 10056
rect 21468 10016 23204 10044
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 28902 10004 28908 10056
rect 28960 10044 28966 10056
rect 30006 10044 30012 10056
rect 28960 10016 30012 10044
rect 28960 10004 28966 10016
rect 30006 10004 30012 10016
rect 30064 10004 30070 10056
rect 30834 10004 30840 10056
rect 30892 10044 30898 10056
rect 34790 10044 34796 10056
rect 30892 10016 34796 10044
rect 30892 10004 30898 10016
rect 34790 10004 34796 10016
rect 34848 10004 34854 10056
rect 36354 10004 36360 10056
rect 36412 10044 36418 10056
rect 38654 10044 38660 10056
rect 36412 10016 38660 10044
rect 36412 10004 36418 10016
rect 38654 10004 38660 10016
rect 38712 10004 38718 10056
rect 38838 10004 38844 10056
rect 38896 10044 38902 10056
rect 41046 10044 41052 10056
rect 38896 10016 41052 10044
rect 38896 10004 38902 10016
rect 41046 10004 41052 10016
rect 41104 10004 41110 10056
rect 25130 9976 25136 9988
rect 15528 9948 17080 9976
rect 17144 9948 25136 9976
rect 15528 9936 15534 9948
rect 11388 9880 14136 9908
rect 11388 9868 11394 9880
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 16482 9908 16488 9920
rect 14516 9880 16488 9908
rect 14516 9868 14522 9880
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 5810 9800 5816 9852
rect 5868 9840 5874 9852
rect 9030 9840 9036 9852
rect 5868 9812 9036 9840
rect 5868 9800 5874 9812
rect 9030 9800 9036 9812
rect 9088 9800 9094 9852
rect 9766 9800 9772 9852
rect 9824 9840 9830 9852
rect 12066 9840 12072 9852
rect 9824 9812 12072 9840
rect 9824 9800 9830 9812
rect 12066 9800 12072 9812
rect 12124 9800 12130 9852
rect 13354 9800 13360 9852
rect 13412 9840 13418 9852
rect 14274 9840 14280 9852
rect 13412 9812 14280 9840
rect 13412 9800 13418 9812
rect 14274 9800 14280 9812
rect 14332 9800 14338 9852
rect 15102 9800 15108 9852
rect 15160 9840 15166 9852
rect 16758 9840 16764 9852
rect 15160 9812 16764 9840
rect 15160 9800 15166 9812
rect 16758 9800 16764 9812
rect 16816 9800 16822 9852
rect 17052 9840 17080 9948
rect 25130 9936 25136 9948
rect 25188 9936 25194 9988
rect 28442 9976 28448 9988
rect 25240 9948 28448 9976
rect 17126 9868 17132 9920
rect 17184 9908 17190 9920
rect 25240 9908 25268 9948
rect 28442 9936 28448 9948
rect 28500 9936 28506 9988
rect 28626 9936 28632 9988
rect 28684 9976 28690 9988
rect 29638 9976 29644 9988
rect 28684 9948 29644 9976
rect 28684 9936 28690 9948
rect 29638 9936 29644 9948
rect 29696 9936 29702 9988
rect 31110 9936 31116 9988
rect 31168 9976 31174 9988
rect 32122 9976 32128 9988
rect 31168 9948 32128 9976
rect 31168 9936 31174 9948
rect 32122 9936 32128 9948
rect 32180 9936 32186 9988
rect 35802 9936 35808 9988
rect 35860 9976 35866 9988
rect 37550 9976 37556 9988
rect 35860 9948 37556 9976
rect 35860 9936 35866 9948
rect 37550 9936 37556 9948
rect 37608 9936 37614 9988
rect 38562 9936 38568 9988
rect 38620 9976 38626 9988
rect 40678 9976 40684 9988
rect 38620 9948 40684 9976
rect 38620 9936 38626 9948
rect 40678 9936 40684 9948
rect 40736 9936 40742 9988
rect 17184 9880 25268 9908
rect 17184 9868 17190 9880
rect 25314 9868 25320 9920
rect 25372 9908 25378 9920
rect 27154 9908 27160 9920
rect 25372 9880 27160 9908
rect 25372 9868 25378 9880
rect 27154 9868 27160 9880
rect 27212 9868 27218 9920
rect 33318 9868 33324 9920
rect 33376 9908 33382 9920
rect 34606 9908 34612 9920
rect 33376 9880 34612 9908
rect 33376 9868 33382 9880
rect 34606 9868 34612 9880
rect 34664 9868 34670 9920
rect 34974 9868 34980 9920
rect 35032 9908 35038 9920
rect 36630 9908 36636 9920
rect 35032 9880 36636 9908
rect 35032 9868 35038 9880
rect 36630 9868 36636 9880
rect 36688 9868 36694 9920
rect 38010 9868 38016 9920
rect 38068 9908 38074 9920
rect 39942 9908 39948 9920
rect 38068 9880 39948 9908
rect 38068 9868 38074 9880
rect 39942 9868 39948 9880
rect 40000 9868 40006 9920
rect 21266 9840 21272 9852
rect 17052 9812 21272 9840
rect 21266 9800 21272 9812
rect 21324 9800 21330 9852
rect 21358 9800 21364 9852
rect 21416 9840 21422 9852
rect 22922 9840 22928 9852
rect 21416 9812 22928 9840
rect 21416 9800 21422 9812
rect 22922 9800 22928 9812
rect 22980 9800 22986 9852
rect 24762 9800 24768 9852
rect 24820 9840 24826 9852
rect 25958 9840 25964 9852
rect 24820 9812 25964 9840
rect 24820 9800 24826 9812
rect 25958 9800 25964 9812
rect 26016 9800 26022 9852
rect 27246 9800 27252 9852
rect 27304 9840 27310 9852
rect 27890 9840 27896 9852
rect 27304 9812 27896 9840
rect 27304 9800 27310 9812
rect 27890 9800 27896 9812
rect 27948 9800 27954 9852
rect 28350 9800 28356 9852
rect 28408 9840 28414 9852
rect 29270 9840 29276 9852
rect 28408 9812 29276 9840
rect 28408 9800 28414 9812
rect 29270 9800 29276 9812
rect 29328 9800 29334 9852
rect 29454 9800 29460 9852
rect 29512 9840 29518 9852
rect 31478 9840 31484 9852
rect 29512 9812 31484 9840
rect 29512 9800 29518 9812
rect 31478 9800 31484 9812
rect 31536 9800 31542 9852
rect 34330 9800 34336 9852
rect 34388 9840 34394 9852
rect 35250 9840 35256 9852
rect 34388 9812 35256 9840
rect 34388 9800 34394 9812
rect 35250 9800 35256 9812
rect 35308 9800 35314 9852
rect 35342 9800 35348 9852
rect 35400 9840 35406 9852
rect 41386 9840 41414 10356
rect 42518 10344 42524 10356
rect 42576 10344 42582 10396
rect 35400 9812 41414 9840
rect 35400 9800 35406 9812
rect 4154 9732 4160 9784
rect 4212 9772 4218 9784
rect 7098 9772 7104 9784
rect 4212 9744 7104 9772
rect 4212 9732 4218 9744
rect 7098 9732 7104 9744
rect 7156 9732 7162 9784
rect 7466 9732 7472 9784
rect 7524 9772 7530 9784
rect 9306 9772 9312 9784
rect 7524 9744 9312 9772
rect 7524 9732 7530 9744
rect 9306 9732 9312 9744
rect 9364 9732 9370 9784
rect 9490 9732 9496 9784
rect 9548 9772 9554 9784
rect 13446 9772 13452 9784
rect 9548 9744 13452 9772
rect 9548 9732 9554 9744
rect 13446 9732 13452 9744
rect 13504 9732 13510 9784
rect 13630 9732 13636 9784
rect 13688 9772 13694 9784
rect 14550 9772 14556 9784
rect 13688 9744 14556 9772
rect 13688 9732 13694 9744
rect 14550 9732 14556 9744
rect 14608 9732 14614 9784
rect 16298 9732 16304 9784
rect 16356 9772 16362 9784
rect 17586 9772 17592 9784
rect 16356 9744 17592 9772
rect 16356 9732 16362 9744
rect 17586 9732 17592 9744
rect 17644 9732 17650 9784
rect 17678 9732 17684 9784
rect 17736 9772 17742 9784
rect 19518 9772 19524 9784
rect 17736 9744 19524 9772
rect 17736 9732 17742 9744
rect 19518 9732 19524 9744
rect 19576 9732 19582 9784
rect 19610 9732 19616 9784
rect 19668 9772 19674 9784
rect 19668 9744 26924 9772
rect 19668 9732 19674 9744
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 7374 9704 7380 9716
rect 6788 9676 7380 9704
rect 6788 9664 6794 9676
rect 7374 9664 7380 9676
rect 7432 9664 7438 9716
rect 8570 9664 8576 9716
rect 8628 9704 8634 9716
rect 11238 9704 11244 9716
rect 8628 9676 11244 9704
rect 8628 9664 8634 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13814 9704 13820 9716
rect 13228 9676 13820 9704
rect 13228 9664 13234 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 17310 9704 17316 9716
rect 16080 9676 17316 9704
rect 16080 9664 16086 9676
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 19150 9664 19156 9716
rect 19208 9704 19214 9716
rect 20622 9704 20628 9716
rect 19208 9676 20628 9704
rect 19208 9664 19214 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 22094 9704 22100 9716
rect 21232 9676 22100 9704
rect 21232 9664 21238 9676
rect 22094 9664 22100 9676
rect 22152 9664 22158 9716
rect 23382 9664 23388 9716
rect 23440 9704 23446 9716
rect 23658 9704 23664 9716
rect 23440 9676 23664 9704
rect 23440 9664 23446 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 23934 9664 23940 9716
rect 23992 9704 23998 9716
rect 25498 9704 25504 9716
rect 23992 9676 25504 9704
rect 23992 9664 23998 9676
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 25590 9664 25596 9716
rect 25648 9704 25654 9716
rect 26510 9704 26516 9716
rect 25648 9676 26516 9704
rect 25648 9664 25654 9676
rect 26510 9664 26516 9676
rect 26568 9664 26574 9716
rect 26896 9704 26924 9744
rect 26970 9732 26976 9784
rect 27028 9772 27034 9784
rect 27982 9772 27988 9784
rect 27028 9744 27988 9772
rect 27028 9732 27034 9744
rect 27982 9732 27988 9744
rect 28040 9732 28046 9784
rect 28074 9732 28080 9784
rect 28132 9772 28138 9784
rect 29086 9772 29092 9784
rect 28132 9744 29092 9772
rect 28132 9732 28138 9744
rect 29086 9732 29092 9744
rect 29144 9732 29150 9784
rect 39114 9732 39120 9784
rect 39172 9772 39178 9784
rect 41690 9772 41696 9784
rect 39172 9744 41696 9772
rect 39172 9732 39178 9744
rect 41690 9732 41696 9744
rect 41748 9732 41754 9784
rect 26896 9676 27476 9704
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 15838 9636 15844 9648
rect 5960 9608 15844 9636
rect 5960 9596 5966 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 16482 9596 16488 9648
rect 16540 9636 16546 9648
rect 27448 9636 27476 9676
rect 27522 9664 27528 9716
rect 27580 9704 27586 9716
rect 29178 9704 29184 9716
rect 27580 9676 29184 9704
rect 27580 9664 27586 9676
rect 29178 9664 29184 9676
rect 29236 9664 29242 9716
rect 32306 9704 32312 9716
rect 31772 9676 32312 9704
rect 31772 9674 31800 9676
rect 31680 9648 31800 9674
rect 32306 9664 32312 9676
rect 32364 9664 32370 9716
rect 32490 9664 32496 9716
rect 32548 9704 32554 9716
rect 33686 9704 33692 9716
rect 32548 9676 33692 9704
rect 32548 9664 32554 9676
rect 33686 9664 33692 9676
rect 33744 9664 33750 9716
rect 34146 9664 34152 9716
rect 34204 9704 34210 9716
rect 35618 9704 35624 9716
rect 34204 9676 35624 9704
rect 34204 9664 34210 9676
rect 35618 9664 35624 9676
rect 35676 9664 35682 9716
rect 37182 9664 37188 9716
rect 37240 9704 37246 9716
rect 39298 9704 39304 9716
rect 37240 9676 39304 9704
rect 37240 9664 37246 9676
rect 39298 9664 39304 9676
rect 39356 9664 39362 9716
rect 39390 9664 39396 9716
rect 39448 9704 39454 9716
rect 40310 9704 40316 9716
rect 39448 9676 40316 9704
rect 39448 9664 39454 9676
rect 40310 9664 40316 9676
rect 40368 9664 40374 9716
rect 28626 9636 28632 9648
rect 16540 9608 27384 9636
rect 27448 9608 28632 9636
rect 16540 9596 16546 9608
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 8478 9568 8484 9580
rect 5316 9540 8484 9568
rect 5316 9528 5322 9540
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 27356 9568 27384 9608
rect 28626 9596 28632 9608
rect 28684 9596 28690 9648
rect 31662 9596 31668 9648
rect 31720 9646 31800 9648
rect 31720 9596 31726 9646
rect 35434 9596 35440 9648
rect 35492 9636 35498 9648
rect 39850 9636 39856 9648
rect 35492 9608 39856 9636
rect 35492 9596 35498 9608
rect 39850 9596 39856 9608
rect 39908 9596 39914 9648
rect 29730 9568 29736 9580
rect 15804 9540 27292 9568
rect 27356 9540 29736 9568
rect 15804 9528 15810 9540
rect 4522 9460 4528 9512
rect 4580 9500 4586 9512
rect 13722 9500 13728 9512
rect 4580 9472 13728 9500
rect 4580 9460 4586 9472
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 16390 9460 16396 9512
rect 16448 9500 16454 9512
rect 26786 9500 26792 9512
rect 16448 9472 26792 9500
rect 16448 9460 16454 9472
rect 26786 9460 26792 9472
rect 26844 9460 26850 9512
rect 27264 9500 27292 9540
rect 29730 9528 29736 9540
rect 29788 9528 29794 9580
rect 31202 9500 31208 9512
rect 27264 9472 31208 9500
rect 31202 9460 31208 9472
rect 31260 9460 31266 9512
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 23290 9432 23296 9444
rect 7064 9404 23296 9432
rect 7064 9392 7070 9404
rect 23290 9392 23296 9404
rect 23348 9392 23354 9444
rect 27430 9432 27436 9444
rect 23400 9404 27436 9432
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 17954 9364 17960 9376
rect 7340 9336 17960 9364
rect 7340 9324 7346 9336
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 23400 9364 23428 9404
rect 27430 9392 27436 9404
rect 27488 9392 27494 9444
rect 31386 9392 31392 9444
rect 31444 9432 31450 9444
rect 32582 9432 32588 9444
rect 31444 9404 32588 9432
rect 31444 9392 31450 9404
rect 32582 9392 32588 9404
rect 32640 9392 32646 9444
rect 21324 9336 23428 9364
rect 21324 9324 21330 9336
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 43622 9364 43628 9376
rect 23900 9336 43628 9364
rect 23900 9324 23906 9336
rect 43622 9324 43628 9336
rect 43680 9324 43686 9376
rect 4338 9256 4344 9308
rect 4396 9296 4402 9308
rect 15562 9296 15568 9308
rect 4396 9268 15568 9296
rect 4396 9256 4402 9268
rect 15562 9256 15568 9268
rect 15620 9256 15626 9308
rect 18138 9256 18144 9308
rect 18196 9296 18202 9308
rect 40494 9296 40500 9308
rect 18196 9268 40500 9296
rect 18196 9256 18202 9268
rect 40494 9256 40500 9268
rect 40552 9256 40558 9308
rect 4706 9188 4712 9240
rect 4764 9228 4770 9240
rect 6914 9228 6920 9240
rect 4764 9200 6920 9228
rect 4764 9188 4770 9200
rect 6914 9188 6920 9200
rect 6972 9188 6978 9240
rect 11882 9188 11888 9240
rect 11940 9228 11946 9240
rect 34146 9228 34152 9240
rect 11940 9200 34152 9228
rect 11940 9188 11946 9200
rect 34146 9188 34152 9200
rect 34204 9188 34210 9240
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 5684 9132 15951 9160
rect 5684 9120 5690 9132
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 5718 9092 5724 9104
rect 3568 9064 5724 9092
rect 3568 9052 3574 9064
rect 5718 9052 5724 9064
rect 5776 9052 5782 9104
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 10962 9092 10968 9104
rect 6236 9064 10968 9092
rect 6236 9052 6242 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 15923 9092 15951 9132
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 35894 9160 35900 9172
rect 16264 9132 35900 9160
rect 16264 9120 16270 9132
rect 35894 9120 35900 9132
rect 35952 9120 35958 9172
rect 18506 9092 18512 9104
rect 11664 9064 12498 9092
rect 15923 9064 18512 9092
rect 11664 9052 11670 9064
rect 7098 8984 7104 9036
rect 7156 9024 7162 9036
rect 12470 9024 12498 9064
rect 18506 9052 18512 9064
rect 18564 9052 18570 9104
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 19668 9064 22094 9092
rect 19668 9052 19674 9064
rect 19426 9024 19432 9036
rect 7156 8996 12434 9024
rect 12470 8996 19432 9024
rect 7156 8984 7162 8996
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 11146 8956 11152 8968
rect 6144 8928 11152 8956
rect 6144 8916 6150 8928
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 4890 8848 4896 8900
rect 4948 8888 4954 8900
rect 8202 8888 8208 8900
rect 4948 8860 8208 8888
rect 4948 8848 4954 8860
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 12406 8888 12434 8996
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 20530 8956 20536 8968
rect 13964 8928 20536 8956
rect 13964 8916 13970 8928
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 22066 8956 22094 9064
rect 26786 9052 26792 9104
rect 26844 9092 26850 9104
rect 28994 9092 29000 9104
rect 26844 9064 29000 9092
rect 26844 9052 26850 9064
rect 28994 9052 29000 9064
rect 29052 9052 29058 9104
rect 30650 9052 30656 9104
rect 30708 9092 30714 9104
rect 35802 9092 35808 9104
rect 30708 9064 35808 9092
rect 30708 9052 30714 9064
rect 35802 9052 35808 9064
rect 35860 9052 35866 9104
rect 26878 8984 26884 9036
rect 26936 9024 26942 9036
rect 41138 9024 41144 9036
rect 26936 8996 41144 9024
rect 26936 8984 26942 8996
rect 41138 8984 41144 8996
rect 41196 8984 41202 9036
rect 29822 8956 29828 8968
rect 22066 8928 29828 8956
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 31662 8916 31668 8968
rect 31720 8956 31726 8968
rect 32122 8956 32128 8968
rect 31720 8928 32128 8956
rect 31720 8916 31726 8928
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 39574 8916 39580 8968
rect 39632 8956 39638 8968
rect 42610 8956 42616 8968
rect 39632 8928 42616 8956
rect 39632 8916 39638 8928
rect 42610 8916 42616 8928
rect 42668 8916 42674 8968
rect 17494 8888 17500 8900
rect 12406 8860 17500 8888
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 21910 8848 21916 8900
rect 21968 8888 21974 8900
rect 23658 8888 23664 8900
rect 21968 8860 23664 8888
rect 21968 8848 21974 8860
rect 23658 8848 23664 8860
rect 23716 8848 23722 8900
rect 24118 8848 24124 8900
rect 24176 8888 24182 8900
rect 34238 8888 34244 8900
rect 24176 8860 34244 8888
rect 24176 8848 24182 8860
rect 34238 8848 34244 8860
rect 34296 8848 34302 8900
rect 35710 8848 35716 8900
rect 35768 8888 35774 8900
rect 42978 8888 42984 8900
rect 35768 8860 42984 8888
rect 35768 8848 35774 8860
rect 42978 8848 42984 8860
rect 43036 8848 43042 8900
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 4798 8820 4804 8832
rect 3292 8792 4804 8820
rect 3292 8780 3298 8792
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 8662 8820 8668 8832
rect 8536 8792 8668 8820
rect 8536 8780 8542 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 11330 8820 11336 8832
rect 9916 8792 11336 8820
rect 9916 8780 9922 8792
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 14090 8820 14096 8832
rect 12584 8792 14096 8820
rect 12584 8780 12590 8792
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 19518 8820 19524 8832
rect 15344 8792 19524 8820
rect 15344 8780 15350 8792
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 22738 8780 22744 8832
rect 22796 8820 22802 8832
rect 28810 8820 28816 8832
rect 22796 8792 28816 8820
rect 22796 8780 22802 8792
rect 28810 8780 28816 8792
rect 28868 8780 28874 8832
rect 30466 8780 30472 8832
rect 30524 8820 30530 8832
rect 42702 8820 42708 8832
rect 30524 8792 42708 8820
rect 30524 8780 30530 8792
rect 42702 8780 42708 8792
rect 42760 8780 42766 8832
rect 1104 8730 43884 8752
rect 1104 8678 2658 8730
rect 2710 8678 2722 8730
rect 2774 8678 2786 8730
rect 2838 8678 2850 8730
rect 2902 8678 2914 8730
rect 2966 8678 2978 8730
rect 3030 8678 8658 8730
rect 8710 8678 8722 8730
rect 8774 8678 8786 8730
rect 8838 8678 8850 8730
rect 8902 8678 8914 8730
rect 8966 8678 8978 8730
rect 9030 8678 14658 8730
rect 14710 8678 14722 8730
rect 14774 8678 14786 8730
rect 14838 8678 14850 8730
rect 14902 8678 14914 8730
rect 14966 8678 14978 8730
rect 15030 8678 20658 8730
rect 20710 8678 20722 8730
rect 20774 8678 20786 8730
rect 20838 8678 20850 8730
rect 20902 8678 20914 8730
rect 20966 8678 20978 8730
rect 21030 8678 26658 8730
rect 26710 8678 26722 8730
rect 26774 8678 26786 8730
rect 26838 8678 26850 8730
rect 26902 8678 26914 8730
rect 26966 8678 26978 8730
rect 27030 8678 32658 8730
rect 32710 8678 32722 8730
rect 32774 8678 32786 8730
rect 32838 8678 32850 8730
rect 32902 8678 32914 8730
rect 32966 8678 32978 8730
rect 33030 8678 38658 8730
rect 38710 8678 38722 8730
rect 38774 8678 38786 8730
rect 38838 8678 38850 8730
rect 38902 8678 38914 8730
rect 38966 8678 38978 8730
rect 39030 8678 43884 8730
rect 1104 8656 43884 8678
rect 3053 8619 3111 8625
rect 3053 8585 3065 8619
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 6270 8616 6276 8628
rect 3467 8588 6276 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3068 8548 3096 8579
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 6696 8588 6745 8616
rect 6696 8576 6702 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 14366 8616 14372 8628
rect 6733 8579 6791 8585
rect 6932 8588 14372 8616
rect 5994 8548 6000 8560
rect 3068 8520 6000 8548
rect 5994 8508 6000 8520
rect 6052 8508 6058 8560
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 2884 8412 2912 8443
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5626 8480 5632 8492
rect 5491 8452 5632 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6086 8480 6092 8492
rect 5859 8452 6092 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6932 8489 6960 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 15102 8616 15108 8628
rect 14875 8588 15108 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 16022 8576 16028 8628
rect 16080 8576 16086 8628
rect 16298 8576 16304 8628
rect 16356 8576 16362 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 17586 8616 17592 8628
rect 16816 8588 17592 8616
rect 16816 8576 16822 8588
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17862 8616 17868 8628
rect 17727 8588 17868 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 17957 8619 18015 8625
rect 17957 8585 17969 8619
rect 18003 8616 18015 8619
rect 18414 8616 18420 8628
rect 18003 8588 18420 8616
rect 18003 8585 18015 8588
rect 17957 8579 18015 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 24118 8616 24124 8628
rect 19484 8588 24124 8616
rect 19484 8576 19490 8588
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 24912 8588 27292 8616
rect 24912 8576 24918 8588
rect 7098 8508 7104 8560
rect 7156 8548 7162 8560
rect 7156 8520 9812 8548
rect 7156 8508 7162 8520
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7760 8452 7972 8480
rect 3326 8412 3332 8424
rect 2884 8384 3332 8412
rect 1673 8375 1731 8381
rect 1688 8276 1716 8375
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 4540 8384 7696 8412
rect 2685 8347 2743 8353
rect 2685 8313 2697 8347
rect 2731 8344 2743 8347
rect 3510 8344 3516 8356
rect 2731 8316 3516 8344
rect 2731 8313 2743 8316
rect 2685 8307 2743 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 4540 8353 4568 8384
rect 7668 8356 7696 8384
rect 4525 8347 4583 8353
rect 4080 8316 4476 8344
rect 4080 8276 4108 8316
rect 1688 8248 4108 8276
rect 4154 8236 4160 8288
rect 4212 8236 4218 8288
rect 4448 8276 4476 8316
rect 4525 8313 4537 8347
rect 4571 8313 4583 8347
rect 5534 8344 5540 8356
rect 4525 8307 4583 8313
rect 4816 8316 5540 8344
rect 4816 8276 4844 8316
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5810 8304 5816 8356
rect 5868 8304 5874 8356
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8344 6055 8347
rect 7101 8347 7159 8353
rect 6043 8316 7052 8344
rect 6043 8313 6055 8316
rect 5997 8307 6055 8313
rect 4448 8248 4844 8276
rect 4890 8236 4896 8288
rect 4948 8236 4954 8288
rect 5258 8236 5264 8288
rect 5316 8236 5322 8288
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 5828 8276 5856 8304
rect 5675 8248 5856 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 6822 8276 6828 8288
rect 6144 8248 6828 8276
rect 6144 8236 6150 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 7024 8276 7052 8316
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7190 8344 7196 8356
rect 7147 8316 7196 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 7432 8316 7481 8344
rect 7432 8304 7438 8316
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 7650 8304 7656 8356
rect 7708 8304 7714 8356
rect 7760 8276 7788 8452
rect 7834 8372 7840 8424
rect 7892 8372 7898 8424
rect 7944 8412 7972 8452
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 8294 8412 8300 8424
rect 7944 8384 8300 8412
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8772 8412 8800 8443
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9784 8489 9812 8520
rect 10778 8508 10784 8560
rect 10836 8548 10842 8560
rect 10873 8551 10931 8557
rect 10873 8548 10885 8551
rect 10836 8520 10885 8548
rect 10836 8508 10842 8520
rect 10873 8517 10885 8520
rect 10919 8517 10931 8551
rect 10873 8511 10931 8517
rect 13722 8508 13728 8560
rect 13780 8548 13786 8560
rect 18598 8548 18604 8560
rect 13780 8520 15148 8548
rect 13780 8508 13786 8520
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9364 8452 9413 8480
rect 9364 8440 9370 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 10410 8440 10416 8492
rect 10468 8440 10474 8492
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11793 8483 11851 8489
rect 11793 8480 11805 8483
rect 11204 8452 11805 8480
rect 11204 8440 11210 8452
rect 11793 8449 11805 8452
rect 11839 8480 11851 8483
rect 13173 8483 13231 8489
rect 11839 8452 12434 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 10594 8412 10600 8424
rect 8772 8384 10600 8412
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 10870 8412 10876 8424
rect 10827 8384 10876 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 7852 8285 7880 8372
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8205 8347 8263 8353
rect 8205 8344 8217 8347
rect 8168 8316 8217 8344
rect 8168 8304 8174 8316
rect 8205 8313 8217 8316
rect 8251 8313 8263 8347
rect 8205 8307 8263 8313
rect 8573 8347 8631 8353
rect 8573 8313 8585 8347
rect 8619 8344 8631 8347
rect 9122 8344 9128 8356
rect 8619 8316 9128 8344
rect 8619 8313 8631 8316
rect 8573 8307 8631 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 9585 8347 9643 8353
rect 9585 8344 9597 8347
rect 9548 8316 9597 8344
rect 9548 8304 9554 8316
rect 9585 8313 9597 8316
rect 9631 8313 9643 8347
rect 9585 8307 9643 8313
rect 9950 8304 9956 8356
rect 10008 8304 10014 8356
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 10704 8344 10732 8375
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11480 8384 11529 8412
rect 11480 8372 11486 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 11054 8344 11060 8356
rect 10704 8316 11060 8344
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 7024 8248 7788 8276
rect 7837 8279 7895 8285
rect 7837 8245 7849 8279
rect 7883 8245 7895 8279
rect 7837 8239 7895 8245
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 11146 8276 11152 8288
rect 8904 8248 11152 8276
rect 8904 8236 8910 8248
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 11241 8279 11299 8285
rect 11241 8245 11253 8279
rect 11287 8276 11299 8279
rect 11330 8276 11336 8288
rect 11287 8248 11336 8276
rect 11287 8245 11299 8248
rect 11241 8239 11299 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12406 8276 12434 8452
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13446 8480 13452 8492
rect 13219 8452 13452 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14366 8480 14372 8492
rect 14139 8452 14372 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 15120 8489 15148 8520
rect 16868 8520 18604 8548
rect 15105 8483 15163 8489
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15746 8440 15752 8492
rect 15804 8440 15810 8492
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16482 8440 16488 8492
rect 16540 8440 16546 8492
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8381 12955 8415
rect 16868 8412 16896 8520
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 22281 8551 22339 8557
rect 18800 8520 22232 8548
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17175 8452 17209 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 12897 8375 12955 8381
rect 14292 8384 16896 8412
rect 16945 8415 17003 8421
rect 12529 8347 12587 8353
rect 12529 8313 12541 8347
rect 12575 8344 12587 8347
rect 12802 8344 12808 8356
rect 12575 8316 12808 8344
rect 12575 8313 12587 8316
rect 12529 8307 12587 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 12710 8276 12716 8288
rect 12406 8248 12716 8276
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 12912 8276 12940 8375
rect 14292 8353 14320 8384
rect 16945 8381 16957 8415
rect 16991 8412 17003 8415
rect 17144 8412 17172 8443
rect 17494 8440 17500 8492
rect 17552 8440 17558 8492
rect 17586 8440 17592 8492
rect 17644 8480 17650 8492
rect 17862 8480 17868 8492
rect 17644 8452 17868 8480
rect 17644 8440 17650 8452
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18138 8440 18144 8492
rect 18196 8440 18202 8492
rect 18800 8489 18828 8520
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 19426 8480 19432 8492
rect 18785 8443 18843 8449
rect 18892 8452 19432 8480
rect 18892 8412 18920 8452
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 20070 8480 20076 8492
rect 19935 8452 20076 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 16991 8384 18920 8412
rect 19061 8415 19119 8421
rect 16991 8381 17003 8384
rect 16945 8375 17003 8381
rect 19061 8381 19073 8415
rect 19107 8381 19119 8415
rect 20165 8415 20223 8421
rect 20165 8412 20177 8415
rect 19061 8375 19119 8381
rect 19536 8384 20177 8412
rect 14277 8347 14335 8353
rect 14277 8313 14289 8347
rect 14323 8313 14335 8347
rect 14277 8307 14335 8313
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 15286 8344 15292 8356
rect 14700 8316 15292 8344
rect 14700 8304 14706 8316
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15565 8347 15623 8353
rect 15565 8313 15577 8347
rect 15611 8344 15623 8347
rect 17034 8344 17040 8356
rect 15611 8316 17040 8344
rect 15611 8313 15623 8316
rect 15565 8307 15623 8313
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17313 8347 17371 8353
rect 17313 8313 17325 8347
rect 17359 8344 17371 8347
rect 17770 8344 17776 8356
rect 17359 8316 17776 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 17770 8304 17776 8316
rect 17828 8304 17834 8356
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 19076 8344 19104 8375
rect 18840 8316 19104 8344
rect 18840 8304 18846 8316
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 19300 8316 19441 8344
rect 19300 8304 19306 8316
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 19429 8307 19487 8313
rect 13722 8276 13728 8288
rect 12912 8248 13728 8276
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 13906 8236 13912 8288
rect 13964 8236 13970 8288
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 17586 8276 17592 8288
rect 14516 8248 17592 8276
rect 14516 8236 14522 8248
rect 17586 8236 17592 8248
rect 17644 8236 17650 8288
rect 18322 8236 18328 8288
rect 18380 8276 18386 8288
rect 18874 8276 18880 8288
rect 18380 8248 18880 8276
rect 18380 8236 18386 8248
rect 18874 8236 18880 8248
rect 18932 8276 18938 8288
rect 19536 8276 19564 8384
rect 20165 8381 20177 8384
rect 20211 8381 20223 8415
rect 20165 8375 20223 8381
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 21361 8415 21419 8421
rect 21361 8412 21373 8415
rect 20772 8384 21373 8412
rect 20772 8372 20778 8384
rect 21361 8381 21373 8384
rect 21407 8412 21419 8415
rect 21726 8412 21732 8424
rect 21407 8384 21732 8412
rect 21407 8381 21419 8384
rect 21361 8375 21419 8381
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 19610 8304 19616 8356
rect 19668 8344 19674 8356
rect 21821 8347 21879 8353
rect 21821 8344 21833 8347
rect 19668 8316 21833 8344
rect 19668 8304 19674 8316
rect 21821 8313 21833 8316
rect 21867 8313 21879 8347
rect 22204 8344 22232 8520
rect 22281 8517 22293 8551
rect 22327 8548 22339 8551
rect 23106 8548 23112 8560
rect 22327 8520 23112 8548
rect 22327 8517 22339 8520
rect 22281 8511 22339 8517
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 24026 8508 24032 8560
rect 24084 8548 24090 8560
rect 24762 8548 24768 8560
rect 24084 8520 24768 8548
rect 24084 8508 24090 8520
rect 24762 8508 24768 8520
rect 24820 8508 24826 8560
rect 26234 8508 26240 8560
rect 26292 8548 26298 8560
rect 26513 8551 26571 8557
rect 26513 8548 26525 8551
rect 26292 8520 26525 8548
rect 26292 8508 26298 8520
rect 26513 8517 26525 8520
rect 26559 8517 26571 8551
rect 26513 8511 26571 8517
rect 22465 8483 22523 8489
rect 22465 8449 22477 8483
rect 22511 8480 22523 8483
rect 22830 8480 22836 8492
rect 22511 8452 22836 8480
rect 22511 8449 22523 8452
rect 22465 8443 22523 8449
rect 22830 8440 22836 8452
rect 22888 8440 22894 8492
rect 23382 8440 23388 8492
rect 23440 8440 23446 8492
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 24302 8480 24308 8492
rect 23716 8452 24308 8480
rect 23716 8440 23722 8452
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 25498 8440 25504 8492
rect 25556 8440 25562 8492
rect 25958 8440 25964 8492
rect 26016 8480 26022 8492
rect 27264 8489 27292 8588
rect 27338 8576 27344 8628
rect 27396 8616 27402 8628
rect 42153 8619 42211 8625
rect 27396 8588 42012 8616
rect 27396 8576 27402 8588
rect 28994 8508 29000 8560
rect 29052 8508 29058 8560
rect 29178 8508 29184 8560
rect 29236 8508 29242 8560
rect 29748 8520 31800 8548
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26016 8452 26985 8480
rect 26016 8440 26022 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 28169 8483 28227 8489
rect 28169 8449 28181 8483
rect 28215 8480 28227 8483
rect 28258 8480 28264 8492
rect 28215 8452 28264 8480
rect 28215 8449 28227 8452
rect 28169 8443 28227 8449
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 22646 8372 22652 8424
rect 22704 8412 22710 8424
rect 22741 8415 22799 8421
rect 22741 8412 22753 8415
rect 22704 8384 22753 8412
rect 22704 8372 22710 8384
rect 22741 8381 22753 8384
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 24394 8372 24400 8424
rect 24452 8372 24458 8424
rect 25222 8372 25228 8424
rect 25280 8412 25286 8424
rect 25777 8415 25835 8421
rect 25777 8412 25789 8415
rect 25280 8384 25789 8412
rect 25280 8372 25286 8384
rect 25777 8381 25789 8384
rect 25823 8381 25835 8415
rect 25777 8375 25835 8381
rect 26697 8415 26755 8421
rect 26697 8381 26709 8415
rect 26743 8412 26755 8415
rect 27338 8412 27344 8424
rect 26743 8384 27344 8412
rect 26743 8381 26755 8384
rect 26697 8375 26755 8381
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 27706 8372 27712 8424
rect 27764 8412 27770 8424
rect 27893 8415 27951 8421
rect 27893 8412 27905 8415
rect 27764 8384 27905 8412
rect 27764 8372 27770 8384
rect 27893 8381 27905 8384
rect 27939 8381 27951 8415
rect 27893 8375 27951 8381
rect 28994 8372 29000 8424
rect 29052 8412 29058 8424
rect 29748 8421 29776 8520
rect 29914 8440 29920 8492
rect 29972 8480 29978 8492
rect 30009 8483 30067 8489
rect 30009 8480 30021 8483
rect 29972 8452 30021 8480
rect 29972 8440 29978 8452
rect 30009 8449 30021 8452
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 30098 8440 30104 8492
rect 30156 8480 30162 8492
rect 30156 8452 30420 8480
rect 30156 8440 30162 8452
rect 29733 8415 29791 8421
rect 29733 8412 29745 8415
rect 29052 8384 29745 8412
rect 29052 8372 29058 8384
rect 29733 8381 29745 8384
rect 29779 8381 29791 8415
rect 29733 8375 29791 8381
rect 23106 8344 23112 8356
rect 22204 8316 23112 8344
rect 21821 8307 21879 8313
rect 23106 8304 23112 8316
rect 23164 8304 23170 8356
rect 23198 8304 23204 8356
rect 23256 8344 23262 8356
rect 23256 8316 23888 8344
rect 23256 8304 23262 8316
rect 18932 8248 19564 8276
rect 18932 8236 18938 8248
rect 19702 8236 19708 8288
rect 19760 8276 19766 8288
rect 22002 8276 22008 8288
rect 19760 8248 22008 8276
rect 19760 8236 19766 8248
rect 22002 8236 22008 8248
rect 22060 8236 22066 8288
rect 22189 8279 22247 8285
rect 22189 8245 22201 8279
rect 22235 8276 22247 8279
rect 22830 8276 22836 8288
rect 22235 8248 22836 8276
rect 22235 8245 22247 8248
rect 22189 8239 22247 8245
rect 22830 8236 22836 8248
rect 22888 8236 22894 8288
rect 23860 8276 23888 8316
rect 25332 8316 25544 8344
rect 25332 8276 25360 8316
rect 23860 8248 25360 8276
rect 25406 8236 25412 8288
rect 25464 8236 25470 8288
rect 25516 8276 25544 8316
rect 26528 8316 26740 8344
rect 26528 8276 26556 8316
rect 25516 8248 26556 8276
rect 26712 8276 26740 8316
rect 26878 8304 26884 8356
rect 26936 8344 26942 8356
rect 28905 8347 28963 8353
rect 26936 8316 27384 8344
rect 26936 8304 26942 8316
rect 27246 8276 27252 8288
rect 26712 8248 27252 8276
rect 27246 8236 27252 8248
rect 27304 8236 27310 8288
rect 27356 8276 27384 8316
rect 28905 8313 28917 8347
rect 28951 8344 28963 8347
rect 29546 8344 29552 8356
rect 28951 8316 29552 8344
rect 28951 8313 28963 8316
rect 28905 8307 28963 8313
rect 29546 8304 29552 8316
rect 29604 8304 29610 8356
rect 30392 8344 30420 8452
rect 30742 8440 30748 8492
rect 30800 8480 30806 8492
rect 30837 8483 30895 8489
rect 30837 8480 30849 8483
rect 30800 8452 30849 8480
rect 30800 8440 30806 8452
rect 30837 8449 30849 8452
rect 30883 8449 30895 8483
rect 30837 8443 30895 8449
rect 31772 8412 31800 8520
rect 32030 8508 32036 8560
rect 32088 8548 32094 8560
rect 32217 8551 32275 8557
rect 32217 8548 32229 8551
rect 32088 8520 32229 8548
rect 32088 8508 32094 8520
rect 32217 8517 32229 8520
rect 32263 8517 32275 8551
rect 32217 8511 32275 8517
rect 33134 8508 33140 8560
rect 33192 8548 33198 8560
rect 33192 8520 33548 8548
rect 33192 8508 33198 8520
rect 31846 8440 31852 8492
rect 31904 8480 31910 8492
rect 31941 8483 31999 8489
rect 31941 8480 31953 8483
rect 31904 8452 31953 8480
rect 31904 8440 31910 8452
rect 31941 8449 31953 8452
rect 31987 8449 31999 8483
rect 31941 8443 31999 8449
rect 33318 8440 33324 8492
rect 33376 8480 33382 8492
rect 33413 8483 33471 8489
rect 33413 8480 33425 8483
rect 33376 8452 33425 8480
rect 33376 8440 33382 8452
rect 33413 8449 33425 8452
rect 33459 8449 33471 8483
rect 33520 8480 33548 8520
rect 33594 8508 33600 8560
rect 33652 8548 33658 8560
rect 34333 8551 34391 8557
rect 34333 8548 34345 8551
rect 33652 8520 34345 8548
rect 33652 8508 33658 8520
rect 34333 8517 34345 8520
rect 34379 8517 34391 8551
rect 40218 8548 40224 8560
rect 34333 8511 34391 8517
rect 38856 8520 40224 8548
rect 33873 8483 33931 8489
rect 33873 8480 33885 8483
rect 33520 8452 33885 8480
rect 33413 8443 33471 8449
rect 33873 8449 33885 8452
rect 33919 8449 33931 8483
rect 33873 8443 33931 8449
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 34701 8483 34759 8489
rect 34701 8449 34713 8483
rect 34747 8480 34759 8483
rect 34790 8480 34796 8492
rect 34747 8452 34796 8480
rect 34747 8449 34759 8452
rect 34701 8443 34759 8449
rect 34790 8440 34796 8452
rect 34848 8440 34854 8492
rect 34882 8440 34888 8492
rect 34940 8480 34946 8492
rect 35621 8483 35679 8489
rect 35621 8480 35633 8483
rect 34940 8452 35633 8480
rect 34940 8440 34946 8452
rect 35621 8449 35633 8452
rect 35667 8449 35679 8483
rect 35621 8443 35679 8449
rect 35894 8440 35900 8492
rect 35952 8440 35958 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 36906 8440 36912 8492
rect 36964 8440 36970 8492
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 38470 8440 38476 8492
rect 38528 8440 38534 8492
rect 38856 8489 38884 8520
rect 40218 8508 40224 8520
rect 40276 8508 40282 8560
rect 41782 8548 41788 8560
rect 40880 8520 41788 8548
rect 38841 8483 38899 8489
rect 38841 8449 38853 8483
rect 38887 8449 38899 8483
rect 38841 8443 38899 8449
rect 38933 8483 38991 8489
rect 38933 8449 38945 8483
rect 38979 8480 38991 8483
rect 39390 8480 39396 8492
rect 38979 8452 39396 8480
rect 38979 8449 38991 8452
rect 38933 8443 38991 8449
rect 39390 8440 39396 8452
rect 39448 8440 39454 8492
rect 39574 8440 39580 8492
rect 39632 8440 39638 8492
rect 40880 8489 40908 8520
rect 41782 8508 41788 8520
rect 41840 8508 41846 8560
rect 40129 8483 40187 8489
rect 40129 8449 40141 8483
rect 40175 8449 40187 8483
rect 40129 8443 40187 8449
rect 40497 8483 40555 8489
rect 40497 8449 40509 8483
rect 40543 8449 40555 8483
rect 40497 8443 40555 8449
rect 40865 8483 40923 8489
rect 40865 8449 40877 8483
rect 40911 8449 40923 8483
rect 40865 8443 40923 8449
rect 41233 8483 41291 8489
rect 41233 8449 41245 8483
rect 41279 8480 41291 8483
rect 41414 8480 41420 8492
rect 41279 8452 41420 8480
rect 41279 8449 41291 8452
rect 41233 8443 41291 8449
rect 32950 8412 32956 8424
rect 31772 8384 32956 8412
rect 32950 8372 32956 8384
rect 33008 8372 33014 8424
rect 33689 8415 33747 8421
rect 33689 8381 33701 8415
rect 33735 8412 33747 8415
rect 33962 8412 33968 8424
rect 33735 8384 33968 8412
rect 33735 8381 33747 8384
rect 33689 8375 33747 8381
rect 33962 8372 33968 8384
rect 34020 8372 34026 8424
rect 34974 8372 34980 8424
rect 35032 8372 35038 8424
rect 35066 8372 35072 8424
rect 35124 8412 35130 8424
rect 37553 8415 37611 8421
rect 37553 8412 37565 8415
rect 35124 8384 37565 8412
rect 35124 8372 35130 8384
rect 37553 8381 37565 8384
rect 37599 8381 37611 8415
rect 37553 8375 37611 8381
rect 32677 8347 32735 8353
rect 32677 8344 32689 8347
rect 30392 8316 32689 8344
rect 32677 8313 32689 8316
rect 32723 8313 32735 8347
rect 32677 8307 32735 8313
rect 33778 8304 33784 8356
rect 33836 8344 33842 8356
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 33836 8316 34069 8344
rect 33836 8304 33842 8316
rect 34057 8313 34069 8316
rect 34103 8313 34115 8347
rect 34057 8307 34115 8313
rect 36630 8304 36636 8356
rect 36688 8304 36694 8356
rect 38194 8304 38200 8356
rect 38252 8344 38258 8356
rect 38289 8347 38347 8353
rect 38289 8344 38301 8347
rect 38252 8316 38301 8344
rect 38252 8304 38258 8316
rect 38289 8313 38301 8316
rect 38335 8313 38347 8347
rect 38289 8307 38347 8313
rect 38654 8304 38660 8356
rect 38712 8304 38718 8356
rect 39114 8304 39120 8356
rect 39172 8304 39178 8356
rect 39298 8304 39304 8356
rect 39356 8344 39362 8356
rect 39393 8347 39451 8353
rect 39393 8344 39405 8347
rect 39356 8316 39405 8344
rect 39356 8304 39362 8316
rect 39393 8313 39405 8316
rect 39439 8313 39451 8347
rect 39393 8307 39451 8313
rect 39942 8304 39948 8356
rect 40000 8304 40006 8356
rect 40034 8304 40040 8356
rect 40092 8304 40098 8356
rect 40144 8344 40172 8443
rect 40512 8412 40540 8443
rect 41414 8440 41420 8452
rect 41472 8440 41478 8492
rect 41598 8440 41604 8492
rect 41656 8440 41662 8492
rect 41984 8489 42012 8588
rect 42153 8585 42165 8619
rect 42199 8616 42211 8619
rect 42794 8616 42800 8628
rect 42199 8588 42800 8616
rect 42199 8585 42211 8588
rect 42153 8579 42211 8585
rect 42794 8576 42800 8588
rect 42852 8576 42858 8628
rect 43438 8576 43444 8628
rect 43496 8576 43502 8628
rect 41969 8483 42027 8489
rect 41969 8449 41981 8483
rect 42015 8449 42027 8483
rect 41969 8443 42027 8449
rect 42702 8440 42708 8492
rect 42760 8480 42766 8492
rect 42797 8483 42855 8489
rect 42797 8480 42809 8483
rect 42760 8452 42809 8480
rect 42760 8440 42766 8452
rect 42797 8449 42809 8452
rect 42843 8480 42855 8483
rect 42889 8483 42947 8489
rect 42889 8480 42901 8483
rect 42843 8452 42901 8480
rect 42843 8449 42855 8452
rect 42797 8443 42855 8449
rect 42889 8449 42901 8452
rect 42935 8449 42947 8483
rect 42889 8443 42947 8449
rect 42978 8440 42984 8492
rect 43036 8480 43042 8492
rect 43257 8483 43315 8489
rect 43257 8480 43269 8483
rect 43036 8452 43269 8480
rect 43036 8440 43042 8452
rect 43257 8449 43269 8452
rect 43303 8449 43315 8483
rect 43257 8443 43315 8449
rect 41506 8412 41512 8424
rect 40512 8384 41512 8412
rect 41506 8372 41512 8384
rect 41564 8372 41570 8424
rect 41322 8344 41328 8356
rect 40144 8316 41328 8344
rect 41322 8304 41328 8316
rect 41380 8304 41386 8356
rect 41417 8347 41475 8353
rect 41417 8313 41429 8347
rect 41463 8344 41475 8347
rect 41690 8344 41696 8356
rect 41463 8316 41696 8344
rect 41463 8313 41475 8316
rect 41417 8307 41475 8313
rect 41690 8304 41696 8316
rect 41748 8304 41754 8356
rect 43070 8304 43076 8356
rect 43128 8304 43134 8356
rect 30650 8276 30656 8288
rect 27356 8248 30656 8276
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 30742 8236 30748 8288
rect 30800 8236 30806 8288
rect 30834 8236 30840 8288
rect 30892 8276 30898 8288
rect 31067 8279 31125 8285
rect 31067 8276 31079 8279
rect 30892 8248 31079 8276
rect 30892 8236 30898 8248
rect 31067 8245 31079 8248
rect 31113 8245 31125 8279
rect 31067 8239 31125 8245
rect 31754 8236 31760 8288
rect 31812 8236 31818 8288
rect 32309 8279 32367 8285
rect 32309 8245 32321 8279
rect 32355 8276 32367 8279
rect 33042 8276 33048 8288
rect 32355 8248 33048 8276
rect 32355 8245 32367 8248
rect 32309 8239 32367 8245
rect 33042 8236 33048 8248
rect 33100 8236 33106 8288
rect 36906 8236 36912 8288
rect 36964 8276 36970 8288
rect 37093 8279 37151 8285
rect 37093 8276 37105 8279
rect 36964 8248 37105 8276
rect 36964 8236 36970 8248
rect 37093 8245 37105 8248
rect 37139 8245 37151 8279
rect 40052 8276 40080 8304
rect 40313 8279 40371 8285
rect 40313 8276 40325 8279
rect 40052 8248 40325 8276
rect 37093 8239 37151 8245
rect 40313 8245 40325 8248
rect 40359 8245 40371 8279
rect 40313 8239 40371 8245
rect 40678 8236 40684 8288
rect 40736 8236 40742 8288
rect 41046 8236 41052 8288
rect 41104 8236 41110 8288
rect 41138 8236 41144 8288
rect 41196 8276 41202 8288
rect 42426 8276 42432 8288
rect 41196 8248 42432 8276
rect 41196 8236 41202 8248
rect 42426 8236 42432 8248
rect 42484 8236 42490 8288
rect 1104 8186 43884 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13918 8186
rect 13970 8134 13982 8186
rect 14034 8134 14046 8186
rect 14098 8134 14110 8186
rect 14162 8134 14174 8186
rect 14226 8134 14238 8186
rect 14290 8134 19918 8186
rect 19970 8134 19982 8186
rect 20034 8134 20046 8186
rect 20098 8134 20110 8186
rect 20162 8134 20174 8186
rect 20226 8134 20238 8186
rect 20290 8134 25918 8186
rect 25970 8134 25982 8186
rect 26034 8134 26046 8186
rect 26098 8134 26110 8186
rect 26162 8134 26174 8186
rect 26226 8134 26238 8186
rect 26290 8134 31918 8186
rect 31970 8134 31982 8186
rect 32034 8134 32046 8186
rect 32098 8134 32110 8186
rect 32162 8134 32174 8186
rect 32226 8134 32238 8186
rect 32290 8134 37918 8186
rect 37970 8134 37982 8186
rect 38034 8134 38046 8186
rect 38098 8134 38110 8186
rect 38162 8134 38174 8186
rect 38226 8134 38238 8186
rect 38290 8134 43884 8186
rect 1104 8112 43884 8134
rect 3050 8032 3056 8084
rect 3108 8032 3114 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 5442 8072 5448 8084
rect 3927 8044 5448 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6086 8032 6092 8084
rect 6144 8032 6150 8084
rect 6454 8032 6460 8084
rect 6512 8032 6518 8084
rect 6564 8044 7420 8072
rect 3605 8007 3663 8013
rect 3605 7973 3617 8007
rect 3651 8004 3663 8007
rect 4062 8004 4068 8016
rect 3651 7976 4068 8004
rect 3651 7973 3663 7976
rect 3605 7967 3663 7973
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 5169 8007 5227 8013
rect 5169 7973 5181 8007
rect 5215 8004 5227 8007
rect 5626 8004 5632 8016
rect 5215 7976 5632 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 5718 7964 5724 8016
rect 5776 8004 5782 8016
rect 6564 8004 6592 8044
rect 5776 7976 6592 8004
rect 7392 8004 7420 8044
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7800 8044 8217 8072
rect 7800 8032 7806 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 8570 8032 8576 8084
rect 8628 8032 8634 8084
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 10318 8072 10324 8084
rect 8812 8044 10324 8072
rect 8812 8032 8818 8044
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 15289 8075 15347 8081
rect 10560 8044 15240 8072
rect 10560 8032 10566 8044
rect 8846 8004 8852 8016
rect 7392 7976 8852 8004
rect 5776 7964 5782 7976
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 10597 8007 10655 8013
rect 10597 7973 10609 8007
rect 10643 7973 10655 8007
rect 10597 7967 10655 7973
rect 13357 8007 13415 8013
rect 13357 7973 13369 8007
rect 13403 7973 13415 8007
rect 13357 7967 13415 7973
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 3786 7936 3792 7948
rect 1719 7908 3792 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 3786 7896 3792 7908
rect 3844 7896 3850 7948
rect 3878 7896 3884 7948
rect 3936 7936 3942 7948
rect 5537 7939 5595 7945
rect 3936 7908 4108 7936
rect 3936 7896 3942 7908
rect 1486 7828 1492 7880
rect 1544 7828 1550 7880
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 2314 7828 2320 7880
rect 2372 7868 2378 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2372 7840 2605 7868
rect 2372 7828 2378 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2958 7828 2964 7880
rect 3016 7828 3022 7880
rect 4080 7877 4108 7908
rect 5537 7905 5549 7939
rect 5583 7936 5595 7939
rect 6086 7936 6092 7948
rect 5583 7908 6092 7936
rect 5583 7905 5595 7908
rect 5537 7899 5595 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6362 7936 6368 7948
rect 6288 7908 6368 7936
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4154 7828 4160 7880
rect 4212 7828 4218 7880
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4396 7840 4445 7868
rect 4396 7828 4402 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 6288 7877 6316 7908
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6733 7939 6791 7945
rect 6733 7936 6745 7939
rect 6472 7908 6745 7936
rect 6273 7871 6331 7877
rect 4764 7840 5856 7868
rect 4764 7828 4770 7840
rect 1670 7760 1676 7812
rect 1728 7800 1734 7812
rect 2225 7803 2283 7809
rect 2225 7800 2237 7803
rect 1728 7772 2237 7800
rect 1728 7760 1734 7772
rect 2225 7769 2237 7772
rect 2271 7769 2283 7803
rect 2225 7763 2283 7769
rect 2406 7760 2412 7812
rect 2464 7760 2470 7812
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 3326 7800 3332 7812
rect 2823 7772 3332 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 3418 7760 3424 7812
rect 3476 7760 3482 7812
rect 5353 7803 5411 7809
rect 5353 7769 5365 7803
rect 5399 7800 5411 7803
rect 5442 7800 5448 7812
rect 5399 7772 5448 7800
rect 5399 7769 5411 7772
rect 5353 7763 5411 7769
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7769 5779 7803
rect 5828 7800 5856 7840
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6472 7800 6500 7908
rect 6733 7905 6745 7908
rect 6779 7905 6791 7939
rect 8938 7936 8944 7948
rect 6733 7899 6791 7905
rect 8266 7908 8944 7936
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 7006 7877 7012 7880
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6604 7840 6653 7868
rect 6604 7828 6610 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6996 7871 7012 7877
rect 6996 7837 7008 7871
rect 6996 7831 7012 7837
rect 7006 7828 7012 7831
rect 7064 7828 7070 7880
rect 8266 7868 8294 7908
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 10612 7936 10640 7967
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 10612 7908 11989 7936
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 13372 7936 13400 7967
rect 14458 7936 14464 7948
rect 13372 7908 14464 7936
rect 11977 7899 12035 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 7208 7840 8294 7868
rect 8389 7871 8447 7877
rect 7208 7800 7236 7840
rect 8389 7837 8401 7871
rect 8435 7868 8447 7871
rect 8478 7868 8484 7880
rect 8435 7840 8484 7868
rect 8435 7837 8447 7840
rect 8389 7831 8447 7837
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8754 7828 8760 7880
rect 8812 7828 8818 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 12250 7877 12256 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 9180 7840 9229 7868
rect 9180 7828 9186 7840
rect 9217 7837 9229 7840
rect 9263 7868 9275 7871
rect 11885 7871 11943 7877
rect 9263 7840 11836 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 5828 7772 7236 7800
rect 5721 7763 5779 7769
rect 1857 7735 1915 7741
rect 1857 7701 1869 7735
rect 1903 7732 1915 7735
rect 5166 7732 5172 7744
rect 1903 7704 5172 7732
rect 1903 7701 1915 7704
rect 1857 7695 1915 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 5736 7732 5764 7763
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 11808 7800 11836 7840
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 11931 7840 12204 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12066 7800 12072 7812
rect 7708 7772 10272 7800
rect 11808 7772 12072 7800
rect 7708 7760 7714 7772
rect 5316 7704 5764 7732
rect 5813 7735 5871 7741
rect 5316 7692 5322 7704
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 6270 7732 6276 7744
rect 5859 7704 6276 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 7006 7732 7012 7744
rect 6512 7704 7012 7732
rect 6512 7692 6518 7704
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8570 7732 8576 7744
rect 8352 7704 8576 7732
rect 8352 7692 8358 7704
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 9953 7735 10011 7741
rect 9953 7701 9965 7735
rect 9999 7732 10011 7735
rect 10134 7732 10140 7744
rect 9999 7704 10140 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10244 7732 10272 7772
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 12176 7800 12204 7840
rect 12244 7831 12256 7877
rect 12308 7868 12314 7880
rect 12308 7840 12344 7868
rect 12250 7828 12256 7831
rect 12308 7828 12314 7840
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 13909 7871 13967 7877
rect 12676 7840 13860 7868
rect 12676 7828 12682 7840
rect 12176 7772 13222 7800
rect 12802 7732 12808 7744
rect 10244 7704 12808 7732
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13194 7732 13222 7772
rect 13262 7760 13268 7812
rect 13320 7800 13326 7812
rect 13832 7800 13860 7840
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 14090 7868 14096 7880
rect 13955 7840 14096 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14826 7828 14832 7880
rect 14884 7828 14890 7880
rect 15102 7828 15108 7880
rect 15160 7828 15166 7880
rect 15212 7800 15240 8044
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 15654 8072 15660 8084
rect 15335 8044 15660 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 18414 8072 18420 8084
rect 17460 8044 18420 8072
rect 17460 8032 17466 8044
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 18877 8075 18935 8081
rect 18877 8072 18889 8075
rect 18748 8044 18889 8072
rect 18748 8032 18754 8044
rect 18877 8041 18889 8044
rect 18923 8041 18935 8075
rect 18877 8035 18935 8041
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 19024 8044 19441 8072
rect 19024 8032 19030 8044
rect 19429 8041 19441 8044
rect 19475 8041 19487 8075
rect 19429 8035 19487 8041
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19613 8075 19671 8081
rect 19613 8072 19625 8075
rect 19576 8044 19625 8072
rect 19576 8032 19582 8044
rect 19613 8041 19625 8044
rect 19659 8041 19671 8075
rect 19613 8035 19671 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22097 8075 22155 8081
rect 22097 8072 22109 8075
rect 21968 8044 22109 8072
rect 21968 8032 21974 8044
rect 22097 8041 22109 8044
rect 22143 8041 22155 8075
rect 22097 8035 22155 8041
rect 22554 8032 22560 8084
rect 22612 8072 22618 8084
rect 22612 8044 23244 8072
rect 22612 8032 22618 8044
rect 16577 8007 16635 8013
rect 16577 7973 16589 8007
rect 16623 8004 16635 8007
rect 16758 8004 16764 8016
rect 16623 7976 16764 8004
rect 16623 7973 16635 7976
rect 16577 7967 16635 7973
rect 16758 7964 16764 7976
rect 16816 7964 16822 8016
rect 17862 7964 17868 8016
rect 17920 7964 17926 8016
rect 17972 7976 19472 8004
rect 15378 7896 15384 7948
rect 15436 7936 15442 7948
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 15436 7908 15577 7936
rect 15436 7896 15442 7908
rect 15565 7905 15577 7908
rect 15611 7905 15623 7939
rect 17972 7936 18000 7976
rect 19444 7948 19472 7976
rect 22186 7964 22192 8016
rect 22244 7964 22250 8016
rect 15565 7899 15623 7905
rect 16132 7908 18000 7936
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 15838 7877 15844 7880
rect 15828 7871 15844 7877
rect 15828 7868 15840 7871
rect 15580 7840 15840 7868
rect 15580 7800 15608 7840
rect 15828 7837 15840 7840
rect 15828 7831 15844 7837
rect 15838 7828 15844 7831
rect 15896 7828 15902 7880
rect 13320 7772 13768 7800
rect 13832 7772 14228 7800
rect 15212 7772 15608 7800
rect 13320 7760 13326 7772
rect 13446 7732 13452 7744
rect 13194 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13740 7741 13768 7772
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7701 13783 7735
rect 13725 7695 13783 7701
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13964 7704 14105 7732
rect 13964 7692 13970 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14200 7732 14228 7772
rect 16132 7732 16160 7908
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18656 7908 19288 7936
rect 18656 7896 18662 7908
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17402 7828 17408 7880
rect 17460 7877 17466 7880
rect 17460 7871 17509 7877
rect 17460 7837 17463 7871
rect 17497 7837 17509 7871
rect 17460 7831 17509 7837
rect 17460 7828 17466 7831
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 18322 7828 18328 7880
rect 18380 7828 18386 7880
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 18966 7868 18972 7880
rect 18555 7840 18972 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19058 7828 19064 7880
rect 19116 7828 19122 7880
rect 19260 7877 19288 7908
rect 19426 7896 19432 7948
rect 19484 7896 19490 7948
rect 19518 7896 19524 7948
rect 19576 7936 19582 7948
rect 20993 7939 21051 7945
rect 19576 7908 20392 7936
rect 19576 7896 19582 7908
rect 19245 7871 19303 7877
rect 19245 7837 19257 7871
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19760 7840 19809 7868
rect 19760 7828 19766 7840
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 20364 7868 20392 7908
rect 20993 7905 21005 7939
rect 21039 7936 21051 7939
rect 21082 7936 21088 7948
rect 21039 7908 21088 7936
rect 21039 7905 21051 7908
rect 20993 7899 21051 7905
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 23216 7936 23244 8044
rect 25796 8044 28994 8072
rect 24136 7976 24808 8004
rect 23293 7939 23351 7945
rect 23293 7936 23305 7939
rect 23216 7908 23305 7936
rect 23293 7905 23305 7908
rect 23339 7905 23351 7939
rect 23293 7899 23351 7905
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 20364 7840 20637 7868
rect 19797 7831 19855 7837
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 21174 7868 21180 7880
rect 20947 7840 21180 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7868 21327 7871
rect 21634 7868 21640 7880
rect 21315 7840 21640 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 21910 7828 21916 7880
rect 21968 7828 21974 7880
rect 22922 7828 22928 7880
rect 22980 7828 22986 7880
rect 23198 7828 23204 7880
rect 23256 7828 23262 7880
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 23569 7871 23627 7877
rect 23569 7868 23581 7871
rect 23532 7840 23581 7868
rect 23532 7828 23538 7840
rect 23569 7837 23581 7840
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 24136 7800 24164 7976
rect 24486 7896 24492 7948
rect 24544 7896 24550 7948
rect 24780 7936 24808 7976
rect 25406 7964 25412 8016
rect 25464 8004 25470 8016
rect 25685 8007 25743 8013
rect 25685 8004 25697 8007
rect 25464 7976 25697 8004
rect 25464 7964 25470 7976
rect 25685 7973 25697 7976
rect 25731 7973 25743 8007
rect 25685 7967 25743 7973
rect 25796 7936 25824 8044
rect 26078 7939 26136 7945
rect 26078 7936 26090 7939
rect 24780 7908 26090 7936
rect 26078 7905 26090 7908
rect 26124 7905 26136 7939
rect 26078 7899 26136 7905
rect 26786 7896 26792 7948
rect 26844 7936 26850 7948
rect 26973 7939 27031 7945
rect 26973 7936 26985 7939
rect 26844 7908 26985 7936
rect 26844 7896 26850 7908
rect 26973 7905 26985 7908
rect 27019 7905 27031 7939
rect 28966 7936 28994 8044
rect 29914 8032 29920 8084
rect 29972 8072 29978 8084
rect 32582 8072 32588 8084
rect 29972 8044 32588 8072
rect 29972 8032 29978 8044
rect 32582 8032 32588 8044
rect 32640 8032 32646 8084
rect 34330 8032 34336 8084
rect 34388 8032 34394 8084
rect 34514 8032 34520 8084
rect 34572 8072 34578 8084
rect 34793 8075 34851 8081
rect 34793 8072 34805 8075
rect 34572 8044 34805 8072
rect 34572 8032 34578 8044
rect 34793 8041 34805 8044
rect 34839 8041 34851 8075
rect 37458 8072 37464 8084
rect 34793 8035 34851 8041
rect 35544 8044 37464 8072
rect 30653 8007 30711 8013
rect 30653 7973 30665 8007
rect 30699 8004 30711 8007
rect 30742 8004 30748 8016
rect 30699 7976 30748 8004
rect 30699 7973 30711 7976
rect 30653 7967 30711 7973
rect 30742 7964 30748 7976
rect 30800 7964 30806 8016
rect 31941 8007 31999 8013
rect 31941 7973 31953 8007
rect 31987 7973 31999 8007
rect 31941 7967 31999 7973
rect 30009 7939 30067 7945
rect 30009 7936 30021 7939
rect 28966 7908 30021 7936
rect 26973 7899 27031 7905
rect 30009 7905 30021 7908
rect 30055 7905 30067 7939
rect 30009 7899 30067 7905
rect 24504 7868 24532 7896
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 24504 7840 24777 7868
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 25038 7828 25044 7880
rect 25096 7828 25102 7880
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7868 25283 7871
rect 25406 7868 25412 7880
rect 25271 7840 25412 7868
rect 25271 7837 25283 7840
rect 25225 7831 25283 7837
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 25958 7828 25964 7880
rect 26016 7828 26022 7880
rect 26234 7828 26240 7880
rect 26292 7828 26298 7880
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27614 7868 27620 7880
rect 27295 7840 27620 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 27706 7828 27712 7880
rect 27764 7868 27770 7880
rect 27893 7871 27951 7877
rect 27893 7868 27905 7871
rect 27764 7840 27905 7868
rect 27764 7828 27770 7840
rect 27893 7837 27905 7840
rect 27939 7837 27951 7871
rect 27893 7831 27951 7837
rect 28166 7828 28172 7880
rect 28224 7828 28230 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 28368 7840 29745 7868
rect 18472 7772 24164 7800
rect 18472 7760 18478 7772
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 24489 7803 24547 7809
rect 24489 7800 24501 7803
rect 24268 7772 24501 7800
rect 24268 7760 24274 7772
rect 24489 7769 24501 7772
rect 24535 7769 24547 7803
rect 24489 7763 24547 7769
rect 24578 7760 24584 7812
rect 24636 7800 24642 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 24636 7772 24685 7800
rect 24636 7760 24642 7772
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 26881 7803 26939 7809
rect 26881 7769 26893 7803
rect 26927 7800 26939 7803
rect 28368 7800 28396 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 26927 7772 28396 7800
rect 26927 7769 26939 7772
rect 26881 7763 26939 7769
rect 29178 7760 29184 7812
rect 29236 7760 29242 7812
rect 14200 7704 16160 7732
rect 16669 7735 16727 7741
rect 14093 7695 14151 7701
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 17402 7732 17408 7744
rect 16715 7704 17408 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 18690 7732 18696 7744
rect 17644 7704 18696 7732
rect 17644 7692 17650 7704
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 19794 7692 19800 7744
rect 19852 7732 19858 7744
rect 19889 7735 19947 7741
rect 19889 7732 19901 7735
rect 19852 7704 19901 7732
rect 19852 7692 19858 7704
rect 19889 7701 19901 7704
rect 19935 7701 19947 7735
rect 19889 7695 19947 7701
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 20438 7732 20444 7744
rect 20036 7704 20444 7732
rect 20036 7692 20042 7704
rect 20438 7692 20444 7704
rect 20496 7732 20502 7744
rect 24949 7735 25007 7741
rect 24949 7732 24961 7735
rect 20496 7704 24961 7732
rect 20496 7692 20502 7704
rect 24949 7701 24961 7704
rect 24995 7732 25007 7735
rect 27062 7732 27068 7744
rect 24995 7704 27068 7732
rect 24995 7701 25007 7704
rect 24949 7695 25007 7701
rect 27062 7692 27068 7704
rect 27120 7692 27126 7744
rect 28905 7735 28963 7741
rect 28905 7701 28917 7735
rect 28951 7732 28963 7735
rect 28994 7732 29000 7744
rect 28951 7704 29000 7732
rect 28951 7701 28963 7704
rect 28905 7695 28963 7701
rect 28994 7692 29000 7704
rect 29052 7692 29058 7744
rect 29089 7735 29147 7741
rect 29089 7701 29101 7735
rect 29135 7732 29147 7735
rect 29362 7732 29368 7744
rect 29135 7704 29368 7732
rect 29135 7701 29147 7704
rect 29089 7695 29147 7701
rect 29362 7692 29368 7704
rect 29420 7692 29426 7744
rect 29454 7692 29460 7744
rect 29512 7732 29518 7744
rect 29549 7735 29607 7741
rect 29549 7732 29561 7735
rect 29512 7704 29561 7732
rect 29512 7692 29518 7704
rect 29549 7701 29561 7704
rect 29595 7701 29607 7735
rect 30024 7732 30052 7899
rect 30926 7896 30932 7948
rect 30984 7896 30990 7948
rect 31205 7939 31263 7945
rect 31205 7905 31217 7939
rect 31251 7936 31263 7939
rect 31956 7936 31984 7967
rect 34698 7964 34704 8016
rect 34756 8004 34762 8016
rect 35161 8007 35219 8013
rect 35161 8004 35173 8007
rect 34756 7976 35173 8004
rect 34756 7964 34762 7976
rect 35161 7973 35173 7976
rect 35207 7973 35219 8007
rect 35161 7967 35219 7973
rect 31251 7908 31984 7936
rect 31251 7905 31263 7908
rect 31205 7899 31263 7905
rect 32950 7896 32956 7948
rect 33008 7896 33014 7948
rect 35544 7945 35572 8044
rect 37458 8032 37464 8044
rect 37516 8032 37522 8084
rect 37550 8032 37556 8084
rect 37608 8032 37614 8084
rect 37826 8032 37832 8084
rect 37884 8072 37890 8084
rect 37921 8075 37979 8081
rect 37921 8072 37933 8075
rect 37884 8044 37933 8072
rect 37884 8032 37890 8044
rect 37921 8041 37933 8044
rect 37967 8041 37979 8075
rect 37921 8035 37979 8041
rect 38657 8075 38715 8081
rect 38657 8041 38669 8075
rect 38703 8072 38715 8075
rect 39206 8072 39212 8084
rect 38703 8044 39212 8072
rect 38703 8041 38715 8044
rect 38657 8035 38715 8041
rect 39206 8032 39212 8044
rect 39264 8032 39270 8084
rect 39393 8075 39451 8081
rect 39393 8041 39405 8075
rect 39439 8072 39451 8075
rect 39758 8072 39764 8084
rect 39439 8044 39764 8072
rect 39439 8041 39451 8044
rect 39393 8035 39451 8041
rect 39758 8032 39764 8044
rect 39816 8032 39822 8084
rect 40126 8032 40132 8084
rect 40184 8072 40190 8084
rect 41049 8075 41107 8081
rect 41049 8072 41061 8075
rect 40184 8044 41061 8072
rect 40184 8032 40190 8044
rect 41049 8041 41061 8044
rect 41095 8041 41107 8075
rect 41049 8035 41107 8041
rect 41506 8032 41512 8084
rect 41564 8032 41570 8084
rect 42705 8075 42763 8081
rect 42705 8041 42717 8075
rect 42751 8072 42763 8075
rect 43162 8072 43168 8084
rect 42751 8044 43168 8072
rect 42751 8041 42763 8044
rect 42705 8035 42763 8041
rect 43162 8032 43168 8044
rect 43220 8032 43226 8084
rect 37182 7964 37188 8016
rect 37240 8004 37246 8016
rect 38197 8007 38255 8013
rect 38197 8004 38209 8007
rect 37240 7976 38209 8004
rect 37240 7964 37246 7976
rect 38197 7973 38209 7976
rect 38243 7973 38255 8007
rect 38197 7967 38255 7973
rect 39117 8007 39175 8013
rect 39117 7973 39129 8007
rect 39163 8004 39175 8007
rect 39482 8004 39488 8016
rect 39163 7976 39488 8004
rect 39163 7973 39175 7976
rect 39117 7967 39175 7973
rect 39482 7964 39488 7976
rect 39540 7964 39546 8016
rect 41322 7964 41328 8016
rect 41380 8004 41386 8016
rect 41690 8004 41696 8016
rect 41380 7976 41696 8004
rect 41380 7964 41386 7976
rect 41690 7964 41696 7976
rect 41748 7964 41754 8016
rect 41969 8007 42027 8013
rect 41969 7973 41981 8007
rect 42015 7973 42027 8007
rect 41969 7967 42027 7973
rect 42337 8007 42395 8013
rect 42337 7973 42349 8007
rect 42383 8004 42395 8007
rect 43346 8004 43352 8016
rect 42383 7976 43352 8004
rect 42383 7973 42395 7976
rect 42337 7967 42395 7973
rect 35529 7939 35587 7945
rect 35529 7936 35541 7939
rect 34164 7908 35541 7936
rect 30190 7828 30196 7880
rect 30248 7828 30254 7880
rect 31018 7828 31024 7880
rect 31076 7877 31082 7880
rect 31076 7871 31104 7877
rect 31092 7837 31104 7871
rect 31076 7831 31104 7837
rect 31076 7828 31082 7831
rect 32674 7828 32680 7880
rect 32732 7828 32738 7880
rect 33042 7828 33048 7880
rect 33100 7828 33106 7880
rect 33318 7828 33324 7880
rect 33376 7828 33382 7880
rect 33410 7828 33416 7880
rect 33468 7868 33474 7880
rect 34164 7868 34192 7908
rect 35529 7905 35541 7908
rect 35575 7905 35587 7939
rect 35529 7899 35587 7905
rect 36173 7939 36231 7945
rect 36173 7905 36185 7939
rect 36219 7936 36231 7939
rect 41984 7936 42012 7967
rect 43346 7964 43352 7976
rect 43404 7964 43410 8016
rect 43530 7936 43536 7948
rect 36219 7908 39528 7936
rect 41984 7908 43536 7936
rect 36219 7905 36231 7908
rect 36173 7899 36231 7905
rect 33468 7840 34192 7868
rect 34517 7871 34575 7877
rect 33468 7828 33474 7840
rect 34517 7837 34529 7871
rect 34563 7868 34575 7871
rect 34790 7868 34796 7880
rect 34563 7840 34796 7868
rect 34563 7837 34575 7840
rect 34517 7831 34575 7837
rect 34790 7828 34796 7840
rect 34848 7828 34854 7880
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7868 35035 7871
rect 35158 7868 35164 7880
rect 35023 7840 35164 7868
rect 35023 7837 35035 7840
rect 34977 7831 35035 7837
rect 35158 7828 35164 7840
rect 35216 7828 35222 7880
rect 35342 7828 35348 7880
rect 35400 7828 35406 7880
rect 35710 7828 35716 7880
rect 35768 7828 35774 7880
rect 36446 7828 36452 7880
rect 36504 7828 36510 7880
rect 36538 7828 36544 7880
rect 36596 7877 36602 7880
rect 36596 7871 36624 7877
rect 36612 7837 36624 7871
rect 36596 7831 36624 7837
rect 36596 7828 36602 7831
rect 36722 7828 36728 7880
rect 36780 7828 36786 7880
rect 37737 7871 37795 7877
rect 37737 7837 37749 7871
rect 37783 7868 37795 7871
rect 37826 7868 37832 7880
rect 37783 7840 37832 7868
rect 37783 7837 37795 7840
rect 37737 7831 37795 7837
rect 37826 7828 37832 7840
rect 37884 7828 37890 7880
rect 38105 7871 38163 7877
rect 38105 7837 38117 7871
rect 38151 7868 38163 7871
rect 38841 7871 38899 7877
rect 38151 7840 38792 7868
rect 38151 7837 38163 7840
rect 38105 7831 38163 7837
rect 32030 7800 32036 7812
rect 31772 7772 32036 7800
rect 31772 7732 31800 7772
rect 32030 7760 32036 7772
rect 32088 7760 32094 7812
rect 32122 7760 32128 7812
rect 32180 7800 32186 7812
rect 35434 7800 35440 7812
rect 32180 7772 35440 7800
rect 32180 7760 32186 7772
rect 35434 7760 35440 7772
rect 35492 7760 35498 7812
rect 37369 7803 37427 7809
rect 37369 7769 37381 7803
rect 37415 7800 37427 7803
rect 38381 7803 38439 7809
rect 38381 7800 38393 7803
rect 37415 7772 38393 7800
rect 37415 7769 37427 7772
rect 37369 7763 37427 7769
rect 38381 7769 38393 7772
rect 38427 7769 38439 7803
rect 38381 7763 38439 7769
rect 30024 7704 31800 7732
rect 31849 7735 31907 7741
rect 29549 7695 29607 7701
rect 31849 7701 31861 7735
rect 31895 7732 31907 7735
rect 32306 7732 32312 7744
rect 31895 7704 32312 7732
rect 31895 7701 31907 7704
rect 31849 7695 31907 7701
rect 32306 7692 32312 7704
rect 32364 7692 32370 7744
rect 32674 7692 32680 7744
rect 32732 7732 32738 7744
rect 33318 7732 33324 7744
rect 32732 7704 33324 7732
rect 32732 7692 32738 7704
rect 33318 7692 33324 7704
rect 33376 7692 33382 7744
rect 33870 7692 33876 7744
rect 33928 7732 33934 7744
rect 34057 7735 34115 7741
rect 34057 7732 34069 7735
rect 33928 7704 34069 7732
rect 33928 7692 33934 7704
rect 34057 7701 34069 7704
rect 34103 7701 34115 7735
rect 34057 7695 34115 7701
rect 34146 7692 34152 7744
rect 34204 7732 34210 7744
rect 36446 7732 36452 7744
rect 34204 7704 36452 7732
rect 34204 7692 34210 7704
rect 36446 7692 36452 7704
rect 36504 7692 36510 7744
rect 38764 7732 38792 7840
rect 38841 7837 38853 7871
rect 38887 7837 38899 7871
rect 38841 7831 38899 7837
rect 38933 7871 38991 7877
rect 38933 7837 38945 7871
rect 38979 7868 38991 7871
rect 39114 7868 39120 7880
rect 38979 7840 39120 7868
rect 38979 7837 38991 7840
rect 38933 7831 38991 7837
rect 38856 7800 38884 7831
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39298 7800 39304 7812
rect 38856 7772 39304 7800
rect 39298 7760 39304 7772
rect 39356 7760 39362 7812
rect 39206 7732 39212 7744
rect 38764 7704 39212 7732
rect 39206 7692 39212 7704
rect 39264 7692 39270 7744
rect 39500 7732 39528 7908
rect 43530 7896 43536 7908
rect 43588 7896 43594 7948
rect 39577 7871 39635 7877
rect 39577 7837 39589 7871
rect 39623 7837 39635 7871
rect 39577 7831 39635 7837
rect 39592 7800 39620 7831
rect 39666 7828 39672 7880
rect 39724 7868 39730 7880
rect 39853 7871 39911 7877
rect 39853 7868 39865 7871
rect 39724 7840 39865 7868
rect 39724 7828 39730 7840
rect 39853 7837 39865 7840
rect 39899 7837 39911 7871
rect 39853 7831 39911 7837
rect 40126 7828 40132 7880
rect 40184 7828 40190 7880
rect 41233 7871 41291 7877
rect 41233 7837 41245 7871
rect 41279 7868 41291 7871
rect 41506 7868 41512 7880
rect 41279 7840 41512 7868
rect 41279 7837 41291 7840
rect 41233 7831 41291 7837
rect 41506 7828 41512 7840
rect 41564 7828 41570 7880
rect 41693 7871 41751 7877
rect 41693 7837 41705 7871
rect 41739 7837 41751 7871
rect 41693 7831 41751 7837
rect 41785 7871 41843 7877
rect 41785 7837 41797 7871
rect 41831 7868 41843 7871
rect 41874 7868 41880 7880
rect 41831 7840 41880 7868
rect 41831 7837 41843 7840
rect 41785 7831 41843 7837
rect 40402 7800 40408 7812
rect 39592 7772 40408 7800
rect 40402 7760 40408 7772
rect 40460 7760 40466 7812
rect 41708 7800 41736 7831
rect 41874 7828 41880 7840
rect 41932 7828 41938 7880
rect 42150 7828 42156 7880
rect 42208 7828 42214 7880
rect 42518 7828 42524 7880
rect 42576 7828 42582 7880
rect 42889 7871 42947 7877
rect 42889 7837 42901 7871
rect 42935 7868 42947 7871
rect 42978 7868 42984 7880
rect 42935 7840 42984 7868
rect 42935 7837 42947 7840
rect 42889 7831 42947 7837
rect 42978 7828 42984 7840
rect 43036 7828 43042 7880
rect 43257 7871 43315 7877
rect 43257 7837 43269 7871
rect 43303 7837 43315 7871
rect 43257 7831 43315 7837
rect 41708 7772 42196 7800
rect 42168 7744 42196 7772
rect 42794 7760 42800 7812
rect 42852 7800 42858 7812
rect 43272 7800 43300 7831
rect 42852 7772 43300 7800
rect 42852 7760 42858 7772
rect 40865 7735 40923 7741
rect 40865 7732 40877 7735
rect 39500 7704 40877 7732
rect 40865 7701 40877 7704
rect 40911 7701 40923 7735
rect 40865 7695 40923 7701
rect 42150 7692 42156 7744
rect 42208 7692 42214 7744
rect 43070 7692 43076 7744
rect 43128 7692 43134 7744
rect 43438 7692 43444 7744
rect 43496 7692 43502 7744
rect 1104 7642 43884 7664
rect 1104 7590 2658 7642
rect 2710 7590 2722 7642
rect 2774 7590 2786 7642
rect 2838 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 8658 7642
rect 8710 7590 8722 7642
rect 8774 7590 8786 7642
rect 8838 7590 8850 7642
rect 8902 7590 8914 7642
rect 8966 7590 8978 7642
rect 9030 7590 14658 7642
rect 14710 7590 14722 7642
rect 14774 7590 14786 7642
rect 14838 7590 14850 7642
rect 14902 7590 14914 7642
rect 14966 7590 14978 7642
rect 15030 7590 20658 7642
rect 20710 7590 20722 7642
rect 20774 7590 20786 7642
rect 20838 7590 20850 7642
rect 20902 7590 20914 7642
rect 20966 7590 20978 7642
rect 21030 7590 26658 7642
rect 26710 7590 26722 7642
rect 26774 7590 26786 7642
rect 26838 7590 26850 7642
rect 26902 7590 26914 7642
rect 26966 7590 26978 7642
rect 27030 7590 32658 7642
rect 32710 7590 32722 7642
rect 32774 7590 32786 7642
rect 32838 7590 32850 7642
rect 32902 7590 32914 7642
rect 32966 7590 32978 7642
rect 33030 7590 38658 7642
rect 38710 7590 38722 7642
rect 38774 7590 38786 7642
rect 38838 7590 38850 7642
rect 38902 7590 38914 7642
rect 38966 7590 38978 7642
rect 39030 7590 43884 7642
rect 1104 7568 43884 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2096 7500 6684 7528
rect 2096 7488 2102 7500
rect 2777 7463 2835 7469
rect 2777 7429 2789 7463
rect 2823 7460 2835 7463
rect 3050 7460 3056 7472
rect 2823 7432 3056 7460
rect 2823 7429 2835 7432
rect 2777 7423 2835 7429
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 3142 7420 3148 7472
rect 3200 7420 3206 7472
rect 3329 7463 3387 7469
rect 3329 7429 3341 7463
rect 3375 7460 3387 7463
rect 6656 7460 6684 7500
rect 6730 7488 6736 7540
rect 6788 7488 6794 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 7834 7528 7840 7540
rect 7147 7500 7840 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8202 7528 8208 7540
rect 7975 7500 8208 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 9306 7528 9312 7540
rect 8343 7500 9312 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 9766 7488 9772 7540
rect 9824 7488 9830 7540
rect 10244 7500 10548 7528
rect 10244 7460 10272 7500
rect 3375 7432 6592 7460
rect 6656 7432 10272 7460
rect 10520 7460 10548 7500
rect 11054 7488 11060 7540
rect 11112 7488 11118 7540
rect 11149 7531 11207 7537
rect 11149 7497 11161 7531
rect 11195 7497 11207 7531
rect 11149 7491 11207 7497
rect 11164 7460 11192 7491
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 12860 7500 15792 7528
rect 12860 7488 12866 7500
rect 10520 7432 11192 7460
rect 11624 7432 14044 7460
rect 3375 7429 3387 7432
rect 3329 7423 3387 7429
rect 2406 7352 2412 7404
rect 2464 7352 2470 7404
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 3234 7392 3240 7404
rect 2639 7364 3240 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 4080 7364 4537 7392
rect 1394 7284 1400 7336
rect 1452 7284 1458 7336
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 1762 7324 1768 7336
rect 1719 7296 1768 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 1302 7216 1308 7268
rect 1360 7256 1366 7268
rect 4080 7256 4108 7364
rect 4525 7361 4537 7364
rect 4571 7392 4583 7395
rect 5350 7392 5356 7404
rect 4571 7364 5356 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5460 7364 5641 7392
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 4212 7296 4261 7324
rect 4212 7284 4218 7296
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 5460 7256 5488 7364
rect 5629 7361 5641 7364
rect 5675 7392 5687 7395
rect 5718 7392 5724 7404
rect 5675 7364 5724 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 5810 7352 5816 7404
rect 5868 7352 5874 7404
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 6012 7324 6040 7355
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6454 7324 6460 7336
rect 5592 7296 6460 7324
rect 5592 7284 5598 7296
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 6564 7324 6592 7432
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7392 6975 7395
rect 7006 7392 7012 7404
rect 6963 7364 7012 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7248 7364 7297 7392
rect 7248 7352 7254 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 7524 7364 7665 7392
rect 7524 7352 7530 7364
rect 7653 7361 7665 7364
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8757 7395 8815 7401
rect 8757 7392 8769 7395
rect 8113 7355 8171 7361
rect 8220 7364 8769 7392
rect 6564 7296 7696 7324
rect 1360 7228 4108 7256
rect 5000 7228 5488 7256
rect 1360 7216 1366 7228
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 5000 7188 5028 7228
rect 2915 7160 5028 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 5132 7160 5273 7188
rect 5132 7148 5138 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 6472 7188 6500 7284
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 7469 7259 7527 7265
rect 7469 7256 7481 7259
rect 7340 7228 7481 7256
rect 7340 7216 7346 7228
rect 7469 7225 7481 7228
rect 7515 7225 7527 7259
rect 7668 7256 7696 7296
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 8128 7324 8156 7355
rect 7800 7296 8156 7324
rect 7800 7284 7806 7296
rect 8220 7256 8248 7364
rect 8757 7361 8769 7364
rect 8803 7392 8815 7395
rect 9122 7392 9128 7404
rect 8803 7364 9128 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9582 7392 9588 7404
rect 9364 7364 9588 7392
rect 9364 7352 9370 7364
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9732 7364 9965 7392
rect 9732 7352 9738 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10226 7392 10232 7404
rect 10091 7364 10232 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8352 7296 8493 7324
rect 8352 7284 8358 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 10060 7324 10088 7355
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10318 7352 10324 7404
rect 10376 7396 10382 7404
rect 10376 7392 10456 7396
rect 11054 7392 11060 7404
rect 10376 7368 11060 7392
rect 10376 7352 10382 7368
rect 10428 7364 11060 7368
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 11330 7352 11336 7404
rect 11388 7352 11394 7404
rect 9272 7296 10088 7324
rect 9272 7284 9278 7296
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 10744 7296 11529 7324
rect 10744 7284 10750 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 7668 7228 8248 7256
rect 9140 7228 10180 7256
rect 7469 7219 7527 7225
rect 6822 7188 6828 7200
rect 6472 7160 6828 7188
rect 5261 7151 5319 7157
rect 6822 7148 6828 7160
rect 6880 7188 6886 7200
rect 9140 7188 9168 7228
rect 6880 7160 9168 7188
rect 9493 7191 9551 7197
rect 6880 7148 6886 7160
rect 9493 7157 9505 7191
rect 9539 7188 9551 7191
rect 9674 7188 9680 7200
rect 9539 7160 9680 7188
rect 9539 7157 9551 7160
rect 9493 7151 9551 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10042 7188 10048 7200
rect 9824 7160 10048 7188
rect 9824 7148 9830 7160
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10152 7188 10180 7228
rect 11624 7188 11652 7432
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 12032 7364 13277 7392
rect 12032 7352 12038 7364
rect 13265 7361 13277 7364
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7361 13691 7395
rect 13633 7355 13691 7361
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13648 7324 13676 7355
rect 13722 7352 13728 7404
rect 13780 7352 13786 7404
rect 14016 7401 14044 7432
rect 14090 7420 14096 7472
rect 14148 7460 14154 7472
rect 15654 7460 15660 7472
rect 14148 7432 15660 7460
rect 14148 7420 14154 7432
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14918 7392 14924 7404
rect 14047 7364 14924 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 15764 7392 15792 7500
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 15988 7500 16313 7528
rect 15988 7488 15994 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 17310 7488 17316 7540
rect 17368 7528 17374 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 17368 7500 17693 7528
rect 17368 7488 17374 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 17681 7491 17739 7497
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18690 7528 18696 7540
rect 18472 7500 18696 7528
rect 18472 7488 18478 7500
rect 18690 7488 18696 7500
rect 18748 7528 18754 7540
rect 19153 7531 19211 7537
rect 19153 7528 19165 7531
rect 18748 7500 19165 7528
rect 18748 7488 18754 7500
rect 19153 7497 19165 7500
rect 19199 7497 19211 7531
rect 19153 7491 19211 7497
rect 19702 7488 19708 7540
rect 19760 7488 19766 7540
rect 23845 7531 23903 7537
rect 23845 7528 23857 7531
rect 21376 7500 23857 7528
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 19794 7460 19800 7472
rect 15896 7432 18092 7460
rect 15896 7420 15902 7432
rect 16390 7392 16396 7404
rect 15427 7364 16396 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16574 7392 16580 7404
rect 16531 7364 16580 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17954 7392 17960 7404
rect 17000 7364 17960 7392
rect 17000 7352 17006 7364
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 18064 7401 18092 7432
rect 19076 7432 19800 7460
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 12860 7296 13676 7324
rect 14384 7296 15117 7324
rect 12860 7284 12866 7296
rect 10152 7160 11652 7188
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 13538 7188 13544 7200
rect 13495 7160 13544 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 14384 7188 14412 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15746 7284 15752 7336
rect 15804 7324 15810 7336
rect 15804 7296 16712 7324
rect 15804 7284 15810 7296
rect 16684 7268 16712 7296
rect 17770 7284 17776 7336
rect 17828 7284 17834 7336
rect 19076 7333 19104 7432
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 20438 7352 20444 7404
rect 20496 7401 20502 7404
rect 20496 7395 20545 7401
rect 20496 7361 20499 7395
rect 20533 7361 20545 7395
rect 21376 7392 21404 7500
rect 23845 7497 23857 7500
rect 23891 7497 23903 7531
rect 23845 7491 23903 7497
rect 24118 7488 24124 7540
rect 24176 7528 24182 7540
rect 24394 7528 24400 7540
rect 24176 7500 24400 7528
rect 24176 7488 24182 7500
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 25133 7531 25191 7537
rect 25133 7497 25145 7531
rect 25179 7528 25191 7531
rect 26234 7528 26240 7540
rect 25179 7500 26240 7528
rect 25179 7497 25191 7500
rect 25133 7491 25191 7497
rect 26234 7488 26240 7500
rect 26292 7488 26298 7540
rect 26344 7500 26740 7528
rect 22646 7460 22652 7472
rect 22296 7432 22652 7460
rect 22296 7401 22324 7432
rect 22646 7420 22652 7432
rect 22704 7460 22710 7472
rect 23198 7460 23204 7472
rect 22704 7432 23204 7460
rect 22704 7420 22710 7432
rect 23198 7420 23204 7432
rect 23256 7420 23262 7472
rect 23400 7432 24256 7460
rect 20496 7355 20545 7361
rect 21284 7364 21404 7392
rect 22281 7395 22339 7401
rect 20496 7352 20502 7355
rect 19061 7327 19119 7333
rect 19061 7293 19073 7327
rect 19107 7293 19119 7327
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 19061 7287 19119 7293
rect 19168 7296 20361 7324
rect 15764 7228 16620 7256
rect 13780 7160 14412 7188
rect 14737 7191 14795 7197
rect 13780 7148 13786 7160
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15764 7188 15792 7228
rect 14783 7160 15792 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16117 7191 16175 7197
rect 16117 7188 16129 7191
rect 15896 7160 16129 7188
rect 15896 7148 15902 7160
rect 16117 7157 16129 7160
rect 16163 7157 16175 7191
rect 16592 7188 16620 7228
rect 16666 7216 16672 7268
rect 16724 7216 16730 7268
rect 19168 7256 19196 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 20625 7327 20683 7333
rect 20625 7293 20637 7327
rect 20671 7324 20683 7327
rect 20990 7324 20996 7336
rect 20671 7296 20996 7324
rect 20671 7293 20683 7296
rect 20625 7287 20683 7293
rect 20990 7284 20996 7296
rect 21048 7324 21054 7336
rect 21284 7324 21312 7364
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22370 7352 22376 7404
rect 22428 7352 22434 7404
rect 23285 7395 23343 7401
rect 23285 7392 23297 7395
rect 22526 7364 23297 7392
rect 21048 7296 21312 7324
rect 21361 7327 21419 7333
rect 21048 7284 21054 7296
rect 21361 7293 21373 7327
rect 21407 7293 21419 7327
rect 21361 7287 21419 7293
rect 20901 7259 20959 7265
rect 18708 7228 19196 7256
rect 19536 7228 20024 7256
rect 18708 7188 18736 7228
rect 16592 7160 18736 7188
rect 18785 7191 18843 7197
rect 16117 7151 16175 7157
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 19536 7188 19564 7228
rect 18831 7160 19564 7188
rect 19613 7191 19671 7197
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 19613 7157 19625 7191
rect 19659 7188 19671 7191
rect 19702 7188 19708 7200
rect 19659 7160 19708 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 19996 7188 20024 7228
rect 20901 7225 20913 7259
rect 20947 7225 20959 7259
rect 20901 7219 20959 7225
rect 20438 7188 20444 7200
rect 19996 7160 20444 7188
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20530 7148 20536 7200
rect 20588 7188 20594 7200
rect 20916 7188 20944 7219
rect 20588 7160 20944 7188
rect 21376 7188 21404 7287
rect 21542 7284 21548 7336
rect 21600 7284 21606 7336
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22526 7324 22554 7364
rect 23285 7361 23297 7364
rect 23331 7392 23343 7395
rect 23400 7392 23428 7432
rect 23331 7364 23428 7392
rect 23331 7361 23343 7364
rect 23285 7355 23343 7361
rect 23566 7352 23572 7404
rect 23624 7352 23630 7404
rect 24026 7401 24032 7404
rect 24020 7355 24032 7401
rect 24026 7352 24032 7355
rect 24084 7352 24090 7404
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24228 7392 24256 7432
rect 24486 7420 24492 7472
rect 24544 7460 24550 7472
rect 26344 7460 26372 7500
rect 24544 7432 26372 7460
rect 24544 7420 24550 7432
rect 26418 7420 26424 7472
rect 26476 7460 26482 7472
rect 26605 7463 26663 7469
rect 26605 7460 26617 7463
rect 26476 7432 26617 7460
rect 26476 7420 26482 7432
rect 26605 7429 26617 7432
rect 26651 7429 26663 7463
rect 26712 7460 26740 7500
rect 27062 7488 27068 7540
rect 27120 7528 27126 7540
rect 31757 7531 31815 7537
rect 27120 7500 31156 7528
rect 27120 7488 27126 7500
rect 26789 7463 26847 7469
rect 26789 7460 26801 7463
rect 26712 7432 26801 7460
rect 26605 7423 26663 7429
rect 26789 7429 26801 7432
rect 26835 7460 26847 7463
rect 27246 7460 27252 7472
rect 26835 7432 27252 7460
rect 26835 7429 26847 7432
rect 26789 7423 26847 7429
rect 27246 7420 27252 7432
rect 27304 7420 27310 7472
rect 27982 7420 27988 7472
rect 28040 7460 28046 7472
rect 28077 7463 28135 7469
rect 28077 7460 28089 7463
rect 28040 7432 28089 7460
rect 28040 7420 28046 7432
rect 28077 7429 28089 7432
rect 28123 7429 28135 7463
rect 28077 7423 28135 7429
rect 24397 7395 24455 7401
rect 24397 7392 24409 7395
rect 24228 7364 24409 7392
rect 24397 7361 24409 7364
rect 24443 7392 24455 7395
rect 25501 7395 25559 7401
rect 25501 7392 25513 7395
rect 24443 7364 25513 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 25501 7361 25513 7364
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 26326 7352 26332 7404
rect 26384 7392 26390 7404
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26384 7364 26985 7392
rect 26384 7352 26390 7364
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 27080 7364 27660 7392
rect 22060 7296 22554 7324
rect 22649 7327 22707 7333
rect 22060 7284 22066 7296
rect 22649 7293 22661 7327
rect 22695 7324 22707 7327
rect 22738 7324 22744 7336
rect 22695 7296 22744 7324
rect 22695 7293 22707 7296
rect 22649 7287 22707 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 25225 7327 25283 7333
rect 25225 7324 25237 7327
rect 24780 7296 25237 7324
rect 22097 7259 22155 7265
rect 22097 7225 22109 7259
rect 22143 7256 22155 7259
rect 22370 7256 22376 7268
rect 22143 7228 22376 7256
rect 22143 7225 22155 7228
rect 22097 7219 22155 7225
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 23477 7259 23535 7265
rect 23477 7225 23489 7259
rect 23523 7256 23535 7259
rect 23842 7256 23848 7268
rect 23523 7228 23848 7256
rect 23523 7225 23535 7228
rect 23477 7219 23535 7225
rect 23842 7216 23848 7228
rect 23900 7216 23906 7268
rect 23753 7191 23811 7197
rect 23753 7188 23765 7191
rect 21376 7160 23765 7188
rect 20588 7148 20594 7160
rect 23753 7157 23765 7160
rect 23799 7188 23811 7191
rect 23934 7188 23940 7200
rect 23799 7160 23940 7188
rect 23799 7157 23811 7160
rect 23753 7151 23811 7157
rect 23934 7148 23940 7160
rect 23992 7148 23998 7200
rect 24210 7148 24216 7200
rect 24268 7188 24274 7200
rect 24780 7188 24808 7296
rect 25225 7293 25237 7296
rect 25271 7293 25283 7327
rect 27080 7324 27108 7364
rect 27632 7336 27660 7364
rect 29546 7352 29552 7404
rect 29604 7352 29610 7404
rect 30374 7352 30380 7404
rect 30432 7352 30438 7404
rect 31018 7392 31024 7404
rect 30484 7364 31024 7392
rect 25225 7287 25283 7293
rect 25976 7296 27108 7324
rect 24268 7160 24808 7188
rect 25240 7188 25268 7287
rect 25314 7188 25320 7200
rect 25240 7160 25320 7188
rect 24268 7148 24274 7160
rect 25314 7148 25320 7160
rect 25372 7148 25378 7200
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 25976 7188 26004 7296
rect 27614 7284 27620 7336
rect 27672 7324 27678 7336
rect 28350 7324 28356 7336
rect 27672 7296 28356 7324
rect 27672 7284 27678 7296
rect 28350 7284 28356 7296
rect 28408 7284 28414 7336
rect 28534 7284 28540 7336
rect 28592 7284 28598 7336
rect 28994 7284 29000 7336
rect 29052 7284 29058 7336
rect 29273 7327 29331 7333
rect 29273 7324 29285 7327
rect 29104 7296 29285 7324
rect 26510 7216 26516 7268
rect 26568 7256 26574 7268
rect 29104 7256 29132 7296
rect 29273 7293 29285 7296
rect 29319 7293 29331 7327
rect 29273 7287 29331 7293
rect 29411 7327 29469 7333
rect 29411 7293 29423 7327
rect 29457 7324 29469 7327
rect 29914 7324 29920 7336
rect 29457 7296 29920 7324
rect 29457 7293 29469 7296
rect 29411 7287 29469 7293
rect 29914 7284 29920 7296
rect 29972 7284 29978 7336
rect 30484 7324 30512 7364
rect 31018 7352 31024 7364
rect 31076 7352 31082 7404
rect 30024 7296 30512 7324
rect 30653 7327 30711 7333
rect 26568 7228 29132 7256
rect 26568 7216 26574 7228
rect 25556 7160 26004 7188
rect 26237 7191 26295 7197
rect 25556 7148 25562 7160
rect 26237 7157 26249 7191
rect 26283 7188 26295 7191
rect 26602 7188 26608 7200
rect 26283 7160 26608 7188
rect 26283 7157 26295 7160
rect 26237 7151 26295 7157
rect 26602 7148 26608 7160
rect 26660 7148 26666 7200
rect 27203 7191 27261 7197
rect 27203 7157 27215 7191
rect 27249 7188 27261 7191
rect 27614 7188 27620 7200
rect 27249 7160 27620 7188
rect 27249 7157 27261 7160
rect 27203 7151 27261 7157
rect 27614 7148 27620 7160
rect 27672 7148 27678 7200
rect 27982 7148 27988 7200
rect 28040 7148 28046 7200
rect 28166 7148 28172 7200
rect 28224 7188 28230 7200
rect 28994 7188 29000 7200
rect 28224 7160 29000 7188
rect 28224 7148 28230 7160
rect 28994 7148 29000 7160
rect 29052 7148 29058 7200
rect 29104 7188 29132 7228
rect 30024 7188 30052 7296
rect 30653 7293 30665 7327
rect 30699 7324 30711 7327
rect 30742 7324 30748 7336
rect 30699 7296 30748 7324
rect 30699 7293 30711 7296
rect 30653 7287 30711 7293
rect 30742 7284 30748 7296
rect 30800 7284 30806 7336
rect 31128 7324 31156 7500
rect 31757 7497 31769 7531
rect 31803 7528 31815 7531
rect 31938 7528 31944 7540
rect 31803 7500 31944 7528
rect 31803 7497 31815 7500
rect 31757 7491 31815 7497
rect 31938 7488 31944 7500
rect 31996 7488 32002 7540
rect 32030 7488 32036 7540
rect 32088 7528 32094 7540
rect 32088 7500 33180 7528
rect 32088 7488 32094 7500
rect 33042 7460 33048 7472
rect 32140 7432 33048 7460
rect 31478 7352 31484 7404
rect 31536 7352 31542 7404
rect 31570 7352 31576 7404
rect 31628 7352 31634 7404
rect 31662 7352 31668 7404
rect 31720 7392 31726 7404
rect 32140 7401 32168 7432
rect 33042 7420 33048 7432
rect 33100 7420 33106 7472
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31720 7364 32137 7392
rect 31720 7352 31726 7364
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 32401 7395 32459 7401
rect 32401 7361 32413 7395
rect 32447 7392 32459 7395
rect 32766 7392 32772 7404
rect 32447 7364 32772 7392
rect 32447 7361 32459 7364
rect 32401 7355 32459 7361
rect 32766 7352 32772 7364
rect 32824 7352 32830 7404
rect 33152 7392 33180 7500
rect 33318 7488 33324 7540
rect 33376 7528 33382 7540
rect 35345 7531 35403 7537
rect 33376 7500 35020 7528
rect 33376 7488 33382 7500
rect 34992 7392 35020 7500
rect 35345 7497 35357 7531
rect 35391 7528 35403 7531
rect 35526 7528 35532 7540
rect 35391 7500 35532 7528
rect 35391 7497 35403 7500
rect 35345 7491 35403 7497
rect 35526 7488 35532 7500
rect 35584 7488 35590 7540
rect 36449 7531 36507 7537
rect 36449 7497 36461 7531
rect 36495 7528 36507 7531
rect 36722 7528 36728 7540
rect 36495 7500 36728 7528
rect 36495 7497 36507 7500
rect 36449 7491 36507 7497
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 36909 7531 36967 7537
rect 36909 7497 36921 7531
rect 36955 7528 36967 7531
rect 36998 7528 37004 7540
rect 36955 7500 37004 7528
rect 36955 7497 36967 7500
rect 36909 7491 36967 7497
rect 36998 7488 37004 7500
rect 37056 7488 37062 7540
rect 39298 7488 39304 7540
rect 39356 7528 39362 7540
rect 39356 7500 40172 7528
rect 39356 7488 39362 7500
rect 35069 7463 35127 7469
rect 35069 7429 35081 7463
rect 35115 7460 35127 7463
rect 35115 7432 37136 7460
rect 35115 7429 35127 7432
rect 35069 7423 35127 7429
rect 35161 7395 35219 7401
rect 35161 7392 35173 7395
rect 33152 7364 33548 7392
rect 34992 7364 35173 7392
rect 31128 7296 31754 7324
rect 30098 7216 30104 7268
rect 30156 7256 30162 7268
rect 31297 7259 31355 7265
rect 31297 7256 31309 7259
rect 30156 7228 31309 7256
rect 30156 7216 30162 7228
rect 31297 7225 31309 7228
rect 31343 7225 31355 7259
rect 31726 7256 31754 7296
rect 33042 7284 33048 7336
rect 33100 7324 33106 7336
rect 33229 7327 33287 7333
rect 33229 7324 33241 7327
rect 33100 7296 33241 7324
rect 33100 7284 33106 7296
rect 33229 7293 33241 7296
rect 33275 7293 33287 7327
rect 33229 7287 33287 7293
rect 33413 7327 33471 7333
rect 33413 7293 33425 7327
rect 33459 7293 33471 7327
rect 33413 7287 33471 7293
rect 33428 7256 33456 7287
rect 31726 7228 32260 7256
rect 31297 7219 31355 7225
rect 29104 7160 30052 7188
rect 30193 7191 30251 7197
rect 30193 7157 30205 7191
rect 30239 7188 30251 7191
rect 30558 7188 30564 7200
rect 30239 7160 30564 7188
rect 30239 7157 30251 7160
rect 30193 7151 30251 7157
rect 30558 7148 30564 7160
rect 30616 7148 30622 7200
rect 30926 7148 30932 7200
rect 30984 7188 30990 7200
rect 32122 7188 32128 7200
rect 30984 7160 32128 7188
rect 30984 7148 30990 7160
rect 32122 7148 32128 7160
rect 32180 7148 32186 7200
rect 32232 7188 32260 7228
rect 32784 7228 33456 7256
rect 33520 7256 33548 7364
rect 35161 7361 35173 7364
rect 35207 7361 35219 7395
rect 35161 7355 35219 7361
rect 35250 7352 35256 7404
rect 35308 7392 35314 7404
rect 35713 7395 35771 7401
rect 35713 7392 35725 7395
rect 35308 7364 35725 7392
rect 35308 7352 35314 7364
rect 35713 7361 35725 7364
rect 35759 7392 35771 7395
rect 35759 7364 36216 7392
rect 35759 7361 35771 7364
rect 35713 7355 35771 7361
rect 33870 7284 33876 7336
rect 33928 7284 33934 7336
rect 34146 7324 34152 7336
rect 33980 7296 34152 7324
rect 33980 7256 34008 7296
rect 34146 7284 34152 7296
rect 34204 7284 34210 7336
rect 34238 7284 34244 7336
rect 34296 7333 34302 7336
rect 34296 7327 34324 7333
rect 34312 7293 34324 7327
rect 34296 7287 34324 7293
rect 34296 7284 34302 7287
rect 34422 7284 34428 7336
rect 34480 7284 34486 7336
rect 35437 7327 35495 7333
rect 35437 7324 35449 7327
rect 34900 7296 35449 7324
rect 34900 7268 34928 7296
rect 35437 7293 35449 7296
rect 35483 7293 35495 7327
rect 36188 7324 36216 7364
rect 36262 7352 36268 7404
rect 36320 7392 36326 7404
rect 37108 7401 37136 7432
rect 36817 7395 36875 7401
rect 36817 7392 36829 7395
rect 36320 7364 36829 7392
rect 36320 7352 36326 7364
rect 36817 7361 36829 7364
rect 36863 7361 36875 7395
rect 36817 7355 36875 7361
rect 37093 7395 37151 7401
rect 37093 7361 37105 7395
rect 37139 7361 37151 7395
rect 37553 7395 37611 7401
rect 37553 7392 37565 7395
rect 37093 7355 37151 7361
rect 37200 7364 37565 7392
rect 37200 7324 37228 7364
rect 37553 7361 37565 7364
rect 37599 7392 37611 7395
rect 38746 7392 38752 7404
rect 37599 7364 38752 7392
rect 37599 7361 37611 7364
rect 37553 7355 37611 7361
rect 38746 7352 38752 7364
rect 38804 7352 38810 7404
rect 39298 7352 39304 7404
rect 39356 7352 39362 7404
rect 39482 7401 39488 7404
rect 39439 7395 39488 7401
rect 39439 7361 39451 7395
rect 39485 7361 39488 7395
rect 39439 7355 39488 7361
rect 39482 7352 39488 7355
rect 39540 7352 39546 7404
rect 36188 7296 37228 7324
rect 35437 7287 35495 7293
rect 37274 7284 37280 7336
rect 37332 7284 37338 7336
rect 38378 7284 38384 7336
rect 38436 7284 38442 7336
rect 38565 7327 38623 7333
rect 38565 7293 38577 7327
rect 38611 7293 38623 7327
rect 38565 7287 38623 7293
rect 39577 7327 39635 7333
rect 39577 7293 39589 7327
rect 39623 7324 39635 7327
rect 39623 7296 39988 7324
rect 39623 7293 39635 7296
rect 39577 7287 39635 7293
rect 33520 7228 34008 7256
rect 32784 7188 32812 7228
rect 34882 7216 34888 7268
rect 34940 7216 34946 7268
rect 36354 7216 36360 7268
rect 36412 7256 36418 7268
rect 36633 7259 36691 7265
rect 36633 7256 36645 7259
rect 36412 7228 36645 7256
rect 36412 7216 36418 7228
rect 36633 7225 36645 7228
rect 36679 7256 36691 7259
rect 37295 7256 37323 7284
rect 38580 7256 38608 7287
rect 38654 7256 38660 7268
rect 36679 7228 37323 7256
rect 37936 7228 38660 7256
rect 36679 7225 36691 7228
rect 36633 7219 36691 7225
rect 32232 7160 32812 7188
rect 33137 7191 33195 7197
rect 33137 7157 33149 7191
rect 33183 7188 33195 7191
rect 34422 7188 34428 7200
rect 33183 7160 34428 7188
rect 33183 7157 33195 7160
rect 33137 7151 33195 7157
rect 34422 7148 34428 7160
rect 34480 7148 34486 7200
rect 35434 7148 35440 7200
rect 35492 7188 35498 7200
rect 37936 7188 37964 7228
rect 38654 7216 38660 7228
rect 38712 7216 38718 7268
rect 39022 7216 39028 7268
rect 39080 7216 39086 7268
rect 35492 7160 37964 7188
rect 38289 7191 38347 7197
rect 35492 7148 35498 7160
rect 38289 7157 38301 7191
rect 38335 7188 38347 7191
rect 39960 7188 39988 7296
rect 40144 7256 40172 7500
rect 40310 7488 40316 7540
rect 40368 7528 40374 7540
rect 40405 7531 40463 7537
rect 40405 7528 40417 7531
rect 40368 7500 40417 7528
rect 40368 7488 40374 7500
rect 40405 7497 40417 7500
rect 40451 7497 40463 7531
rect 40405 7491 40463 7497
rect 40678 7488 40684 7540
rect 40736 7488 40742 7540
rect 41782 7488 41788 7540
rect 41840 7528 41846 7540
rect 42061 7531 42119 7537
rect 42061 7528 42073 7531
rect 41840 7500 42073 7528
rect 41840 7488 41846 7500
rect 42061 7497 42073 7500
rect 42107 7497 42119 7531
rect 42061 7491 42119 7497
rect 42705 7531 42763 7537
rect 42705 7497 42717 7531
rect 42751 7528 42763 7531
rect 42886 7528 42892 7540
rect 42751 7500 42892 7528
rect 42751 7497 42763 7500
rect 42705 7491 42763 7497
rect 42886 7488 42892 7500
rect 42944 7488 42950 7540
rect 43073 7531 43131 7537
rect 43073 7497 43085 7531
rect 43119 7528 43131 7531
rect 43254 7528 43260 7540
rect 43119 7500 43260 7528
rect 43119 7497 43131 7500
rect 43073 7491 43131 7497
rect 43254 7488 43260 7500
rect 43312 7488 43318 7540
rect 40221 7463 40279 7469
rect 40221 7429 40233 7463
rect 40267 7460 40279 7463
rect 40267 7432 40908 7460
rect 40267 7429 40279 7432
rect 40221 7423 40279 7429
rect 40880 7401 40908 7432
rect 40589 7395 40647 7401
rect 40589 7361 40601 7395
rect 40635 7361 40647 7395
rect 40589 7355 40647 7361
rect 40865 7395 40923 7401
rect 40865 7361 40877 7395
rect 40911 7361 40923 7395
rect 40865 7355 40923 7361
rect 40604 7324 40632 7355
rect 42242 7352 42248 7404
rect 42300 7352 42306 7404
rect 42426 7352 42432 7404
rect 42484 7392 42490 7404
rect 42521 7395 42579 7401
rect 42521 7392 42533 7395
rect 42484 7364 42533 7392
rect 42484 7352 42490 7364
rect 42521 7361 42533 7364
rect 42567 7361 42579 7395
rect 42521 7355 42579 7361
rect 42886 7352 42892 7404
rect 42944 7352 42950 7404
rect 43257 7395 43315 7401
rect 43257 7361 43269 7395
rect 43303 7361 43315 7395
rect 43257 7355 43315 7361
rect 42334 7324 42340 7336
rect 40604 7296 42340 7324
rect 42334 7284 42340 7296
rect 42392 7284 42398 7336
rect 41966 7256 41972 7268
rect 40144 7228 41972 7256
rect 41966 7216 41972 7228
rect 42024 7216 42030 7268
rect 42058 7216 42064 7268
rect 42116 7256 42122 7268
rect 43272 7256 43300 7355
rect 42116 7228 43300 7256
rect 42116 7216 42122 7228
rect 38335 7160 39988 7188
rect 38335 7157 38347 7160
rect 38289 7151 38347 7157
rect 43438 7148 43444 7200
rect 43496 7148 43502 7200
rect 1104 7098 43884 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13918 7098
rect 13970 7046 13982 7098
rect 14034 7046 14046 7098
rect 14098 7046 14110 7098
rect 14162 7046 14174 7098
rect 14226 7046 14238 7098
rect 14290 7046 19918 7098
rect 19970 7046 19982 7098
rect 20034 7046 20046 7098
rect 20098 7046 20110 7098
rect 20162 7046 20174 7098
rect 20226 7046 20238 7098
rect 20290 7046 25918 7098
rect 25970 7046 25982 7098
rect 26034 7046 26046 7098
rect 26098 7046 26110 7098
rect 26162 7046 26174 7098
rect 26226 7046 26238 7098
rect 26290 7046 31918 7098
rect 31970 7046 31982 7098
rect 32034 7046 32046 7098
rect 32098 7046 32110 7098
rect 32162 7046 32174 7098
rect 32226 7046 32238 7098
rect 32290 7046 37918 7098
rect 37970 7046 37982 7098
rect 38034 7046 38046 7098
rect 38098 7046 38110 7098
rect 38162 7046 38174 7098
rect 38226 7046 38238 7098
rect 38290 7046 43884 7098
rect 1104 7024 43884 7046
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 7834 6984 7840 6996
rect 6052 6956 7840 6984
rect 6052 6944 6058 6956
rect 7834 6944 7840 6956
rect 7892 6984 7898 6996
rect 10226 6984 10232 6996
rect 7892 6956 10232 6984
rect 7892 6944 7898 6956
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 10410 6984 10416 6996
rect 10336 6956 10416 6984
rect 3970 6876 3976 6928
rect 4028 6876 4034 6928
rect 4890 6876 4896 6928
rect 4948 6876 4954 6928
rect 5074 6876 5080 6928
rect 5132 6876 5138 6928
rect 10336 6916 10364 6956
rect 10410 6944 10416 6956
rect 10468 6984 10474 6996
rect 12618 6984 12624 6996
rect 10468 6956 12624 6984
rect 10468 6944 10474 6956
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 13446 6944 13452 6996
rect 13504 6944 13510 6996
rect 19334 6984 19340 6996
rect 13556 6956 19340 6984
rect 10152 6888 10364 6916
rect 1394 6808 1400 6860
rect 1452 6808 1458 6860
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 4338 6848 4344 6860
rect 3007 6820 4344 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4908 6848 4936 6876
rect 4479 6820 4936 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 5350 6848 5356 6860
rect 5224 6820 5356 6848
rect 5224 6808 5230 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5534 6857 5540 6860
rect 5491 6851 5540 6857
rect 5491 6817 5503 6851
rect 5537 6817 5540 6851
rect 5491 6811 5540 6817
rect 5534 6808 5540 6811
rect 5592 6808 5598 6860
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 7742 6848 7748 6860
rect 7340 6820 7748 6848
rect 7340 6808 7346 6820
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 9306 6848 9312 6860
rect 8312 6820 9312 6848
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1719 6752 2268 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2240 6724 2268 6752
rect 2314 6740 2320 6792
rect 2372 6740 2378 6792
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3050 6780 3056 6792
rect 2823 6752 3056 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3292 6752 3801 6780
rect 3292 6740 3298 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 4614 6740 4620 6792
rect 4672 6740 4678 6792
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 2222 6672 2228 6724
rect 2280 6712 2286 6724
rect 3145 6715 3203 6721
rect 3145 6712 3157 6715
rect 2280 6684 3157 6712
rect 2280 6672 2286 6684
rect 3145 6681 3157 6684
rect 3191 6681 3203 6715
rect 3145 6675 3203 6681
rect 3329 6715 3387 6721
rect 3329 6681 3341 6715
rect 3375 6712 3387 6715
rect 4062 6712 4068 6724
rect 3375 6684 4068 6712
rect 3375 6681 3387 6684
rect 3329 6675 3387 6681
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 3160 6644 3188 6675
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 6748 6712 6776 6743
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 6880 6752 8033 6780
rect 6880 6740 6886 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8312 6780 8340 6820
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9836 6851 9894 6857
rect 9836 6817 9848 6851
rect 9882 6848 9894 6851
rect 10152 6848 10180 6888
rect 12158 6876 12164 6928
rect 12216 6876 12222 6928
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 13556 6916 13584 6956
rect 19334 6944 19340 6956
rect 19392 6944 19398 6996
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 27982 6984 27988 6996
rect 19484 6956 27988 6984
rect 19484 6944 19490 6956
rect 27982 6944 27988 6956
rect 28040 6944 28046 6996
rect 28350 6944 28356 6996
rect 28408 6984 28414 6996
rect 30926 6984 30932 6996
rect 28408 6956 30932 6984
rect 28408 6944 28414 6956
rect 30926 6944 30932 6956
rect 30984 6944 30990 6996
rect 31018 6944 31024 6996
rect 31076 6984 31082 6996
rect 32030 6984 32036 6996
rect 31076 6956 32036 6984
rect 31076 6944 31082 6956
rect 32030 6944 32036 6956
rect 32088 6944 32094 6996
rect 32214 6944 32220 6996
rect 32272 6984 32278 6996
rect 32582 6984 32588 6996
rect 32272 6956 32588 6984
rect 32272 6944 32278 6956
rect 32582 6944 32588 6956
rect 32640 6944 32646 6996
rect 33042 6984 33048 6996
rect 32692 6956 33048 6984
rect 12768 6888 13584 6916
rect 12768 6876 12774 6888
rect 18506 6876 18512 6928
rect 18564 6916 18570 6928
rect 19058 6916 19064 6928
rect 18564 6888 19064 6916
rect 18564 6876 18570 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 25409 6919 25467 6925
rect 20364 6888 21588 6916
rect 9882 6820 10180 6848
rect 9882 6817 9894 6820
rect 9836 6811 9894 6817
rect 10226 6808 10232 6860
rect 10284 6808 10290 6860
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10965 6851 11023 6857
rect 10965 6848 10977 6851
rect 10376 6820 10977 6848
rect 10376 6808 10382 6820
rect 10965 6817 10977 6820
rect 11011 6817 11023 6851
rect 10965 6811 11023 6817
rect 8168 6752 8340 6780
rect 8168 6740 8174 6752
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 10560 6752 10701 6780
rect 10560 6740 10566 6752
rect 10689 6749 10701 6752
rect 10735 6780 10747 6783
rect 10778 6780 10784 6792
rect 10735 6752 10784 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6780 10931 6783
rect 11146 6780 11152 6792
rect 10919 6752 11152 6780
rect 10919 6749 10931 6752
rect 10873 6743 10931 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11514 6780 11520 6792
rect 11287 6752 11520 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 12176 6789 12204 6876
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14240 6820 14688 6848
rect 14240 6808 14246 6820
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 14274 6780 14280 6792
rect 13955 6752 14280 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 14660 6789 14688 6820
rect 17678 6808 17684 6860
rect 17736 6808 17742 6860
rect 20364 6848 20392 6888
rect 18432 6820 20392 6848
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14918 6740 14924 6792
rect 14976 6740 14982 6792
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 16850 6780 16856 6792
rect 16807 6752 16856 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 8294 6712 8300 6724
rect 6104 6684 8300 6712
rect 6104 6644 6132 6684
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8772 6684 9260 6712
rect 3160 6616 6132 6644
rect 6273 6647 6331 6653
rect 6273 6613 6285 6647
rect 6319 6644 6331 6647
rect 6362 6644 6368 6656
rect 6319 6616 6368 6644
rect 6319 6613 6331 6616
rect 6273 6607 6331 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 7282 6644 7288 6656
rect 6512 6616 7288 6644
rect 6512 6604 6518 6616
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 8202 6644 8208 6656
rect 7515 6616 8208 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8772 6653 8800 6684
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 9033 6647 9091 6653
rect 9033 6613 9045 6647
rect 9079 6644 9091 6647
rect 9122 6644 9128 6656
rect 9079 6616 9128 6644
rect 9079 6613 9091 6616
rect 9033 6607 9091 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9232 6644 9260 6684
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 16500 6712 16528 6743
rect 16850 6740 16856 6752
rect 16908 6780 16914 6792
rect 17310 6780 17316 6792
rect 16908 6752 17316 6780
rect 16908 6740 16914 6752
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17402 6740 17408 6792
rect 17460 6740 17466 6792
rect 17770 6740 17776 6792
rect 17828 6740 17834 6792
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 18012 6752 18061 6780
rect 18012 6740 18018 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18322 6712 18328 6724
rect 11112 6684 18328 6712
rect 11112 6672 11118 6684
rect 18322 6672 18328 6684
rect 18380 6672 18386 6724
rect 10226 6644 10232 6656
rect 9232 6616 10232 6644
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 11977 6647 12035 6653
rect 11977 6613 11989 6647
rect 12023 6644 12035 6647
rect 12066 6644 12072 6656
rect 12023 6616 12072 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 14734 6644 14740 6656
rect 14415 6616 14740 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 15746 6604 15752 6656
rect 15804 6604 15810 6656
rect 17218 6604 17224 6656
rect 17276 6604 17282 6656
rect 17310 6604 17316 6656
rect 17368 6644 17374 6656
rect 18432 6644 18460 6820
rect 20438 6808 20444 6860
rect 20496 6808 20502 6860
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 20990 6848 20996 6860
rect 20947 6820 20996 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19150 6780 19156 6792
rect 19107 6752 19156 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 19886 6740 19892 6792
rect 19944 6740 19950 6792
rect 19978 6740 19984 6792
rect 20036 6789 20042 6792
rect 20036 6783 20085 6789
rect 20036 6749 20039 6783
rect 20073 6749 20085 6783
rect 20036 6743 20085 6749
rect 20036 6740 20042 6743
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 21085 6783 21143 6789
rect 21085 6749 21097 6783
rect 21131 6780 21143 6783
rect 21358 6780 21364 6792
rect 21131 6752 21364 6780
rect 21131 6749 21143 6752
rect 21085 6743 21143 6749
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 21560 6712 21588 6888
rect 25409 6885 25421 6919
rect 25455 6885 25467 6919
rect 25409 6879 25467 6885
rect 28537 6919 28595 6925
rect 28537 6885 28549 6919
rect 28583 6885 28595 6919
rect 28537 6879 28595 6885
rect 22462 6808 22468 6860
rect 22520 6808 22526 6860
rect 23106 6808 23112 6860
rect 23164 6848 23170 6860
rect 24210 6848 24216 6860
rect 23164 6820 24216 6848
rect 23164 6808 23170 6820
rect 24210 6808 24216 6820
rect 24268 6848 24274 6860
rect 24397 6851 24455 6857
rect 24397 6848 24409 6851
rect 24268 6820 24409 6848
rect 24268 6808 24274 6820
rect 24397 6817 24409 6820
rect 24443 6817 24455 6851
rect 25424 6848 25452 6879
rect 26145 6851 26203 6857
rect 26145 6848 26157 6851
rect 25424 6820 26157 6848
rect 24397 6811 24455 6817
rect 26145 6817 26157 6820
rect 26191 6817 26203 6851
rect 26145 6811 26203 6817
rect 26234 6808 26240 6860
rect 26292 6848 26298 6860
rect 27522 6848 27528 6860
rect 26292 6820 27528 6848
rect 26292 6808 26298 6820
rect 27522 6808 27528 6820
rect 27580 6808 27586 6860
rect 28552 6848 28580 6879
rect 28626 6876 28632 6928
rect 28684 6876 28690 6928
rect 28994 6876 29000 6928
rect 29052 6916 29058 6928
rect 29052 6888 29868 6916
rect 29052 6876 29058 6888
rect 29362 6848 29368 6860
rect 28552 6820 29368 6848
rect 29362 6808 29368 6820
rect 29420 6808 29426 6860
rect 29840 6848 29868 6888
rect 31570 6876 31576 6928
rect 31628 6916 31634 6928
rect 32692 6916 32720 6956
rect 33042 6944 33048 6956
rect 33100 6984 33106 6996
rect 33410 6984 33416 6996
rect 33100 6956 33416 6984
rect 33100 6944 33106 6956
rect 33410 6944 33416 6956
rect 33468 6944 33474 6996
rect 34238 6944 34244 6996
rect 34296 6984 34302 6996
rect 36538 6984 36544 6996
rect 34296 6956 36544 6984
rect 34296 6944 34302 6956
rect 31628 6888 32720 6916
rect 31628 6876 31634 6888
rect 34146 6876 34152 6928
rect 34204 6876 34210 6928
rect 35820 6916 35848 6956
rect 36538 6944 36544 6956
rect 36596 6944 36602 6996
rect 36998 6944 37004 6996
rect 37056 6984 37062 6996
rect 37458 6984 37464 6996
rect 37056 6956 37464 6984
rect 37056 6944 37062 6956
rect 37458 6944 37464 6956
rect 37516 6944 37522 6996
rect 38562 6984 38568 6996
rect 37844 6956 38568 6984
rect 35820 6888 35940 6916
rect 29840 6820 30144 6848
rect 21910 6740 21916 6792
rect 21968 6740 21974 6792
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22204 6712 22232 6743
rect 22738 6740 22744 6792
rect 22796 6740 22802 6792
rect 24670 6740 24676 6792
rect 24728 6740 24734 6792
rect 25498 6740 25504 6792
rect 25556 6740 25562 6792
rect 25590 6740 25596 6792
rect 25648 6780 25654 6792
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25648 6752 25697 6780
rect 25648 6740 25654 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 26418 6740 26424 6792
rect 26476 6740 26482 6792
rect 26510 6740 26516 6792
rect 26568 6789 26574 6792
rect 26568 6783 26596 6789
rect 26584 6749 26596 6783
rect 26568 6743 26596 6749
rect 26568 6740 26574 6743
rect 26694 6740 26700 6792
rect 26752 6740 26758 6792
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6780 27859 6783
rect 28074 6780 28080 6792
rect 27847 6752 28080 6780
rect 27847 6749 27859 6752
rect 27801 6743 27859 6749
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 28813 6783 28871 6789
rect 28813 6749 28825 6783
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 28905 6783 28963 6789
rect 28905 6749 28917 6783
rect 28951 6749 28963 6783
rect 28905 6743 28963 6749
rect 29181 6783 29239 6789
rect 29181 6749 29193 6783
rect 29227 6780 29239 6783
rect 29270 6780 29276 6792
rect 29227 6752 29276 6780
rect 29227 6749 29239 6752
rect 29181 6743 29239 6749
rect 23014 6712 23020 6724
rect 18800 6684 19472 6712
rect 21560 6684 23020 6712
rect 18800 6653 18828 6684
rect 17368 6616 18460 6644
rect 18785 6647 18843 6653
rect 17368 6604 17374 6616
rect 18785 6613 18797 6647
rect 18831 6613 18843 6647
rect 18785 6607 18843 6613
rect 18874 6604 18880 6656
rect 18932 6604 18938 6656
rect 19245 6647 19303 6653
rect 19245 6613 19257 6647
rect 19291 6644 19303 6647
rect 19334 6644 19340 6656
rect 19291 6616 19340 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19444 6644 19472 6684
rect 23014 6672 23020 6684
rect 23072 6672 23078 6724
rect 23106 6672 23112 6724
rect 23164 6712 23170 6724
rect 23164 6684 23612 6712
rect 23164 6672 23170 6684
rect 19886 6644 19892 6656
rect 19444 6616 19892 6644
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 20162 6604 20168 6656
rect 20220 6644 20226 6656
rect 20438 6644 20444 6656
rect 20220 6616 20444 6644
rect 20220 6604 20226 6616
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 20588 6616 21189 6644
rect 20588 6604 20594 6616
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 23198 6644 23204 6656
rect 21784 6616 23204 6644
rect 21784 6604 21790 6616
rect 23198 6604 23204 6616
rect 23256 6604 23262 6656
rect 23474 6604 23480 6656
rect 23532 6604 23538 6656
rect 23584 6644 23612 6684
rect 23658 6672 23664 6724
rect 23716 6712 23722 6724
rect 24688 6712 24716 6740
rect 25608 6712 25636 6740
rect 23716 6684 24716 6712
rect 24780 6684 25636 6712
rect 27341 6715 27399 6721
rect 23716 6672 23722 6684
rect 23934 6644 23940 6656
rect 23584 6616 23940 6644
rect 23934 6604 23940 6616
rect 23992 6644 23998 6656
rect 24780 6644 24808 6684
rect 27341 6681 27353 6715
rect 27387 6712 27399 6715
rect 28828 6712 28856 6743
rect 27387 6684 28856 6712
rect 27387 6681 27399 6684
rect 27341 6675 27399 6681
rect 23992 6616 24808 6644
rect 23992 6604 23998 6616
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 26418 6644 26424 6656
rect 25004 6616 26424 6644
rect 25004 6604 25010 6616
rect 26418 6604 26424 6616
rect 26476 6604 26482 6656
rect 27798 6604 27804 6656
rect 27856 6644 27862 6656
rect 28920 6644 28948 6743
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 29638 6740 29644 6792
rect 29696 6780 29702 6792
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 29696 6752 29745 6780
rect 29696 6740 29702 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 30006 6740 30012 6792
rect 30064 6740 30070 6792
rect 30116 6789 30144 6820
rect 31386 6808 31392 6860
rect 31444 6848 31450 6860
rect 31444 6820 31984 6848
rect 31444 6808 31450 6820
rect 30101 6783 30159 6789
rect 30101 6749 30113 6783
rect 30147 6780 30159 6783
rect 30282 6780 30288 6792
rect 30147 6752 30288 6780
rect 30147 6749 30159 6752
rect 30101 6743 30159 6749
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 30374 6740 30380 6792
rect 30432 6740 30438 6792
rect 30558 6740 30564 6792
rect 30616 6740 30622 6792
rect 30653 6783 30711 6789
rect 30653 6749 30665 6783
rect 30699 6780 30711 6783
rect 30834 6780 30840 6792
rect 30699 6752 30840 6780
rect 30699 6749 30711 6752
rect 30653 6743 30711 6749
rect 30834 6740 30840 6752
rect 30892 6740 30898 6792
rect 30926 6740 30932 6792
rect 30984 6740 30990 6792
rect 31294 6740 31300 6792
rect 31352 6780 31358 6792
rect 31956 6789 31984 6820
rect 32582 6808 32588 6860
rect 32640 6808 32646 6860
rect 33686 6808 33692 6860
rect 33744 6808 33750 6860
rect 31941 6783 31999 6789
rect 31352 6752 31892 6780
rect 31352 6740 31358 6752
rect 28994 6672 29000 6724
rect 29052 6712 29058 6724
rect 30392 6712 30420 6740
rect 29052 6684 29868 6712
rect 29052 6672 29058 6684
rect 27856 6616 28948 6644
rect 29089 6647 29147 6653
rect 27856 6604 27862 6616
rect 29089 6613 29101 6647
rect 29135 6644 29147 6647
rect 29178 6644 29184 6656
rect 29135 6616 29184 6644
rect 29135 6613 29147 6616
rect 29089 6607 29147 6613
rect 29178 6604 29184 6616
rect 29236 6604 29242 6656
rect 29270 6604 29276 6656
rect 29328 6644 29334 6656
rect 29365 6647 29423 6653
rect 29365 6644 29377 6647
rect 29328 6616 29377 6644
rect 29328 6604 29334 6616
rect 29365 6613 29377 6616
rect 29411 6613 29423 6647
rect 29365 6607 29423 6613
rect 29546 6604 29552 6656
rect 29604 6604 29610 6656
rect 29840 6653 29868 6684
rect 30300 6684 30420 6712
rect 30300 6653 30328 6684
rect 31386 6672 31392 6724
rect 31444 6712 31450 6724
rect 31864 6712 31892 6752
rect 31941 6749 31953 6783
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 32217 6783 32275 6789
rect 32217 6749 32229 6783
rect 32263 6780 32275 6783
rect 32306 6780 32312 6792
rect 32263 6752 32312 6780
rect 32263 6749 32275 6752
rect 32217 6743 32275 6749
rect 32306 6740 32312 6752
rect 32364 6740 32370 6792
rect 32490 6740 32496 6792
rect 32548 6740 32554 6792
rect 32861 6783 32919 6789
rect 32861 6749 32873 6783
rect 32907 6749 32919 6783
rect 32861 6743 32919 6749
rect 32876 6712 32904 6743
rect 33226 6740 33232 6792
rect 33284 6780 33290 6792
rect 33965 6783 34023 6789
rect 33965 6780 33977 6783
rect 33284 6752 33977 6780
rect 33284 6740 33290 6752
rect 33965 6749 33977 6752
rect 34011 6749 34023 6783
rect 34164 6780 34192 6876
rect 34606 6808 34612 6860
rect 34664 6848 34670 6860
rect 35912 6857 35940 6888
rect 37550 6876 37556 6928
rect 37608 6916 37614 6928
rect 37737 6919 37795 6925
rect 37737 6916 37749 6919
rect 37608 6888 37749 6916
rect 37608 6876 37614 6888
rect 37737 6885 37749 6888
rect 37783 6885 37795 6919
rect 37737 6879 37795 6885
rect 34701 6851 34759 6857
rect 34701 6848 34713 6851
rect 34664 6820 34713 6848
rect 34664 6808 34670 6820
rect 34701 6817 34713 6820
rect 34747 6817 34759 6851
rect 34701 6811 34759 6817
rect 35897 6851 35955 6857
rect 35897 6817 35909 6851
rect 35943 6817 35955 6851
rect 35897 6811 35955 6817
rect 36078 6808 36084 6860
rect 36136 6808 36142 6860
rect 36538 6808 36544 6860
rect 36596 6808 36602 6860
rect 36630 6808 36636 6860
rect 36688 6848 36694 6860
rect 36998 6857 37004 6860
rect 36817 6851 36875 6857
rect 36817 6848 36829 6851
rect 36688 6820 36829 6848
rect 36688 6808 36694 6820
rect 36817 6817 36829 6820
rect 36863 6817 36875 6851
rect 36817 6811 36875 6817
rect 36955 6851 37004 6857
rect 36955 6817 36967 6851
rect 37001 6817 37004 6851
rect 36955 6811 37004 6817
rect 36998 6808 37004 6811
rect 37056 6808 37062 6860
rect 37274 6808 37280 6860
rect 37332 6848 37338 6860
rect 37844 6857 37872 6956
rect 38562 6944 38568 6956
rect 38620 6944 38626 6996
rect 38841 6987 38899 6993
rect 38841 6953 38853 6987
rect 38887 6984 38899 6987
rect 39022 6984 39028 6996
rect 38887 6956 39028 6984
rect 38887 6953 38899 6956
rect 38841 6947 38899 6953
rect 39022 6944 39028 6956
rect 39080 6944 39086 6996
rect 39206 6944 39212 6996
rect 39264 6984 39270 6996
rect 41138 6984 41144 6996
rect 39264 6956 41144 6984
rect 39264 6944 39270 6956
rect 41138 6944 41144 6956
rect 41196 6944 41202 6996
rect 42058 6984 42064 6996
rect 41386 6956 42064 6984
rect 39393 6919 39451 6925
rect 38672 6888 39344 6916
rect 37829 6851 37887 6857
rect 37829 6848 37841 6851
rect 37332 6820 37841 6848
rect 37332 6808 37338 6820
rect 37829 6817 37841 6820
rect 37875 6817 37887 6851
rect 38672 6848 38700 6888
rect 37829 6811 37887 6817
rect 38488 6820 38700 6848
rect 34977 6783 35035 6789
rect 34977 6780 34989 6783
rect 34164 6752 34989 6780
rect 33965 6743 34023 6749
rect 34977 6749 34989 6752
rect 35023 6749 35035 6783
rect 35802 6756 35808 6808
rect 35860 6756 35866 6808
rect 34977 6743 35035 6749
rect 37090 6740 37096 6792
rect 37148 6740 37154 6792
rect 37734 6740 37740 6792
rect 37792 6780 37798 6792
rect 38105 6783 38163 6789
rect 38105 6780 38117 6783
rect 37792 6752 38117 6780
rect 37792 6740 37798 6752
rect 38105 6749 38117 6752
rect 38151 6780 38163 6783
rect 38488 6780 38516 6820
rect 38746 6808 38752 6860
rect 38804 6848 38810 6860
rect 38804 6820 39252 6848
rect 38804 6808 38810 6820
rect 38151 6752 38516 6780
rect 38151 6749 38163 6752
rect 38105 6743 38163 6749
rect 38562 6740 38568 6792
rect 38620 6780 38626 6792
rect 39224 6789 39252 6820
rect 39117 6783 39175 6789
rect 39117 6780 39129 6783
rect 38620 6752 39129 6780
rect 38620 6740 38626 6752
rect 39117 6749 39129 6752
rect 39163 6749 39175 6783
rect 39117 6743 39175 6749
rect 39209 6783 39267 6789
rect 39209 6749 39221 6783
rect 39255 6749 39267 6783
rect 39316 6780 39344 6888
rect 39393 6885 39405 6919
rect 39439 6885 39451 6919
rect 39393 6879 39451 6885
rect 39669 6919 39727 6925
rect 39669 6885 39681 6919
rect 39715 6885 39727 6919
rect 39669 6879 39727 6885
rect 39408 6848 39436 6879
rect 39408 6820 39620 6848
rect 39485 6783 39543 6789
rect 39485 6780 39497 6783
rect 39316 6752 39497 6780
rect 39209 6743 39267 6749
rect 39485 6749 39497 6752
rect 39531 6749 39543 6783
rect 39485 6743 39543 6749
rect 31444 6684 31800 6712
rect 31864 6684 32076 6712
rect 32876 6684 33272 6712
rect 31444 6672 31450 6684
rect 29825 6647 29883 6653
rect 29825 6613 29837 6647
rect 29871 6613 29883 6647
rect 29825 6607 29883 6613
rect 30285 6647 30343 6653
rect 30285 6613 30297 6647
rect 30331 6613 30343 6647
rect 30285 6607 30343 6613
rect 30377 6647 30435 6653
rect 30377 6613 30389 6647
rect 30423 6644 30435 6647
rect 30558 6644 30564 6656
rect 30423 6616 30564 6644
rect 30423 6613 30435 6616
rect 30377 6607 30435 6613
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 31478 6604 31484 6656
rect 31536 6644 31542 6656
rect 31772 6653 31800 6684
rect 32048 6653 32076 6684
rect 33244 6656 33272 6684
rect 33686 6672 33692 6724
rect 33744 6712 33750 6724
rect 35066 6712 35072 6724
rect 33744 6684 35072 6712
rect 33744 6672 33750 6684
rect 35066 6672 35072 6684
rect 35124 6672 35130 6724
rect 35342 6672 35348 6724
rect 35400 6712 35406 6724
rect 35400 6684 36124 6712
rect 35400 6672 35406 6684
rect 31665 6647 31723 6653
rect 31665 6644 31677 6647
rect 31536 6616 31677 6644
rect 31536 6604 31542 6616
rect 31665 6613 31677 6616
rect 31711 6613 31723 6647
rect 31665 6607 31723 6613
rect 31757 6647 31815 6653
rect 31757 6613 31769 6647
rect 31803 6613 31815 6647
rect 31757 6607 31815 6613
rect 32033 6647 32091 6653
rect 32033 6613 32045 6647
rect 32079 6613 32091 6647
rect 32033 6607 32091 6613
rect 32306 6604 32312 6656
rect 32364 6604 32370 6656
rect 32490 6604 32496 6656
rect 32548 6644 32554 6656
rect 32674 6644 32680 6656
rect 32548 6616 32680 6644
rect 32548 6604 32554 6616
rect 32674 6604 32680 6616
rect 32732 6604 32738 6656
rect 33226 6604 33232 6656
rect 33284 6604 33290 6656
rect 33502 6604 33508 6656
rect 33560 6644 33566 6656
rect 33597 6647 33655 6653
rect 33597 6644 33609 6647
rect 33560 6616 33609 6644
rect 33560 6604 33566 6616
rect 33597 6613 33609 6616
rect 33643 6613 33655 6647
rect 33597 6607 33655 6613
rect 34514 6604 34520 6656
rect 34572 6644 34578 6656
rect 35250 6644 35256 6656
rect 34572 6616 35256 6644
rect 34572 6604 34578 6616
rect 35250 6604 35256 6616
rect 35308 6604 35314 6656
rect 35618 6604 35624 6656
rect 35676 6604 35682 6656
rect 36096 6644 36124 6684
rect 37568 6684 38976 6712
rect 37568 6644 37596 6684
rect 36096 6616 37596 6644
rect 37642 6604 37648 6656
rect 37700 6644 37706 6656
rect 38746 6644 38752 6656
rect 37700 6616 38752 6644
rect 37700 6604 37706 6616
rect 38746 6604 38752 6616
rect 38804 6604 38810 6656
rect 38948 6653 38976 6684
rect 38933 6647 38991 6653
rect 38933 6613 38945 6647
rect 38979 6613 38991 6647
rect 39500 6644 39528 6743
rect 39592 6712 39620 6820
rect 39684 6780 39712 6879
rect 39850 6876 39856 6928
rect 39908 6916 39914 6928
rect 41386 6916 41414 6956
rect 42058 6944 42064 6956
rect 42116 6944 42122 6996
rect 42334 6944 42340 6996
rect 42392 6944 42398 6996
rect 39908 6888 41414 6916
rect 39908 6876 39914 6888
rect 39758 6808 39764 6860
rect 39816 6848 39822 6860
rect 41874 6848 41880 6860
rect 39816 6820 41880 6848
rect 39816 6808 39822 6820
rect 41874 6808 41880 6820
rect 41932 6808 41938 6860
rect 39684 6752 41414 6780
rect 41386 6712 41414 6752
rect 41690 6740 41696 6792
rect 41748 6780 41754 6792
rect 42521 6783 42579 6789
rect 42521 6780 42533 6783
rect 41748 6752 42533 6780
rect 41748 6740 41754 6752
rect 42521 6749 42533 6752
rect 42567 6749 42579 6783
rect 42521 6743 42579 6749
rect 42702 6740 42708 6792
rect 42760 6740 42766 6792
rect 43165 6783 43223 6789
rect 43165 6749 43177 6783
rect 43211 6780 43223 6783
rect 43257 6783 43315 6789
rect 43257 6780 43269 6783
rect 43211 6752 43269 6780
rect 43211 6749 43223 6752
rect 43165 6743 43223 6749
rect 43257 6749 43269 6752
rect 43303 6749 43315 6783
rect 43257 6743 43315 6749
rect 42978 6712 42984 6724
rect 39592 6684 40448 6712
rect 41386 6684 42984 6712
rect 40126 6644 40132 6656
rect 39500 6616 40132 6644
rect 38933 6607 38991 6613
rect 40126 6604 40132 6616
rect 40184 6604 40190 6656
rect 40420 6644 40448 6684
rect 42978 6672 42984 6684
rect 43036 6672 43042 6724
rect 43070 6672 43076 6724
rect 43128 6672 43134 6724
rect 42794 6644 42800 6656
rect 40420 6616 42800 6644
rect 42794 6604 42800 6616
rect 42852 6604 42858 6656
rect 42886 6604 42892 6656
rect 42944 6604 42950 6656
rect 43438 6604 43444 6656
rect 43496 6604 43502 6656
rect 1104 6554 43884 6576
rect 1104 6502 2658 6554
rect 2710 6502 2722 6554
rect 2774 6502 2786 6554
rect 2838 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 8658 6554
rect 8710 6502 8722 6554
rect 8774 6502 8786 6554
rect 8838 6502 8850 6554
rect 8902 6502 8914 6554
rect 8966 6502 8978 6554
rect 9030 6502 14658 6554
rect 14710 6502 14722 6554
rect 14774 6502 14786 6554
rect 14838 6502 14850 6554
rect 14902 6502 14914 6554
rect 14966 6502 14978 6554
rect 15030 6502 20658 6554
rect 20710 6502 20722 6554
rect 20774 6502 20786 6554
rect 20838 6502 20850 6554
rect 20902 6502 20914 6554
rect 20966 6502 20978 6554
rect 21030 6502 26658 6554
rect 26710 6502 26722 6554
rect 26774 6502 26786 6554
rect 26838 6502 26850 6554
rect 26902 6502 26914 6554
rect 26966 6502 26978 6554
rect 27030 6502 32658 6554
rect 32710 6502 32722 6554
rect 32774 6502 32786 6554
rect 32838 6502 32850 6554
rect 32902 6502 32914 6554
rect 32966 6502 32978 6554
rect 33030 6502 38658 6554
rect 38710 6502 38722 6554
rect 38774 6502 38786 6554
rect 38838 6502 38850 6554
rect 38902 6502 38914 6554
rect 38966 6502 38978 6554
rect 39030 6502 43884 6554
rect 1104 6480 43884 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3418 6440 3424 6452
rect 2832 6412 3424 6440
rect 2832 6400 2838 6412
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 5810 6440 5816 6452
rect 3660 6412 5816 6440
rect 3660 6400 3666 6412
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 5960 6412 6561 6440
rect 5960 6400 5966 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6696 6412 6745 6440
rect 6696 6400 6702 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 8754 6440 8760 6452
rect 6733 6403 6791 6409
rect 6932 6412 8760 6440
rect 6454 6372 6460 6384
rect 5184 6344 6460 6372
rect 5184 6316 5212 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 1670 6304 1676 6316
rect 1535 6276 1676 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 2958 6304 2964 6316
rect 1820 6276 2964 6304
rect 1820 6264 1826 6276
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2464 6208 2605 6236
rect 2464 6196 2470 6208
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 2774 6196 2780 6248
rect 2832 6196 2838 6248
rect 3510 6230 3516 6282
rect 3568 6230 3574 6282
rect 3602 6264 3608 6316
rect 3660 6314 3666 6316
rect 3660 6313 3673 6314
rect 3660 6307 3688 6313
rect 3676 6273 3688 6307
rect 3660 6267 3688 6273
rect 3660 6264 3666 6267
rect 3786 6264 3792 6316
rect 3844 6264 3850 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 4479 6276 4537 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 5718 6304 5724 6316
rect 5491 6276 5724 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6932 6313 6960 6412
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9309 6443 9367 6449
rect 9309 6440 9321 6443
rect 9272 6412 9321 6440
rect 9272 6400 9278 6412
rect 9309 6409 9321 6412
rect 9355 6409 9367 6443
rect 9309 6403 9367 6409
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 9950 6440 9956 6452
rect 9640 6412 9956 6440
rect 9640 6400 9646 6412
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10502 6440 10508 6452
rect 10100 6412 10508 6440
rect 10100 6400 10106 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 13630 6440 13636 6452
rect 13495 6412 13636 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13814 6400 13820 6452
rect 13872 6400 13878 6452
rect 18874 6440 18880 6452
rect 14016 6412 18880 6440
rect 9140 6372 9168 6400
rect 10226 6372 10232 6384
rect 9140 6344 10232 6372
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10520 6372 10548 6400
rect 14016 6372 14044 6412
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19242 6400 19248 6452
rect 19300 6400 19306 6452
rect 20346 6440 20352 6452
rect 19444 6412 20352 6440
rect 10520 6344 14044 6372
rect 14274 6332 14280 6384
rect 14332 6332 14338 6384
rect 14918 6332 14924 6384
rect 14976 6372 14982 6384
rect 17034 6372 17040 6384
rect 14976 6344 17040 6372
rect 14976 6332 14982 6344
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 17310 6332 17316 6384
rect 17368 6372 17374 6384
rect 17678 6372 17684 6384
rect 17368 6344 17684 6372
rect 17368 6332 17374 6344
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 17770 6332 17776 6384
rect 17828 6372 17834 6384
rect 18046 6372 18052 6384
rect 17828 6344 18052 6372
rect 17828 6332 17834 6344
rect 18046 6332 18052 6344
rect 18104 6372 18110 6384
rect 18782 6372 18788 6384
rect 18104 6344 18788 6372
rect 18104 6332 18110 6344
rect 18782 6332 18788 6344
rect 18840 6332 18846 6384
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7650 6264 7656 6316
rect 7708 6264 7714 6316
rect 7926 6264 7932 6316
rect 7984 6264 7990 6316
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 9033 6307 9091 6313
rect 8711 6276 8984 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 3513 6205 3525 6230
rect 3559 6205 3571 6230
rect 3513 6199 3571 6205
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 7791 6239 7849 6245
rect 7791 6236 7803 6239
rect 5868 6208 7803 6236
rect 5868 6196 5874 6208
rect 7791 6205 7803 6208
rect 7837 6236 7849 6239
rect 7837 6208 8156 6236
rect 7837 6205 7849 6208
rect 7791 6199 7849 6205
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3237 6171 3295 6177
rect 3237 6168 3249 6171
rect 3108 6140 3249 6168
rect 3108 6128 3114 6140
rect 3237 6137 3249 6140
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 4522 6128 4528 6180
rect 4580 6168 4586 6180
rect 4709 6171 4767 6177
rect 4709 6168 4721 6171
rect 4580 6140 4721 6168
rect 4580 6128 4586 6140
rect 4709 6137 4721 6140
rect 4755 6137 4767 6171
rect 4709 6131 4767 6137
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6100 2559 6103
rect 3326 6100 3332 6112
rect 2547 6072 3332 6100
rect 2547 6069 2559 6072
rect 2501 6063 2559 6069
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 6362 6100 6368 6112
rect 6227 6072 6368 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7834 6100 7840 6112
rect 7055 6072 7840 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8128 6100 8156 6208
rect 8202 6196 8208 6248
rect 8260 6196 8266 6248
rect 8294 6196 8300 6248
rect 8352 6196 8358 6248
rect 8846 6196 8852 6248
rect 8904 6196 8910 6248
rect 8956 6236 8984 6276
rect 9033 6273 9045 6307
rect 9079 6304 9091 6307
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 9079 6276 9137 6304
rect 9079 6273 9091 6276
rect 9033 6267 9091 6273
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 10686 6304 10692 6316
rect 9815 6276 10692 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 11077 6307 11135 6313
rect 11077 6273 11089 6307
rect 11123 6304 11135 6307
rect 11238 6304 11244 6316
rect 11123 6276 11244 6304
rect 11123 6273 11135 6276
rect 11077 6267 11135 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 13633 6307 13691 6313
rect 13633 6304 13645 6307
rect 13596 6276 13645 6304
rect 13596 6264 13602 6276
rect 13633 6273 13645 6276
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14001 6307 14059 6313
rect 14001 6304 14013 6307
rect 13872 6276 14013 6304
rect 13872 6264 13878 6276
rect 14001 6273 14013 6276
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 14182 6264 14188 6316
rect 14240 6304 14246 6316
rect 17586 6304 17592 6316
rect 14240 6276 17592 6304
rect 14240 6264 14246 6276
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17696 6304 17724 6332
rect 19444 6313 19472 6412
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 23658 6440 23664 6452
rect 20496 6412 23664 6440
rect 20496 6400 20502 6412
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 23750 6400 23756 6452
rect 23808 6400 23814 6452
rect 23860 6412 24992 6440
rect 19518 6332 19524 6384
rect 19576 6372 19582 6384
rect 19978 6372 19984 6384
rect 19576 6344 19984 6372
rect 19576 6332 19582 6344
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 22922 6332 22928 6384
rect 22980 6372 22986 6384
rect 23860 6372 23888 6412
rect 22980 6344 23888 6372
rect 24029 6375 24087 6381
rect 22980 6332 22986 6344
rect 24029 6341 24041 6375
rect 24075 6372 24087 6375
rect 24397 6375 24455 6381
rect 24397 6372 24409 6375
rect 24075 6344 24409 6372
rect 24075 6341 24087 6344
rect 24029 6335 24087 6341
rect 24397 6341 24409 6344
rect 24443 6341 24455 6375
rect 24397 6335 24455 6341
rect 24581 6375 24639 6381
rect 24581 6341 24593 6375
rect 24627 6372 24639 6375
rect 24854 6372 24860 6384
rect 24627 6344 24860 6372
rect 24627 6341 24639 6344
rect 24581 6335 24639 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 24964 6372 24992 6412
rect 25038 6400 25044 6452
rect 25096 6440 25102 6452
rect 26510 6440 26516 6452
rect 25096 6412 26516 6440
rect 25096 6400 25102 6412
rect 26510 6400 26516 6412
rect 26568 6440 26574 6452
rect 29914 6440 29920 6452
rect 26568 6412 29920 6440
rect 26568 6400 26574 6412
rect 29914 6400 29920 6412
rect 29972 6440 29978 6452
rect 31386 6440 31392 6452
rect 29972 6412 31392 6440
rect 29972 6400 29978 6412
rect 31386 6400 31392 6412
rect 31444 6400 31450 6452
rect 31665 6443 31723 6449
rect 31665 6409 31677 6443
rect 31711 6440 31723 6443
rect 36909 6443 36967 6449
rect 31711 6412 35020 6440
rect 31711 6409 31723 6412
rect 31665 6403 31723 6409
rect 27154 6372 27160 6384
rect 24964 6344 25452 6372
rect 17865 6307 17923 6313
rect 17865 6304 17877 6307
rect 17696 6276 17877 6304
rect 17865 6273 17877 6276
rect 17911 6273 17923 6307
rect 19429 6307 19487 6313
rect 17865 6267 17923 6273
rect 18248 6276 19196 6304
rect 10042 6236 10048 6248
rect 8956 6208 10048 6236
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6205 11391 6239
rect 11333 6199 11391 6205
rect 8312 6168 8340 6196
rect 11348 6168 11376 6199
rect 11514 6196 11520 6248
rect 11572 6236 11578 6248
rect 16942 6236 16948 6248
rect 11572 6208 16948 6236
rect 11572 6196 11578 6208
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 8312 6140 10456 6168
rect 11348 6140 15577 6168
rect 8938 6100 8944 6112
rect 8128 6072 8944 6100
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6100 9091 6103
rect 9214 6100 9220 6112
rect 9079 6072 9220 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 9582 6060 9588 6112
rect 9640 6060 9646 6112
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 9916 6072 9965 6100
rect 9916 6060 9922 6072
rect 9953 6069 9965 6072
rect 9999 6069 10011 6103
rect 10428 6100 10456 6140
rect 15565 6137 15577 6140
rect 15611 6137 15623 6171
rect 15565 6131 15623 6137
rect 11514 6100 11520 6112
rect 10428 6072 11520 6100
rect 9953 6063 10011 6069
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12618 6100 12624 6112
rect 11848 6072 12624 6100
rect 11848 6060 11854 6072
rect 12618 6060 12624 6072
rect 12676 6100 12682 6112
rect 17310 6100 17316 6112
rect 12676 6072 17316 6100
rect 12676 6060 12682 6072
rect 17310 6060 17316 6072
rect 17368 6060 17374 6112
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 18248 6100 18276 6276
rect 19168 6248 19196 6276
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19610 6264 19616 6316
rect 19668 6264 19674 6316
rect 19702 6264 19708 6316
rect 19760 6264 19766 6316
rect 19794 6264 19800 6316
rect 19852 6264 19858 6316
rect 20714 6264 20720 6316
rect 20772 6264 20778 6316
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6304 21879 6307
rect 21910 6304 21916 6316
rect 21867 6276 21916 6304
rect 21867 6273 21879 6276
rect 21821 6267 21879 6273
rect 21910 6264 21916 6276
rect 21968 6264 21974 6316
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 23474 6264 23480 6316
rect 23532 6304 23538 6316
rect 23750 6304 23756 6316
rect 23532 6276 23756 6304
rect 23532 6264 23538 6276
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 23934 6264 23940 6316
rect 23992 6264 23998 6316
rect 24118 6264 24124 6316
rect 24176 6264 24182 6316
rect 24305 6307 24363 6313
rect 24305 6273 24317 6307
rect 24351 6273 24363 6307
rect 24305 6267 24363 6273
rect 18322 6196 18328 6248
rect 18380 6236 18386 6248
rect 18380 6208 19104 6236
rect 18380 6196 18386 6208
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 18969 6171 19027 6177
rect 18969 6168 18981 6171
rect 18840 6140 18981 6168
rect 18840 6128 18846 6140
rect 18969 6137 18981 6140
rect 19015 6137 19027 6171
rect 19076 6168 19104 6208
rect 19150 6196 19156 6248
rect 19208 6236 19214 6248
rect 19628 6236 19656 6264
rect 19208 6208 19656 6236
rect 19208 6196 19214 6208
rect 19978 6196 19984 6248
rect 20036 6196 20042 6248
rect 20346 6196 20352 6248
rect 20404 6196 20410 6248
rect 20898 6245 20904 6248
rect 20855 6239 20904 6245
rect 20855 6205 20867 6239
rect 20901 6205 20904 6239
rect 20855 6199 20904 6205
rect 20898 6196 20904 6199
rect 20956 6196 20962 6248
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6236 21051 6239
rect 21174 6236 21180 6248
rect 21039 6208 21180 6236
rect 21039 6205 21051 6208
rect 20993 6199 21051 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 22738 6236 22744 6248
rect 21692 6208 22744 6236
rect 21692 6196 21698 6208
rect 22738 6196 22744 6208
rect 22796 6196 22802 6248
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6236 23627 6239
rect 24320 6236 24348 6267
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 25424 6313 25452 6344
rect 26344 6344 27160 6372
rect 24765 6307 24823 6313
rect 24765 6304 24777 6307
rect 24728 6276 24777 6304
rect 24728 6264 24734 6276
rect 24765 6273 24777 6276
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 25409 6307 25467 6313
rect 25409 6273 25421 6307
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 26237 6307 26295 6313
rect 26237 6273 26249 6307
rect 26283 6304 26295 6307
rect 26344 6304 26372 6344
rect 27154 6332 27160 6344
rect 27212 6332 27218 6384
rect 27522 6332 27528 6384
rect 27580 6372 27586 6384
rect 30742 6372 30748 6384
rect 27580 6344 28212 6372
rect 27580 6332 27586 6344
rect 28184 6316 28212 6344
rect 30024 6344 30748 6372
rect 26283 6276 26372 6304
rect 26283 6273 26295 6276
rect 26237 6267 26295 6273
rect 26418 6264 26424 6316
rect 26476 6304 26482 6316
rect 26605 6307 26663 6313
rect 26605 6304 26617 6307
rect 26476 6276 26617 6304
rect 26476 6264 26482 6276
rect 26605 6273 26617 6276
rect 26651 6304 26663 6307
rect 27430 6304 27436 6316
rect 26651 6276 27436 6304
rect 26651 6273 26663 6276
rect 26605 6267 26663 6273
rect 27430 6264 27436 6276
rect 27488 6264 27494 6316
rect 27614 6264 27620 6316
rect 27672 6304 27678 6316
rect 27709 6307 27767 6313
rect 27709 6304 27721 6307
rect 27672 6276 27721 6304
rect 27672 6264 27678 6276
rect 27709 6273 27721 6276
rect 27755 6273 27767 6307
rect 27709 6267 27767 6273
rect 27982 6264 27988 6316
rect 28040 6264 28046 6316
rect 28166 6264 28172 6316
rect 28224 6264 28230 6316
rect 28350 6264 28356 6316
rect 28408 6264 28414 6316
rect 29362 6264 29368 6316
rect 29420 6264 29426 6316
rect 23615 6208 24348 6236
rect 23615 6205 23627 6208
rect 23569 6199 23627 6205
rect 24394 6196 24400 6248
rect 24452 6236 24458 6248
rect 25130 6236 25136 6248
rect 24452 6208 25136 6236
rect 24452 6196 24458 6208
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 26970 6236 26976 6248
rect 26160 6208 26976 6236
rect 20364 6168 20392 6196
rect 19076 6140 20392 6168
rect 20441 6171 20499 6177
rect 18969 6131 19027 6137
rect 20441 6137 20453 6171
rect 20487 6137 20499 6171
rect 22186 6168 22192 6180
rect 20441 6131 20499 6137
rect 21376 6140 22192 6168
rect 17460 6072 18276 6100
rect 17460 6060 17466 6072
rect 18598 6060 18604 6112
rect 18656 6060 18662 6112
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 19521 6103 19579 6109
rect 19521 6100 19533 6103
rect 18748 6072 19533 6100
rect 18748 6060 18754 6072
rect 19521 6069 19533 6072
rect 19567 6069 19579 6103
rect 19521 6063 19579 6069
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 19978 6100 19984 6112
rect 19668 6072 19984 6100
rect 19668 6060 19674 6072
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 20456 6100 20484 6131
rect 20714 6100 20720 6112
rect 20456 6072 20720 6100
rect 20714 6060 20720 6072
rect 20772 6100 20778 6112
rect 21376 6100 21404 6140
rect 22186 6128 22192 6140
rect 22244 6168 22250 6180
rect 23658 6168 23664 6180
rect 22244 6140 23664 6168
rect 22244 6128 22250 6140
rect 23658 6128 23664 6140
rect 23716 6128 23722 6180
rect 26160 6177 26188 6208
rect 26970 6196 26976 6208
rect 27028 6196 27034 6248
rect 29089 6239 29147 6245
rect 29089 6236 29101 6239
rect 28368 6208 29101 6236
rect 28368 6180 28396 6208
rect 29089 6205 29101 6208
rect 29135 6205 29147 6239
rect 29089 6199 29147 6205
rect 29227 6239 29285 6245
rect 29227 6205 29239 6239
rect 29273 6236 29285 6239
rect 30024 6236 30052 6344
rect 30742 6332 30748 6344
rect 30800 6372 30806 6384
rect 31570 6372 31576 6384
rect 30800 6344 31576 6372
rect 30800 6332 30806 6344
rect 31570 6332 31576 6344
rect 31628 6332 31634 6384
rect 32401 6375 32459 6381
rect 31680 6344 32352 6372
rect 31680 6316 31708 6344
rect 30282 6264 30288 6316
rect 30340 6304 30346 6316
rect 30377 6307 30435 6313
rect 30377 6304 30389 6307
rect 30340 6276 30389 6304
rect 30340 6264 30346 6276
rect 30377 6273 30389 6276
rect 30423 6273 30435 6307
rect 30377 6267 30435 6273
rect 30650 6264 30656 6316
rect 30708 6304 30714 6316
rect 31205 6307 31263 6313
rect 31205 6304 31217 6307
rect 30708 6276 31217 6304
rect 30708 6264 30714 6276
rect 31205 6273 31217 6276
rect 31251 6273 31263 6307
rect 31205 6267 31263 6273
rect 31294 6264 31300 6316
rect 31352 6304 31358 6316
rect 31481 6307 31539 6313
rect 31481 6304 31493 6307
rect 31352 6276 31493 6304
rect 31352 6264 31358 6276
rect 31481 6273 31493 6276
rect 31527 6273 31539 6307
rect 31481 6267 31539 6273
rect 31662 6264 31668 6316
rect 31720 6264 31726 6316
rect 31754 6264 31760 6316
rect 31812 6264 31818 6316
rect 31846 6264 31852 6316
rect 31904 6304 31910 6316
rect 32217 6307 32275 6313
rect 32217 6304 32229 6307
rect 31904 6276 32229 6304
rect 31904 6264 31910 6276
rect 32217 6273 32229 6276
rect 32263 6273 32275 6307
rect 32324 6304 32352 6344
rect 32401 6341 32413 6375
rect 32447 6372 32459 6375
rect 32766 6372 32772 6384
rect 32447 6344 32772 6372
rect 32447 6341 32459 6344
rect 32401 6335 32459 6341
rect 32766 6332 32772 6344
rect 32824 6332 32830 6384
rect 34992 6372 35020 6412
rect 36909 6409 36921 6443
rect 36955 6440 36967 6443
rect 37090 6440 37096 6452
rect 36955 6412 37096 6440
rect 36955 6409 36967 6412
rect 36909 6403 36967 6409
rect 37090 6400 37096 6412
rect 37148 6400 37154 6452
rect 37182 6400 37188 6452
rect 37240 6440 37246 6452
rect 39758 6440 39764 6452
rect 37240 6412 39764 6440
rect 37240 6400 37246 6412
rect 39758 6400 39764 6412
rect 39816 6400 39822 6452
rect 40494 6400 40500 6452
rect 40552 6400 40558 6452
rect 42610 6400 42616 6452
rect 42668 6400 42674 6452
rect 43438 6400 43444 6452
rect 43496 6400 43502 6452
rect 34992 6344 36584 6372
rect 32324 6276 32536 6304
rect 32217 6267 32275 6273
rect 29273 6208 30052 6236
rect 30101 6239 30159 6245
rect 29273 6205 29285 6208
rect 29227 6199 29285 6205
rect 30101 6205 30113 6239
rect 30147 6205 30159 6239
rect 31864 6236 31892 6264
rect 30101 6199 30159 6205
rect 30760 6208 31892 6236
rect 26145 6171 26203 6177
rect 26145 6137 26157 6171
rect 26191 6137 26203 6171
rect 26145 6131 26203 6137
rect 26421 6171 26479 6177
rect 26421 6137 26433 6171
rect 26467 6168 26479 6171
rect 26467 6140 27292 6168
rect 26467 6137 26479 6140
rect 26421 6131 26479 6137
rect 20772 6072 21404 6100
rect 20772 6060 20778 6072
rect 21634 6060 21640 6112
rect 21692 6060 21698 6112
rect 21910 6060 21916 6112
rect 21968 6100 21974 6112
rect 22005 6103 22063 6109
rect 22005 6100 22017 6103
rect 21968 6072 22017 6100
rect 21968 6060 21974 6072
rect 22005 6069 22017 6072
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 22281 6103 22339 6109
rect 22281 6069 22293 6103
rect 22327 6100 22339 6103
rect 22922 6100 22928 6112
rect 22327 6072 22928 6100
rect 22327 6069 22339 6072
rect 22281 6063 22339 6069
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 23014 6060 23020 6112
rect 23072 6100 23078 6112
rect 26326 6100 26332 6112
rect 23072 6072 26332 6100
rect 23072 6060 23078 6072
rect 26326 6060 26332 6072
rect 26384 6100 26390 6112
rect 26694 6100 26700 6112
rect 26384 6072 26700 6100
rect 26384 6060 26390 6072
rect 26694 6060 26700 6072
rect 26752 6060 26758 6112
rect 26786 6060 26792 6112
rect 26844 6100 26850 6112
rect 26973 6103 27031 6109
rect 26973 6100 26985 6103
rect 26844 6072 26985 6100
rect 26844 6060 26850 6072
rect 26973 6069 26985 6072
rect 27019 6069 27031 6103
rect 27264 6100 27292 6140
rect 28350 6128 28356 6180
rect 28408 6128 28414 6180
rect 28810 6128 28816 6180
rect 28868 6128 28874 6180
rect 29914 6128 29920 6180
rect 29972 6168 29978 6180
rect 30116 6168 30144 6199
rect 29972 6140 30144 6168
rect 29972 6128 29978 6140
rect 29362 6100 29368 6112
rect 27264 6072 29368 6100
rect 26973 6063 27031 6069
rect 29362 6060 29368 6072
rect 29420 6060 29426 6112
rect 29730 6060 29736 6112
rect 29788 6100 29794 6112
rect 30009 6103 30067 6109
rect 30009 6100 30021 6103
rect 29788 6072 30021 6100
rect 29788 6060 29794 6072
rect 30009 6069 30021 6072
rect 30055 6069 30067 6103
rect 30116 6100 30144 6140
rect 30760 6100 30788 6208
rect 32030 6196 32036 6248
rect 32088 6236 32094 6248
rect 32508 6236 32536 6276
rect 32582 6264 32588 6316
rect 32640 6304 32646 6316
rect 32677 6307 32735 6313
rect 32677 6304 32689 6307
rect 32640 6276 32689 6304
rect 32640 6264 32646 6276
rect 32677 6273 32689 6276
rect 32723 6273 32735 6307
rect 32677 6267 32735 6273
rect 32858 6264 32864 6316
rect 32916 6264 32922 6316
rect 35066 6264 35072 6316
rect 35124 6304 35130 6316
rect 35529 6307 35587 6313
rect 35529 6304 35541 6307
rect 35124 6276 35541 6304
rect 35124 6264 35130 6276
rect 35529 6273 35541 6276
rect 35575 6304 35587 6307
rect 35618 6304 35624 6316
rect 35575 6276 35624 6304
rect 35575 6273 35587 6276
rect 35529 6267 35587 6273
rect 35618 6264 35624 6276
rect 35676 6264 35682 6316
rect 35805 6307 35863 6313
rect 35805 6273 35817 6307
rect 35851 6304 35863 6307
rect 36078 6304 36084 6316
rect 35851 6276 36084 6304
rect 35851 6273 35863 6276
rect 35805 6267 35863 6273
rect 36078 6264 36084 6276
rect 36136 6264 36142 6316
rect 36173 6307 36231 6313
rect 36173 6273 36185 6307
rect 36219 6304 36231 6307
rect 36446 6304 36452 6316
rect 36219 6276 36452 6304
rect 36219 6273 36231 6276
rect 36173 6267 36231 6273
rect 36446 6264 36452 6276
rect 36504 6264 36510 6316
rect 32088 6208 32352 6236
rect 32508 6208 32812 6236
rect 32088 6196 32094 6208
rect 30834 6128 30840 6180
rect 30892 6168 30898 6180
rect 31570 6168 31576 6180
rect 30892 6140 31576 6168
rect 30892 6128 30898 6140
rect 31570 6128 31576 6140
rect 31628 6168 31634 6180
rect 31941 6171 31999 6177
rect 31628 6140 31892 6168
rect 31628 6128 31634 6140
rect 30116 6072 30788 6100
rect 31113 6103 31171 6109
rect 30009 6063 30067 6069
rect 31113 6069 31125 6103
rect 31159 6100 31171 6103
rect 31294 6100 31300 6112
rect 31159 6072 31300 6100
rect 31159 6069 31171 6072
rect 31113 6063 31171 6069
rect 31294 6060 31300 6072
rect 31352 6060 31358 6112
rect 31386 6060 31392 6112
rect 31444 6060 31450 6112
rect 31864 6100 31892 6140
rect 31941 6137 31953 6171
rect 31987 6168 31999 6171
rect 32214 6168 32220 6180
rect 31987 6140 32220 6168
rect 31987 6137 31999 6140
rect 31941 6131 31999 6137
rect 32214 6128 32220 6140
rect 32272 6128 32278 6180
rect 32324 6168 32352 6208
rect 32493 6171 32551 6177
rect 32493 6168 32505 6171
rect 32324 6140 32505 6168
rect 32493 6137 32505 6140
rect 32539 6137 32551 6171
rect 32784 6168 32812 6208
rect 32950 6196 32956 6248
rect 33008 6236 33014 6248
rect 33045 6239 33103 6245
rect 33045 6236 33057 6239
rect 33008 6208 33057 6236
rect 33008 6196 33014 6208
rect 33045 6205 33057 6208
rect 33091 6205 33103 6239
rect 33045 6199 33103 6205
rect 33502 6196 33508 6248
rect 33560 6196 33566 6248
rect 33781 6239 33839 6245
rect 33781 6236 33793 6239
rect 33612 6208 33793 6236
rect 33410 6168 33416 6180
rect 32784 6140 33416 6168
rect 32493 6131 32551 6137
rect 33410 6128 33416 6140
rect 33468 6168 33474 6180
rect 33612 6168 33640 6208
rect 33781 6205 33793 6208
rect 33827 6205 33839 6239
rect 33781 6199 33839 6205
rect 33870 6196 33876 6248
rect 33928 6245 33934 6248
rect 33928 6239 33956 6245
rect 33944 6205 33956 6239
rect 33928 6199 33956 6205
rect 33928 6196 33934 6199
rect 34054 6196 34060 6248
rect 34112 6196 34118 6248
rect 35894 6196 35900 6248
rect 35952 6196 35958 6248
rect 36556 6236 36584 6344
rect 37734 6264 37740 6316
rect 37792 6264 37798 6316
rect 38378 6264 38384 6316
rect 38436 6304 38442 6316
rect 38565 6307 38623 6313
rect 38565 6304 38577 6307
rect 38436 6276 38577 6304
rect 38436 6264 38442 6276
rect 38565 6273 38577 6276
rect 38611 6273 38623 6307
rect 38565 6267 38623 6273
rect 38654 6264 38660 6316
rect 38712 6304 38718 6316
rect 38749 6307 38807 6313
rect 38749 6304 38761 6307
rect 38712 6276 38761 6304
rect 38712 6264 38718 6276
rect 38749 6273 38761 6276
rect 38795 6273 38807 6307
rect 38749 6267 38807 6273
rect 39574 6264 39580 6316
rect 39632 6313 39638 6316
rect 39632 6307 39660 6313
rect 39648 6273 39660 6307
rect 39632 6267 39660 6273
rect 40405 6307 40463 6313
rect 40405 6273 40417 6307
rect 40451 6304 40463 6307
rect 40681 6307 40739 6313
rect 40681 6304 40693 6307
rect 40451 6276 40693 6304
rect 40451 6273 40463 6276
rect 40405 6267 40463 6273
rect 40681 6273 40693 6276
rect 40727 6273 40739 6307
rect 40681 6267 40739 6273
rect 39632 6264 39638 6267
rect 42794 6264 42800 6316
rect 42852 6264 42858 6316
rect 42889 6307 42947 6313
rect 42889 6273 42901 6307
rect 42935 6273 42947 6307
rect 42889 6267 42947 6273
rect 43257 6307 43315 6313
rect 43257 6273 43269 6307
rect 43303 6304 43315 6307
rect 43346 6304 43352 6316
rect 43303 6276 43352 6304
rect 43303 6273 43315 6276
rect 43257 6267 43315 6273
rect 37182 6236 37188 6248
rect 36556 6208 37188 6236
rect 37182 6196 37188 6208
rect 37240 6196 37246 6248
rect 37458 6196 37464 6248
rect 37516 6196 37522 6248
rect 39298 6236 39304 6248
rect 38672 6208 39304 6236
rect 34606 6168 34612 6180
rect 33468 6140 33640 6168
rect 33468 6128 33474 6140
rect 32309 6103 32367 6109
rect 32309 6100 32321 6103
rect 31864 6072 32321 6100
rect 32309 6069 32321 6072
rect 32355 6069 32367 6103
rect 33612 6100 33640 6140
rect 34440 6140 34612 6168
rect 34440 6100 34468 6140
rect 34606 6128 34612 6140
rect 34664 6128 34670 6180
rect 38672 6168 38700 6208
rect 39298 6196 39304 6208
rect 39356 6236 39362 6248
rect 39485 6239 39543 6245
rect 39485 6236 39497 6239
rect 39356 6208 39497 6236
rect 39356 6196 39362 6208
rect 39485 6205 39497 6208
rect 39531 6205 39543 6239
rect 39485 6199 39543 6205
rect 39758 6196 39764 6248
rect 39816 6196 39822 6248
rect 39942 6196 39948 6248
rect 40000 6236 40006 6248
rect 42904 6236 42932 6267
rect 43346 6264 43352 6276
rect 43404 6264 43410 6316
rect 40000 6208 42932 6236
rect 40000 6196 40006 6208
rect 38120 6140 38700 6168
rect 33612 6072 34468 6100
rect 32309 6063 32367 6069
rect 34514 6060 34520 6112
rect 34572 6100 34578 6112
rect 34701 6103 34759 6109
rect 34701 6100 34713 6103
rect 34572 6072 34713 6100
rect 34572 6060 34578 6072
rect 34701 6069 34713 6072
rect 34747 6069 34759 6103
rect 34701 6063 34759 6069
rect 34793 6103 34851 6109
rect 34793 6069 34805 6103
rect 34839 6100 34851 6103
rect 34882 6100 34888 6112
rect 34839 6072 34888 6100
rect 34839 6069 34851 6072
rect 34793 6063 34851 6069
rect 34882 6060 34888 6072
rect 34940 6060 34946 6112
rect 35526 6060 35532 6112
rect 35584 6100 35590 6112
rect 36262 6100 36268 6112
rect 35584 6072 36268 6100
rect 35584 6060 35590 6072
rect 36262 6060 36268 6072
rect 36320 6060 36326 6112
rect 36630 6060 36636 6112
rect 36688 6100 36694 6112
rect 38120 6100 38148 6140
rect 39206 6128 39212 6180
rect 39264 6128 39270 6180
rect 36688 6072 38148 6100
rect 38473 6103 38531 6109
rect 36688 6060 36694 6072
rect 38473 6069 38485 6103
rect 38519 6100 38531 6103
rect 39758 6100 39764 6112
rect 38519 6072 39764 6100
rect 38519 6069 38531 6072
rect 38473 6063 38531 6069
rect 39758 6060 39764 6072
rect 39816 6060 39822 6112
rect 43070 6060 43076 6112
rect 43128 6060 43134 6112
rect 1104 6010 43884 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13918 6010
rect 13970 5958 13982 6010
rect 14034 5958 14046 6010
rect 14098 5958 14110 6010
rect 14162 5958 14174 6010
rect 14226 5958 14238 6010
rect 14290 5958 19918 6010
rect 19970 5958 19982 6010
rect 20034 5958 20046 6010
rect 20098 5958 20110 6010
rect 20162 5958 20174 6010
rect 20226 5958 20238 6010
rect 20290 5958 25918 6010
rect 25970 5958 25982 6010
rect 26034 5958 26046 6010
rect 26098 5958 26110 6010
rect 26162 5958 26174 6010
rect 26226 5958 26238 6010
rect 26290 5958 31918 6010
rect 31970 5958 31982 6010
rect 32034 5958 32046 6010
rect 32098 5958 32110 6010
rect 32162 5958 32174 6010
rect 32226 5958 32238 6010
rect 32290 5958 37918 6010
rect 37970 5958 37982 6010
rect 38034 5958 38046 6010
rect 38098 5958 38110 6010
rect 38162 5958 38174 6010
rect 38226 5958 38238 6010
rect 38290 5958 43884 6010
rect 1104 5936 43884 5958
rect 3050 5856 3056 5908
rect 3108 5856 3114 5908
rect 4430 5856 4436 5908
rect 4488 5856 4494 5908
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 5442 5896 5448 5908
rect 4672 5868 5448 5896
rect 4672 5856 4678 5868
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 6972 5868 7328 5896
rect 6972 5856 6978 5868
rect 3418 5788 3424 5840
rect 3476 5788 3482 5840
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 5408 5800 5948 5828
rect 5408 5788 5414 5800
rect 1762 5720 1768 5772
rect 1820 5760 1826 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1820 5732 2053 5760
rect 1820 5720 1826 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 4522 5760 4528 5772
rect 3292 5732 4528 5760
rect 3292 5720 3298 5732
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4614 5720 4620 5772
rect 4672 5720 4678 5772
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 5810 5760 5816 5772
rect 5767 5732 5816 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 5920 5769 5948 5800
rect 6362 5788 6368 5840
rect 6420 5788 6426 5840
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 5905 5723 5963 5729
rect 5994 5720 6000 5772
rect 6052 5720 6058 5772
rect 6730 5720 6736 5772
rect 6788 5769 6794 5772
rect 6788 5763 6837 5769
rect 6788 5729 6791 5763
rect 6825 5729 6837 5763
rect 7300 5760 7328 5868
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7616 5868 7941 5896
rect 7616 5856 7622 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 11974 5896 11980 5908
rect 8812 5868 11980 5896
rect 8812 5856 8818 5868
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12584 5868 12909 5896
rect 12584 5856 12590 5868
rect 12897 5865 12909 5868
rect 12943 5896 12955 5899
rect 13170 5896 13176 5908
rect 12943 5868 13176 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 13354 5856 13360 5908
rect 13412 5856 13418 5908
rect 13633 5899 13691 5905
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 13722 5896 13728 5908
rect 13679 5868 13728 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 13722 5856 13728 5868
rect 13780 5896 13786 5908
rect 14182 5896 14188 5908
rect 13780 5868 14188 5896
rect 13780 5856 13786 5868
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14366 5856 14372 5908
rect 14424 5896 14430 5908
rect 15105 5899 15163 5905
rect 15105 5896 15117 5899
rect 14424 5868 15117 5896
rect 14424 5856 14430 5868
rect 15105 5865 15117 5868
rect 15151 5865 15163 5899
rect 15105 5859 15163 5865
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15252 5868 16252 5896
rect 15252 5856 15258 5868
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 7432 5800 7696 5828
rect 7432 5788 7438 5800
rect 7668 5760 7696 5800
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 7837 5831 7895 5837
rect 7837 5828 7849 5831
rect 7800 5800 7849 5828
rect 7800 5788 7806 5800
rect 7837 5797 7849 5800
rect 7883 5797 7895 5831
rect 7837 5791 7895 5797
rect 8018 5788 8024 5840
rect 8076 5828 8082 5840
rect 8662 5828 8668 5840
rect 8076 5800 8668 5828
rect 8076 5788 8082 5800
rect 8662 5788 8668 5800
rect 8720 5788 8726 5840
rect 10134 5788 10140 5840
rect 10192 5788 10198 5840
rect 12066 5788 12072 5840
rect 12124 5788 12130 5840
rect 14829 5831 14887 5837
rect 12544 5800 14780 5828
rect 9585 5763 9643 5769
rect 9585 5760 9597 5763
rect 7300 5732 7512 5760
rect 7668 5732 9597 5760
rect 6788 5723 6837 5729
rect 6788 5720 6794 5723
rect 1486 5652 1492 5704
rect 1544 5652 1550 5704
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4304 5664 4353 5692
rect 4304 5652 4310 5664
rect 4341 5661 4353 5664
rect 4387 5692 4399 5695
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4387 5688 4568 5692
rect 4724 5688 4905 5692
rect 4387 5664 4905 5688
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4540 5660 4752 5664
rect 4893 5661 4905 5664
rect 4939 5692 4951 5695
rect 5534 5692 5540 5704
rect 4939 5664 5540 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 6012 5692 6040 5720
rect 5920 5664 6040 5692
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 2556 5596 3249 5624
rect 2556 5584 2562 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3237 5587 3295 5593
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 3881 5627 3939 5633
rect 3881 5624 3893 5627
rect 3476 5596 3893 5624
rect 3476 5584 3482 5596
rect 3881 5593 3893 5596
rect 3927 5593 3939 5627
rect 3881 5587 3939 5593
rect 4065 5627 4123 5633
rect 4065 5593 4077 5627
rect 4111 5624 4123 5627
rect 5920 5624 5948 5664
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 4111 5596 5948 5624
rect 4111 5593 4123 5596
rect 4065 5587 4123 5593
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 3510 5556 3516 5568
rect 1627 5528 3516 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 3602 5516 3608 5568
rect 3660 5556 3666 5568
rect 4706 5556 4712 5568
rect 3660 5528 4712 5556
rect 3660 5516 3666 5528
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5629 5559 5687 5565
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 6822 5556 6828 5568
rect 5675 5528 6828 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7484 5556 7512 5732
rect 9585 5729 9597 5732
rect 9631 5729 9643 5763
rect 9585 5723 9643 5729
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5760 9919 5763
rect 10042 5760 10048 5772
rect 9907 5732 10048 5760
rect 9907 5729 9919 5732
rect 9861 5723 9919 5729
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10778 5720 10784 5772
rect 10836 5720 10842 5772
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 12544 5769 12572 5800
rect 11676 5763 11734 5769
rect 11676 5760 11688 5763
rect 11204 5732 11688 5760
rect 11204 5720 11210 5732
rect 11676 5729 11688 5732
rect 11722 5760 11734 5763
rect 12529 5763 12587 5769
rect 11722 5732 12388 5760
rect 11722 5729 11734 5732
rect 11676 5723 11734 5729
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7607 5664 7665 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 9766 5701 9772 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7984 5664 8125 5692
rect 7984 5652 7990 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8435 5664 8953 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9744 5695 9772 5701
rect 9744 5661 9756 5695
rect 9744 5655 9772 5661
rect 9766 5652 9772 5655
rect 9824 5652 9830 5704
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 10612 5624 10640 5655
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 12360 5692 12388 5732
rect 12529 5729 12541 5763
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 12710 5720 12716 5772
rect 12768 5720 12774 5772
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13096 5732 13553 5760
rect 13096 5704 13124 5732
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 14277 5763 14335 5769
rect 14277 5729 14289 5763
rect 14323 5760 14335 5763
rect 14366 5760 14372 5772
rect 14323 5732 14372 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 14752 5760 14780 5800
rect 14829 5797 14841 5831
rect 14875 5828 14887 5831
rect 15286 5828 15292 5840
rect 14875 5800 15292 5828
rect 14875 5797 14887 5800
rect 14829 5791 14887 5797
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 15378 5760 15384 5772
rect 14752 5732 15384 5760
rect 15378 5720 15384 5732
rect 15436 5760 15442 5772
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 15436 5732 16037 5760
rect 15436 5720 15442 5732
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16224 5760 16252 5868
rect 16316 5868 18368 5896
rect 16316 5837 16344 5868
rect 16301 5831 16359 5837
rect 16301 5797 16313 5831
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 17402 5828 17408 5840
rect 16448 5800 17408 5828
rect 16448 5788 16454 5800
rect 16960 5769 16988 5800
rect 17402 5788 17408 5800
rect 17460 5788 17466 5840
rect 16945 5763 17003 5769
rect 16224 5732 16804 5760
rect 16025 5723 16083 5729
rect 12360 5664 12572 5692
rect 12544 5624 12572 5664
rect 13078 5652 13084 5704
rect 13136 5652 13142 5704
rect 13170 5652 13176 5704
rect 13228 5652 13234 5704
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 14461 5695 14519 5701
rect 13504 5664 14412 5692
rect 13504 5652 13510 5664
rect 13354 5624 13360 5636
rect 8628 5596 8892 5624
rect 10612 5596 11008 5624
rect 12544 5596 13360 5624
rect 8628 5584 8634 5596
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7484 5528 8217 5556
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 8386 5516 8392 5568
rect 8444 5556 8450 5568
rect 8665 5559 8723 5565
rect 8665 5556 8677 5559
rect 8444 5528 8677 5556
rect 8444 5516 8450 5528
rect 8665 5525 8677 5528
rect 8711 5525 8723 5559
rect 8864 5556 8892 5596
rect 9490 5556 9496 5568
rect 8864 5528 9496 5556
rect 8665 5519 8723 5525
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 10870 5516 10876 5568
rect 10928 5516 10934 5568
rect 10980 5556 11008 5596
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 13722 5584 13728 5636
rect 13780 5584 13786 5636
rect 14384 5633 14412 5664
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 14918 5692 14924 5704
rect 14507 5664 14924 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 15746 5652 15752 5704
rect 15804 5652 15810 5704
rect 15930 5701 15936 5704
rect 15908 5695 15936 5701
rect 15908 5661 15920 5695
rect 15908 5655 15936 5661
rect 15930 5652 15936 5655
rect 15988 5652 15994 5704
rect 16776 5701 16804 5732
rect 16945 5729 16957 5763
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17586 5692 17592 5704
rect 17451 5664 17592 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 14369 5627 14427 5633
rect 14369 5593 14381 5627
rect 14415 5593 14427 5627
rect 16776 5624 16804 5655
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 17770 5692 17776 5704
rect 17727 5664 17776 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18340 5692 18368 5868
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 18877 5899 18935 5905
rect 18877 5896 18889 5899
rect 18656 5868 18889 5896
rect 18656 5856 18662 5868
rect 18877 5865 18889 5868
rect 18923 5896 18935 5899
rect 19058 5896 19064 5908
rect 18923 5868 19064 5896
rect 18923 5865 18935 5868
rect 18877 5859 18935 5865
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 19242 5856 19248 5908
rect 19300 5856 19306 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 19978 5896 19984 5908
rect 19668 5868 19984 5896
rect 19668 5856 19674 5868
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20714 5896 20720 5908
rect 20312 5868 20720 5896
rect 20312 5856 20318 5868
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 21542 5896 21548 5908
rect 20956 5868 21548 5896
rect 20956 5856 20962 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 23569 5899 23627 5905
rect 23569 5896 23581 5899
rect 21692 5868 23581 5896
rect 21692 5856 21698 5868
rect 23569 5865 23581 5868
rect 23615 5865 23627 5899
rect 23569 5859 23627 5865
rect 23934 5856 23940 5908
rect 23992 5856 23998 5908
rect 24118 5856 24124 5908
rect 24176 5896 24182 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 24176 5868 24409 5896
rect 24176 5856 24182 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 29178 5896 29184 5908
rect 24397 5859 24455 5865
rect 26068 5868 29184 5896
rect 18417 5831 18475 5837
rect 18417 5797 18429 5831
rect 18463 5828 18475 5831
rect 20346 5828 20352 5840
rect 18463 5800 18552 5828
rect 18463 5797 18475 5800
rect 18417 5791 18475 5797
rect 18524 5769 18552 5800
rect 18892 5800 20352 5828
rect 18509 5763 18567 5769
rect 18509 5729 18521 5763
rect 18555 5729 18567 5763
rect 18892 5760 18920 5800
rect 20346 5788 20352 5800
rect 20404 5788 20410 5840
rect 20438 5788 20444 5840
rect 20496 5788 20502 5840
rect 24578 5828 24584 5840
rect 21560 5800 24584 5828
rect 18509 5723 18567 5729
rect 18616 5732 18920 5760
rect 18984 5732 19932 5760
rect 18616 5692 18644 5732
rect 18984 5692 19012 5732
rect 18340 5664 18644 5692
rect 18800 5664 19012 5692
rect 18800 5624 18828 5664
rect 19334 5652 19340 5704
rect 19392 5688 19398 5704
rect 19429 5695 19487 5701
rect 19429 5688 19441 5695
rect 19392 5661 19441 5688
rect 19475 5661 19487 5695
rect 19392 5660 19487 5661
rect 19392 5652 19398 5660
rect 19429 5655 19487 5660
rect 19610 5652 19616 5704
rect 19668 5692 19674 5704
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19668 5664 19717 5692
rect 19668 5652 19674 5664
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19794 5652 19800 5704
rect 19852 5652 19858 5704
rect 19904 5692 19932 5732
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 21560 5760 21588 5800
rect 24578 5788 24584 5800
rect 24636 5788 24642 5840
rect 20036 5732 21588 5760
rect 21637 5763 21695 5769
rect 20036 5720 20042 5732
rect 21637 5729 21649 5763
rect 21683 5760 21695 5763
rect 22097 5763 22155 5769
rect 22097 5760 22109 5763
rect 21683 5732 22109 5760
rect 21683 5729 21695 5732
rect 21637 5723 21695 5729
rect 22097 5729 22109 5732
rect 22143 5729 22155 5763
rect 22097 5723 22155 5729
rect 23477 5763 23535 5769
rect 23477 5729 23489 5763
rect 23523 5760 23535 5763
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 23523 5732 24961 5760
rect 23523 5729 23535 5732
rect 23477 5723 23535 5729
rect 24949 5729 24961 5732
rect 24995 5760 25007 5763
rect 25317 5763 25375 5769
rect 25317 5760 25329 5763
rect 24995 5732 25329 5760
rect 24995 5729 25007 5732
rect 24949 5723 25007 5729
rect 25317 5729 25329 5732
rect 25363 5729 25375 5763
rect 25317 5723 25375 5729
rect 25682 5720 25688 5772
rect 25740 5760 25746 5772
rect 26068 5769 26096 5868
rect 29178 5856 29184 5868
rect 29236 5896 29242 5908
rect 30190 5896 30196 5908
rect 29236 5868 30196 5896
rect 29236 5856 29242 5868
rect 30190 5856 30196 5868
rect 30248 5856 30254 5908
rect 30282 5856 30288 5908
rect 30340 5896 30346 5908
rect 31018 5896 31024 5908
rect 30340 5868 31024 5896
rect 30340 5856 30346 5868
rect 31018 5856 31024 5868
rect 31076 5896 31082 5908
rect 32950 5896 32956 5908
rect 31076 5868 32956 5896
rect 31076 5856 31082 5868
rect 32950 5856 32956 5868
rect 33008 5856 33014 5908
rect 33689 5899 33747 5905
rect 33689 5865 33701 5899
rect 33735 5896 33747 5899
rect 34054 5896 34060 5908
rect 33735 5868 34060 5896
rect 33735 5865 33747 5868
rect 33689 5859 33747 5865
rect 34054 5856 34060 5868
rect 34112 5856 34118 5908
rect 34330 5856 34336 5908
rect 34388 5856 34394 5908
rect 34698 5856 34704 5908
rect 34756 5856 34762 5908
rect 35084 5868 36492 5896
rect 26602 5828 26608 5840
rect 26252 5800 26608 5828
rect 26252 5772 26280 5800
rect 26602 5788 26608 5800
rect 26660 5788 26666 5840
rect 27798 5788 27804 5840
rect 27856 5828 27862 5840
rect 29914 5828 29920 5840
rect 27856 5800 29920 5828
rect 27856 5788 27862 5800
rect 29914 5788 29920 5800
rect 29972 5788 29978 5840
rect 31294 5788 31300 5840
rect 31352 5828 31358 5840
rect 31389 5831 31447 5837
rect 31389 5828 31401 5831
rect 31352 5800 31401 5828
rect 31352 5788 31358 5800
rect 31389 5797 31401 5800
rect 31435 5797 31447 5831
rect 31389 5791 31447 5797
rect 33965 5831 34023 5837
rect 33965 5797 33977 5831
rect 34011 5828 34023 5831
rect 35084 5828 35112 5868
rect 34011 5800 35112 5828
rect 36464 5828 36492 5868
rect 36538 5856 36544 5908
rect 36596 5896 36602 5908
rect 36817 5899 36875 5905
rect 36817 5896 36829 5899
rect 36596 5868 36829 5896
rect 36596 5856 36602 5868
rect 36817 5865 36829 5868
rect 36863 5865 36875 5899
rect 36817 5859 36875 5865
rect 37366 5856 37372 5908
rect 37424 5856 37430 5908
rect 37458 5856 37464 5908
rect 37516 5896 37522 5908
rect 38105 5899 38163 5905
rect 37516 5868 38056 5896
rect 37516 5856 37522 5868
rect 37642 5828 37648 5840
rect 36464 5800 37648 5828
rect 34011 5797 34023 5800
rect 33965 5791 34023 5797
rect 37642 5788 37648 5800
rect 37700 5788 37706 5840
rect 38028 5828 38056 5868
rect 38105 5865 38117 5899
rect 38151 5896 38163 5899
rect 38151 5868 39160 5896
rect 38151 5865 38163 5868
rect 38105 5859 38163 5865
rect 39132 5828 39160 5868
rect 39206 5856 39212 5908
rect 39264 5856 39270 5908
rect 42886 5828 42892 5840
rect 38028 5800 38240 5828
rect 39132 5800 42892 5828
rect 38212 5772 38240 5800
rect 42886 5788 42892 5800
rect 42944 5788 42950 5840
rect 43438 5788 43444 5840
rect 43496 5788 43502 5840
rect 26053 5763 26111 5769
rect 26053 5760 26065 5763
rect 25740 5732 26065 5760
rect 25740 5720 25746 5732
rect 26053 5729 26065 5732
rect 26099 5729 26111 5763
rect 26053 5723 26111 5729
rect 26234 5720 26240 5772
rect 26292 5720 26298 5772
rect 26326 5720 26332 5772
rect 26384 5760 26390 5772
rect 26697 5763 26755 5769
rect 26697 5760 26709 5763
rect 26384 5732 26709 5760
rect 26384 5720 26390 5732
rect 26697 5729 26709 5732
rect 26743 5729 26755 5763
rect 26697 5723 26755 5729
rect 27111 5763 27169 5769
rect 27111 5729 27123 5763
rect 27157 5760 27169 5763
rect 27157 5732 27844 5760
rect 27157 5729 27169 5732
rect 27111 5723 27169 5729
rect 19904 5664 20024 5692
rect 16776 5596 18828 5624
rect 14369 5587 14427 5593
rect 18874 5584 18880 5636
rect 18932 5584 18938 5636
rect 18966 5584 18972 5636
rect 19024 5624 19030 5636
rect 19024 5596 19104 5624
rect 19024 5584 19030 5596
rect 15470 5556 15476 5568
rect 10980 5528 15476 5556
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 16482 5556 16488 5568
rect 15712 5528 16488 5556
rect 15712 5516 15718 5528
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 18417 5559 18475 5565
rect 18417 5525 18429 5559
rect 18463 5556 18475 5559
rect 18782 5556 18788 5568
rect 18463 5528 18788 5556
rect 18463 5525 18475 5528
rect 18417 5519 18475 5525
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 19076 5565 19104 5596
rect 19150 5584 19156 5636
rect 19208 5624 19214 5636
rect 19208 5596 19748 5624
rect 19208 5584 19214 5596
rect 19720 5568 19748 5596
rect 19061 5559 19119 5565
rect 19061 5525 19073 5559
rect 19107 5525 19119 5559
rect 19061 5519 19119 5525
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19521 5559 19579 5565
rect 19521 5556 19533 5559
rect 19392 5528 19533 5556
rect 19392 5516 19398 5528
rect 19521 5525 19533 5528
rect 19567 5525 19579 5559
rect 19521 5519 19579 5525
rect 19702 5516 19708 5568
rect 19760 5516 19766 5568
rect 19996 5556 20024 5664
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 20898 5701 20904 5704
rect 20855 5695 20904 5701
rect 20855 5661 20867 5695
rect 20901 5661 20904 5695
rect 20855 5655 20904 5661
rect 20898 5652 20904 5655
rect 20956 5652 20962 5704
rect 20990 5652 20996 5704
rect 21048 5652 21054 5704
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 21542 5584 21548 5636
rect 21600 5624 21606 5636
rect 21928 5624 21956 5655
rect 22186 5652 22192 5704
rect 22244 5652 22250 5704
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 24820 5664 24869 5692
rect 24820 5652 24826 5664
rect 24857 5661 24869 5664
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 25225 5695 25283 5701
rect 25225 5661 25237 5695
rect 25271 5661 25283 5695
rect 25225 5655 25283 5661
rect 21600 5596 21956 5624
rect 21600 5584 21606 5596
rect 23842 5584 23848 5636
rect 23900 5624 23906 5636
rect 25240 5624 25268 5655
rect 25590 5652 25596 5704
rect 25648 5692 25654 5704
rect 25958 5692 25964 5704
rect 25648 5664 25964 5692
rect 25648 5652 25654 5664
rect 25958 5652 25964 5664
rect 26016 5652 26022 5704
rect 26988 5652 26994 5704
rect 27046 5652 27052 5704
rect 27246 5652 27252 5704
rect 27304 5652 27310 5704
rect 27816 5692 27844 5732
rect 27890 5720 27896 5772
rect 27948 5760 27954 5772
rect 27985 5763 28043 5769
rect 27985 5760 27997 5763
rect 27948 5732 27997 5760
rect 27948 5720 27954 5732
rect 27985 5729 27997 5732
rect 28031 5729 28043 5763
rect 27985 5723 28043 5729
rect 28166 5720 28172 5772
rect 28224 5760 28230 5772
rect 28224 5732 30696 5760
rect 28224 5720 28230 5732
rect 28261 5695 28319 5701
rect 27816 5664 28028 5692
rect 28000 5636 28028 5664
rect 28261 5661 28273 5695
rect 28307 5692 28319 5695
rect 28350 5692 28356 5704
rect 28307 5664 28356 5692
rect 28307 5661 28319 5664
rect 28261 5655 28319 5661
rect 28350 5652 28356 5664
rect 28408 5652 28414 5704
rect 29730 5652 29736 5704
rect 29788 5652 29794 5704
rect 30668 5692 30696 5732
rect 30742 5720 30748 5772
rect 30800 5720 30806 5772
rect 31478 5720 31484 5772
rect 31536 5760 31542 5772
rect 31941 5763 31999 5769
rect 31941 5760 31953 5763
rect 31536 5732 31953 5760
rect 31536 5720 31542 5732
rect 31941 5729 31953 5732
rect 31987 5729 31999 5763
rect 31941 5723 31999 5729
rect 32674 5720 32680 5772
rect 32732 5720 32738 5772
rect 36446 5720 36452 5772
rect 36504 5760 36510 5772
rect 36504 5732 38056 5760
rect 36504 5720 36510 5732
rect 30926 5692 30932 5704
rect 30668 5664 30932 5692
rect 30926 5652 30932 5664
rect 30984 5652 30990 5704
rect 31662 5652 31668 5704
rect 31720 5652 31726 5704
rect 31754 5652 31760 5704
rect 31812 5701 31818 5704
rect 31812 5695 31840 5701
rect 31828 5661 31840 5695
rect 31812 5655 31840 5661
rect 32953 5695 33011 5701
rect 32953 5661 32965 5695
rect 32999 5692 33011 5695
rect 33042 5692 33048 5704
rect 32999 5664 33048 5692
rect 32999 5661 33011 5664
rect 32953 5655 33011 5661
rect 31812 5652 31818 5655
rect 33042 5652 33048 5664
rect 33100 5692 33106 5704
rect 33781 5695 33839 5701
rect 33781 5692 33793 5695
rect 33100 5664 33793 5692
rect 33100 5652 33106 5664
rect 33781 5661 33793 5664
rect 33827 5661 33839 5695
rect 33781 5655 33839 5661
rect 34514 5652 34520 5704
rect 34572 5652 34578 5704
rect 35434 5652 35440 5704
rect 35492 5652 35498 5704
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5661 35771 5695
rect 35713 5655 35771 5661
rect 35805 5695 35863 5701
rect 35805 5661 35817 5695
rect 35851 5692 35863 5695
rect 35986 5692 35992 5704
rect 35851 5664 35992 5692
rect 35851 5661 35863 5664
rect 35805 5655 35863 5661
rect 26234 5624 26240 5636
rect 23900 5596 24808 5624
rect 23900 5584 23906 5596
rect 21634 5556 21640 5568
rect 19996 5528 21640 5556
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 21729 5559 21787 5565
rect 21729 5525 21741 5559
rect 21775 5556 21787 5559
rect 22002 5556 22008 5568
rect 21775 5528 22008 5556
rect 21775 5525 21787 5528
rect 21729 5519 21787 5525
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 24780 5565 24808 5596
rect 24872 5596 25268 5624
rect 25516 5596 26240 5624
rect 24872 5568 24900 5596
rect 24765 5559 24823 5565
rect 24765 5525 24777 5559
rect 24811 5525 24823 5559
rect 24765 5519 24823 5525
rect 24854 5516 24860 5568
rect 24912 5516 24918 5568
rect 25038 5516 25044 5568
rect 25096 5556 25102 5568
rect 25516 5556 25544 5596
rect 26234 5584 26240 5596
rect 26292 5584 26298 5636
rect 27982 5584 27988 5636
rect 28040 5624 28046 5636
rect 29362 5624 29368 5636
rect 28040 5596 29368 5624
rect 28040 5584 28046 5596
rect 29362 5584 29368 5596
rect 29420 5584 29426 5636
rect 33152 5596 35388 5624
rect 25096 5528 25544 5556
rect 25096 5516 25102 5528
rect 25590 5516 25596 5568
rect 25648 5556 25654 5568
rect 27798 5556 27804 5568
rect 25648 5528 27804 5556
rect 25648 5516 25654 5528
rect 27798 5516 27804 5528
rect 27856 5516 27862 5568
rect 27893 5559 27951 5565
rect 27893 5525 27905 5559
rect 27939 5556 27951 5559
rect 28258 5556 28264 5568
rect 27939 5528 28264 5556
rect 27939 5525 27951 5528
rect 27893 5519 27951 5525
rect 28258 5516 28264 5528
rect 28316 5516 28322 5568
rect 29178 5516 29184 5568
rect 29236 5556 29242 5568
rect 29549 5559 29607 5565
rect 29549 5556 29561 5559
rect 29236 5528 29561 5556
rect 29236 5516 29242 5528
rect 29549 5525 29561 5528
rect 29595 5525 29607 5559
rect 29549 5519 29607 5525
rect 30742 5516 30748 5568
rect 30800 5556 30806 5568
rect 31386 5556 31392 5568
rect 30800 5528 31392 5556
rect 30800 5516 30806 5528
rect 31386 5516 31392 5528
rect 31444 5516 31450 5568
rect 31938 5516 31944 5568
rect 31996 5556 32002 5568
rect 32585 5559 32643 5565
rect 32585 5556 32597 5559
rect 31996 5528 32597 5556
rect 31996 5516 32002 5528
rect 32585 5525 32597 5528
rect 32631 5525 32643 5559
rect 32585 5519 32643 5525
rect 32766 5516 32772 5568
rect 32824 5556 32830 5568
rect 33152 5556 33180 5596
rect 32824 5528 33180 5556
rect 35360 5556 35388 5596
rect 35728 5556 35756 5655
rect 35986 5652 35992 5664
rect 36044 5652 36050 5704
rect 36081 5695 36139 5701
rect 36081 5661 36093 5695
rect 36127 5692 36139 5695
rect 36127 5664 37504 5692
rect 36127 5661 36139 5664
rect 36081 5655 36139 5661
rect 37476 5636 37504 5664
rect 37550 5652 37556 5704
rect 37608 5652 37614 5704
rect 37921 5695 37979 5701
rect 37921 5661 37933 5695
rect 37967 5661 37979 5695
rect 38028 5692 38056 5732
rect 38194 5720 38200 5772
rect 38252 5720 38258 5772
rect 43530 5760 43536 5772
rect 43180 5732 43536 5760
rect 38473 5695 38531 5701
rect 38473 5692 38485 5695
rect 38028 5664 38485 5692
rect 37921 5655 37979 5661
rect 38473 5661 38485 5664
rect 38519 5692 38531 5695
rect 39206 5692 39212 5704
rect 38519 5664 39212 5692
rect 38519 5661 38531 5664
rect 38473 5655 38531 5661
rect 37458 5584 37464 5636
rect 37516 5624 37522 5636
rect 37734 5624 37740 5636
rect 37516 5596 37740 5624
rect 37516 5584 37522 5596
rect 37734 5584 37740 5596
rect 37792 5624 37798 5636
rect 37936 5624 37964 5655
rect 39206 5652 39212 5664
rect 39264 5692 39270 5704
rect 39301 5695 39359 5701
rect 39301 5692 39313 5695
rect 39264 5664 39313 5692
rect 39264 5652 39270 5664
rect 39301 5661 39313 5664
rect 39347 5661 39359 5695
rect 39301 5655 39359 5661
rect 40218 5652 40224 5704
rect 40276 5692 40282 5704
rect 41874 5692 41880 5704
rect 40276 5664 41880 5692
rect 40276 5652 40282 5664
rect 41874 5652 41880 5664
rect 41932 5652 41938 5704
rect 42889 5695 42947 5701
rect 42889 5661 42901 5695
rect 42935 5692 42947 5695
rect 43180 5692 43208 5732
rect 43530 5720 43536 5732
rect 43588 5720 43594 5772
rect 42935 5664 43208 5692
rect 43257 5695 43315 5701
rect 42935 5661 42947 5664
rect 42889 5655 42947 5661
rect 43257 5661 43269 5695
rect 43303 5661 43315 5695
rect 43257 5655 43315 5661
rect 37792 5596 37964 5624
rect 37792 5584 37798 5596
rect 38194 5584 38200 5636
rect 38252 5624 38258 5636
rect 38252 5596 39344 5624
rect 38252 5584 38258 5596
rect 39316 5568 39344 5596
rect 39666 5584 39672 5636
rect 39724 5624 39730 5636
rect 43272 5624 43300 5655
rect 39724 5596 43300 5624
rect 39724 5584 39730 5596
rect 36078 5556 36084 5568
rect 35360 5528 36084 5556
rect 32824 5516 32830 5528
rect 36078 5516 36084 5528
rect 36136 5516 36142 5568
rect 39298 5516 39304 5568
rect 39356 5516 39362 5568
rect 39485 5559 39543 5565
rect 39485 5525 39497 5559
rect 39531 5556 39543 5559
rect 42978 5556 42984 5568
rect 39531 5528 42984 5556
rect 39531 5525 39543 5528
rect 39485 5519 39543 5525
rect 42978 5516 42984 5528
rect 43036 5516 43042 5568
rect 43070 5516 43076 5568
rect 43128 5516 43134 5568
rect 1104 5466 43884 5488
rect 1104 5414 2658 5466
rect 2710 5414 2722 5466
rect 2774 5414 2786 5466
rect 2838 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 8658 5466
rect 8710 5414 8722 5466
rect 8774 5414 8786 5466
rect 8838 5414 8850 5466
rect 8902 5414 8914 5466
rect 8966 5414 8978 5466
rect 9030 5414 14658 5466
rect 14710 5414 14722 5466
rect 14774 5414 14786 5466
rect 14838 5414 14850 5466
rect 14902 5414 14914 5466
rect 14966 5414 14978 5466
rect 15030 5414 20658 5466
rect 20710 5414 20722 5466
rect 20774 5414 20786 5466
rect 20838 5414 20850 5466
rect 20902 5414 20914 5466
rect 20966 5414 20978 5466
rect 21030 5414 26658 5466
rect 26710 5414 26722 5466
rect 26774 5414 26786 5466
rect 26838 5414 26850 5466
rect 26902 5414 26914 5466
rect 26966 5414 26978 5466
rect 27030 5414 32658 5466
rect 32710 5414 32722 5466
rect 32774 5414 32786 5466
rect 32838 5414 32850 5466
rect 32902 5414 32914 5466
rect 32966 5414 32978 5466
rect 33030 5414 38658 5466
rect 38710 5414 38722 5466
rect 38774 5414 38786 5466
rect 38838 5414 38850 5466
rect 38902 5414 38914 5466
rect 38966 5414 38978 5466
rect 39030 5414 43884 5466
rect 1104 5392 43884 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 2774 5352 2780 5364
rect 1627 5324 2780 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 4798 5352 4804 5364
rect 2976 5324 4804 5352
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1578 5216 1584 5228
rect 1443 5188 1584 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2498 5176 2504 5228
rect 2556 5216 2562 5228
rect 2777 5219 2835 5225
rect 2777 5216 2789 5219
rect 2556 5188 2789 5216
rect 2556 5176 2562 5188
rect 2777 5185 2789 5188
rect 2823 5216 2835 5219
rect 2976 5216 3004 5324
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5460 5324 6684 5352
rect 4522 5244 4528 5296
rect 4580 5284 4586 5296
rect 5460 5284 5488 5324
rect 6454 5284 6460 5296
rect 4580 5256 5488 5284
rect 6380 5256 6460 5284
rect 4580 5244 4586 5256
rect 2823 5188 3004 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 3878 5225 3884 5228
rect 3835 5219 3884 5225
rect 3835 5185 3847 5219
rect 3881 5185 3884 5219
rect 3835 5179 3884 5185
rect 3878 5176 3884 5179
rect 3936 5176 3942 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 4982 5216 4988 5228
rect 4847 5188 4988 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5166 5216 5172 5228
rect 5123 5188 5172 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 6380 5225 6408 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6656 5225 6684 5324
rect 7098 5312 7104 5364
rect 7156 5312 7162 5364
rect 7377 5355 7435 5361
rect 7377 5321 7389 5355
rect 7423 5352 7435 5355
rect 7650 5352 7656 5364
rect 7423 5324 7656 5352
rect 7423 5321 7435 5324
rect 7377 5315 7435 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8662 5352 8668 5364
rect 8128 5324 8668 5352
rect 7116 5284 7144 5312
rect 7116 5256 7604 5284
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 6687 5188 7052 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 2961 5151 3019 5157
rect 2740 5120 2912 5148
rect 2740 5108 2746 5120
rect 2884 5080 2912 5120
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3050 5148 3056 5160
rect 3007 5120 3056 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4019 5120 4384 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 3142 5080 3148 5092
rect 2884 5052 3148 5080
rect 3142 5040 3148 5052
rect 3200 5040 3206 5092
rect 3418 5040 3424 5092
rect 3476 5040 3482 5092
rect 1673 5015 1731 5021
rect 1673 4981 1685 5015
rect 1719 5012 1731 5015
rect 4356 5012 4384 5120
rect 1719 4984 4384 5012
rect 1719 4981 1731 4984
rect 1673 4975 1731 4981
rect 4614 4972 4620 5024
rect 4672 4972 4678 5024
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 6454 5012 6460 5024
rect 5859 4984 6460 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 7024 5012 7052 5188
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7156 5188 7481 5216
rect 7156 5176 7162 5188
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7576 5080 7604 5256
rect 8128 5225 8156 5324
rect 8662 5312 8668 5324
rect 8720 5352 8726 5364
rect 8720 5324 9628 5352
rect 8720 5312 8726 5324
rect 9600 5284 9628 5324
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 10008 5324 10057 5352
rect 10008 5312 10014 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 11333 5355 11391 5361
rect 10376 5324 10916 5352
rect 10376 5312 10382 5324
rect 10778 5284 10784 5296
rect 9600 5256 10784 5284
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 10888 5284 10916 5324
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11514 5352 11520 5364
rect 11379 5324 11520 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 12710 5352 12716 5364
rect 11716 5324 12716 5352
rect 11606 5284 11612 5296
rect 10888 5256 11612 5284
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 9122 5176 9128 5228
rect 9180 5176 9186 5228
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 11054 5216 11060 5228
rect 10643 5188 11060 5216
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 11716 5216 11744 5324
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13044 5324 13829 5352
rect 13044 5312 13050 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 17218 5352 17224 5364
rect 13817 5315 13875 5321
rect 14108 5324 17224 5352
rect 11563 5188 11744 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 12710 5176 12716 5228
rect 12768 5176 12774 5228
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 13906 5216 13912 5228
rect 13688 5188 13912 5216
rect 13688 5176 13694 5188
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14108 5216 14136 5324
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 18233 5355 18291 5361
rect 17644 5324 18184 5352
rect 17644 5312 17650 5324
rect 14182 5244 14188 5296
rect 14240 5244 14246 5296
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16540 5256 18092 5284
rect 16540 5244 16546 5256
rect 14047 5188 14136 5216
rect 14369 5219 14427 5225
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 15010 5216 15016 5228
rect 14415 5188 15016 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15838 5176 15844 5228
rect 15896 5176 15902 5228
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16850 5216 16856 5228
rect 16715 5188 16856 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 18064 5225 18092 5256
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5185 18107 5219
rect 18156 5216 18184 5324
rect 18233 5321 18245 5355
rect 18279 5352 18291 5355
rect 19242 5352 19248 5364
rect 18279 5324 19248 5352
rect 18279 5321 18291 5324
rect 18233 5315 18291 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 21637 5355 21695 5361
rect 19659 5324 21496 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 18325 5287 18383 5293
rect 18325 5253 18337 5287
rect 18371 5284 18383 5287
rect 19061 5287 19119 5293
rect 19061 5284 19073 5287
rect 18371 5256 19073 5284
rect 18371 5253 18383 5256
rect 18325 5247 18383 5253
rect 19061 5253 19073 5256
rect 19107 5253 19119 5287
rect 19426 5284 19432 5296
rect 19061 5247 19119 5253
rect 19352 5256 19432 5284
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18156 5188 18429 5216
rect 18049 5179 18107 5185
rect 18417 5185 18429 5188
rect 18463 5185 18475 5219
rect 18417 5179 18475 5185
rect 7926 5108 7932 5160
rect 7984 5108 7990 5160
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8352 5120 8861 5148
rect 8352 5108 8358 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 8987 5151 9045 5157
rect 8987 5117 8999 5151
rect 9033 5148 9045 5151
rect 9306 5148 9312 5160
rect 9033 5120 9312 5148
rect 9033 5117 9045 5120
rect 8987 5111 9045 5117
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 11701 5151 11759 5157
rect 11701 5117 11713 5151
rect 11747 5117 11759 5151
rect 11701 5111 11759 5117
rect 7653 5083 7711 5089
rect 7653 5080 7665 5083
rect 7576 5052 7665 5080
rect 7653 5049 7665 5052
rect 7699 5049 7711 5083
rect 7653 5043 7711 5049
rect 8570 5040 8576 5092
rect 8628 5040 8634 5092
rect 10318 5080 10324 5092
rect 9508 5052 10324 5080
rect 9508 5012 9536 5052
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 7024 4984 9536 5012
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 10778 5012 10784 5024
rect 9815 4984 10784 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11716 5012 11744 5111
rect 11790 5108 11796 5160
rect 11848 5148 11854 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 11848 5120 12449 5148
rect 11848 5108 11854 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12575 5151 12633 5157
rect 12575 5117 12587 5151
rect 12621 5148 12633 5151
rect 13354 5148 13360 5160
rect 12621 5120 13360 5148
rect 12621 5117 12633 5120
rect 12575 5111 12633 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 14458 5148 14464 5160
rect 13556 5120 14464 5148
rect 11882 5040 11888 5092
rect 11940 5080 11946 5092
rect 12161 5083 12219 5089
rect 12161 5080 12173 5083
rect 11940 5052 12173 5080
rect 11940 5040 11946 5052
rect 12161 5049 12173 5052
rect 12207 5049 12219 5083
rect 13556 5080 13584 5120
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 14642 5108 14648 5160
rect 14700 5108 14706 5160
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 15194 5148 15200 5160
rect 14875 5120 15200 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15436 5120 15577 5148
rect 15436 5108 15442 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 15654 5108 15660 5160
rect 15712 5157 15718 5160
rect 15712 5151 15761 5157
rect 15712 5117 15715 5151
rect 15749 5148 15761 5151
rect 16022 5148 16028 5160
rect 15749 5120 16028 5148
rect 15749 5117 15761 5120
rect 15712 5111 15761 5117
rect 15712 5108 15718 5111
rect 16022 5108 16028 5120
rect 16080 5108 16086 5160
rect 17957 5151 18015 5157
rect 17957 5117 17969 5151
rect 18003 5117 18015 5151
rect 18064 5148 18092 5179
rect 18506 5176 18512 5228
rect 18564 5176 18570 5228
rect 18598 5176 18604 5228
rect 18656 5176 18662 5228
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 18966 5216 18972 5228
rect 18831 5188 18972 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19352 5225 19380 5256
rect 19426 5244 19432 5256
rect 19484 5284 19490 5296
rect 19794 5284 19800 5296
rect 19484 5256 19800 5284
rect 19484 5244 19490 5256
rect 19794 5244 19800 5256
rect 19852 5244 19858 5296
rect 19978 5244 19984 5296
rect 20036 5244 20042 5296
rect 21468 5284 21496 5324
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 22094 5352 22100 5364
rect 21683 5324 22100 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 22094 5312 22100 5324
rect 22152 5312 22158 5364
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22511 5355 22569 5361
rect 22511 5352 22523 5355
rect 22244 5324 22523 5352
rect 22244 5312 22250 5324
rect 22511 5321 22523 5324
rect 22557 5321 22569 5355
rect 22511 5315 22569 5321
rect 23290 5312 23296 5364
rect 23348 5352 23354 5364
rect 23934 5352 23940 5364
rect 23348 5324 23940 5352
rect 23348 5312 23354 5324
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 24762 5312 24768 5364
rect 24820 5312 24826 5364
rect 25498 5312 25504 5364
rect 25556 5352 25562 5364
rect 30466 5352 30472 5364
rect 25556 5324 30472 5352
rect 25556 5312 25562 5324
rect 30466 5312 30472 5324
rect 30524 5312 30530 5364
rect 30745 5355 30803 5361
rect 30745 5321 30757 5355
rect 30791 5352 30803 5355
rect 31202 5352 31208 5364
rect 30791 5324 31208 5352
rect 30791 5321 30803 5324
rect 30745 5315 30803 5321
rect 31202 5312 31208 5324
rect 31260 5312 31266 5364
rect 31754 5312 31760 5364
rect 31812 5312 31818 5364
rect 35618 5352 35624 5364
rect 31864 5324 35624 5352
rect 25593 5287 25651 5293
rect 21468 5256 22416 5284
rect 19337 5219 19395 5225
rect 19337 5185 19349 5219
rect 19383 5185 19395 5219
rect 19337 5179 19395 5185
rect 19521 5219 19579 5225
rect 19521 5185 19533 5219
rect 19567 5215 19579 5219
rect 19567 5187 19656 5215
rect 19567 5185 19579 5187
rect 19521 5179 19579 5185
rect 18877 5151 18935 5157
rect 18877 5148 18889 5151
rect 18064 5120 18889 5148
rect 17957 5111 18015 5117
rect 18877 5117 18889 5120
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 12161 5043 12219 5049
rect 13280 5052 13584 5080
rect 13633 5083 13691 5089
rect 13280 5012 13308 5052
rect 13633 5049 13645 5083
rect 13679 5080 13691 5083
rect 13722 5080 13728 5092
rect 13679 5052 13728 5080
rect 13679 5049 13691 5052
rect 13633 5043 13691 5049
rect 13722 5040 13728 5052
rect 13780 5080 13786 5092
rect 13780 5052 14412 5080
rect 13780 5040 13786 5052
rect 11716 4984 13308 5012
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 13446 5012 13452 5024
rect 13403 4984 13452 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 14277 5015 14335 5021
rect 14277 5012 14289 5015
rect 13964 4984 14289 5012
rect 13964 4972 13970 4984
rect 14277 4981 14289 4984
rect 14323 4981 14335 5015
rect 14384 5012 14412 5052
rect 14734 5040 14740 5092
rect 14792 5080 14798 5092
rect 15289 5083 15347 5089
rect 15289 5080 15301 5083
rect 14792 5052 15301 5080
rect 14792 5040 14798 5052
rect 15289 5049 15301 5052
rect 15335 5049 15347 5083
rect 15289 5043 15347 5049
rect 17681 5083 17739 5089
rect 17681 5049 17693 5083
rect 17727 5080 17739 5083
rect 17972 5080 18000 5111
rect 19058 5108 19064 5160
rect 19116 5108 19122 5160
rect 19150 5108 19156 5160
rect 19208 5148 19214 5160
rect 19628 5148 19656 5187
rect 19702 5176 19708 5228
rect 19760 5216 19766 5228
rect 19996 5216 20024 5244
rect 19760 5188 19932 5216
rect 19996 5188 20208 5216
rect 19760 5176 19766 5188
rect 19208 5140 19380 5148
rect 19444 5140 19656 5148
rect 19208 5120 19656 5140
rect 19208 5108 19214 5120
rect 19352 5112 19472 5120
rect 18969 5083 19027 5089
rect 18969 5080 18981 5083
rect 17727 5052 17908 5080
rect 17972 5052 18981 5080
rect 17727 5049 17739 5052
rect 17681 5043 17739 5049
rect 15194 5012 15200 5024
rect 14384 4984 15200 5012
rect 14277 4975 14335 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 16264 4984 16497 5012
rect 16264 4972 16270 4984
rect 16485 4981 16497 4984
rect 16531 4981 16543 5015
rect 16485 4975 16543 4981
rect 17770 4972 17776 5024
rect 17828 4972 17834 5024
rect 17880 5012 17908 5052
rect 18969 5049 18981 5052
rect 19015 5049 19027 5083
rect 18969 5043 19027 5049
rect 18690 5012 18696 5024
rect 17880 4984 18696 5012
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19245 5015 19303 5021
rect 19245 5012 19257 5015
rect 18840 4984 19257 5012
rect 18840 4972 18846 4984
rect 19245 4981 19257 4984
rect 19291 4981 19303 5015
rect 19628 5012 19656 5120
rect 19794 5108 19800 5160
rect 19852 5108 19858 5160
rect 19904 5148 19932 5188
rect 19981 5151 20039 5157
rect 19981 5148 19993 5151
rect 19904 5120 19993 5148
rect 19981 5117 19993 5120
rect 20027 5148 20039 5151
rect 20070 5148 20076 5160
rect 20027 5120 20076 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 20180 5148 20208 5188
rect 22002 5176 22008 5228
rect 22060 5176 22066 5228
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 22388 5225 22416 5256
rect 25593 5253 25605 5287
rect 25639 5284 25651 5287
rect 25774 5284 25780 5296
rect 25639 5256 25780 5284
rect 25639 5253 25651 5256
rect 25593 5247 25651 5253
rect 25774 5244 25780 5256
rect 25832 5244 25838 5296
rect 25958 5244 25964 5296
rect 26016 5284 26022 5296
rect 26016 5256 26740 5284
rect 26016 5244 26022 5256
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5185 22431 5219
rect 22582 5219 22640 5225
rect 22582 5216 22594 5219
rect 22373 5179 22431 5185
rect 22572 5185 22594 5216
rect 22628 5185 22640 5219
rect 22572 5179 22640 5185
rect 20441 5151 20499 5157
rect 20441 5148 20453 5151
rect 20180 5120 20453 5148
rect 20441 5117 20453 5120
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 20714 5108 20720 5160
rect 20772 5108 20778 5160
rect 20898 5157 20904 5160
rect 20855 5151 20904 5157
rect 20855 5117 20867 5151
rect 20901 5117 20904 5151
rect 20855 5111 20904 5117
rect 20898 5108 20904 5111
rect 20956 5108 20962 5160
rect 20993 5151 21051 5157
rect 20993 5117 21005 5151
rect 21039 5148 21051 5151
rect 21174 5148 21180 5160
rect 21039 5120 21180 5148
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 21174 5108 21180 5120
rect 21232 5148 21238 5160
rect 21818 5148 21824 5160
rect 21232 5120 21824 5148
rect 21232 5108 21238 5120
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 22204 5148 22232 5179
rect 22462 5148 22468 5160
rect 22204 5120 22468 5148
rect 22462 5108 22468 5120
rect 22520 5108 22526 5160
rect 19702 5040 19708 5092
rect 19760 5080 19766 5092
rect 20530 5080 20536 5092
rect 19760 5052 20536 5080
rect 19760 5040 19766 5052
rect 20530 5040 20536 5052
rect 20588 5040 20594 5092
rect 21450 5040 21456 5092
rect 21508 5080 21514 5092
rect 21508 5052 21864 5080
rect 21508 5040 21514 5052
rect 21542 5012 21548 5024
rect 19628 4984 21548 5012
rect 19245 4975 19303 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 21836 5021 21864 5052
rect 22186 5040 22192 5092
rect 22244 5080 22250 5092
rect 22572 5080 22600 5179
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23934 5176 23940 5228
rect 23992 5225 23998 5228
rect 23992 5219 24020 5225
rect 24008 5185 24020 5219
rect 23992 5179 24020 5185
rect 23992 5176 23998 5179
rect 24118 5176 24124 5228
rect 24176 5176 24182 5228
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5215 25743 5219
rect 26602 5216 26608 5228
rect 25792 5215 26608 5216
rect 25731 5188 26608 5215
rect 25731 5187 25820 5188
rect 25731 5185 25743 5187
rect 25685 5179 25743 5185
rect 26602 5176 26608 5188
rect 26660 5176 26666 5228
rect 26712 5216 26740 5256
rect 27080 5256 28994 5284
rect 26970 5216 26976 5228
rect 26712 5188 26976 5216
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 22738 5108 22744 5160
rect 22796 5148 22802 5160
rect 23109 5151 23167 5157
rect 23109 5148 23121 5151
rect 22796 5120 23121 5148
rect 22796 5108 22802 5120
rect 23109 5117 23121 5120
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 22244 5052 22600 5080
rect 23124 5080 23152 5111
rect 23290 5108 23296 5160
rect 23348 5148 23354 5160
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 23348 5120 23857 5148
rect 23348 5108 23354 5120
rect 23845 5117 23857 5120
rect 23891 5148 23903 5151
rect 24486 5148 24492 5160
rect 23891 5120 24492 5148
rect 23891 5117 23903 5120
rect 23845 5111 23903 5117
rect 24486 5108 24492 5120
rect 24544 5108 24550 5160
rect 25317 5151 25375 5157
rect 25317 5117 25329 5151
rect 25363 5148 25375 5151
rect 25590 5148 25596 5160
rect 25363 5120 25596 5148
rect 25363 5117 25375 5120
rect 25317 5111 25375 5117
rect 25590 5108 25596 5120
rect 25648 5108 25654 5160
rect 25866 5108 25872 5160
rect 25924 5148 25930 5160
rect 27080 5148 27108 5256
rect 27338 5176 27344 5228
rect 27396 5216 27402 5228
rect 27709 5219 27767 5225
rect 27709 5216 27721 5219
rect 27396 5188 27721 5216
rect 27396 5176 27402 5188
rect 27705 5187 27721 5188
rect 27709 5185 27721 5187
rect 27755 5185 27767 5219
rect 27709 5179 27767 5185
rect 28258 5176 28264 5228
rect 28316 5176 28322 5228
rect 28966 5216 28994 5256
rect 30558 5244 30564 5296
rect 30616 5284 30622 5296
rect 31864 5284 31892 5324
rect 35618 5312 35624 5324
rect 35676 5312 35682 5364
rect 43162 5352 43168 5364
rect 36556 5324 43168 5352
rect 30616 5256 31892 5284
rect 30616 5244 30622 5256
rect 32030 5244 32036 5296
rect 32088 5284 32094 5296
rect 32088 5256 33732 5284
rect 32088 5244 32094 5256
rect 33704 5228 33732 5256
rect 35710 5244 35716 5296
rect 35768 5284 35774 5296
rect 36556 5284 36584 5324
rect 43162 5312 43168 5324
rect 43220 5312 43226 5364
rect 43438 5312 43444 5364
rect 43496 5312 43502 5364
rect 35768 5256 36584 5284
rect 35768 5244 35774 5256
rect 36630 5244 36636 5296
rect 36688 5284 36694 5296
rect 42702 5284 42708 5296
rect 36688 5256 42708 5284
rect 36688 5244 36694 5256
rect 42702 5244 42708 5256
rect 42760 5244 42766 5296
rect 28966 5188 29132 5216
rect 25924 5120 27108 5148
rect 27985 5151 28043 5157
rect 25924 5108 25930 5120
rect 27985 5117 27997 5151
rect 28031 5117 28043 5151
rect 27985 5111 28043 5117
rect 23569 5083 23627 5089
rect 23124 5052 23428 5080
rect 22244 5040 22250 5052
rect 21821 5015 21879 5021
rect 21821 4981 21833 5015
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 21910 4972 21916 5024
rect 21968 5012 21974 5024
rect 23290 5012 23296 5024
rect 21968 4984 23296 5012
rect 21968 4972 21974 4984
rect 23290 4972 23296 4984
rect 23348 4972 23354 5024
rect 23400 5012 23428 5052
rect 23569 5049 23581 5083
rect 23615 5080 23627 5083
rect 23658 5080 23664 5092
rect 23615 5052 23664 5080
rect 23615 5049 23627 5052
rect 23569 5043 23627 5049
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 25222 5040 25228 5092
rect 25280 5080 25286 5092
rect 26329 5083 26387 5089
rect 26329 5080 26341 5083
rect 25280 5052 26341 5080
rect 25280 5040 25286 5052
rect 26329 5049 26341 5052
rect 26375 5080 26387 5083
rect 26375 5052 27016 5080
rect 26375 5049 26387 5052
rect 26329 5043 26387 5049
rect 26988 5024 27016 5052
rect 24026 5012 24032 5024
rect 23400 4984 24032 5012
rect 24026 4972 24032 4984
rect 24084 4972 24090 5024
rect 25314 4972 25320 5024
rect 25372 4972 25378 5024
rect 25409 5015 25467 5021
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 25777 5015 25835 5021
rect 25777 5012 25789 5015
rect 25455 4984 25789 5012
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 25777 4981 25789 4984
rect 25823 4981 25835 5015
rect 25777 4975 25835 4981
rect 25961 5015 26019 5021
rect 25961 4981 25973 5015
rect 26007 5012 26019 5015
rect 26418 5012 26424 5024
rect 26007 4984 26424 5012
rect 26007 4981 26019 4984
rect 25961 4975 26019 4981
rect 26418 4972 26424 4984
rect 26476 4972 26482 5024
rect 26970 4972 26976 5024
rect 27028 4972 27034 5024
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 27890 5012 27896 5024
rect 27580 4984 27896 5012
rect 27580 4972 27586 4984
rect 27890 4972 27896 4984
rect 27948 5012 27954 5024
rect 28000 5012 28028 5111
rect 28626 5108 28632 5160
rect 28684 5148 28690 5160
rect 28813 5151 28871 5157
rect 28813 5148 28825 5151
rect 28684 5120 28825 5148
rect 28684 5108 28690 5120
rect 28813 5117 28825 5120
rect 28859 5117 28871 5151
rect 28813 5111 28871 5117
rect 28902 5108 28908 5160
rect 28960 5148 28966 5160
rect 28997 5151 29055 5157
rect 28997 5148 29009 5151
rect 28960 5120 29009 5148
rect 28960 5108 28966 5120
rect 28997 5117 29009 5120
rect 29043 5117 29055 5151
rect 29104 5148 29132 5188
rect 29730 5176 29736 5228
rect 29788 5176 29794 5228
rect 30006 5176 30012 5228
rect 30064 5176 30070 5228
rect 30653 5219 30711 5225
rect 30653 5185 30665 5219
rect 30699 5216 30711 5219
rect 30929 5219 30987 5225
rect 30929 5216 30941 5219
rect 30699 5188 30941 5216
rect 30699 5185 30711 5188
rect 30653 5179 30711 5185
rect 30929 5185 30941 5188
rect 30975 5185 30987 5219
rect 30929 5179 30987 5185
rect 31938 5176 31944 5228
rect 31996 5176 32002 5228
rect 32398 5176 32404 5228
rect 32456 5176 32462 5228
rect 33318 5176 33324 5228
rect 33376 5216 33382 5228
rect 33413 5219 33471 5225
rect 33413 5216 33425 5219
rect 33376 5188 33425 5216
rect 33376 5176 33382 5188
rect 33413 5185 33425 5188
rect 33459 5185 33471 5219
rect 33413 5179 33471 5185
rect 33686 5176 33692 5228
rect 33744 5176 33750 5228
rect 34606 5176 34612 5228
rect 34664 5176 34670 5228
rect 34882 5176 34888 5228
rect 34940 5176 34946 5228
rect 35529 5219 35587 5225
rect 35529 5185 35541 5219
rect 35575 5216 35587 5219
rect 35805 5219 35863 5225
rect 35805 5216 35817 5219
rect 35575 5188 35817 5216
rect 35575 5185 35587 5188
rect 35529 5179 35587 5185
rect 35805 5185 35817 5188
rect 35851 5185 35863 5219
rect 35805 5179 35863 5185
rect 36078 5176 36084 5228
rect 36136 5176 36142 5228
rect 36357 5219 36415 5225
rect 36357 5185 36369 5219
rect 36403 5216 36415 5219
rect 36446 5216 36452 5228
rect 36403 5188 36452 5216
rect 36403 5185 36415 5188
rect 36357 5179 36415 5185
rect 36446 5176 36452 5188
rect 36504 5176 36510 5228
rect 37458 5176 37464 5228
rect 37516 5216 37522 5228
rect 37553 5219 37611 5225
rect 37553 5216 37565 5219
rect 37516 5188 37565 5216
rect 37516 5176 37522 5188
rect 37553 5185 37565 5188
rect 37599 5185 37611 5219
rect 37553 5179 37611 5185
rect 39206 5176 39212 5228
rect 39264 5176 39270 5228
rect 42886 5176 42892 5228
rect 42944 5176 42950 5228
rect 43254 5176 43260 5228
rect 43312 5176 43318 5228
rect 29850 5151 29908 5157
rect 29850 5148 29862 5151
rect 29104 5120 29862 5148
rect 28997 5111 29055 5117
rect 29850 5117 29862 5120
rect 29896 5148 29908 5151
rect 30558 5148 30564 5160
rect 29896 5120 30564 5148
rect 29896 5117 29908 5120
rect 29850 5111 29908 5117
rect 30558 5108 30564 5120
rect 30616 5108 30622 5160
rect 31570 5108 31576 5160
rect 31628 5148 31634 5160
rect 32125 5151 32183 5157
rect 32125 5148 32137 5151
rect 31628 5120 32137 5148
rect 31628 5108 31634 5120
rect 32125 5117 32137 5120
rect 32171 5117 32183 5151
rect 32125 5111 32183 5117
rect 33873 5151 33931 5157
rect 33873 5117 33885 5151
rect 33919 5117 33931 5151
rect 33873 5111 33931 5117
rect 34333 5151 34391 5157
rect 34333 5117 34345 5151
rect 34379 5117 34391 5151
rect 34333 5111 34391 5117
rect 28534 5040 28540 5092
rect 28592 5080 28598 5092
rect 28920 5080 28948 5108
rect 28592 5052 28948 5080
rect 28592 5040 28598 5052
rect 29454 5040 29460 5092
rect 29512 5040 29518 5092
rect 30926 5040 30932 5092
rect 30984 5080 30990 5092
rect 31294 5080 31300 5092
rect 30984 5052 31300 5080
rect 30984 5040 30990 5052
rect 31294 5040 31300 5052
rect 31352 5040 31358 5092
rect 33888 5080 33916 5111
rect 32784 5052 33916 5080
rect 34348 5080 34376 5111
rect 34422 5108 34428 5160
rect 34480 5148 34486 5160
rect 34747 5151 34805 5157
rect 34747 5148 34759 5151
rect 34480 5120 34759 5148
rect 34480 5108 34486 5120
rect 34747 5117 34759 5120
rect 34793 5148 34805 5151
rect 34793 5120 35756 5148
rect 34793 5117 34805 5120
rect 34747 5111 34805 5117
rect 34348 5052 34468 5080
rect 27948 4984 28028 5012
rect 27948 4972 27954 4984
rect 28074 4972 28080 5024
rect 28132 4972 28138 5024
rect 28166 4972 28172 5024
rect 28224 5012 28230 5024
rect 29178 5012 29184 5024
rect 28224 4984 29184 5012
rect 28224 4972 28230 4984
rect 29178 4972 29184 4984
rect 29236 4972 29242 5024
rect 31478 4972 31484 5024
rect 31536 5012 31542 5024
rect 32784 5012 32812 5052
rect 31536 4984 32812 5012
rect 31536 4972 31542 4984
rect 33042 4972 33048 5024
rect 33100 5012 33106 5024
rect 33137 5015 33195 5021
rect 33137 5012 33149 5015
rect 33100 4984 33149 5012
rect 33100 4972 33106 4984
rect 33137 4981 33149 4984
rect 33183 4981 33195 5015
rect 33137 4975 33195 4981
rect 33229 5015 33287 5021
rect 33229 4981 33241 5015
rect 33275 5012 33287 5015
rect 33686 5012 33692 5024
rect 33275 4984 33692 5012
rect 33275 4981 33287 4984
rect 33229 4975 33287 4981
rect 33686 4972 33692 4984
rect 33744 4972 33750 5024
rect 34440 5012 34468 5052
rect 34698 5012 34704 5024
rect 34440 4984 34704 5012
rect 34698 4972 34704 4984
rect 34756 4972 34762 5024
rect 35250 4972 35256 5024
rect 35308 5012 35314 5024
rect 35621 5015 35679 5021
rect 35621 5012 35633 5015
rect 35308 4984 35633 5012
rect 35308 4972 35314 4984
rect 35621 4981 35633 4984
rect 35667 4981 35679 5015
rect 35728 5012 35756 5120
rect 37182 5108 37188 5160
rect 37240 5148 37246 5160
rect 37277 5151 37335 5157
rect 37277 5148 37289 5151
rect 37240 5120 37289 5148
rect 37240 5108 37246 5120
rect 37277 5117 37289 5120
rect 37323 5117 37335 5151
rect 37277 5111 37335 5117
rect 39485 5151 39543 5157
rect 39485 5117 39497 5151
rect 39531 5117 39543 5151
rect 39485 5111 39543 5117
rect 36906 5080 36912 5092
rect 36740 5052 36912 5080
rect 36740 5012 36768 5052
rect 36906 5040 36912 5052
rect 36964 5040 36970 5092
rect 38470 5040 38476 5092
rect 38528 5040 38534 5092
rect 35728 4984 36768 5012
rect 35621 4975 35679 4981
rect 36814 4972 36820 5024
rect 36872 5012 36878 5024
rect 37093 5015 37151 5021
rect 37093 5012 37105 5015
rect 36872 4984 37105 5012
rect 36872 4972 36878 4984
rect 37093 4981 37105 4984
rect 37139 4981 37151 5015
rect 37093 4975 37151 4981
rect 37366 4972 37372 5024
rect 37424 5012 37430 5024
rect 38289 5015 38347 5021
rect 38289 5012 38301 5015
rect 37424 4984 38301 5012
rect 37424 4972 37430 4984
rect 38289 4981 38301 4984
rect 38335 4981 38347 5015
rect 38289 4975 38347 4981
rect 38654 4972 38660 5024
rect 38712 5012 38718 5024
rect 39500 5012 39528 5111
rect 38712 4984 39528 5012
rect 38712 4972 38718 4984
rect 43070 4972 43076 5024
rect 43128 4972 43134 5024
rect 1104 4922 43884 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13918 4922
rect 13970 4870 13982 4922
rect 14034 4870 14046 4922
rect 14098 4870 14110 4922
rect 14162 4870 14174 4922
rect 14226 4870 14238 4922
rect 14290 4870 19918 4922
rect 19970 4870 19982 4922
rect 20034 4870 20046 4922
rect 20098 4870 20110 4922
rect 20162 4870 20174 4922
rect 20226 4870 20238 4922
rect 20290 4870 25918 4922
rect 25970 4870 25982 4922
rect 26034 4870 26046 4922
rect 26098 4870 26110 4922
rect 26162 4870 26174 4922
rect 26226 4870 26238 4922
rect 26290 4870 31918 4922
rect 31970 4870 31982 4922
rect 32034 4870 32046 4922
rect 32098 4870 32110 4922
rect 32162 4870 32174 4922
rect 32226 4870 32238 4922
rect 32290 4870 37918 4922
rect 37970 4870 37982 4922
rect 38034 4870 38046 4922
rect 38098 4870 38110 4922
rect 38162 4870 38174 4922
rect 38226 4870 38238 4922
rect 38290 4870 43884 4922
rect 1104 4848 43884 4870
rect 3418 4768 3424 4820
rect 3476 4768 3482 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3752 4780 7052 4808
rect 3752 4768 3758 4780
rect 5905 4743 5963 4749
rect 5905 4740 5917 4743
rect 5736 4712 5917 4740
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 3602 4672 3608 4684
rect 3384 4644 3608 4672
rect 3384 4632 3390 4644
rect 3602 4632 3608 4644
rect 3660 4672 3666 4684
rect 3789 4675 3847 4681
rect 3789 4672 3801 4675
rect 3660 4644 3801 4672
rect 3660 4632 3666 4644
rect 3789 4641 3801 4644
rect 3835 4641 3847 4675
rect 3789 4635 3847 4641
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 4856 4644 5457 4672
rect 4856 4632 4862 4644
rect 5445 4641 5457 4644
rect 5491 4672 5503 4675
rect 5534 4672 5540 4684
rect 5491 4644 5540 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5736 4672 5764 4712
rect 5905 4709 5917 4712
rect 5951 4709 5963 4743
rect 5905 4703 5963 4709
rect 5644 4644 5764 4672
rect 1394 4564 1400 4616
rect 1452 4604 1458 4616
rect 1489 4607 1547 4613
rect 1489 4604 1501 4607
rect 1452 4576 1501 4604
rect 1452 4564 1458 4576
rect 1489 4573 1501 4576
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1857 4607 1915 4613
rect 1857 4604 1869 4607
rect 1728 4576 1869 4604
rect 1728 4564 1734 4576
rect 1857 4573 1869 4576
rect 1903 4573 1915 4607
rect 1857 4567 1915 4573
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 2590 4604 2596 4616
rect 2455 4576 2596 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2774 4604 2780 4616
rect 2731 4576 2780 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 2774 4564 2780 4576
rect 2832 4604 2838 4616
rect 3050 4604 3056 4616
rect 2832 4576 3056 4604
rect 2832 4564 2838 4576
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3896 4576 4077 4604
rect 2038 4496 2044 4548
rect 2096 4496 2102 4548
rect 3142 4496 3148 4548
rect 3200 4536 3206 4548
rect 3896 4536 3924 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5644 4604 5672 4644
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 5868 4644 6193 4672
rect 5868 4632 5874 4644
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 6454 4632 6460 4684
rect 6512 4632 6518 4684
rect 5261 4567 5319 4573
rect 5368 4576 5672 4604
rect 3200 4508 3924 4536
rect 3200 4496 3206 4508
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4468 1639 4471
rect 2498 4468 2504 4480
rect 1627 4440 2504 4468
rect 1627 4437 1639 4440
rect 1581 4431 1639 4437
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 4798 4428 4804 4480
rect 4856 4428 4862 4480
rect 5074 4428 5080 4480
rect 5132 4428 5138 4480
rect 5276 4468 5304 4567
rect 5368 4548 5396 4576
rect 6270 4564 6276 4616
rect 6328 4613 6334 4616
rect 6328 4607 6356 4613
rect 6344 4573 6356 4607
rect 7024 4604 7052 4780
rect 7098 4768 7104 4820
rect 7156 4768 7162 4820
rect 7760 4780 8524 4808
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 7760 4681 7788 4780
rect 8496 4740 8524 4780
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 8757 4811 8815 4817
rect 8757 4808 8769 4811
rect 8628 4780 8769 4808
rect 8628 4768 8634 4780
rect 8757 4777 8769 4780
rect 8803 4777 8815 4811
rect 8757 4771 8815 4777
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 9122 4808 9128 4820
rect 8987 4780 9128 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 11425 4811 11483 4817
rect 9364 4780 11376 4808
rect 9364 4768 9370 4780
rect 9030 4740 9036 4752
rect 8496 4712 9036 4740
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 11348 4740 11376 4780
rect 11425 4777 11437 4811
rect 11471 4808 11483 4811
rect 12710 4808 12716 4820
rect 11471 4780 12716 4808
rect 11471 4777 11483 4780
rect 11425 4771 11483 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 12986 4768 12992 4820
rect 13044 4768 13050 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14366 4808 14372 4820
rect 14139 4780 14372 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14734 4808 14740 4820
rect 14476 4780 14740 4808
rect 11790 4740 11796 4752
rect 11348 4712 11796 4740
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 13004 4740 13032 4768
rect 12912 4712 13032 4740
rect 13909 4743 13967 4749
rect 7745 4675 7803 4681
rect 7745 4672 7757 4675
rect 7616 4644 7757 4672
rect 7616 4632 7622 4644
rect 7745 4641 7757 4644
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 9950 4632 9956 4684
rect 10008 4672 10014 4684
rect 10318 4672 10324 4684
rect 10008 4644 10324 4672
rect 10008 4632 10014 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 12802 4672 12808 4684
rect 12544 4644 12808 4672
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7024 4576 8033 4604
rect 6328 4567 6356 4573
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 6328 4564 6334 4567
rect 5350 4496 5356 4548
rect 5408 4496 5414 4548
rect 7190 4496 7196 4548
rect 7248 4536 7254 4548
rect 7469 4539 7527 4545
rect 7469 4536 7481 4539
rect 7248 4508 7481 4536
rect 7248 4496 7254 4508
rect 7469 4505 7481 4508
rect 7515 4536 7527 4539
rect 7742 4536 7748 4548
rect 7515 4508 7748 4536
rect 7515 4505 7527 4508
rect 7469 4499 7527 4505
rect 7742 4496 7748 4508
rect 7800 4496 7806 4548
rect 8036 4536 8064 4567
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9732 4576 9774 4604
rect 9732 4564 9738 4576
rect 10410 4564 10416 4616
rect 10468 4564 10474 4616
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11480 4576 11805 4604
rect 11480 4564 11486 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 10137 4539 10195 4545
rect 8036 4508 9674 4536
rect 6730 4468 6736 4480
rect 5276 4440 6736 4468
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7558 4428 7564 4480
rect 7616 4428 7622 4480
rect 9646 4468 9674 4508
rect 10137 4505 10149 4539
rect 10183 4536 10195 4539
rect 11146 4536 11152 4548
rect 10183 4508 11152 4536
rect 10183 4505 10195 4508
rect 10137 4499 10195 4505
rect 10152 4468 10180 4499
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11808 4536 11836 4567
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 12544 4604 12572 4644
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 12912 4681 12940 4712
rect 13909 4709 13921 4743
rect 13955 4740 13967 4743
rect 14476 4740 14504 4780
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 14884 4780 15056 4808
rect 14884 4768 14890 4780
rect 13955 4712 14504 4740
rect 15028 4740 15056 4780
rect 15102 4768 15108 4820
rect 15160 4808 15166 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15160 4780 15945 4808
rect 15160 4768 15166 4780
rect 15933 4777 15945 4780
rect 15979 4777 15991 4811
rect 16850 4808 16856 4820
rect 15933 4771 15991 4777
rect 16500 4780 16856 4808
rect 15197 4743 15255 4749
rect 15028 4712 15148 4740
rect 13955 4709 13967 4712
rect 13909 4703 13967 4709
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4641 12955 4675
rect 15120 4672 15148 4712
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 15378 4740 15384 4752
rect 15243 4712 15384 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 15473 4743 15531 4749
rect 15473 4709 15485 4743
rect 15519 4740 15531 4743
rect 15562 4740 15568 4752
rect 15519 4712 15568 4740
rect 15519 4709 15531 4712
rect 15473 4703 15531 4709
rect 15562 4700 15568 4712
rect 15620 4700 15626 4752
rect 16390 4672 16396 4684
rect 15120 4644 16396 4672
rect 12897 4635 12955 4641
rect 15580 4616 15608 4644
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 16500 4681 16528 4780
rect 16850 4768 16856 4780
rect 16908 4808 16914 4820
rect 17310 4808 17316 4820
rect 16908 4780 17316 4808
rect 16908 4768 16914 4780
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 17494 4768 17500 4820
rect 17552 4768 17558 4820
rect 18046 4768 18052 4820
rect 18104 4768 18110 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 19150 4808 19156 4820
rect 18380 4780 19156 4808
rect 18380 4768 18386 4780
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4777 19671 4811
rect 20898 4808 20904 4820
rect 19613 4771 19671 4777
rect 19720 4780 20904 4808
rect 17586 4700 17592 4752
rect 17644 4740 17650 4752
rect 17773 4743 17831 4749
rect 17773 4740 17785 4743
rect 17644 4712 17785 4740
rect 17644 4700 17650 4712
rect 17773 4709 17785 4712
rect 17819 4709 17831 4743
rect 18064 4740 18092 4768
rect 17773 4703 17831 4709
rect 18039 4712 18092 4740
rect 18233 4743 18291 4749
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4641 16543 4675
rect 18039 4672 18067 4712
rect 18233 4709 18245 4743
rect 18279 4740 18291 4743
rect 18414 4740 18420 4752
rect 18279 4712 18420 4740
rect 18279 4709 18291 4712
rect 18233 4703 18291 4709
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 19242 4700 19248 4752
rect 19300 4700 19306 4752
rect 18095 4675 18153 4681
rect 18095 4672 18107 4675
rect 18039 4644 18107 4672
rect 16485 4635 16543 4641
rect 18095 4641 18107 4644
rect 18141 4641 18153 4675
rect 18095 4635 18153 4641
rect 18598 4632 18604 4684
rect 18656 4672 18662 4684
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 18656 4644 18705 4672
rect 18656 4632 18662 4644
rect 18693 4641 18705 4644
rect 18739 4641 18751 4675
rect 18693 4635 18751 4641
rect 18782 4632 18788 4684
rect 18840 4672 18846 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 18840 4644 19533 4672
rect 18840 4632 18846 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 12176 4576 12572 4604
rect 12176 4536 12204 4576
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 13173 4607 13231 4613
rect 13173 4604 13185 4607
rect 12676 4576 13185 4604
rect 12676 4564 12682 4576
rect 13173 4573 13185 4576
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14366 4604 14372 4616
rect 14148 4576 14372 4604
rect 14148 4564 14154 4576
rect 14366 4564 14372 4576
rect 14424 4604 14430 4616
rect 14829 4607 14887 4613
rect 14829 4604 14841 4607
rect 14424 4576 14841 4604
rect 14424 4564 14430 4576
rect 14829 4573 14841 4576
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14976 4576 15117 4604
rect 14976 4564 14982 4576
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15286 4564 15292 4616
rect 15344 4604 15350 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 15344 4576 15393 4604
rect 15344 4564 15350 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 15562 4564 15568 4616
rect 15620 4564 15626 4616
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16206 4604 16212 4616
rect 16163 4576 16212 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 16776 4536 16804 4567
rect 17678 4564 17684 4616
rect 17736 4564 17742 4616
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 18008 4607 18066 4613
rect 18008 4573 18020 4607
rect 18054 4604 18066 4607
rect 19058 4604 19064 4616
rect 18054 4576 19064 4604
rect 18054 4573 18066 4576
rect 18008 4567 18066 4573
rect 11808 4508 12204 4536
rect 12248 4508 16804 4536
rect 17880 4536 17908 4567
rect 19058 4564 19064 4576
rect 19116 4604 19122 4616
rect 19628 4604 19656 4771
rect 19116 4576 19656 4604
rect 19116 4564 19122 4576
rect 18782 4536 18788 4548
rect 17880 4508 18788 4536
rect 9646 4440 10180 4468
rect 10226 4428 10232 4480
rect 10284 4428 10290 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 12248 4468 12276 4508
rect 18782 4496 18788 4508
rect 18840 4496 18846 4548
rect 19720 4536 19748 4780
rect 20898 4768 20904 4780
rect 20956 4808 20962 4820
rect 22002 4808 22008 4820
rect 20956 4780 22008 4808
rect 20956 4768 20962 4780
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22189 4811 22247 4817
rect 22189 4808 22201 4811
rect 22152 4780 22201 4808
rect 22152 4768 22158 4780
rect 22189 4777 22201 4780
rect 22235 4777 22247 4811
rect 22189 4771 22247 4777
rect 22278 4768 22284 4820
rect 22336 4808 22342 4820
rect 25041 4811 25099 4817
rect 22336 4780 23612 4808
rect 22336 4768 22342 4780
rect 19812 4712 20668 4740
rect 19812 4613 19840 4712
rect 20073 4675 20131 4681
rect 20073 4641 20085 4675
rect 20119 4672 20131 4675
rect 20254 4672 20260 4684
rect 20119 4644 20260 4672
rect 20119 4641 20131 4644
rect 20073 4635 20131 4641
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 20530 4632 20536 4684
rect 20588 4632 20594 4684
rect 20640 4672 20668 4712
rect 21542 4700 21548 4752
rect 21600 4700 21606 4752
rect 21726 4700 21732 4752
rect 21784 4740 21790 4752
rect 22296 4740 22324 4768
rect 23584 4749 23612 4780
rect 25041 4777 25053 4811
rect 25087 4808 25099 4811
rect 25317 4811 25375 4817
rect 25317 4808 25329 4811
rect 25087 4780 25329 4808
rect 25087 4777 25099 4780
rect 25041 4771 25099 4777
rect 25317 4777 25329 4780
rect 25363 4808 25375 4811
rect 26050 4808 26056 4820
rect 25363 4780 26056 4808
rect 25363 4777 25375 4780
rect 25317 4771 25375 4777
rect 26050 4768 26056 4780
rect 26108 4808 26114 4820
rect 26418 4808 26424 4820
rect 26108 4780 26424 4808
rect 26108 4768 26114 4780
rect 26418 4768 26424 4780
rect 26476 4768 26482 4820
rect 26605 4811 26663 4817
rect 26605 4777 26617 4811
rect 26651 4808 26663 4811
rect 26970 4808 26976 4820
rect 26651 4780 26976 4808
rect 26651 4777 26663 4780
rect 26605 4771 26663 4777
rect 26970 4768 26976 4780
rect 27028 4808 27034 4820
rect 27798 4808 27804 4820
rect 27028 4780 27804 4808
rect 27028 4768 27034 4780
rect 27798 4768 27804 4780
rect 27856 4768 27862 4820
rect 29273 4811 29331 4817
rect 28000 4780 29224 4808
rect 21784 4712 22324 4740
rect 23569 4743 23627 4749
rect 21784 4700 21790 4712
rect 23569 4709 23581 4743
rect 23615 4709 23627 4743
rect 23569 4703 23627 4709
rect 20806 4672 20812 4684
rect 20640 4644 20812 4672
rect 20806 4632 20812 4644
rect 20864 4672 20870 4684
rect 21560 4672 21588 4700
rect 20864 4644 21588 4672
rect 20864 4632 20870 4644
rect 21634 4632 21640 4684
rect 21692 4672 21698 4684
rect 23198 4681 23204 4684
rect 23017 4675 23075 4681
rect 23017 4672 23029 4675
rect 21692 4644 23029 4672
rect 21692 4632 21698 4644
rect 23017 4641 23029 4644
rect 23063 4641 23075 4675
rect 23017 4635 23075 4641
rect 23176 4675 23204 4681
rect 23176 4641 23188 4675
rect 23176 4635 23204 4641
rect 23198 4632 23204 4635
rect 23256 4632 23262 4684
rect 23290 4632 23296 4684
rect 23348 4632 23354 4684
rect 27801 4675 27859 4681
rect 26418 4621 26424 4673
rect 26476 4621 26482 4673
rect 27801 4641 27813 4675
rect 27847 4672 27859 4675
rect 27890 4672 27896 4684
rect 27847 4644 27896 4672
rect 27847 4641 27859 4644
rect 27801 4635 27859 4641
rect 27890 4632 27896 4644
rect 27948 4632 27954 4684
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4573 19855 4607
rect 19797 4567 19855 4573
rect 19886 4564 19892 4616
rect 19944 4564 19950 4616
rect 20898 4564 20904 4616
rect 20956 4613 20962 4616
rect 20956 4607 20984 4613
rect 20972 4573 20984 4607
rect 20956 4567 20984 4573
rect 20956 4564 20962 4567
rect 21082 4564 21088 4616
rect 21140 4564 21146 4616
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 21652 4576 22017 4604
rect 21652 4536 21680 4576
rect 22005 4573 22017 4576
rect 22051 4604 22063 4607
rect 22186 4604 22192 4616
rect 22051 4576 22192 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 24026 4564 24032 4616
rect 24084 4564 24090 4616
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 24673 4607 24731 4613
rect 24673 4573 24685 4607
rect 24719 4604 24731 4607
rect 24762 4604 24768 4616
rect 24719 4576 24768 4604
rect 24719 4573 24731 4576
rect 24673 4567 24731 4573
rect 18892 4508 19748 4536
rect 21560 4508 21680 4536
rect 11112 4440 12276 4468
rect 12805 4471 12863 4477
rect 11112 4428 11118 4440
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 13354 4468 13360 4480
rect 12851 4440 13360 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14550 4468 14556 4480
rect 13780 4440 14556 4468
rect 13780 4428 13786 4440
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 18601 4471 18659 4477
rect 18601 4468 18613 4471
rect 15528 4440 18613 4468
rect 15528 4428 15534 4440
rect 18601 4437 18613 4440
rect 18647 4468 18659 4471
rect 18892 4468 18920 4508
rect 18647 4440 18920 4468
rect 18647 4437 18659 4440
rect 18601 4431 18659 4437
rect 19058 4428 19064 4480
rect 19116 4468 19122 4480
rect 21560 4468 21588 4508
rect 21818 4496 21824 4548
rect 21876 4496 21882 4548
rect 24228 4536 24256 4567
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 25041 4607 25099 4613
rect 25041 4573 25053 4607
rect 25087 4604 25099 4607
rect 25222 4604 25228 4616
rect 25087 4576 25228 4604
rect 25087 4573 25099 4576
rect 25041 4567 25099 4573
rect 25222 4564 25228 4576
rect 25280 4604 25286 4616
rect 25406 4604 25412 4616
rect 25280 4576 25412 4604
rect 25280 4564 25286 4576
rect 25406 4564 25412 4576
rect 25464 4564 25470 4616
rect 25958 4564 25964 4616
rect 26016 4604 26022 4616
rect 26053 4607 26111 4613
rect 26053 4604 26065 4607
rect 26016 4576 26065 4604
rect 26016 4564 26022 4576
rect 26053 4573 26065 4576
rect 26099 4573 26111 4607
rect 26053 4567 26111 4573
rect 26326 4564 26332 4616
rect 26384 4564 26390 4616
rect 26694 4564 26700 4616
rect 26752 4564 26758 4616
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27525 4607 27583 4613
rect 27525 4604 27537 4607
rect 27488 4576 27537 4604
rect 27488 4564 27494 4576
rect 27525 4573 27537 4576
rect 27571 4573 27583 4607
rect 27525 4567 27583 4573
rect 27614 4564 27620 4616
rect 27672 4604 27678 4616
rect 28000 4604 28028 4780
rect 29196 4740 29224 4780
rect 29273 4777 29285 4811
rect 29319 4808 29331 4811
rect 30006 4808 30012 4820
rect 29319 4780 30012 4808
rect 29319 4777 29331 4780
rect 29273 4771 29331 4777
rect 30006 4768 30012 4780
rect 30064 4768 30070 4820
rect 30558 4808 30564 4820
rect 30208 4780 30564 4808
rect 29730 4740 29736 4752
rect 29196 4712 29736 4740
rect 29730 4700 29736 4712
rect 29788 4740 29794 4752
rect 30208 4749 30236 4780
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 31386 4768 31392 4820
rect 31444 4808 31450 4820
rect 32582 4808 32588 4820
rect 31444 4780 32588 4808
rect 31444 4768 31450 4780
rect 32582 4768 32588 4780
rect 32640 4808 32646 4820
rect 32640 4780 33088 4808
rect 32640 4768 32646 4780
rect 30193 4743 30251 4749
rect 29788 4712 29868 4740
rect 29788 4700 29794 4712
rect 28258 4632 28264 4684
rect 28316 4632 28322 4684
rect 28902 4632 28908 4684
rect 28960 4672 28966 4684
rect 29840 4672 29868 4712
rect 30193 4709 30205 4743
rect 30239 4709 30251 4743
rect 30193 4703 30251 4709
rect 30650 4681 30656 4684
rect 30469 4675 30527 4681
rect 30469 4672 30481 4675
rect 28960 4644 29776 4672
rect 29840 4644 30481 4672
rect 28960 4632 28966 4644
rect 27672 4576 28028 4604
rect 27672 4564 27678 4576
rect 28534 4564 28540 4616
rect 28592 4564 28598 4616
rect 28626 4564 28632 4616
rect 28684 4604 28690 4616
rect 29748 4613 29776 4644
rect 30469 4641 30481 4644
rect 30515 4641 30527 4675
rect 30469 4635 30527 4641
rect 30607 4675 30656 4681
rect 30607 4641 30619 4675
rect 30653 4641 30656 4675
rect 30607 4635 30656 4641
rect 30650 4632 30656 4635
rect 30708 4672 30714 4684
rect 31665 4675 31723 4681
rect 31665 4672 31677 4675
rect 30708 4644 31677 4672
rect 30708 4632 30714 4644
rect 31665 4641 31677 4644
rect 31711 4641 31723 4675
rect 31665 4635 31723 4641
rect 31754 4632 31760 4684
rect 31812 4672 31818 4684
rect 32125 4675 32183 4681
rect 32125 4672 32137 4675
rect 31812 4644 32137 4672
rect 31812 4632 31818 4644
rect 32125 4641 32137 4644
rect 32171 4641 32183 4675
rect 32125 4635 32183 4641
rect 32398 4632 32404 4684
rect 32456 4632 32462 4684
rect 33060 4672 33088 4780
rect 33318 4768 33324 4820
rect 33376 4768 33382 4820
rect 34054 4768 34060 4820
rect 34112 4808 34118 4820
rect 36630 4808 36636 4820
rect 34112 4780 36636 4808
rect 34112 4768 34118 4780
rect 36630 4768 36636 4780
rect 36688 4768 36694 4820
rect 39485 4811 39543 4817
rect 39485 4808 39497 4811
rect 36740 4780 39497 4808
rect 35066 4700 35072 4752
rect 35124 4700 35130 4752
rect 36538 4700 36544 4752
rect 36596 4740 36602 4752
rect 36740 4740 36768 4780
rect 39485 4777 39497 4780
rect 39531 4777 39543 4811
rect 39485 4771 39543 4777
rect 39758 4768 39764 4820
rect 39816 4808 39822 4820
rect 42886 4808 42892 4820
rect 39816 4780 42892 4808
rect 39816 4768 39822 4780
rect 42886 4768 42892 4780
rect 42944 4768 42950 4820
rect 36596 4712 36768 4740
rect 36596 4700 36602 4712
rect 36814 4700 36820 4752
rect 36872 4700 36878 4752
rect 43438 4700 43444 4752
rect 43496 4700 43502 4752
rect 37210 4675 37268 4681
rect 37210 4672 37222 4675
rect 33060 4644 37222 4672
rect 37210 4641 37222 4644
rect 37256 4641 37268 4675
rect 37210 4635 37268 4641
rect 37366 4632 37372 4684
rect 37424 4632 37430 4684
rect 37550 4632 37556 4684
rect 37608 4672 37614 4684
rect 37608 4644 37964 4672
rect 37608 4632 37614 4644
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 28684 4576 29561 4604
rect 28684 4564 28690 4576
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 29733 4607 29791 4613
rect 29733 4573 29745 4607
rect 29779 4573 29791 4607
rect 29733 4567 29791 4573
rect 28902 4536 28908 4548
rect 24228 4508 28908 4536
rect 19116 4440 21588 4468
rect 21729 4471 21787 4477
rect 19116 4428 19122 4440
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 22094 4468 22100 4480
rect 21775 4440 22100 4468
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 22370 4428 22376 4480
rect 22428 4428 22434 4480
rect 22922 4428 22928 4480
rect 22980 4468 22986 4480
rect 24228 4468 24256 4508
rect 28902 4496 28908 4508
rect 28960 4496 28966 4548
rect 22980 4440 24256 4468
rect 22980 4428 22986 4440
rect 25222 4428 25228 4480
rect 25280 4428 25286 4480
rect 25590 4428 25596 4480
rect 25648 4468 25654 4480
rect 25958 4468 25964 4480
rect 25648 4440 25964 4468
rect 25648 4428 25654 4440
rect 25958 4428 25964 4440
rect 26016 4428 26022 4480
rect 26418 4428 26424 4480
rect 26476 4428 26482 4480
rect 26694 4428 26700 4480
rect 26752 4468 26758 4480
rect 26789 4471 26847 4477
rect 26789 4468 26801 4471
rect 26752 4440 26801 4468
rect 26752 4428 26758 4440
rect 26789 4437 26801 4440
rect 26835 4437 26847 4471
rect 29564 4468 29592 4567
rect 30742 4564 30748 4616
rect 30800 4564 30806 4616
rect 31478 4564 31484 4616
rect 31536 4564 31542 4616
rect 32582 4613 32588 4616
rect 32539 4607 32588 4613
rect 32539 4573 32551 4607
rect 32585 4573 32588 4607
rect 32539 4567 32588 4573
rect 32582 4564 32588 4567
rect 32640 4564 32646 4616
rect 32674 4564 32680 4616
rect 32732 4564 32738 4616
rect 34057 4607 34115 4613
rect 34057 4573 34069 4607
rect 34103 4604 34115 4607
rect 34146 4604 34152 4616
rect 34103 4576 34152 4604
rect 34103 4573 34115 4576
rect 34057 4567 34115 4573
rect 34146 4564 34152 4576
rect 34204 4564 34210 4616
rect 35253 4607 35311 4613
rect 35253 4573 35265 4607
rect 35299 4604 35311 4607
rect 36078 4604 36084 4616
rect 35299 4576 36084 4604
rect 35299 4573 35311 4576
rect 35253 4567 35311 4573
rect 36078 4564 36084 4576
rect 36136 4564 36142 4616
rect 36173 4607 36231 4613
rect 36173 4573 36185 4607
rect 36219 4573 36231 4607
rect 36173 4567 36231 4573
rect 31294 4496 31300 4548
rect 31352 4536 31358 4548
rect 31352 4508 31708 4536
rect 31352 4496 31358 4508
rect 30466 4468 30472 4480
rect 29564 4440 30472 4468
rect 26789 4431 26847 4437
rect 30466 4428 30472 4440
rect 30524 4428 30530 4480
rect 30650 4428 30656 4480
rect 30708 4468 30714 4480
rect 31389 4471 31447 4477
rect 31389 4468 31401 4471
rect 30708 4440 31401 4468
rect 30708 4428 30714 4440
rect 31389 4437 31401 4440
rect 31435 4437 31447 4471
rect 31680 4468 31708 4508
rect 34238 4496 34244 4548
rect 34296 4496 34302 4548
rect 32950 4468 32956 4480
rect 31680 4440 32956 4468
rect 31389 4431 31447 4437
rect 32950 4428 32956 4440
rect 33008 4428 33014 4480
rect 33502 4428 33508 4480
rect 33560 4468 33566 4480
rect 36188 4468 36216 4567
rect 36354 4564 36360 4616
rect 36412 4564 36418 4616
rect 37090 4564 37096 4616
rect 37148 4564 37154 4616
rect 37936 4604 37964 4644
rect 38378 4632 38384 4684
rect 38436 4672 38442 4684
rect 38473 4675 38531 4681
rect 38473 4672 38485 4675
rect 38436 4644 38485 4672
rect 38436 4632 38442 4644
rect 38473 4641 38485 4644
rect 38519 4641 38531 4675
rect 38473 4635 38531 4641
rect 38488 4604 38516 4635
rect 38654 4604 38660 4616
rect 37936 4576 38424 4604
rect 38488 4576 38660 4604
rect 38013 4539 38071 4545
rect 38013 4505 38025 4539
rect 38059 4536 38071 4539
rect 38289 4539 38347 4545
rect 38289 4536 38301 4539
rect 38059 4508 38301 4536
rect 38059 4505 38071 4508
rect 38013 4499 38071 4505
rect 38289 4505 38301 4508
rect 38335 4505 38347 4539
rect 38396 4536 38424 4576
rect 38654 4564 38660 4576
rect 38712 4564 38718 4616
rect 38749 4607 38807 4613
rect 38749 4573 38761 4607
rect 38795 4573 38807 4607
rect 38749 4567 38807 4573
rect 38764 4536 38792 4567
rect 42794 4564 42800 4616
rect 42852 4604 42858 4616
rect 42889 4607 42947 4613
rect 42889 4604 42901 4607
rect 42852 4576 42901 4604
rect 42852 4564 42858 4576
rect 42889 4573 42901 4576
rect 42935 4573 42947 4607
rect 42889 4567 42947 4573
rect 43162 4564 43168 4616
rect 43220 4604 43226 4616
rect 43257 4607 43315 4613
rect 43257 4604 43269 4607
rect 43220 4576 43269 4604
rect 43220 4564 43226 4576
rect 43257 4573 43269 4576
rect 43303 4573 43315 4607
rect 43257 4567 43315 4573
rect 38396 4508 38792 4536
rect 38289 4499 38347 4505
rect 36630 4468 36636 4480
rect 33560 4440 36636 4468
rect 33560 4428 33566 4440
rect 36630 4428 36636 4440
rect 36688 4428 36694 4480
rect 37274 4428 37280 4480
rect 37332 4468 37338 4480
rect 38197 4471 38255 4477
rect 38197 4468 38209 4471
rect 37332 4440 38209 4468
rect 37332 4428 37338 4440
rect 38197 4437 38209 4440
rect 38243 4437 38255 4471
rect 38197 4431 38255 4437
rect 43070 4428 43076 4480
rect 43128 4428 43134 4480
rect 1104 4378 43884 4400
rect 1104 4326 2658 4378
rect 2710 4326 2722 4378
rect 2774 4326 2786 4378
rect 2838 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 8658 4378
rect 8710 4326 8722 4378
rect 8774 4326 8786 4378
rect 8838 4326 8850 4378
rect 8902 4326 8914 4378
rect 8966 4326 8978 4378
rect 9030 4326 14658 4378
rect 14710 4326 14722 4378
rect 14774 4326 14786 4378
rect 14838 4326 14850 4378
rect 14902 4326 14914 4378
rect 14966 4326 14978 4378
rect 15030 4326 20658 4378
rect 20710 4326 20722 4378
rect 20774 4326 20786 4378
rect 20838 4326 20850 4378
rect 20902 4326 20914 4378
rect 20966 4326 20978 4378
rect 21030 4326 26658 4378
rect 26710 4326 26722 4378
rect 26774 4326 26786 4378
rect 26838 4326 26850 4378
rect 26902 4326 26914 4378
rect 26966 4326 26978 4378
rect 27030 4326 32658 4378
rect 32710 4326 32722 4378
rect 32774 4326 32786 4378
rect 32838 4326 32850 4378
rect 32902 4326 32914 4378
rect 32966 4326 32978 4378
rect 33030 4326 38658 4378
rect 38710 4326 38722 4378
rect 38774 4326 38786 4378
rect 38838 4326 38850 4378
rect 38902 4326 38914 4378
rect 38966 4326 38978 4378
rect 39030 4326 43884 4378
rect 1104 4304 43884 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2685 4267 2743 4273
rect 2685 4264 2697 4267
rect 2464 4236 2697 4264
rect 2464 4224 2470 4236
rect 2685 4233 2697 4236
rect 2731 4264 2743 4267
rect 3142 4264 3148 4276
rect 2731 4236 3148 4264
rect 2731 4233 2743 4236
rect 2685 4227 2743 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 5166 4264 5172 4276
rect 3436 4236 5172 4264
rect 1486 4156 1492 4208
rect 1544 4156 1550 4208
rect 1854 4156 1860 4208
rect 1912 4156 1918 4208
rect 2222 4156 2228 4208
rect 2280 4156 2286 4208
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4196 2927 4199
rect 3050 4196 3056 4208
rect 2915 4168 3056 4196
rect 2915 4165 2927 4168
rect 2869 4159 2927 4165
rect 3050 4156 3056 4168
rect 3108 4196 3114 4208
rect 3436 4196 3464 4236
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5813 4267 5871 4273
rect 5813 4264 5825 4267
rect 5408 4236 5825 4264
rect 5408 4224 5414 4236
rect 5813 4233 5825 4236
rect 5859 4233 5871 4267
rect 5813 4227 5871 4233
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 6638 4264 6644 4276
rect 5960 4236 6644 4264
rect 5960 4224 5966 4236
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 8386 4224 8392 4276
rect 8444 4224 8450 4276
rect 13262 4264 13268 4276
rect 8588 4236 13268 4264
rect 3108 4168 3464 4196
rect 3108 4156 3114 4168
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4097 2559 4131
rect 2501 4091 2559 4097
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3326 4128 3332 4140
rect 3191 4100 3332 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 2516 4060 2544 4091
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 3436 4137 3464 4168
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 4890 4196 4896 4208
rect 4488 4168 4896 4196
rect 4488 4156 4494 4168
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 5000 4168 5212 4196
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4614 4128 4620 4140
rect 4295 4100 4620 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5000 4128 5028 4168
rect 4724 4100 5028 4128
rect 4724 4060 4752 4100
rect 5074 4088 5080 4140
rect 5132 4088 5138 4140
rect 5184 4128 5212 4168
rect 7282 4128 7288 4140
rect 5184 4100 7288 4128
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 8404 4128 8432 4224
rect 8588 4205 8616 4236
rect 13262 4224 13268 4236
rect 13320 4264 13326 4276
rect 13906 4264 13912 4276
rect 13320 4236 13912 4264
rect 13320 4224 13326 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 16666 4224 16672 4276
rect 16724 4264 16730 4276
rect 18601 4267 18659 4273
rect 18601 4264 18613 4267
rect 16724 4236 18613 4264
rect 16724 4224 16730 4236
rect 18601 4233 18613 4236
rect 18647 4233 18659 4267
rect 18601 4227 18659 4233
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 19058 4264 19064 4276
rect 18748 4236 19064 4264
rect 18748 4224 18754 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 19242 4224 19248 4276
rect 19300 4264 19306 4276
rect 21637 4267 21695 4273
rect 19300 4236 21588 4264
rect 19300 4224 19306 4236
rect 8573 4199 8631 4205
rect 8573 4165 8585 4199
rect 8619 4165 8631 4199
rect 8573 4159 8631 4165
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 21560 4196 21588 4236
rect 21637 4233 21649 4267
rect 21683 4264 21695 4267
rect 21818 4264 21824 4276
rect 21683 4236 21824 4264
rect 21683 4233 21695 4236
rect 21637 4227 21695 4233
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 22189 4267 22247 4273
rect 22189 4233 22201 4267
rect 22235 4264 22247 4267
rect 22370 4264 22376 4276
rect 22235 4236 22376 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 22557 4267 22615 4273
rect 22557 4264 22569 4267
rect 22520 4236 22569 4264
rect 22520 4224 22526 4236
rect 22557 4233 22569 4236
rect 22603 4233 22615 4267
rect 25130 4264 25136 4276
rect 22557 4227 22615 4233
rect 23124 4236 25136 4264
rect 23124 4196 23152 4236
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 25961 4267 26019 4273
rect 25961 4264 25973 4267
rect 25280 4236 25973 4264
rect 25280 4224 25286 4236
rect 25961 4233 25973 4236
rect 26007 4233 26019 4267
rect 25961 4227 26019 4233
rect 26145 4267 26203 4273
rect 26145 4233 26157 4267
rect 26191 4264 26203 4267
rect 26326 4264 26332 4276
rect 26191 4236 26332 4264
rect 26191 4233 26203 4236
rect 26145 4227 26203 4233
rect 26326 4224 26332 4236
rect 26384 4224 26390 4276
rect 27062 4224 27068 4276
rect 27120 4264 27126 4276
rect 27433 4267 27491 4273
rect 27433 4264 27445 4267
rect 27120 4236 27445 4264
rect 27120 4224 27126 4236
rect 27433 4233 27445 4236
rect 27479 4233 27491 4267
rect 27433 4227 27491 4233
rect 28166 4224 28172 4276
rect 28224 4264 28230 4276
rect 29273 4267 29331 4273
rect 28224 4236 28672 4264
rect 28224 4224 28230 4236
rect 10928 4168 12296 4196
rect 21560 4168 23152 4196
rect 10928 4156 10934 4168
rect 9766 4137 9772 4140
rect 9723 4131 9772 4137
rect 8404 4100 8984 4128
rect 8956 4072 8984 4100
rect 9723 4097 9735 4131
rect 9769 4097 9772 4131
rect 9723 4091 9772 4097
rect 9766 4088 9772 4091
rect 9824 4088 9830 4140
rect 9858 4088 9864 4140
rect 9916 4088 9922 4140
rect 10778 4088 10784 4140
rect 10836 4088 10842 4140
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 1544 4032 2544 4060
rect 4172 4032 4752 4060
rect 4801 4063 4859 4069
rect 1544 4020 1550 4032
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 3050 3992 3056 4004
rect 2087 3964 3056 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 4172 4001 4200 4032
rect 4801 4029 4813 4063
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3961 4215 3995
rect 4157 3955 4215 3961
rect 4430 3952 4436 4004
rect 4488 3952 4494 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1762 3924 1768 3936
rect 1627 3896 1768 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 1762 3884 1768 3896
rect 1820 3884 1826 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 2590 3924 2596 3936
rect 2363 3896 2596 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 2682 3884 2688 3936
rect 2740 3884 2746 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 3878 3924 3884 3936
rect 3007 3896 3884 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4816 3924 4844 4023
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 7742 4060 7748 4072
rect 5500 4032 7748 4060
rect 5500 4020 5506 4032
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8628 4032 8677 4060
rect 8628 4020 8634 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 8846 4020 8852 4072
rect 8904 4020 8910 4072
rect 8938 4020 8944 4072
rect 8996 4020 9002 4072
rect 9398 4060 9404 4072
rect 9232 4032 9404 4060
rect 9232 3992 9260 4032
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 10042 4060 10048 4072
rect 9631 4032 10048 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 11072 4060 11100 4091
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11790 4128 11796 4140
rect 11204 4100 11796 4128
rect 11204 4088 11210 4100
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 12268 4137 12296 4168
rect 25314 4156 25320 4208
rect 25372 4196 25378 4208
rect 25372 4168 25824 4196
rect 25372 4156 25378 4168
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4097 12311 4131
rect 12253 4091 12311 4097
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4128 12771 4131
rect 13078 4128 13084 4140
rect 12759 4100 13084 4128
rect 12759 4097 12771 4100
rect 12713 4091 12771 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13630 4088 13636 4140
rect 13688 4088 13694 4140
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 15654 4128 15660 4140
rect 14599 4100 15660 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 16850 4088 16856 4140
rect 16908 4088 16914 4140
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4128 18567 4131
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18555 4100 18797 4128
rect 18555 4097 18567 4100
rect 18509 4091 18567 4097
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19024 4100 20024 4128
rect 19024 4088 19030 4100
rect 10551 4032 11100 4060
rect 12897 4063 12955 4069
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 12897 4029 12909 4063
rect 12943 4060 12955 4063
rect 12943 4032 13222 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 7208 3964 9260 3992
rect 7208 3924 7236 3964
rect 9306 3952 9312 4004
rect 9364 3952 9370 4004
rect 12158 3992 12164 4004
rect 10520 3964 12164 3992
rect 4816 3896 7236 3924
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 10520 3924 10548 3964
rect 12158 3952 12164 3964
rect 12216 3952 12222 4004
rect 7331 3896 10548 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 10873 3927 10931 3933
rect 10873 3893 10885 3927
rect 10919 3924 10931 3927
rect 10962 3924 10968 3936
rect 10919 3896 10968 3924
rect 10919 3893 10931 3896
rect 10873 3887 10931 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 11882 3924 11888 3936
rect 11572 3896 11888 3924
rect 11572 3884 11578 3896
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 12032 3896 12081 3924
rect 12032 3884 12038 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 13194 3924 13222 4032
rect 13354 4020 13360 4072
rect 13412 4020 13418 4072
rect 13750 4063 13808 4069
rect 13750 4060 13762 4063
rect 13464 4032 13762 4060
rect 13262 3952 13268 4004
rect 13320 3992 13326 4004
rect 13464 3992 13492 4032
rect 13750 4029 13762 4032
rect 13796 4029 13808 4063
rect 13750 4023 13808 4029
rect 13906 4020 13912 4072
rect 13964 4020 13970 4072
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 14516 4032 16681 4060
rect 14516 4020 14522 4032
rect 16669 4029 16681 4032
rect 16715 4060 16727 4063
rect 16758 4060 16764 4072
rect 16715 4032 16764 4060
rect 16715 4029 16727 4032
rect 16669 4023 16727 4029
rect 16758 4020 16764 4032
rect 16816 4020 16822 4072
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17589 4063 17647 4069
rect 17589 4060 17601 4063
rect 17313 4023 17371 4029
rect 17420 4032 17601 4060
rect 13320 3964 13492 3992
rect 13320 3952 13326 3964
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 14792 3964 16436 3992
rect 14792 3952 14798 3964
rect 15562 3924 15568 3936
rect 13194 3896 15568 3924
rect 12069 3887 12127 3893
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 16408 3924 16436 3964
rect 16482 3952 16488 4004
rect 16540 3992 16546 4004
rect 17328 3992 17356 4023
rect 16540 3964 17356 3992
rect 16540 3952 16546 3964
rect 17420 3924 17448 4032
rect 17589 4029 17601 4032
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17678 4020 17684 4072
rect 17736 4069 17742 4072
rect 19996 4069 20024 4100
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4128 22983 4131
rect 23014 4128 23020 4140
rect 22971 4100 23020 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 24118 4088 24124 4140
rect 24176 4088 24182 4140
rect 25225 4131 25283 4137
rect 25225 4128 25237 4131
rect 25056 4100 25237 4128
rect 17736 4063 17764 4069
rect 17752 4029 17764 4063
rect 17736 4023 17764 4029
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4029 19855 4063
rect 19797 4023 19855 4029
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20530 4060 20536 4072
rect 20027 4032 20536 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 17736 4020 17742 4023
rect 18506 3924 18512 3936
rect 16408 3896 18512 3924
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 19812 3924 19840 4023
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 20714 4020 20720 4072
rect 20772 4020 20778 4072
rect 20898 4069 20904 4072
rect 20855 4063 20904 4069
rect 20855 4029 20867 4063
rect 20901 4029 20904 4063
rect 20855 4023 20904 4029
rect 20898 4020 20904 4023
rect 20956 4020 20962 4072
rect 20990 4020 20996 4072
rect 21048 4060 21054 4072
rect 21634 4060 21640 4072
rect 21048 4032 21640 4060
rect 21048 4020 21054 4032
rect 21634 4020 21640 4032
rect 21692 4020 21698 4072
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22186 4060 22192 4072
rect 22051 4032 22192 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22186 4020 22192 4032
rect 22244 4020 22250 4072
rect 22830 4020 22836 4072
rect 22888 4060 22894 4072
rect 23109 4063 23167 4069
rect 23109 4060 23121 4063
rect 22888 4032 23121 4060
rect 22888 4020 22894 4032
rect 23109 4029 23121 4032
rect 23155 4060 23167 4063
rect 23198 4060 23204 4072
rect 23155 4032 23204 4060
rect 23155 4029 23167 4032
rect 23109 4023 23167 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23569 4063 23627 4069
rect 23569 4029 23581 4063
rect 23615 4060 23627 4063
rect 23658 4060 23664 4072
rect 23615 4032 23664 4060
rect 23615 4029 23627 4032
rect 23569 4023 23627 4029
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 23842 4020 23848 4072
rect 23900 4020 23906 4072
rect 23983 4063 24041 4069
rect 23983 4029 23995 4063
rect 24029 4060 24041 4063
rect 24302 4060 24308 4072
rect 24029 4032 24308 4060
rect 24029 4029 24041 4032
rect 23983 4023 24041 4029
rect 24302 4020 24308 4032
rect 24360 4060 24366 4072
rect 24360 4032 24624 4060
rect 24360 4020 24366 4032
rect 20438 3952 20444 4004
rect 20496 3952 20502 4004
rect 21450 3952 21456 4004
rect 21508 3992 21514 4004
rect 23474 3992 23480 4004
rect 21508 3964 23480 3992
rect 21508 3952 21514 3964
rect 23474 3952 23480 3964
rect 23532 3952 23538 4004
rect 24596 3992 24624 4032
rect 24670 4020 24676 4072
rect 24728 4060 24734 4072
rect 24765 4063 24823 4069
rect 24765 4060 24777 4063
rect 24728 4032 24777 4060
rect 24728 4020 24734 4032
rect 24765 4029 24777 4032
rect 24811 4029 24823 4063
rect 24765 4023 24823 4029
rect 25056 3992 25084 4100
rect 25225 4097 25237 4100
rect 25271 4097 25283 4131
rect 25225 4091 25283 4097
rect 25406 4088 25412 4140
rect 25464 4088 25470 4140
rect 25796 4137 25824 4168
rect 25866 4156 25872 4208
rect 25924 4196 25930 4208
rect 25924 4168 27384 4196
rect 25924 4156 25930 4168
rect 25781 4131 25839 4137
rect 25781 4097 25793 4131
rect 25827 4097 25839 4131
rect 25958 4128 25964 4140
rect 25781 4091 25839 4097
rect 25884 4100 25964 4128
rect 25884 4069 25912 4100
rect 25958 4088 25964 4100
rect 26016 4088 26022 4140
rect 26050 4088 26056 4140
rect 26108 4128 26114 4140
rect 27356 4137 27384 4168
rect 28442 4156 28448 4208
rect 28500 4196 28506 4208
rect 28500 4168 28580 4196
rect 28500 4156 28506 4168
rect 26630 4131 26688 4137
rect 26630 4128 26642 4131
rect 26108 4100 26642 4128
rect 26108 4088 26114 4100
rect 26630 4097 26642 4100
rect 26676 4097 26688 4131
rect 26630 4091 26688 4097
rect 27341 4131 27399 4137
rect 27341 4097 27353 4131
rect 27387 4128 27399 4131
rect 27387 4100 27568 4128
rect 27387 4097 27399 4100
rect 27341 4091 27399 4097
rect 27540 4072 27568 4100
rect 28258 4088 28264 4140
rect 28316 4088 28322 4140
rect 28552 4137 28580 4168
rect 28537 4131 28595 4137
rect 28537 4097 28549 4131
rect 28583 4097 28595 4131
rect 28644 4128 28672 4236
rect 29273 4233 29285 4267
rect 29319 4264 29331 4267
rect 29454 4264 29460 4276
rect 29319 4236 29460 4264
rect 29319 4233 29331 4236
rect 29273 4227 29331 4233
rect 29454 4224 29460 4236
rect 29512 4224 29518 4276
rect 29822 4224 29828 4276
rect 29880 4264 29886 4276
rect 30469 4267 30527 4273
rect 30469 4264 30481 4267
rect 29880 4236 30481 4264
rect 29880 4224 29886 4236
rect 30469 4233 30481 4236
rect 30515 4233 30527 4267
rect 30469 4227 30527 4233
rect 31478 4224 31484 4276
rect 31536 4264 31542 4276
rect 32766 4264 32772 4276
rect 31536 4236 32772 4264
rect 31536 4224 31542 4236
rect 32766 4224 32772 4236
rect 32824 4224 32830 4276
rect 33134 4224 33140 4276
rect 33192 4264 33198 4276
rect 33192 4236 34192 4264
rect 33192 4224 33198 4236
rect 28718 4156 28724 4208
rect 28776 4196 28782 4208
rect 31662 4196 31668 4208
rect 28776 4168 31668 4196
rect 28776 4156 28782 4168
rect 31662 4156 31668 4168
rect 31720 4156 31726 4208
rect 30466 4128 30472 4140
rect 28644 4100 30472 4128
rect 28537 4091 28595 4097
rect 30466 4088 30472 4100
rect 30524 4088 30530 4140
rect 30650 4088 30656 4140
rect 30708 4088 30714 4140
rect 31018 4088 31024 4140
rect 31076 4128 31082 4140
rect 32214 4128 32220 4140
rect 31076 4100 32220 4128
rect 31076 4088 31082 4100
rect 32214 4088 32220 4100
rect 32272 4128 32278 4140
rect 32401 4131 32459 4137
rect 32401 4128 32413 4131
rect 32272 4100 32413 4128
rect 32272 4088 32278 4100
rect 32401 4097 32413 4100
rect 32447 4097 32459 4131
rect 32401 4091 32459 4097
rect 32582 4088 32588 4140
rect 32640 4088 32646 4140
rect 33410 4088 33416 4140
rect 33468 4137 33474 4140
rect 33468 4131 33496 4137
rect 33484 4097 33496 4131
rect 34164 4128 34192 4236
rect 34238 4224 34244 4276
rect 34296 4224 34302 4276
rect 34514 4224 34520 4276
rect 34572 4264 34578 4276
rect 39758 4264 39764 4276
rect 34572 4236 39764 4264
rect 34572 4224 34578 4236
rect 39758 4224 39764 4236
rect 39816 4224 39822 4276
rect 36170 4156 36176 4208
rect 36228 4156 36234 4208
rect 39482 4156 39488 4208
rect 39540 4156 39546 4208
rect 39574 4156 39580 4208
rect 39632 4196 39638 4208
rect 42150 4196 42156 4208
rect 39632 4168 42156 4196
rect 39632 4156 39638 4168
rect 42150 4156 42156 4168
rect 42208 4156 42214 4208
rect 34164 4100 34652 4128
rect 33468 4091 33496 4097
rect 33468 4088 33474 4091
rect 25317 4063 25375 4069
rect 25317 4029 25329 4063
rect 25363 4060 25375 4063
rect 25869 4063 25927 4069
rect 25363 4032 25824 4060
rect 25363 4029 25375 4032
rect 25317 4023 25375 4029
rect 24596 3964 25084 3992
rect 25590 3952 25596 4004
rect 25648 3952 25654 4004
rect 25796 3992 25824 4032
rect 25869 4029 25881 4063
rect 25915 4029 25927 4063
rect 25869 4023 25927 4029
rect 26237 4063 26295 4069
rect 26237 4029 26249 4063
rect 26283 4029 26295 4063
rect 26237 4023 26295 4029
rect 26252 3992 26280 4023
rect 27522 4020 27528 4072
rect 27580 4020 27586 4072
rect 27617 4063 27675 4069
rect 27617 4029 27629 4063
rect 27663 4060 27675 4063
rect 27798 4060 27804 4072
rect 27663 4032 27804 4060
rect 27663 4029 27675 4032
rect 27617 4023 27675 4029
rect 27798 4020 27804 4032
rect 27856 4020 27862 4072
rect 28966 4032 32996 4060
rect 25796 3964 26280 3992
rect 26786 3952 26792 4004
rect 26844 3992 26850 4004
rect 27982 3992 27988 4004
rect 26844 3964 27988 3992
rect 26844 3952 26850 3964
rect 27982 3952 27988 3964
rect 28040 3952 28046 4004
rect 28966 3992 28994 4032
rect 28920 3964 28994 3992
rect 23014 3924 23020 3936
rect 19812 3896 23020 3924
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 26234 3884 26240 3936
rect 26292 3924 26298 3936
rect 26559 3927 26617 3933
rect 26559 3924 26571 3927
rect 26292 3896 26571 3924
rect 26292 3884 26298 3896
rect 26559 3893 26571 3896
rect 26605 3893 26617 3927
rect 26559 3887 26617 3893
rect 26973 3927 27031 3933
rect 26973 3893 26985 3927
rect 27019 3924 27031 3927
rect 27338 3924 27344 3936
rect 27019 3896 27344 3924
rect 27019 3893 27031 3896
rect 26973 3887 27031 3893
rect 27338 3884 27344 3896
rect 27396 3884 27402 3936
rect 27430 3884 27436 3936
rect 27488 3924 27494 3936
rect 28920 3924 28948 3964
rect 32214 3952 32220 4004
rect 32272 3992 32278 4004
rect 32582 3992 32588 4004
rect 32272 3964 32588 3992
rect 32272 3952 32278 3964
rect 32582 3952 32588 3964
rect 32640 3952 32646 4004
rect 32968 3992 32996 4032
rect 33042 4020 33048 4072
rect 33100 4020 33106 4072
rect 33134 4020 33140 4072
rect 33192 4060 33198 4072
rect 33321 4063 33379 4069
rect 33321 4060 33333 4063
rect 33192 4032 33333 4060
rect 33192 4020 33198 4032
rect 33321 4029 33333 4032
rect 33367 4029 33379 4063
rect 33321 4023 33379 4029
rect 33594 4020 33600 4072
rect 33652 4020 33658 4072
rect 34330 4020 34336 4072
rect 34388 4020 34394 4072
rect 34517 4063 34575 4069
rect 34517 4029 34529 4063
rect 34563 4029 34575 4063
rect 34624 4060 34652 4100
rect 35342 4088 35348 4140
rect 35400 4137 35406 4140
rect 35400 4131 35428 4137
rect 35416 4097 35428 4131
rect 36188 4128 36216 4156
rect 36909 4131 36967 4137
rect 36909 4128 36921 4131
rect 36188 4100 36921 4128
rect 35400 4091 35428 4097
rect 36909 4097 36921 4100
rect 36955 4128 36967 4131
rect 37182 4128 37188 4140
rect 36955 4100 37188 4128
rect 36955 4097 36967 4100
rect 36909 4091 36967 4097
rect 35400 4088 35406 4091
rect 37182 4088 37188 4100
rect 37240 4088 37246 4140
rect 38381 4131 38439 4137
rect 38381 4097 38393 4131
rect 38427 4128 38439 4131
rect 38473 4131 38531 4137
rect 38473 4128 38485 4131
rect 38427 4100 38485 4128
rect 38427 4097 38439 4100
rect 38381 4091 38439 4097
rect 38473 4097 38485 4100
rect 38519 4097 38531 4131
rect 38473 4091 38531 4097
rect 38746 4088 38752 4140
rect 38804 4128 38810 4140
rect 39025 4131 39083 4137
rect 39025 4128 39037 4131
rect 38804 4100 39037 4128
rect 38804 4088 38810 4100
rect 39025 4097 39037 4100
rect 39071 4128 39083 4131
rect 39500 4128 39528 4156
rect 39071 4100 39528 4128
rect 39071 4097 39083 4100
rect 39025 4091 39083 4097
rect 42058 4088 42064 4140
rect 42116 4128 42122 4140
rect 42245 4131 42303 4137
rect 42245 4128 42257 4131
rect 42116 4100 42257 4128
rect 42116 4088 42122 4100
rect 42245 4097 42257 4100
rect 42291 4097 42303 4131
rect 42245 4091 42303 4097
rect 42610 4088 42616 4140
rect 42668 4088 42674 4140
rect 42889 4131 42947 4137
rect 42889 4097 42901 4131
rect 42935 4097 42947 4131
rect 42889 4091 42947 4097
rect 35253 4063 35311 4069
rect 35253 4060 35265 4063
rect 34624 4032 35265 4060
rect 34517 4023 34575 4029
rect 35253 4029 35265 4032
rect 35299 4029 35311 4063
rect 35253 4023 35311 4029
rect 33152 3992 33180 4020
rect 32968 3964 33180 3992
rect 27488 3896 28948 3924
rect 27488 3884 27494 3896
rect 30466 3884 30472 3936
rect 30524 3924 30530 3936
rect 34532 3924 34560 4023
rect 35526 4020 35532 4072
rect 35584 4020 35590 4072
rect 36078 4020 36084 4072
rect 36136 4060 36142 4072
rect 36173 4063 36231 4069
rect 36173 4060 36185 4063
rect 36136 4032 36185 4060
rect 36136 4020 36142 4032
rect 36173 4029 36185 4032
rect 36219 4029 36231 4063
rect 36173 4023 36231 4029
rect 36262 4020 36268 4072
rect 36320 4060 36326 4072
rect 39206 4060 39212 4072
rect 36320 4032 39212 4060
rect 36320 4020 36326 4032
rect 39206 4020 39212 4032
rect 39264 4020 39270 4072
rect 39482 4020 39488 4072
rect 39540 4060 39546 4072
rect 42904 4060 42932 4091
rect 42978 4088 42984 4140
rect 43036 4128 43042 4140
rect 43257 4131 43315 4137
rect 43257 4128 43269 4131
rect 43036 4100 43269 4128
rect 43036 4088 43042 4100
rect 43257 4097 43269 4100
rect 43303 4097 43315 4131
rect 43257 4091 43315 4097
rect 39540 4032 42932 4060
rect 39540 4020 39546 4032
rect 34974 3952 34980 4004
rect 35032 3952 35038 4004
rect 36722 3952 36728 4004
rect 36780 3952 36786 4004
rect 38841 3995 38899 4001
rect 38841 3992 38853 3995
rect 36832 3964 38853 3992
rect 30524 3896 34560 3924
rect 30524 3884 30530 3896
rect 34790 3884 34796 3936
rect 34848 3924 34854 3936
rect 36832 3924 36860 3964
rect 38841 3961 38853 3964
rect 38887 3961 38899 3995
rect 38841 3955 38899 3961
rect 41966 3952 41972 4004
rect 42024 3992 42030 4004
rect 42061 3995 42119 4001
rect 42061 3992 42073 3995
rect 42024 3964 42073 3992
rect 42024 3952 42030 3964
rect 42061 3961 42073 3964
rect 42107 3961 42119 3995
rect 42061 3955 42119 3961
rect 43438 3952 43444 4004
rect 43496 3952 43502 4004
rect 34848 3896 36860 3924
rect 34848 3884 34854 3896
rect 37826 3884 37832 3936
rect 37884 3924 37890 3936
rect 38289 3927 38347 3933
rect 38289 3924 38301 3927
rect 37884 3896 38301 3924
rect 37884 3884 37890 3896
rect 38289 3893 38301 3896
rect 38335 3893 38347 3927
rect 38289 3887 38347 3893
rect 38657 3927 38715 3933
rect 38657 3893 38669 3927
rect 38703 3924 38715 3927
rect 38746 3924 38752 3936
rect 38703 3896 38752 3924
rect 38703 3893 38715 3896
rect 38657 3887 38715 3893
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 41782 3884 41788 3936
rect 41840 3924 41846 3936
rect 42429 3927 42487 3933
rect 42429 3924 42441 3927
rect 41840 3896 42441 3924
rect 41840 3884 41846 3896
rect 42429 3893 42441 3896
rect 42475 3893 42487 3927
rect 42429 3887 42487 3893
rect 43070 3884 43076 3936
rect 43128 3884 43134 3936
rect 1104 3834 43884 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13918 3834
rect 13970 3782 13982 3834
rect 14034 3782 14046 3834
rect 14098 3782 14110 3834
rect 14162 3782 14174 3834
rect 14226 3782 14238 3834
rect 14290 3782 19918 3834
rect 19970 3782 19982 3834
rect 20034 3782 20046 3834
rect 20098 3782 20110 3834
rect 20162 3782 20174 3834
rect 20226 3782 20238 3834
rect 20290 3782 25918 3834
rect 25970 3782 25982 3834
rect 26034 3782 26046 3834
rect 26098 3782 26110 3834
rect 26162 3782 26174 3834
rect 26226 3782 26238 3834
rect 26290 3782 31918 3834
rect 31970 3782 31982 3834
rect 32034 3782 32046 3834
rect 32098 3782 32110 3834
rect 32162 3782 32174 3834
rect 32226 3782 32238 3834
rect 32290 3782 37918 3834
rect 37970 3782 37982 3834
rect 38034 3782 38046 3834
rect 38098 3782 38110 3834
rect 38162 3782 38174 3834
rect 38226 3782 38238 3834
rect 38290 3782 43884 3834
rect 1104 3760 43884 3782
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 2958 3720 2964 3732
rect 1820 3692 2964 3720
rect 1820 3680 1826 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 6638 3720 6644 3732
rect 3108 3692 6644 3720
rect 3108 3680 3114 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7524 3692 7849 3720
rect 7524 3680 7530 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 9048 3692 9674 3720
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3652 2835 3655
rect 3694 3652 3700 3664
rect 2823 3624 3700 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 4062 3612 4068 3664
rect 4120 3652 4126 3664
rect 4430 3652 4436 3664
rect 4120 3624 4436 3652
rect 4120 3612 4126 3624
rect 4430 3612 4436 3624
rect 4488 3612 4494 3664
rect 5813 3655 5871 3661
rect 5813 3621 5825 3655
rect 5859 3621 5871 3655
rect 9048 3652 9076 3692
rect 5813 3615 5871 3621
rect 7024 3624 7512 3652
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 4614 3584 4620 3596
rect 2455 3556 4620 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 4801 3587 4859 3593
rect 4801 3584 4813 3587
rect 4764 3556 4813 3584
rect 4764 3544 4770 3556
rect 4801 3553 4813 3556
rect 4847 3553 4859 3587
rect 5828 3584 5856 3615
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 5828 3556 6561 3584
rect 4801 3547 4859 3553
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 6708 3587 6766 3593
rect 6708 3553 6720 3587
rect 6754 3584 6766 3587
rect 7024 3584 7052 3624
rect 6754 3556 7052 3584
rect 7101 3587 7159 3593
rect 6754 3553 6766 3556
rect 6708 3547 6766 3553
rect 7101 3553 7113 3587
rect 7147 3584 7159 3587
rect 7374 3584 7380 3596
rect 7147 3556 7380 3584
rect 7147 3553 7159 3556
rect 7101 3547 7159 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 1489 3519 1547 3525
rect 1489 3516 1501 3519
rect 1452 3488 1501 3516
rect 1452 3476 1458 3488
rect 1489 3485 1501 3488
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2740 3488 3249 3516
rect 2740 3476 2746 3488
rect 3237 3485 3249 3488
rect 3283 3516 3295 3519
rect 5074 3516 5080 3528
rect 3283 3488 5080 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 7484 3516 7512 3624
rect 7576 3624 9076 3652
rect 9646 3652 9674 3692
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9916 3692 9965 3720
rect 9916 3680 9922 3692
rect 9953 3689 9965 3692
rect 9999 3689 10011 3723
rect 9953 3683 10011 3689
rect 10336 3692 11468 3720
rect 10336 3652 10364 3692
rect 9646 3624 10364 3652
rect 7576 3593 7604 3624
rect 10410 3612 10416 3664
rect 10468 3652 10474 3664
rect 11440 3652 11468 3692
rect 11514 3680 11520 3732
rect 11572 3680 11578 3732
rect 11716 3692 12756 3720
rect 11716 3652 11744 3692
rect 10468 3624 10548 3652
rect 11440 3624 11744 3652
rect 12728 3652 12756 3692
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 12860 3692 13369 3720
rect 12860 3680 12866 3692
rect 13357 3689 13369 3692
rect 13403 3720 13415 3723
rect 13722 3720 13728 3732
rect 13403 3692 13728 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13872 3692 14105 3720
rect 13872 3680 13878 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 16485 3723 16543 3729
rect 14093 3683 14151 3689
rect 15028 3692 16436 3720
rect 15028 3652 15056 3692
rect 12728 3624 15056 3652
rect 10468 3612 10474 3624
rect 7561 3587 7619 3593
rect 7561 3553 7573 3587
rect 7607 3553 7619 3587
rect 7834 3584 7840 3596
rect 7561 3547 7619 3553
rect 7668 3556 7840 3584
rect 7668 3516 7696 3556
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8570 3584 8576 3596
rect 8352 3556 8576 3584
rect 8352 3544 8358 3556
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8938 3544 8944 3596
rect 8996 3544 9002 3596
rect 9766 3584 9772 3596
rect 9508 3556 9772 3584
rect 7484 3488 7696 3516
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 7926 3516 7932 3528
rect 7800 3488 7932 3516
rect 7800 3476 7806 3488
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 8021 3479 8079 3485
rect 8588 3488 9229 3516
rect 1854 3408 1860 3460
rect 1912 3408 1918 3460
rect 2222 3408 2228 3460
rect 2280 3408 2286 3460
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 2593 3451 2651 3457
rect 2593 3448 2605 3451
rect 2464 3420 2605 3448
rect 2464 3408 2470 3420
rect 2593 3417 2605 3420
rect 2639 3417 2651 3451
rect 2593 3411 2651 3417
rect 3421 3451 3479 3457
rect 3421 3417 3433 3451
rect 3467 3448 3479 3451
rect 3970 3448 3976 3460
rect 3467 3420 3976 3448
rect 3467 3417 3479 3420
rect 3421 3411 3479 3417
rect 3970 3408 3976 3420
rect 4028 3408 4034 3460
rect 8036 3448 8064 3479
rect 8588 3457 8616 3488
rect 9217 3485 9229 3488
rect 9263 3516 9275 3519
rect 9508 3516 9536 3556
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10520 3593 10548 3624
rect 15102 3612 15108 3664
rect 15160 3652 15166 3664
rect 16408 3652 16436 3692
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 17862 3720 17868 3732
rect 16531 3692 17868 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18012 3692 18276 3720
rect 18012 3680 18018 3692
rect 17494 3652 17500 3664
rect 15160 3624 15516 3652
rect 16408 3624 17500 3652
rect 15160 3612 15166 3624
rect 15488 3596 15516 3624
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 18248 3652 18276 3692
rect 18322 3680 18328 3732
rect 18380 3720 18386 3732
rect 18380 3692 20576 3720
rect 18380 3680 18386 3692
rect 19242 3652 19248 3664
rect 18248 3624 19248 3652
rect 19242 3612 19248 3624
rect 19300 3612 19306 3664
rect 19334 3612 19340 3664
rect 19392 3612 19398 3664
rect 10505 3587 10563 3593
rect 10244 3556 10456 3584
rect 10244 3516 10272 3556
rect 9263 3488 9536 3516
rect 9600 3488 10272 3516
rect 10321 3519 10379 3525
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 7760 3420 8064 3448
rect 8573 3451 8631 3457
rect 1578 3340 1584 3392
rect 1636 3340 1642 3392
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 1949 3383 2007 3389
rect 1949 3380 1961 3383
rect 1728 3352 1961 3380
rect 1728 3340 1734 3352
rect 1949 3349 1961 3352
rect 1995 3349 2007 3383
rect 1949 3343 2007 3349
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 7760 3380 7788 3420
rect 8573 3417 8585 3451
rect 8619 3417 8631 3451
rect 8573 3411 8631 3417
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 9490 3448 9496 3460
rect 8803 3420 9496 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 5951 3352 7788 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8588 3380 8616 3411
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 8076 3352 8616 3380
rect 8076 3340 8082 3352
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9600 3380 9628 3488
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 8904 3352 9628 3380
rect 8904 3340 8910 3352
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 9732 3352 10149 3380
rect 9732 3340 9738 3352
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 10336 3380 10364 3479
rect 10428 3448 10456 3556
rect 10505 3553 10517 3587
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 11606 3544 11612 3596
rect 11664 3544 11670 3596
rect 12268 3556 15240 3584
rect 10778 3476 10784 3528
rect 10836 3476 10842 3528
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 10928 3488 11897 3516
rect 10928 3476 10934 3488
rect 11885 3485 11897 3488
rect 11931 3516 11943 3519
rect 12268 3516 12296 3556
rect 13173 3519 13231 3525
rect 11931 3488 12296 3516
rect 12728 3488 13124 3516
rect 11931 3485 11943 3488
rect 11885 3479 11943 3485
rect 12728 3448 12756 3488
rect 10428 3420 12756 3448
rect 12805 3451 12863 3457
rect 12805 3417 12817 3451
rect 12851 3417 12863 3451
rect 13096 3448 13124 3488
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 13262 3516 13268 3528
rect 13219 3488 13268 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13688 3488 13737 3516
rect 13688 3476 13694 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 14642 3476 14648 3528
rect 14700 3476 14706 3528
rect 14458 3448 14464 3460
rect 13096 3420 14464 3448
rect 12805 3411 12863 3417
rect 11330 3380 11336 3392
rect 10336 3352 11336 3380
rect 10137 3343 10195 3349
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 12526 3340 12532 3392
rect 12584 3380 12590 3392
rect 12621 3383 12679 3389
rect 12621 3380 12633 3383
rect 12584 3352 12633 3380
rect 12584 3340 12590 3352
rect 12621 3349 12633 3352
rect 12667 3349 12679 3383
rect 12621 3343 12679 3349
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 12820 3380 12848 3411
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 14829 3451 14887 3457
rect 14829 3417 14841 3451
rect 14875 3448 14887 3451
rect 15102 3448 15108 3460
rect 14875 3420 15108 3448
rect 14875 3417 14887 3420
rect 14829 3411 14887 3417
rect 15102 3408 15108 3420
rect 15160 3408 15166 3460
rect 15212 3448 15240 3556
rect 15470 3544 15476 3596
rect 15528 3544 15534 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 19484 3556 19625 3584
rect 19484 3544 19490 3556
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 20548 3584 20576 3692
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 24302 3720 24308 3732
rect 20956 3692 24308 3720
rect 20956 3680 20962 3692
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25188 3692 26280 3720
rect 25188 3680 25194 3692
rect 20625 3655 20683 3661
rect 20625 3621 20637 3655
rect 20671 3652 20683 3655
rect 20990 3652 20996 3664
rect 20671 3624 20996 3652
rect 20671 3621 20683 3624
rect 20625 3615 20683 3621
rect 20990 3612 20996 3624
rect 21048 3612 21054 3664
rect 21836 3624 22508 3652
rect 21358 3584 21364 3596
rect 20548 3556 21364 3584
rect 19613 3547 19671 3553
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 21836 3528 21864 3624
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 15712 3488 15761 3516
rect 15712 3476 15718 3488
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17494 3516 17500 3528
rect 17276 3488 17500 3516
rect 17276 3476 17282 3488
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17678 3476 17684 3528
rect 17736 3516 17742 3528
rect 17773 3519 17831 3525
rect 17773 3516 17785 3519
rect 17736 3488 17785 3516
rect 17736 3476 17742 3488
rect 17773 3485 17785 3488
rect 17819 3485 17831 3519
rect 17773 3479 17831 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 19334 3516 19340 3528
rect 18196 3488 19340 3516
rect 18196 3476 18202 3488
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19518 3476 19524 3528
rect 19576 3476 19582 3528
rect 19886 3476 19892 3528
rect 19944 3516 19950 3528
rect 20530 3516 20536 3528
rect 19944 3488 20536 3516
rect 19944 3476 19950 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 21818 3476 21824 3528
rect 21876 3476 21882 3528
rect 19794 3448 19800 3460
rect 15212 3420 19800 3448
rect 19794 3408 19800 3420
rect 19852 3408 19858 3460
rect 20898 3408 20904 3460
rect 20956 3448 20962 3460
rect 21174 3448 21180 3460
rect 20956 3420 21180 3448
rect 20956 3408 20962 3420
rect 21174 3408 21180 3420
rect 21232 3448 21238 3460
rect 22480 3448 22508 3624
rect 23474 3612 23480 3664
rect 23532 3652 23538 3664
rect 25038 3652 25044 3664
rect 23532 3624 25044 3652
rect 23532 3612 23538 3624
rect 25038 3612 25044 3624
rect 25096 3652 25102 3664
rect 26252 3652 26280 3692
rect 26326 3680 26332 3732
rect 26384 3720 26390 3732
rect 26384 3692 27568 3720
rect 26384 3680 26390 3692
rect 25096 3624 25912 3652
rect 26252 3624 26464 3652
rect 25096 3612 25102 3624
rect 25884 3596 25912 3624
rect 22646 3544 22652 3596
rect 22704 3544 22710 3596
rect 25682 3544 25688 3596
rect 25740 3544 25746 3596
rect 25866 3544 25872 3596
rect 25924 3544 25930 3596
rect 26326 3544 26332 3596
rect 26384 3544 26390 3596
rect 26436 3584 26464 3624
rect 26602 3584 26608 3596
rect 26436 3556 26608 3584
rect 26602 3544 26608 3556
rect 26660 3544 26666 3596
rect 26786 3593 26792 3596
rect 26743 3587 26792 3593
rect 26743 3553 26755 3587
rect 26789 3553 26792 3587
rect 26743 3547 26792 3553
rect 26786 3544 26792 3547
rect 26844 3544 26850 3596
rect 26878 3544 26884 3596
rect 26936 3544 26942 3596
rect 27062 3544 27068 3596
rect 27120 3584 27126 3596
rect 27120 3556 27476 3584
rect 27120 3544 27126 3556
rect 22925 3519 22983 3525
rect 22925 3485 22937 3519
rect 22971 3485 22983 3519
rect 23842 3516 23848 3528
rect 22925 3479 22983 3485
rect 23584 3488 23848 3516
rect 22940 3448 22968 3479
rect 21232 3420 22416 3448
rect 22480 3420 22968 3448
rect 21232 3408 21238 3420
rect 12768 3352 12848 3380
rect 12897 3383 12955 3389
rect 12768 3340 12774 3352
rect 12897 3349 12909 3383
rect 12943 3380 12955 3383
rect 12986 3380 12992 3392
rect 12943 3352 12992 3380
rect 12943 3349 12955 3352
rect 12897 3343 12955 3349
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 13354 3340 13360 3392
rect 13412 3340 13418 3392
rect 13538 3340 13544 3392
rect 13596 3340 13602 3392
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 13998 3380 14004 3392
rect 13688 3352 14004 3380
rect 13688 3340 13694 3352
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 15654 3380 15660 3392
rect 14240 3352 15660 3380
rect 14240 3340 14246 3352
rect 15654 3340 15660 3352
rect 15712 3380 15718 3392
rect 16758 3380 16764 3392
rect 15712 3352 16764 3380
rect 15712 3340 15718 3352
rect 16758 3340 16764 3352
rect 16816 3380 16822 3392
rect 17862 3380 17868 3392
rect 16816 3352 17868 3380
rect 16816 3340 16822 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 18196 3352 18521 3380
rect 18196 3340 18202 3352
rect 18509 3349 18521 3352
rect 18555 3349 18567 3383
rect 18509 3343 18567 3349
rect 20438 3340 20444 3392
rect 20496 3380 20502 3392
rect 21450 3380 21456 3392
rect 20496 3352 21456 3380
rect 20496 3340 20502 3352
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 22002 3340 22008 3392
rect 22060 3340 22066 3392
rect 22388 3380 22416 3420
rect 23584 3380 23612 3488
rect 23842 3476 23848 3488
rect 23900 3476 23906 3528
rect 24949 3519 25007 3525
rect 24949 3485 24961 3519
rect 24995 3516 25007 3519
rect 25222 3516 25228 3528
rect 24995 3488 25228 3516
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 27448 3448 27476 3556
rect 27540 3516 27568 3692
rect 28258 3680 28264 3732
rect 28316 3720 28322 3732
rect 29273 3723 29331 3729
rect 28316 3692 28994 3720
rect 28316 3680 28322 3692
rect 28258 3544 28264 3596
rect 28316 3544 28322 3596
rect 28966 3584 28994 3692
rect 29273 3689 29285 3723
rect 29319 3720 29331 3723
rect 29319 3692 30236 3720
rect 29319 3689 29331 3692
rect 29273 3683 29331 3689
rect 30208 3652 30236 3692
rect 30558 3680 30564 3732
rect 30616 3680 30622 3732
rect 31110 3680 31116 3732
rect 31168 3720 31174 3732
rect 32585 3723 32643 3729
rect 31168 3692 32536 3720
rect 31168 3680 31174 3692
rect 30742 3652 30748 3664
rect 30208 3624 30748 3652
rect 30742 3612 30748 3624
rect 30800 3612 30806 3664
rect 29549 3587 29607 3593
rect 29549 3584 29561 3587
rect 28966 3556 29561 3584
rect 29549 3553 29561 3556
rect 29595 3553 29607 3587
rect 29549 3547 29607 3553
rect 31570 3544 31576 3596
rect 31628 3544 31634 3596
rect 32508 3584 32536 3692
rect 32585 3689 32597 3723
rect 32631 3720 32643 3723
rect 33594 3720 33600 3732
rect 32631 3692 33600 3720
rect 32631 3689 32643 3692
rect 32585 3683 32643 3689
rect 33594 3680 33600 3692
rect 33652 3680 33658 3732
rect 34974 3680 34980 3732
rect 35032 3720 35038 3732
rect 35253 3723 35311 3729
rect 35253 3720 35265 3723
rect 35032 3692 35265 3720
rect 35032 3680 35038 3692
rect 35253 3689 35265 3692
rect 35299 3689 35311 3723
rect 35253 3683 35311 3689
rect 35526 3680 35532 3732
rect 35584 3720 35590 3732
rect 38289 3723 38347 3729
rect 38289 3720 38301 3723
rect 35584 3692 38301 3720
rect 35584 3680 35590 3692
rect 38289 3689 38301 3692
rect 38335 3689 38347 3723
rect 38289 3683 38347 3689
rect 41506 3680 41512 3732
rect 41564 3720 41570 3732
rect 42061 3723 42119 3729
rect 42061 3720 42073 3723
rect 41564 3692 42073 3720
rect 41564 3680 41570 3692
rect 42061 3689 42073 3692
rect 42107 3689 42119 3723
rect 42061 3683 42119 3689
rect 38470 3612 38476 3664
rect 38528 3652 38534 3664
rect 38746 3652 38752 3664
rect 38528 3624 38752 3652
rect 38528 3612 38534 3624
rect 38746 3612 38752 3624
rect 38804 3612 38810 3664
rect 41414 3612 41420 3664
rect 41472 3652 41478 3664
rect 42613 3655 42671 3661
rect 42613 3652 42625 3655
rect 41472 3624 42625 3652
rect 41472 3612 41478 3624
rect 42613 3621 42625 3624
rect 42659 3621 42671 3655
rect 42613 3615 42671 3621
rect 43438 3612 43444 3664
rect 43496 3612 43502 3664
rect 32677 3587 32735 3593
rect 32677 3584 32689 3587
rect 32508 3556 32689 3584
rect 32677 3553 32689 3556
rect 32723 3553 32735 3587
rect 35066 3584 35072 3596
rect 32677 3547 32735 3553
rect 34808 3556 35072 3584
rect 28442 3516 28448 3528
rect 27540 3488 28448 3516
rect 28442 3476 28448 3488
rect 28500 3516 28506 3528
rect 28537 3519 28595 3525
rect 28537 3516 28549 3519
rect 28500 3488 28549 3516
rect 28500 3476 28506 3488
rect 28537 3485 28549 3488
rect 28583 3485 28595 3519
rect 28537 3479 28595 3485
rect 28626 3476 28632 3528
rect 28684 3516 28690 3528
rect 29454 3516 29460 3528
rect 28684 3488 29460 3516
rect 28684 3476 28690 3488
rect 29454 3476 29460 3488
rect 29512 3476 29518 3528
rect 29825 3519 29883 3525
rect 29825 3485 29837 3519
rect 29871 3516 29883 3519
rect 29871 3485 29893 3516
rect 29825 3479 29893 3485
rect 29730 3448 29736 3460
rect 23676 3420 25912 3448
rect 27448 3420 29736 3448
rect 23676 3389 23704 3420
rect 22388 3352 23612 3380
rect 23661 3383 23719 3389
rect 23661 3349 23673 3383
rect 23707 3349 23719 3383
rect 23661 3343 23719 3349
rect 25038 3340 25044 3392
rect 25096 3380 25102 3392
rect 25133 3383 25191 3389
rect 25133 3380 25145 3383
rect 25096 3352 25145 3380
rect 25096 3340 25102 3352
rect 25133 3349 25145 3352
rect 25179 3349 25191 3383
rect 25884 3380 25912 3420
rect 29730 3408 29736 3420
rect 29788 3408 29794 3460
rect 29865 3448 29893 3479
rect 31846 3476 31852 3528
rect 31904 3476 31910 3528
rect 32950 3476 32956 3528
rect 33008 3476 33014 3528
rect 34808 3516 34836 3556
rect 35066 3544 35072 3556
rect 35124 3584 35130 3596
rect 35124 3556 35664 3584
rect 35124 3544 35130 3556
rect 33060 3488 34836 3516
rect 30098 3448 30104 3460
rect 29865 3420 30104 3448
rect 30098 3408 30104 3420
rect 30156 3408 30162 3460
rect 32306 3448 32312 3460
rect 30392 3420 32312 3448
rect 27154 3380 27160 3392
rect 25884 3352 27160 3380
rect 25133 3343 25191 3349
rect 27154 3340 27160 3352
rect 27212 3340 27218 3392
rect 27338 3340 27344 3392
rect 27396 3380 27402 3392
rect 27525 3383 27583 3389
rect 27525 3380 27537 3383
rect 27396 3352 27537 3380
rect 27396 3340 27402 3352
rect 27525 3349 27537 3352
rect 27571 3349 27583 3383
rect 27525 3343 27583 3349
rect 28534 3340 28540 3392
rect 28592 3380 28598 3392
rect 30392 3380 30420 3420
rect 32306 3408 32312 3420
rect 32364 3408 32370 3460
rect 33060 3448 33088 3488
rect 34882 3476 34888 3528
rect 34940 3476 34946 3528
rect 32968 3420 33088 3448
rect 28592 3352 30420 3380
rect 28592 3340 28598 3352
rect 30466 3340 30472 3392
rect 30524 3380 30530 3392
rect 32968 3380 32996 3420
rect 33410 3408 33416 3460
rect 33468 3448 33474 3460
rect 33870 3448 33876 3460
rect 33468 3420 33876 3448
rect 33468 3408 33474 3420
rect 33870 3408 33876 3420
rect 33928 3408 33934 3460
rect 35636 3448 35664 3556
rect 36262 3544 36268 3596
rect 36320 3584 36326 3596
rect 37277 3587 37335 3593
rect 37277 3584 37289 3587
rect 36320 3556 37289 3584
rect 36320 3544 36326 3556
rect 37277 3553 37289 3556
rect 37323 3553 37335 3587
rect 37277 3547 37335 3553
rect 37844 3556 42932 3584
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 35989 3519 36047 3525
rect 35989 3516 36001 3519
rect 35952 3488 36001 3516
rect 35952 3476 35958 3488
rect 35989 3485 36001 3488
rect 36035 3485 36047 3519
rect 35989 3479 36047 3485
rect 36538 3476 36544 3528
rect 36596 3516 36602 3528
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 36596 3488 37565 3516
rect 36596 3476 36602 3488
rect 37553 3485 37565 3488
rect 37599 3485 37611 3519
rect 37553 3479 37611 3485
rect 37642 3476 37648 3528
rect 37700 3516 37706 3528
rect 37844 3516 37872 3556
rect 37700 3488 37872 3516
rect 37700 3476 37706 3488
rect 38286 3476 38292 3528
rect 38344 3516 38350 3528
rect 38381 3519 38439 3525
rect 38381 3516 38393 3519
rect 38344 3488 38393 3516
rect 38344 3476 38350 3488
rect 38381 3485 38393 3488
rect 38427 3485 38439 3519
rect 39117 3519 39175 3525
rect 38381 3479 38439 3485
rect 38672 3488 39068 3516
rect 36354 3448 36360 3460
rect 35636 3420 36360 3448
rect 36354 3408 36360 3420
rect 36412 3408 36418 3460
rect 37734 3408 37740 3460
rect 37792 3448 37798 3460
rect 38672 3448 38700 3488
rect 37792 3420 38700 3448
rect 37792 3408 37798 3420
rect 38746 3408 38752 3460
rect 38804 3408 38810 3460
rect 30524 3352 32996 3380
rect 30524 3340 30530 3352
rect 33042 3340 33048 3392
rect 33100 3380 33106 3392
rect 33689 3383 33747 3389
rect 33689 3380 33701 3383
rect 33100 3352 33701 3380
rect 33100 3340 33106 3352
rect 33689 3349 33701 3352
rect 33735 3349 33747 3383
rect 33689 3343 33747 3349
rect 34698 3340 34704 3392
rect 34756 3340 34762 3392
rect 35158 3340 35164 3392
rect 35216 3380 35222 3392
rect 38933 3383 38991 3389
rect 38933 3380 38945 3383
rect 35216 3352 38945 3380
rect 35216 3340 35222 3352
rect 38933 3349 38945 3352
rect 38979 3349 38991 3383
rect 39040 3380 39068 3488
rect 39117 3485 39129 3519
rect 39163 3516 39175 3519
rect 39298 3516 39304 3528
rect 39163 3488 39304 3516
rect 39163 3485 39175 3488
rect 39117 3479 39175 3485
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 42245 3519 42303 3525
rect 42245 3485 42257 3519
rect 42291 3485 42303 3519
rect 42245 3479 42303 3485
rect 39206 3408 39212 3460
rect 39264 3448 39270 3460
rect 41966 3448 41972 3460
rect 39264 3420 41972 3448
rect 39264 3408 39270 3420
rect 41966 3408 41972 3420
rect 42024 3408 42030 3460
rect 42260 3448 42288 3479
rect 42518 3476 42524 3528
rect 42576 3476 42582 3528
rect 42904 3525 42932 3556
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3485 42855 3519
rect 42797 3479 42855 3485
rect 42889 3519 42947 3525
rect 42889 3485 42901 3519
rect 42935 3485 42947 3519
rect 42889 3479 42947 3485
rect 42702 3448 42708 3460
rect 42260 3420 42708 3448
rect 42702 3408 42708 3420
rect 42760 3408 42766 3460
rect 42812 3448 42840 3479
rect 43254 3476 43260 3528
rect 43312 3476 43318 3528
rect 42812 3420 43300 3448
rect 43272 3392 43300 3420
rect 42337 3383 42395 3389
rect 42337 3380 42349 3383
rect 39040 3352 42349 3380
rect 38933 3343 38991 3349
rect 42337 3349 42349 3352
rect 42383 3349 42395 3383
rect 42337 3343 42395 3349
rect 43070 3340 43076 3392
rect 43128 3340 43134 3392
rect 43254 3340 43260 3392
rect 43312 3340 43318 3392
rect 1104 3290 43884 3312
rect 1104 3238 2658 3290
rect 2710 3238 2722 3290
rect 2774 3238 2786 3290
rect 2838 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 8658 3290
rect 8710 3238 8722 3290
rect 8774 3238 8786 3290
rect 8838 3238 8850 3290
rect 8902 3238 8914 3290
rect 8966 3238 8978 3290
rect 9030 3238 14658 3290
rect 14710 3238 14722 3290
rect 14774 3238 14786 3290
rect 14838 3238 14850 3290
rect 14902 3238 14914 3290
rect 14966 3238 14978 3290
rect 15030 3238 20658 3290
rect 20710 3238 20722 3290
rect 20774 3238 20786 3290
rect 20838 3238 20850 3290
rect 20902 3238 20914 3290
rect 20966 3238 20978 3290
rect 21030 3238 26658 3290
rect 26710 3238 26722 3290
rect 26774 3238 26786 3290
rect 26838 3238 26850 3290
rect 26902 3238 26914 3290
rect 26966 3238 26978 3290
rect 27030 3238 32658 3290
rect 32710 3238 32722 3290
rect 32774 3238 32786 3290
rect 32838 3238 32850 3290
rect 32902 3238 32914 3290
rect 32966 3238 32978 3290
rect 33030 3238 38658 3290
rect 38710 3238 38722 3290
rect 38774 3238 38786 3290
rect 38838 3238 38850 3290
rect 38902 3238 38914 3290
rect 38966 3238 38978 3290
rect 39030 3238 43884 3290
rect 1104 3216 43884 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 6178 3176 6184 3188
rect 2915 3148 6184 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 7742 3136 7748 3188
rect 7800 3136 7806 3188
rect 13357 3179 13415 3185
rect 8128 3148 13216 3176
rect 2774 3068 2780 3120
rect 2832 3068 2838 3120
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 7760 3108 7788 3136
rect 8018 3108 8024 3120
rect 3108 3080 8024 3108
rect 3108 3068 3114 3080
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 2314 3000 2320 3052
rect 2372 3000 2378 3052
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 8128 3049 8156 3148
rect 10778 3108 10784 3120
rect 9692 3080 10784 3108
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 5224 3012 6653 3040
rect 5224 3000 5230 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 8113 3043 8171 3049
rect 7791 3012 8064 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 1394 2932 1400 2984
rect 1452 2932 1458 2984
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2941 1731 2975
rect 1673 2935 1731 2941
rect 1688 2836 1716 2935
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 6362 2972 6368 2984
rect 4764 2944 6368 2972
rect 4764 2932 4770 2944
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7892 2944 7941 2972
rect 7892 2932 7898 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 8036 2972 8064 3012
rect 8113 3009 8125 3043
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8294 2972 8300 2984
rect 8036 2944 8300 2972
rect 7929 2935 7987 2941
rect 8294 2932 8300 2944
rect 8352 2932 8358 2984
rect 8662 2932 8668 2984
rect 8720 2972 8726 2984
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 8720 2944 8861 2972
rect 8720 2932 8726 2944
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 8938 2932 8944 2984
rect 8996 2981 9002 2984
rect 8996 2975 9024 2981
rect 9012 2941 9024 2975
rect 8996 2935 9024 2941
rect 8996 2932 9002 2935
rect 9122 2932 9128 2984
rect 9180 2932 9186 2984
rect 2498 2864 2504 2916
rect 2556 2864 2562 2916
rect 7484 2876 8524 2904
rect 7484 2836 7512 2876
rect 1688 2808 7512 2836
rect 7561 2839 7619 2845
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 7834 2836 7840 2848
rect 7607 2808 7840 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 8496 2836 8524 2876
rect 8570 2864 8576 2916
rect 8628 2864 8634 2916
rect 9692 2836 9720 3080
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3040 10287 3043
rect 10502 3040 10508 3052
rect 10275 3012 10508 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10612 3049 10640 3080
rect 10778 3068 10784 3080
rect 10836 3068 10842 3120
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 10686 3000 10692 3052
rect 10744 3040 10750 3052
rect 11716 3049 11744 3148
rect 13188 3108 13216 3148
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 14274 3176 14280 3188
rect 13403 3148 14280 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14921 3179 14979 3185
rect 14921 3145 14933 3179
rect 14967 3176 14979 3179
rect 15930 3176 15936 3188
rect 14967 3148 15936 3176
rect 14967 3145 14979 3148
rect 14921 3139 14979 3145
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16482 3136 16488 3188
rect 16540 3136 16546 3188
rect 16850 3136 16856 3188
rect 16908 3136 16914 3188
rect 17218 3136 17224 3188
rect 17276 3136 17282 3188
rect 17497 3179 17555 3185
rect 17497 3145 17509 3179
rect 17543 3176 17555 3179
rect 19518 3176 19524 3188
rect 17543 3148 19524 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 19794 3136 19800 3188
rect 19852 3176 19858 3188
rect 25961 3179 26019 3185
rect 19852 3148 25268 3176
rect 19852 3136 19858 3148
rect 13630 3108 13636 3120
rect 13188 3080 13636 3108
rect 13630 3068 13636 3080
rect 13688 3068 13694 3120
rect 13814 3108 13820 3120
rect 13740 3080 13820 3108
rect 12618 3049 12624 3052
rect 11701 3043 11759 3049
rect 10744 3012 11652 3040
rect 10744 3000 10750 3012
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 10042 2972 10048 2984
rect 9815 2944 10048 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10318 2932 10324 2984
rect 10376 2932 10382 2984
rect 11514 2932 11520 2984
rect 11572 2932 11578 2984
rect 11624 2972 11652 3012
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12575 3043 12624 3049
rect 12575 3009 12587 3043
rect 12621 3009 12624 3043
rect 12575 3003 12624 3009
rect 12618 3000 12624 3003
rect 12676 3000 12682 3052
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 13740 3049 13768 3080
rect 13814 3068 13820 3080
rect 13872 3108 13878 3120
rect 14458 3108 14464 3120
rect 13872 3080 14464 3108
rect 13872 3068 13878 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 22097 3111 22155 3117
rect 22097 3077 22109 3111
rect 22143 3108 22155 3111
rect 22646 3108 22652 3120
rect 22143 3080 22652 3108
rect 22143 3077 22155 3080
rect 22097 3071 22155 3077
rect 22646 3068 22652 3080
rect 22704 3108 22710 3120
rect 22704 3080 23244 3108
rect 22704 3068 22710 3080
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 13412 3012 13461 3040
rect 13412 3000 13418 3012
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14056 3012 14933 3040
rect 14056 3000 14062 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15059 3012 15240 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11624 2944 12449 2972
rect 11333 2907 11391 2913
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 12161 2907 12219 2913
rect 12161 2904 12173 2907
rect 11379 2876 12173 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 12161 2873 12173 2876
rect 12207 2873 12219 2907
rect 12161 2867 12219 2873
rect 8496 2808 9720 2836
rect 10045 2839 10103 2845
rect 10045 2805 10057 2839
rect 10091 2836 10103 2839
rect 10134 2836 10140 2848
rect 10091 2808 10140 2836
rect 10091 2805 10103 2808
rect 10045 2799 10103 2805
rect 10134 2796 10140 2808
rect 10192 2796 10198 2848
rect 12268 2836 12296 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12710 2932 12716 2984
rect 12768 2932 12774 2984
rect 15028 2972 15056 3003
rect 14384 2944 15056 2972
rect 15105 2975 15163 2981
rect 14384 2836 14412 2944
rect 15105 2941 15117 2975
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 14461 2907 14519 2913
rect 14461 2873 14473 2907
rect 14507 2904 14519 2907
rect 15120 2904 15148 2935
rect 14507 2876 15148 2904
rect 14507 2873 14519 2876
rect 14461 2867 14519 2873
rect 12268 2808 14412 2836
rect 14550 2796 14556 2848
rect 14608 2796 14614 2848
rect 15212 2836 15240 3012
rect 15470 3000 15476 3052
rect 15528 3000 15534 3052
rect 15746 3000 15752 3052
rect 15804 3040 15810 3052
rect 15804 3012 16712 3040
rect 15804 3000 15810 3012
rect 16684 2972 16712 3012
rect 16758 3000 16764 3052
rect 16816 3000 16822 3052
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 17144 2972 17172 3003
rect 18138 3000 18144 3052
rect 18196 3000 18202 3052
rect 18322 3049 18328 3052
rect 18300 3043 18328 3049
rect 18300 3009 18312 3043
rect 18300 3003 18328 3009
rect 18322 3000 18328 3003
rect 18380 3000 18386 3052
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 19208 3012 19625 3040
rect 19208 3000 19214 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 20438 3000 20444 3052
rect 20496 3049 20502 3052
rect 20496 3043 20524 3049
rect 20512 3009 20524 3043
rect 20496 3003 20524 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 21545 3043 21603 3049
rect 21545 3040 21557 3043
rect 21315 3012 21557 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 21545 3009 21557 3012
rect 21591 3009 21603 3043
rect 21545 3003 21603 3009
rect 20496 3000 20502 3003
rect 21910 3000 21916 3052
rect 21968 3000 21974 3052
rect 22922 3000 22928 3052
rect 22980 3000 22986 3052
rect 23216 3049 23244 3080
rect 23860 3080 24992 3108
rect 23201 3043 23259 3049
rect 23201 3009 23213 3043
rect 23247 3040 23259 3043
rect 23293 3043 23351 3049
rect 23293 3040 23305 3043
rect 23247 3012 23305 3040
rect 23247 3009 23259 3012
rect 23201 3003 23259 3009
rect 23293 3009 23305 3012
rect 23339 3009 23351 3043
rect 23293 3003 23351 3009
rect 23566 3000 23572 3052
rect 23624 3040 23630 3052
rect 23860 3049 23888 3080
rect 24964 3052 24992 3080
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23624 3012 23857 3040
rect 23624 3000 23630 3012
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23845 3003 23903 3009
rect 24118 3000 24124 3052
rect 24176 3000 24182 3052
rect 24946 3000 24952 3052
rect 25004 3000 25010 3052
rect 25240 3049 25268 3148
rect 25961 3145 25973 3179
rect 26007 3176 26019 3179
rect 26418 3176 26424 3188
rect 26007 3148 26424 3176
rect 26007 3145 26019 3148
rect 25961 3139 26019 3145
rect 26418 3136 26424 3148
rect 26476 3136 26482 3188
rect 27154 3136 27160 3188
rect 27212 3176 27218 3188
rect 28810 3176 28816 3188
rect 27212 3148 28816 3176
rect 27212 3136 27218 3148
rect 28810 3136 28816 3148
rect 28868 3136 28874 3188
rect 30282 3136 30288 3188
rect 30340 3136 30346 3188
rect 31481 3179 31539 3185
rect 31481 3145 31493 3179
rect 31527 3176 31539 3179
rect 32490 3176 32496 3188
rect 31527 3148 32496 3176
rect 31527 3145 31539 3148
rect 31481 3139 31539 3145
rect 32490 3136 32496 3148
rect 32548 3136 32554 3188
rect 34882 3136 34888 3188
rect 34940 3176 34946 3188
rect 36173 3179 36231 3185
rect 36173 3176 36185 3179
rect 34940 3148 36185 3176
rect 34940 3136 34946 3148
rect 36173 3145 36185 3148
rect 36219 3145 36231 3179
rect 36173 3139 36231 3145
rect 36354 3136 36360 3188
rect 36412 3176 36418 3188
rect 38470 3176 38476 3188
rect 36412 3148 38476 3176
rect 36412 3136 36418 3148
rect 38470 3136 38476 3148
rect 38528 3136 38534 3188
rect 38565 3179 38623 3185
rect 38565 3145 38577 3179
rect 38611 3145 38623 3179
rect 38565 3139 38623 3145
rect 38933 3179 38991 3185
rect 38933 3145 38945 3179
rect 38979 3176 38991 3179
rect 39114 3176 39120 3188
rect 38979 3148 39120 3176
rect 38979 3145 38991 3148
rect 38933 3139 38991 3145
rect 25866 3068 25872 3120
rect 25924 3108 25930 3120
rect 25924 3080 27568 3108
rect 25924 3068 25930 3080
rect 25225 3043 25283 3049
rect 25225 3009 25237 3043
rect 25271 3009 25283 3043
rect 25225 3003 25283 3009
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 17586 2972 17592 2984
rect 16684 2944 17592 2972
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 17954 2972 17960 2984
rect 17788 2944 17960 2972
rect 17788 2904 17816 2944
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 19337 2975 19395 2981
rect 18472 2944 18644 2972
rect 18472 2932 18478 2944
rect 16132 2876 17816 2904
rect 16132 2836 16160 2876
rect 15212 2808 16160 2836
rect 18616 2836 18644 2944
rect 19337 2941 19349 2975
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 18690 2864 18696 2916
rect 18748 2864 18754 2916
rect 19352 2904 19380 2935
rect 19426 2932 19432 2984
rect 19484 2932 19490 2984
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 20346 2972 20352 2984
rect 19852 2944 20352 2972
rect 19852 2932 19858 2944
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 20625 2975 20683 2981
rect 20625 2941 20637 2975
rect 20671 2972 20683 2975
rect 21358 2972 21364 2984
rect 20671 2944 21364 2972
rect 20671 2941 20683 2944
rect 20625 2935 20683 2941
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 26068 2972 26096 3003
rect 27338 3000 27344 3052
rect 27396 3000 27402 3052
rect 27540 3049 27568 3080
rect 29454 3068 29460 3120
rect 29512 3108 29518 3120
rect 31846 3108 31852 3120
rect 29512 3080 31852 3108
rect 29512 3068 29518 3080
rect 31846 3068 31852 3080
rect 31904 3068 31910 3120
rect 38580 3108 38608 3139
rect 39114 3136 39120 3148
rect 39172 3136 39178 3188
rect 40402 3136 40408 3188
rect 40460 3136 40466 3188
rect 41138 3136 41144 3188
rect 41196 3136 41202 3188
rect 41598 3136 41604 3188
rect 41656 3136 41662 3188
rect 41785 3179 41843 3185
rect 41785 3145 41797 3179
rect 41831 3176 41843 3179
rect 41874 3176 41880 3188
rect 41831 3148 41880 3176
rect 41831 3145 41843 3148
rect 41785 3139 41843 3145
rect 41874 3136 41880 3148
rect 41932 3136 41938 3188
rect 41966 3136 41972 3188
rect 42024 3176 42030 3188
rect 42024 3148 43300 3176
rect 42024 3136 42030 3148
rect 39390 3108 39396 3120
rect 38580 3080 39396 3108
rect 39390 3068 39396 3080
rect 39448 3068 39454 3120
rect 39500 3080 42564 3108
rect 27525 3043 27583 3049
rect 27525 3009 27537 3043
rect 27571 3009 27583 3043
rect 27525 3003 27583 3009
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 27709 3043 27767 3049
rect 27709 3040 27721 3043
rect 27672 3012 27721 3040
rect 27672 3000 27678 3012
rect 27709 3009 27721 3012
rect 27755 3009 27767 3043
rect 27709 3003 27767 3009
rect 28534 3000 28540 3052
rect 28592 3049 28598 3052
rect 28592 3043 28620 3049
rect 28608 3009 28620 3043
rect 28592 3003 28620 3009
rect 29365 3043 29423 3049
rect 29365 3009 29377 3043
rect 29411 3040 29423 3043
rect 29641 3043 29699 3049
rect 29641 3040 29653 3043
rect 29411 3012 29653 3040
rect 29411 3009 29423 3012
rect 29365 3003 29423 3009
rect 29641 3009 29653 3012
rect 29687 3009 29699 3043
rect 29641 3003 29699 3009
rect 28592 3000 28598 3003
rect 30098 3000 30104 3052
rect 30156 3000 30162 3052
rect 30466 3000 30472 3052
rect 30524 3000 30530 3052
rect 30742 3000 30748 3052
rect 30800 3000 30806 3052
rect 32398 3000 32404 3052
rect 32456 3000 32462 3052
rect 32582 3000 32588 3052
rect 32640 3000 32646 3052
rect 33318 3000 33324 3052
rect 33376 3000 33382 3052
rect 33594 3000 33600 3052
rect 33652 3000 33658 3052
rect 34238 3000 34244 3052
rect 34296 3040 34302 3052
rect 34333 3043 34391 3049
rect 34333 3040 34345 3043
rect 34296 3012 34345 3040
rect 34296 3000 34302 3012
rect 34333 3009 34345 3012
rect 34379 3009 34391 3043
rect 34333 3003 34391 3009
rect 34422 3000 34428 3052
rect 34480 3040 34486 3052
rect 34517 3043 34575 3049
rect 34517 3040 34529 3043
rect 34480 3012 34529 3040
rect 34480 3000 34486 3012
rect 34517 3009 34529 3012
rect 34563 3009 34575 3043
rect 34517 3003 34575 3009
rect 35250 3000 35256 3052
rect 35308 3000 35314 3052
rect 38378 3000 38384 3052
rect 38436 3000 38442 3052
rect 38749 3043 38807 3049
rect 38749 3009 38761 3043
rect 38795 3040 38807 3043
rect 39114 3040 39120 3052
rect 38795 3012 39120 3040
rect 38795 3009 38807 3012
rect 38749 3003 38807 3009
rect 39114 3000 39120 3012
rect 39172 3000 39178 3052
rect 39500 3040 39528 3080
rect 39224 3012 39528 3040
rect 26418 2972 26424 2984
rect 26068 2944 26424 2972
rect 26418 2932 26424 2944
rect 26476 2932 26482 2984
rect 28442 2972 28448 2984
rect 27586 2944 28448 2972
rect 19610 2904 19616 2916
rect 19352 2876 19616 2904
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 20073 2907 20131 2913
rect 20073 2873 20085 2907
rect 20119 2873 20131 2907
rect 20073 2867 20131 2873
rect 22189 2907 22247 2913
rect 22189 2873 22201 2907
rect 22235 2904 22247 2907
rect 22278 2904 22284 2916
rect 22235 2876 22284 2904
rect 22235 2873 22247 2876
rect 22189 2867 22247 2873
rect 19794 2836 19800 2848
rect 18616 2808 19800 2836
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 20088 2836 20116 2867
rect 22278 2864 22284 2876
rect 22336 2864 22342 2916
rect 23124 2876 23704 2904
rect 20346 2836 20352 2848
rect 20088 2808 20352 2836
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 21140 2808 21373 2836
rect 21140 2796 21146 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 21361 2799 21419 2805
rect 21450 2796 21456 2848
rect 21508 2836 21514 2848
rect 23124 2836 23152 2876
rect 21508 2808 23152 2836
rect 23477 2839 23535 2845
rect 21508 2796 21514 2808
rect 23477 2805 23489 2839
rect 23523 2836 23535 2839
rect 23566 2836 23572 2848
rect 23523 2808 23572 2836
rect 23523 2805 23535 2808
rect 23477 2799 23535 2805
rect 23566 2796 23572 2808
rect 23624 2796 23630 2848
rect 23676 2836 23704 2876
rect 24854 2864 24860 2916
rect 24912 2864 24918 2916
rect 26237 2907 26295 2913
rect 26237 2873 26249 2907
rect 26283 2904 26295 2907
rect 26510 2904 26516 2916
rect 26283 2876 26516 2904
rect 26283 2873 26295 2876
rect 26237 2867 26295 2873
rect 26510 2864 26516 2876
rect 26568 2864 26574 2916
rect 27154 2864 27160 2916
rect 27212 2864 27218 2916
rect 27586 2836 27614 2944
rect 28442 2932 28448 2944
rect 28500 2932 28506 2984
rect 28718 2932 28724 2984
rect 28776 2932 28782 2984
rect 33042 2932 33048 2984
rect 33100 2932 33106 2984
rect 33410 2932 33416 2984
rect 33468 2981 33474 2984
rect 33468 2975 33496 2981
rect 33484 2941 33496 2975
rect 33468 2935 33496 2941
rect 33468 2932 33474 2935
rect 35342 2932 35348 2984
rect 35400 2981 35406 2984
rect 35400 2975 35428 2981
rect 35416 2941 35428 2975
rect 35400 2935 35428 2941
rect 35400 2932 35406 2935
rect 35526 2932 35532 2984
rect 35584 2932 35590 2984
rect 37182 2932 37188 2984
rect 37240 2972 37246 2984
rect 39224 2972 39252 3012
rect 40586 3000 40592 3052
rect 40644 3000 40650 3052
rect 41322 3000 41328 3052
rect 41380 3000 41386 3052
rect 41414 3000 41420 3052
rect 41472 3000 41478 3052
rect 41966 3000 41972 3052
rect 42024 3000 42030 3052
rect 42242 3000 42248 3052
rect 42300 3000 42306 3052
rect 42536 3049 42564 3080
rect 43272 3049 43300 3148
rect 43438 3136 43444 3188
rect 43496 3136 43502 3188
rect 42521 3043 42579 3049
rect 42521 3009 42533 3043
rect 42567 3009 42579 3043
rect 42521 3003 42579 3009
rect 42889 3043 42947 3049
rect 42889 3009 42901 3043
rect 42935 3009 42947 3043
rect 42889 3003 42947 3009
rect 43257 3043 43315 3049
rect 43257 3009 43269 3043
rect 43303 3009 43315 3043
rect 43257 3003 43315 3009
rect 37240 2944 39252 2972
rect 37240 2932 37246 2944
rect 39390 2932 39396 2984
rect 39448 2972 39454 2984
rect 42904 2972 42932 3003
rect 39448 2944 42932 2972
rect 39448 2932 39454 2944
rect 28166 2864 28172 2916
rect 28224 2864 28230 2916
rect 34072 2876 34652 2904
rect 23676 2808 27614 2836
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 29178 2836 29184 2848
rect 27764 2808 29184 2836
rect 27764 2796 27770 2808
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 29454 2796 29460 2848
rect 29512 2796 29518 2848
rect 29730 2796 29736 2848
rect 29788 2836 29794 2848
rect 33962 2836 33968 2848
rect 29788 2808 33968 2836
rect 29788 2796 29794 2808
rect 33962 2796 33968 2808
rect 34020 2836 34026 2848
rect 34072 2836 34100 2876
rect 34020 2808 34100 2836
rect 34020 2796 34026 2808
rect 34146 2796 34152 2848
rect 34204 2836 34210 2848
rect 34241 2839 34299 2845
rect 34241 2836 34253 2839
rect 34204 2808 34253 2836
rect 34204 2796 34210 2808
rect 34241 2805 34253 2808
rect 34287 2805 34299 2839
rect 34624 2836 34652 2876
rect 34698 2864 34704 2916
rect 34756 2904 34762 2916
rect 34977 2907 35035 2913
rect 34977 2904 34989 2907
rect 34756 2876 34989 2904
rect 34756 2864 34762 2876
rect 34977 2873 34989 2876
rect 35023 2873 35035 2907
rect 34977 2867 35035 2873
rect 36998 2864 37004 2916
rect 37056 2904 37062 2916
rect 40954 2904 40960 2916
rect 37056 2876 40960 2904
rect 37056 2864 37062 2876
rect 40954 2864 40960 2876
rect 41012 2864 41018 2916
rect 42705 2907 42763 2913
rect 42705 2873 42717 2907
rect 42751 2904 42763 2907
rect 42886 2904 42892 2916
rect 42751 2876 42892 2904
rect 42751 2873 42763 2876
rect 42705 2867 42763 2873
rect 42886 2864 42892 2876
rect 42944 2864 42950 2916
rect 38286 2836 38292 2848
rect 34624 2808 38292 2836
rect 34241 2799 34299 2805
rect 38286 2796 38292 2808
rect 38344 2796 38350 2848
rect 38562 2796 38568 2848
rect 38620 2836 38626 2848
rect 42061 2839 42119 2845
rect 42061 2836 42073 2839
rect 38620 2808 42073 2836
rect 38620 2796 38626 2808
rect 42061 2805 42073 2808
rect 42107 2805 42119 2839
rect 42061 2799 42119 2805
rect 43070 2796 43076 2848
rect 43128 2796 43134 2848
rect 1104 2746 43884 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13918 2746
rect 13970 2694 13982 2746
rect 14034 2694 14046 2746
rect 14098 2694 14110 2746
rect 14162 2694 14174 2746
rect 14226 2694 14238 2746
rect 14290 2694 19918 2746
rect 19970 2694 19982 2746
rect 20034 2694 20046 2746
rect 20098 2694 20110 2746
rect 20162 2694 20174 2746
rect 20226 2694 20238 2746
rect 20290 2694 25918 2746
rect 25970 2694 25982 2746
rect 26034 2694 26046 2746
rect 26098 2694 26110 2746
rect 26162 2694 26174 2746
rect 26226 2694 26238 2746
rect 26290 2694 31918 2746
rect 31970 2694 31982 2746
rect 32034 2694 32046 2746
rect 32098 2694 32110 2746
rect 32162 2694 32174 2746
rect 32226 2694 32238 2746
rect 32290 2694 37918 2746
rect 37970 2694 37982 2746
rect 38034 2694 38046 2746
rect 38098 2694 38110 2746
rect 38162 2694 38174 2746
rect 38226 2694 38238 2746
rect 38290 2694 43884 2746
rect 1104 2672 43884 2694
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 7190 2632 7196 2644
rect 3467 2604 7196 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 8481 2635 8539 2641
rect 7423 2604 8248 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 5537 2567 5595 2573
rect 5537 2533 5549 2567
rect 5583 2564 5595 2567
rect 5902 2564 5908 2576
rect 5583 2536 5908 2564
rect 5583 2533 5595 2536
rect 5537 2527 5595 2533
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 8220 2564 8248 2604
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8570 2632 8576 2644
rect 8527 2604 8576 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 8941 2635 8999 2641
rect 8941 2601 8953 2635
rect 8987 2632 8999 2635
rect 9306 2632 9312 2644
rect 8987 2604 9312 2632
rect 8987 2601 8999 2604
rect 8941 2595 8999 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 9916 2604 10241 2632
rect 9916 2592 9922 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 11333 2635 11391 2641
rect 10376 2604 11284 2632
rect 10376 2592 10382 2604
rect 9122 2564 9128 2576
rect 8220 2536 9128 2564
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 1673 2499 1731 2505
rect 1673 2496 1685 2499
rect 1360 2468 1685 2496
rect 1360 2456 1366 2468
rect 1673 2465 1685 2468
rect 1719 2465 1731 2499
rect 1673 2459 1731 2465
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 3234 2496 3240 2508
rect 2639 2468 3240 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 5776 2468 6377 2496
rect 5776 2456 5782 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 1394 2388 1400 2440
rect 1452 2388 1458 2440
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 1820 2400 2329 2428
rect 1820 2388 1826 2400
rect 2317 2397 2329 2400
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 3326 2320 3332 2372
rect 3384 2320 3390 2372
rect 5718 2320 5724 2372
rect 5776 2320 5782 2372
rect 6380 2360 6408 2459
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 7432 2468 7481 2496
rect 7432 2456 7438 2468
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 11256 2496 11284 2604
rect 11333 2601 11345 2635
rect 11379 2632 11391 2635
rect 12529 2635 12587 2641
rect 11379 2604 12480 2632
rect 11379 2601 11391 2604
rect 11333 2595 11391 2601
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11256 2468 11529 2496
rect 7469 2459 7527 2465
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 12452 2496 12480 2604
rect 12529 2601 12541 2635
rect 12575 2632 12587 2635
rect 12710 2632 12716 2644
rect 12575 2604 12716 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 18601 2635 18659 2641
rect 14016 2604 17264 2632
rect 12618 2524 12624 2576
rect 12676 2564 12682 2576
rect 14016 2564 14044 2604
rect 12676 2536 14044 2564
rect 12676 2524 12682 2536
rect 14090 2524 14096 2576
rect 14148 2564 14154 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 14148 2536 14565 2564
rect 14148 2524 14154 2536
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 14553 2527 14611 2533
rect 12452 2468 16574 2496
rect 11517 2459 11575 2465
rect 6638 2388 6644 2440
rect 6696 2428 6702 2440
rect 6696 2400 7512 2428
rect 6696 2388 6702 2400
rect 7374 2360 7380 2372
rect 6380 2332 7380 2360
rect 7374 2320 7380 2332
rect 7432 2320 7438 2372
rect 7484 2360 7512 2400
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 9677 2431 9735 2437
rect 9677 2428 9689 2431
rect 7852 2400 9689 2428
rect 7852 2360 7880 2400
rect 9677 2397 9689 2400
rect 9723 2428 9735 2431
rect 9766 2428 9772 2440
rect 9723 2400 9772 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 9953 2431 10011 2437
rect 9953 2397 9965 2431
rect 9999 2397 10011 2431
rect 10045 2431 10103 2437
rect 10045 2430 10057 2431
rect 10091 2430 10103 2431
rect 10321 2431 10379 2437
rect 9953 2391 10011 2397
rect 7484 2332 7880 2360
rect 9398 2320 9404 2372
rect 9456 2360 9462 2372
rect 9968 2360 9996 2391
rect 10042 2378 10048 2430
rect 10100 2378 10106 2430
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 9456 2332 9996 2360
rect 10336 2360 10364 2391
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2428 11851 2431
rect 12434 2428 12440 2440
rect 11839 2400 12440 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 14550 2428 14556 2440
rect 13771 2400 14556 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 11606 2360 11612 2372
rect 10336 2332 11612 2360
rect 9456 2320 9462 2332
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3568 2264 3893 2292
rect 3568 2252 3574 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 3881 2255 3939 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4580 2264 4721 2292
rect 4580 2252 4586 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6914 2292 6920 2304
rect 6043 2264 6920 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7282 2252 7288 2304
rect 7340 2292 7346 2304
rect 12636 2292 12664 2391
rect 12710 2320 12716 2372
rect 12768 2360 12774 2372
rect 13004 2360 13032 2391
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 12768 2332 13032 2360
rect 14185 2363 14243 2369
rect 12768 2320 12774 2332
rect 14185 2329 14197 2363
rect 14231 2329 14243 2363
rect 14185 2323 14243 2329
rect 7340 2264 12664 2292
rect 7340 2252 7346 2264
rect 12802 2252 12808 2304
rect 12860 2252 12866 2304
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 13538 2252 13544 2304
rect 13596 2252 13602 2304
rect 14200 2292 14228 2323
rect 14366 2320 14372 2372
rect 14424 2320 14430 2372
rect 14752 2360 14780 2391
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 16546 2428 16574 2468
rect 17236 2437 17264 2604
rect 18601 2601 18613 2635
rect 18647 2632 18659 2635
rect 18690 2632 18696 2644
rect 18647 2604 18696 2632
rect 18647 2601 18659 2604
rect 18601 2595 18659 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 18782 2592 18788 2644
rect 18840 2632 18846 2644
rect 20257 2635 20315 2641
rect 18840 2604 20208 2632
rect 18840 2592 18846 2604
rect 20180 2564 20208 2604
rect 20257 2601 20269 2635
rect 20303 2632 20315 2635
rect 20346 2632 20352 2644
rect 20303 2604 20352 2632
rect 20303 2601 20315 2604
rect 20257 2595 20315 2601
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 21266 2632 21272 2644
rect 20456 2604 21272 2632
rect 20456 2564 20484 2604
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 21358 2592 21364 2644
rect 21416 2592 21422 2644
rect 23385 2635 23443 2641
rect 22204 2604 23060 2632
rect 20180 2536 20484 2564
rect 20346 2456 20352 2508
rect 20404 2456 20410 2508
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16546 2400 16681 2428
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 17862 2388 17868 2440
rect 17920 2388 17926 2440
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 17494 2360 17500 2372
rect 14752 2332 17500 2360
rect 17494 2320 17500 2332
rect 17552 2320 17558 2372
rect 17604 2360 17632 2388
rect 19260 2360 19288 2391
rect 19518 2388 19524 2440
rect 19576 2428 19582 2440
rect 19576 2400 20484 2428
rect 19576 2388 19582 2400
rect 20346 2360 20352 2372
rect 17604 2332 20352 2360
rect 20346 2320 20352 2332
rect 20404 2320 20410 2372
rect 20456 2360 20484 2400
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20588 2400 20637 2428
rect 20588 2388 20594 2400
rect 20625 2397 20637 2400
rect 20671 2428 20683 2431
rect 22204 2428 22232 2604
rect 23032 2564 23060 2604
rect 23385 2601 23397 2635
rect 23431 2632 23443 2635
rect 24026 2632 24032 2644
rect 23431 2604 24032 2632
rect 23431 2601 23443 2604
rect 23385 2595 23443 2601
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 25961 2635 26019 2641
rect 24228 2604 25636 2632
rect 24228 2564 24256 2604
rect 23032 2536 24256 2564
rect 22370 2456 22376 2508
rect 22428 2456 22434 2508
rect 24946 2456 24952 2508
rect 25004 2456 25010 2508
rect 20671 2400 22232 2428
rect 22281 2431 22339 2437
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 22281 2397 22293 2431
rect 22327 2428 22339 2431
rect 22649 2431 22707 2437
rect 22327 2400 22508 2428
rect 22327 2397 22339 2400
rect 22281 2391 22339 2397
rect 22480 2372 22508 2400
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 20456 2332 22232 2360
rect 14458 2292 14464 2304
rect 14200 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 15286 2252 15292 2304
rect 15344 2292 15350 2304
rect 15473 2295 15531 2301
rect 15473 2292 15485 2295
rect 15344 2264 15485 2292
rect 15344 2252 15350 2264
rect 15473 2261 15485 2264
rect 15519 2261 15531 2295
rect 15473 2255 15531 2261
rect 16574 2252 16580 2304
rect 16632 2292 16638 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16632 2264 16865 2292
rect 16632 2252 16638 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2292 17463 2295
rect 17678 2292 17684 2304
rect 17451 2264 17684 2292
rect 17451 2261 17463 2264
rect 17405 2255 17463 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 18104 2264 22109 2292
rect 18104 2252 18110 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22204 2292 22232 2332
rect 22462 2320 22468 2372
rect 22520 2320 22526 2372
rect 22664 2304 22692 2391
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 25608 2428 25636 2604
rect 25961 2601 25973 2635
rect 26007 2632 26019 2635
rect 26326 2632 26332 2644
rect 26007 2604 26332 2632
rect 26007 2601 26019 2604
rect 25961 2595 26019 2601
rect 26326 2592 26332 2604
rect 26384 2592 26390 2644
rect 28166 2592 28172 2644
rect 28224 2592 28230 2644
rect 28718 2632 28724 2644
rect 28368 2604 28724 2632
rect 28077 2567 28135 2573
rect 28077 2533 28089 2567
rect 28123 2564 28135 2567
rect 28368 2564 28396 2604
rect 28718 2592 28724 2604
rect 28776 2592 28782 2644
rect 28810 2592 28816 2644
rect 28868 2632 28874 2644
rect 30098 2632 30104 2644
rect 28868 2604 30104 2632
rect 28868 2592 28874 2604
rect 30098 2592 30104 2604
rect 30156 2632 30162 2644
rect 31389 2635 31447 2641
rect 30156 2604 31064 2632
rect 30156 2592 30162 2604
rect 28123 2536 28396 2564
rect 28123 2533 28135 2536
rect 28077 2527 28135 2533
rect 25774 2456 25780 2508
rect 25832 2496 25838 2508
rect 27062 2496 27068 2508
rect 25832 2468 27068 2496
rect 25832 2456 25838 2468
rect 27062 2456 27068 2468
rect 27120 2456 27126 2508
rect 29178 2456 29184 2508
rect 29236 2496 29242 2508
rect 30374 2496 30380 2508
rect 29236 2468 30380 2496
rect 29236 2456 29242 2468
rect 30374 2456 30380 2468
rect 30432 2456 30438 2508
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 25608 2400 27353 2428
rect 27341 2397 27353 2400
rect 27387 2428 27399 2431
rect 28810 2428 28816 2440
rect 27387 2400 28816 2428
rect 27387 2397 27399 2400
rect 27341 2391 27399 2397
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 28902 2388 28908 2440
rect 28960 2388 28966 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 29104 2400 30665 2428
rect 22922 2320 22928 2372
rect 22980 2360 22986 2372
rect 26418 2360 26424 2372
rect 22980 2332 26424 2360
rect 22980 2320 22986 2332
rect 26418 2320 26424 2332
rect 26476 2360 26482 2372
rect 28920 2360 28948 2388
rect 26476 2332 28948 2360
rect 26476 2320 26482 2332
rect 22554 2292 22560 2304
rect 22204 2264 22560 2292
rect 22097 2255 22155 2261
rect 22554 2252 22560 2264
rect 22612 2252 22618 2304
rect 22646 2252 22652 2304
rect 22704 2292 22710 2304
rect 29104 2292 29132 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 31036 2360 31064 2604
rect 31389 2601 31401 2635
rect 31435 2632 31447 2635
rect 31662 2632 31668 2644
rect 31435 2604 31668 2632
rect 31435 2601 31447 2604
rect 31389 2595 31447 2601
rect 31662 2592 31668 2604
rect 31720 2592 31726 2644
rect 33137 2635 33195 2641
rect 33137 2601 33149 2635
rect 33183 2632 33195 2635
rect 33502 2632 33508 2644
rect 33183 2604 33508 2632
rect 33183 2601 33195 2604
rect 33137 2595 33195 2601
rect 33502 2592 33508 2604
rect 33560 2592 33566 2644
rect 34698 2592 34704 2644
rect 34756 2592 34762 2644
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 35805 2635 35863 2641
rect 35805 2632 35817 2635
rect 35676 2604 35817 2632
rect 35676 2592 35682 2604
rect 35805 2601 35817 2604
rect 35851 2601 35863 2635
rect 35805 2595 35863 2601
rect 42153 2567 42211 2573
rect 42153 2533 42165 2567
rect 42199 2564 42211 2567
rect 42794 2564 42800 2576
rect 42199 2536 42800 2564
rect 42199 2533 42211 2536
rect 42153 2527 42211 2533
rect 42794 2524 42800 2536
rect 42852 2524 42858 2576
rect 43438 2524 43444 2576
rect 43496 2524 43502 2576
rect 31110 2456 31116 2508
rect 31168 2496 31174 2508
rect 32122 2496 32128 2508
rect 31168 2468 32128 2496
rect 31168 2456 31174 2468
rect 32122 2456 32128 2468
rect 32180 2456 32186 2508
rect 33778 2456 33784 2508
rect 33836 2496 33842 2508
rect 33836 2468 34468 2496
rect 33836 2456 33842 2468
rect 34440 2440 34468 2468
rect 39298 2456 39304 2508
rect 39356 2496 39362 2508
rect 39356 2468 42932 2496
rect 39356 2456 39362 2468
rect 32401 2431 32459 2437
rect 32401 2397 32413 2431
rect 32447 2397 32459 2431
rect 32401 2391 32459 2397
rect 32416 2360 32444 2391
rect 34146 2388 34152 2440
rect 34204 2388 34210 2440
rect 34422 2388 34428 2440
rect 34480 2428 34486 2440
rect 35342 2428 35348 2440
rect 34480 2400 35348 2428
rect 34480 2388 34486 2400
rect 35342 2388 35348 2400
rect 35400 2388 35406 2440
rect 35434 2388 35440 2440
rect 35492 2388 35498 2440
rect 35713 2431 35771 2437
rect 35713 2397 35725 2431
rect 35759 2428 35771 2431
rect 35986 2428 35992 2440
rect 35759 2400 35992 2428
rect 35759 2397 35771 2400
rect 35713 2391 35771 2397
rect 35728 2360 35756 2391
rect 35986 2388 35992 2400
rect 36044 2388 36050 2440
rect 36538 2388 36544 2440
rect 36596 2388 36602 2440
rect 42904 2437 42932 2468
rect 36817 2431 36875 2437
rect 36817 2397 36829 2431
rect 36863 2397 36875 2431
rect 36817 2391 36875 2397
rect 41969 2431 42027 2437
rect 41969 2397 41981 2431
rect 42015 2397 42027 2431
rect 41969 2391 42027 2397
rect 42521 2431 42579 2437
rect 42521 2397 42533 2431
rect 42567 2397 42579 2431
rect 42521 2391 42579 2397
rect 42889 2431 42947 2437
rect 42889 2397 42901 2431
rect 42935 2397 42947 2431
rect 42889 2391 42947 2397
rect 43257 2431 43315 2437
rect 43257 2397 43269 2431
rect 43303 2428 43315 2431
rect 43303 2400 43944 2428
rect 43303 2397 43315 2400
rect 43257 2391 43315 2397
rect 31036 2332 32444 2360
rect 33888 2332 35756 2360
rect 36004 2360 36032 2388
rect 36832 2360 36860 2391
rect 36004 2332 36860 2360
rect 22704 2264 29132 2292
rect 22704 2252 22710 2264
rect 32122 2252 32128 2304
rect 32180 2292 32186 2304
rect 33888 2292 33916 2332
rect 36906 2320 36912 2372
rect 36964 2360 36970 2372
rect 41984 2360 42012 2391
rect 36964 2332 42012 2360
rect 36964 2320 36970 2332
rect 32180 2264 33916 2292
rect 32180 2252 32186 2264
rect 33962 2252 33968 2304
rect 34020 2252 34026 2304
rect 39482 2252 39488 2304
rect 39540 2292 39546 2304
rect 42536 2292 42564 2391
rect 39540 2264 42564 2292
rect 42705 2295 42763 2301
rect 39540 2252 39546 2264
rect 42705 2261 42717 2295
rect 42751 2292 42763 2295
rect 42886 2292 42892 2304
rect 42751 2264 42892 2292
rect 42751 2261 42763 2264
rect 42705 2255 42763 2261
rect 42886 2252 42892 2264
rect 42944 2252 42950 2304
rect 43070 2252 43076 2304
rect 43128 2252 43134 2304
rect 1104 2202 43884 2224
rect 1104 2150 2658 2202
rect 2710 2150 2722 2202
rect 2774 2150 2786 2202
rect 2838 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 8658 2202
rect 8710 2150 8722 2202
rect 8774 2150 8786 2202
rect 8838 2150 8850 2202
rect 8902 2150 8914 2202
rect 8966 2150 8978 2202
rect 9030 2150 14658 2202
rect 14710 2150 14722 2202
rect 14774 2150 14786 2202
rect 14838 2150 14850 2202
rect 14902 2150 14914 2202
rect 14966 2150 14978 2202
rect 15030 2150 20658 2202
rect 20710 2150 20722 2202
rect 20774 2150 20786 2202
rect 20838 2150 20850 2202
rect 20902 2150 20914 2202
rect 20966 2150 20978 2202
rect 21030 2150 26658 2202
rect 26710 2150 26722 2202
rect 26774 2150 26786 2202
rect 26838 2150 26850 2202
rect 26902 2150 26914 2202
rect 26966 2150 26978 2202
rect 27030 2150 32658 2202
rect 32710 2150 32722 2202
rect 32774 2150 32786 2202
rect 32838 2150 32850 2202
rect 32902 2150 32914 2202
rect 32966 2150 32978 2202
rect 33030 2150 38658 2202
rect 38710 2150 38722 2202
rect 38774 2150 38786 2202
rect 38838 2150 38850 2202
rect 38902 2150 38914 2202
rect 38966 2150 38978 2202
rect 39030 2150 43884 2202
rect 1104 2128 43884 2150
rect 9858 2048 9864 2100
rect 9916 2088 9922 2100
rect 13170 2088 13176 2100
rect 9916 2060 13176 2088
rect 9916 2048 9922 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 17494 2048 17500 2100
rect 17552 2088 17558 2100
rect 19150 2088 19156 2100
rect 17552 2060 19156 2088
rect 17552 2048 17558 2060
rect 19150 2048 19156 2060
rect 19208 2048 19214 2100
rect 19426 2048 19432 2100
rect 19484 2088 19490 2100
rect 30006 2088 30012 2100
rect 19484 2060 30012 2088
rect 19484 2048 19490 2060
rect 30006 2048 30012 2060
rect 30064 2048 30070 2100
rect 32766 2048 32772 2100
rect 32824 2088 32830 2100
rect 35802 2088 35808 2100
rect 32824 2060 35808 2088
rect 32824 2048 32830 2060
rect 35802 2048 35808 2060
rect 35860 2048 35866 2100
rect 4798 1980 4804 2032
rect 4856 2020 4862 2032
rect 11330 2020 11336 2032
rect 4856 1992 11336 2020
rect 4856 1980 4862 1992
rect 11330 1980 11336 1992
rect 11388 1980 11394 2032
rect 15654 1980 15660 2032
rect 15712 2020 15718 2032
rect 15712 1992 26924 2020
rect 15712 1980 15718 1992
rect 4062 1912 4068 1964
rect 4120 1952 4126 1964
rect 11146 1952 11152 1964
rect 4120 1924 11152 1952
rect 4120 1912 4126 1924
rect 11146 1912 11152 1924
rect 11204 1912 11210 1964
rect 13538 1952 13544 1964
rect 11624 1924 13544 1952
rect 9766 1844 9772 1896
rect 9824 1884 9830 1896
rect 10594 1884 10600 1896
rect 9824 1856 10600 1884
rect 9824 1844 9830 1856
rect 10594 1844 10600 1856
rect 10652 1844 10658 1896
rect 5166 1776 5172 1828
rect 5224 1816 5230 1828
rect 11624 1816 11652 1924
rect 13538 1912 13544 1924
rect 13596 1912 13602 1964
rect 15470 1912 15476 1964
rect 15528 1952 15534 1964
rect 21082 1952 21088 1964
rect 15528 1924 21088 1952
rect 15528 1912 15534 1924
rect 21082 1912 21088 1924
rect 21140 1912 21146 1964
rect 11790 1844 11796 1896
rect 11848 1884 11854 1896
rect 19978 1884 19984 1896
rect 11848 1856 19984 1884
rect 11848 1844 11854 1856
rect 19978 1844 19984 1856
rect 20036 1844 20042 1896
rect 24394 1884 24400 1896
rect 20088 1856 24400 1884
rect 5224 1788 11652 1816
rect 5224 1776 5230 1788
rect 13078 1776 13084 1828
rect 13136 1816 13142 1828
rect 20088 1816 20116 1856
rect 24394 1844 24400 1856
rect 24452 1844 24458 1896
rect 26896 1884 26924 1992
rect 28994 1980 29000 2032
rect 29052 2020 29058 2032
rect 29052 1992 32996 2020
rect 29052 1980 29058 1992
rect 29086 1912 29092 1964
rect 29144 1952 29150 1964
rect 32968 1952 32996 1992
rect 33042 1980 33048 2032
rect 33100 2020 33106 2032
rect 36906 2020 36912 2032
rect 33100 1992 36912 2020
rect 33100 1980 33106 1992
rect 36906 1980 36912 1992
rect 36964 1980 36970 2032
rect 37826 1952 37832 1964
rect 29144 1924 32812 1952
rect 32968 1924 37832 1952
rect 29144 1912 29150 1924
rect 26896 1856 31754 1884
rect 13136 1788 20116 1816
rect 13136 1776 13142 1788
rect 20162 1776 20168 1828
rect 20220 1816 20226 1828
rect 24578 1816 24584 1828
rect 20220 1788 24584 1816
rect 20220 1776 20226 1788
rect 24578 1776 24584 1788
rect 24636 1776 24642 1828
rect 31726 1816 31754 1856
rect 32784 1816 32812 1924
rect 37826 1912 37832 1924
rect 37884 1912 37890 1964
rect 39390 1816 39396 1828
rect 31726 1788 32444 1816
rect 32784 1788 39396 1816
rect 6546 1708 6552 1760
rect 6604 1748 6610 1760
rect 13446 1748 13452 1760
rect 6604 1720 13452 1748
rect 6604 1708 6610 1720
rect 13446 1708 13452 1720
rect 13504 1708 13510 1760
rect 17034 1708 17040 1760
rect 17092 1748 17098 1760
rect 32306 1748 32312 1760
rect 17092 1720 32312 1748
rect 17092 1708 17098 1720
rect 32306 1708 32312 1720
rect 32364 1708 32370 1760
rect 32416 1748 32444 1788
rect 39390 1776 39396 1788
rect 39448 1776 39454 1828
rect 32416 1720 35848 1748
rect 9398 1640 9404 1692
rect 9456 1680 9462 1692
rect 17586 1680 17592 1692
rect 9456 1652 17592 1680
rect 9456 1640 9462 1652
rect 17586 1640 17592 1652
rect 17644 1640 17650 1692
rect 17770 1640 17776 1692
rect 17828 1680 17834 1692
rect 22646 1680 22652 1692
rect 17828 1652 22652 1680
rect 17828 1640 17834 1652
rect 22646 1640 22652 1652
rect 22704 1640 22710 1692
rect 25038 1640 25044 1692
rect 25096 1680 25102 1692
rect 35710 1680 35716 1692
rect 25096 1652 35716 1680
rect 25096 1640 25102 1652
rect 35710 1640 35716 1652
rect 35768 1640 35774 1692
rect 35820 1680 35848 1720
rect 35894 1708 35900 1760
rect 35952 1748 35958 1760
rect 39666 1748 39672 1760
rect 35952 1720 39672 1748
rect 35952 1708 35958 1720
rect 39666 1708 39672 1720
rect 39724 1708 39730 1760
rect 37090 1680 37096 1692
rect 35820 1652 37096 1680
rect 37090 1640 37096 1652
rect 37148 1640 37154 1692
rect 40034 1640 40040 1692
rect 40092 1680 40098 1692
rect 41966 1680 41972 1692
rect 40092 1652 41972 1680
rect 40092 1640 40098 1652
rect 41966 1640 41972 1652
rect 42024 1640 42030 1692
rect 5534 1572 5540 1624
rect 5592 1612 5598 1624
rect 5592 1584 13860 1612
rect 5592 1572 5598 1584
rect 1670 1504 1676 1556
rect 1728 1544 1734 1556
rect 12342 1544 12348 1556
rect 1728 1516 12348 1544
rect 1728 1504 1734 1516
rect 12342 1504 12348 1516
rect 12400 1504 12406 1556
rect 13832 1544 13860 1584
rect 14458 1572 14464 1624
rect 14516 1612 14522 1624
rect 17402 1612 17408 1624
rect 14516 1584 17408 1612
rect 14516 1572 14522 1584
rect 17402 1572 17408 1584
rect 17460 1572 17466 1624
rect 22002 1572 22008 1624
rect 22060 1612 22066 1624
rect 43916 1612 43944 2400
rect 22060 1584 43944 1612
rect 22060 1572 22066 1584
rect 16206 1544 16212 1556
rect 13832 1516 16212 1544
rect 16206 1504 16212 1516
rect 16264 1504 16270 1556
rect 25222 1544 25228 1556
rect 19306 1516 25228 1544
rect 10594 1436 10600 1488
rect 10652 1476 10658 1488
rect 19306 1476 19334 1516
rect 25222 1504 25228 1516
rect 25280 1504 25286 1556
rect 32030 1504 32036 1556
rect 32088 1544 32094 1556
rect 34054 1544 34060 1556
rect 32088 1516 34060 1544
rect 32088 1504 32094 1516
rect 34054 1504 34060 1516
rect 34112 1504 34118 1556
rect 39114 1544 39120 1556
rect 34532 1516 39120 1544
rect 10652 1448 19334 1476
rect 10652 1436 10658 1448
rect 19610 1436 19616 1488
rect 19668 1476 19674 1488
rect 19668 1448 22048 1476
rect 19668 1436 19674 1448
rect 22020 1408 22048 1448
rect 22094 1436 22100 1488
rect 22152 1476 22158 1488
rect 34422 1476 34428 1488
rect 22152 1448 34428 1476
rect 22152 1436 22158 1448
rect 34422 1436 34428 1448
rect 34480 1436 34486 1488
rect 28350 1408 28356 1420
rect 19352 1380 20760 1408
rect 22020 1380 28356 1408
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 9950 1340 9956 1352
rect 5040 1312 9956 1340
rect 5040 1300 5046 1312
rect 9950 1300 9956 1312
rect 10008 1300 10014 1352
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 4430 1232 4436 1284
rect 4488 1272 4494 1284
rect 11716 1272 11744 1300
rect 4488 1244 11744 1272
rect 4488 1232 4494 1244
rect 15102 1232 15108 1284
rect 15160 1272 15166 1284
rect 19352 1272 19380 1380
rect 20732 1340 20760 1380
rect 28350 1368 28356 1380
rect 28408 1368 28414 1420
rect 34532 1408 34560 1516
rect 39114 1504 39120 1516
rect 39172 1504 39178 1556
rect 37274 1436 37280 1488
rect 37332 1476 37338 1488
rect 42242 1476 42248 1488
rect 37332 1448 42248 1476
rect 37332 1436 37338 1448
rect 42242 1436 42248 1448
rect 42300 1436 42306 1488
rect 40586 1408 40592 1420
rect 34348 1380 34560 1408
rect 34624 1380 40592 1408
rect 20732 1312 31984 1340
rect 15160 1244 19380 1272
rect 15160 1232 15166 1244
rect 20070 1232 20076 1284
rect 20128 1272 20134 1284
rect 21910 1272 21916 1284
rect 20128 1244 21916 1272
rect 20128 1232 20134 1244
rect 21910 1232 21916 1244
rect 21968 1232 21974 1284
rect 22002 1232 22008 1284
rect 22060 1272 22066 1284
rect 28074 1272 28080 1284
rect 22060 1244 28080 1272
rect 22060 1232 22066 1244
rect 28074 1232 28080 1244
rect 28132 1232 28138 1284
rect 11698 1164 11704 1216
rect 11756 1204 11762 1216
rect 12802 1204 12808 1216
rect 11756 1176 12808 1204
rect 11756 1164 11762 1176
rect 12802 1164 12808 1176
rect 12860 1164 12866 1216
rect 19150 1164 19156 1216
rect 19208 1204 19214 1216
rect 23750 1204 23756 1216
rect 19208 1176 23756 1204
rect 19208 1164 19214 1176
rect 23750 1164 23756 1176
rect 23808 1164 23814 1216
rect 4614 1096 4620 1148
rect 4672 1136 4678 1148
rect 23474 1136 23480 1148
rect 4672 1108 23480 1136
rect 4672 1096 4678 1108
rect 23474 1096 23480 1108
rect 23532 1096 23538 1148
rect 30834 1136 30840 1148
rect 23584 1108 30840 1136
rect 8478 1028 8484 1080
rect 8536 1068 8542 1080
rect 15470 1068 15476 1080
rect 8536 1040 15476 1068
rect 8536 1028 8542 1040
rect 15470 1028 15476 1040
rect 15528 1028 15534 1080
rect 15562 1028 15568 1080
rect 15620 1068 15626 1080
rect 23584 1068 23612 1108
rect 30834 1096 30840 1108
rect 30892 1096 30898 1148
rect 31956 1136 31984 1312
rect 33318 1232 33324 1284
rect 33376 1272 33382 1284
rect 34348 1272 34376 1380
rect 34422 1300 34428 1352
rect 34480 1340 34486 1352
rect 34624 1340 34652 1380
rect 40586 1368 40592 1380
rect 40644 1368 40650 1420
rect 34480 1312 34652 1340
rect 34480 1300 34486 1312
rect 40402 1300 40408 1352
rect 40460 1340 40466 1352
rect 41414 1340 41420 1352
rect 40460 1312 41420 1340
rect 40460 1300 40466 1312
rect 41414 1300 41420 1312
rect 41472 1300 41478 1352
rect 33376 1244 34376 1272
rect 33376 1232 33382 1244
rect 39206 1232 39212 1284
rect 39264 1272 39270 1284
rect 43254 1272 43260 1284
rect 39264 1244 43260 1272
rect 39264 1232 39270 1244
rect 43254 1232 43260 1244
rect 43312 1232 43318 1284
rect 38010 1164 38016 1216
rect 38068 1204 38074 1216
rect 42150 1204 42156 1216
rect 38068 1176 42156 1204
rect 38068 1164 38074 1176
rect 42150 1164 42156 1176
rect 42208 1164 42214 1216
rect 35894 1136 35900 1148
rect 31956 1108 35900 1136
rect 35894 1096 35900 1108
rect 35952 1096 35958 1148
rect 36814 1096 36820 1148
rect 36872 1136 36878 1148
rect 39574 1136 39580 1148
rect 36872 1108 39580 1136
rect 36872 1096 36878 1108
rect 39574 1096 39580 1108
rect 39632 1096 39638 1148
rect 15620 1040 23612 1068
rect 15620 1028 15626 1040
rect 23658 1028 23664 1080
rect 23716 1068 23722 1080
rect 28994 1068 29000 1080
rect 23716 1040 29000 1068
rect 23716 1028 23722 1040
rect 28994 1028 29000 1040
rect 29052 1028 29058 1080
rect 29638 1028 29644 1080
rect 29696 1068 29702 1080
rect 38378 1068 38384 1080
rect 29696 1040 38384 1068
rect 29696 1028 29702 1040
rect 38378 1028 38384 1040
rect 38436 1028 38442 1080
rect 6270 960 6276 1012
rect 6328 1000 6334 1012
rect 27430 1000 27436 1012
rect 6328 972 27436 1000
rect 6328 960 6334 972
rect 27430 960 27436 972
rect 27488 960 27494 1012
rect 11514 892 11520 944
rect 11572 932 11578 944
rect 29546 932 29552 944
rect 11572 904 29552 932
rect 11572 892 11578 904
rect 29546 892 29552 904
rect 29604 892 29610 944
rect 13722 824 13728 876
rect 13780 864 13786 876
rect 26234 864 26240 876
rect 13780 836 26240 864
rect 13780 824 13786 836
rect 26234 824 26240 836
rect 26292 824 26298 876
rect 6086 756 6092 808
rect 6144 796 6150 808
rect 39298 796 39304 808
rect 6144 768 39304 796
rect 6144 756 6150 768
rect 39298 756 39304 768
rect 39356 756 39362 808
rect 1578 688 1584 740
rect 1636 728 1642 740
rect 37458 728 37464 740
rect 1636 700 37464 728
rect 1636 688 1642 700
rect 37458 688 37464 700
rect 37516 688 37522 740
rect 2498 620 2504 672
rect 2556 660 2562 672
rect 36446 660 36452 672
rect 2556 632 36452 660
rect 2556 620 2562 632
rect 36446 620 36452 632
rect 36504 620 36510 672
rect 10778 552 10784 604
rect 10836 592 10842 604
rect 21818 592 21824 604
rect 10836 564 21824 592
rect 10836 552 10842 564
rect 21818 552 21824 564
rect 21876 552 21882 604
rect 23474 552 23480 604
rect 23532 592 23538 604
rect 33134 592 33140 604
rect 23532 564 33140 592
rect 23532 552 23538 564
rect 33134 552 33140 564
rect 33192 552 33198 604
rect 3786 484 3792 536
rect 3844 524 3850 536
rect 14458 524 14464 536
rect 3844 496 14464 524
rect 3844 484 3850 496
rect 14458 484 14464 496
rect 14516 484 14522 536
rect 16666 484 16672 536
rect 16724 524 16730 536
rect 22002 524 22008 536
rect 16724 496 22008 524
rect 16724 484 16730 496
rect 22002 484 22008 496
rect 22060 484 22066 536
rect 35710 484 35716 536
rect 35768 524 35774 536
rect 42610 524 42616 536
rect 35768 496 42616 524
rect 35768 484 35774 496
rect 42610 484 42616 496
rect 42668 484 42674 536
rect 4890 416 4896 468
rect 4948 456 4954 468
rect 19058 456 19064 468
rect 4948 428 19064 456
rect 4948 416 4954 428
rect 19058 416 19064 428
rect 19116 416 19122 468
rect 7098 348 7104 400
rect 7156 388 7162 400
rect 15562 388 15568 400
rect 7156 360 15568 388
rect 7156 348 7162 360
rect 15562 348 15568 360
rect 15620 348 15626 400
rect 30926 348 30932 400
rect 30984 388 30990 400
rect 42058 388 42064 400
rect 30984 360 42064 388
rect 30984 348 30990 360
rect 42058 348 42064 360
rect 42116 348 42122 400
rect 28534 280 28540 332
rect 28592 320 28598 332
rect 40034 320 40040 332
rect 28592 292 40040 320
rect 28592 280 28598 292
rect 40034 280 40040 292
rect 40092 280 40098 332
rect 24946 212 24952 264
rect 25004 252 25010 264
rect 37274 252 37280 264
rect 25004 224 37280 252
rect 25004 212 25010 224
rect 37274 212 37280 224
rect 37332 212 37338 264
rect 27338 144 27344 196
rect 27396 184 27402 196
rect 41322 184 41328 196
rect 27396 156 41328 184
rect 27396 144 27402 156
rect 41322 144 41328 156
rect 41380 144 41386 196
rect 15194 76 15200 128
rect 15252 116 15258 128
rect 21174 116 21180 128
rect 15252 88 21180 116
rect 15252 76 15258 88
rect 21174 76 21180 88
rect 21232 76 21238 128
rect 26142 76 26148 128
rect 26200 116 26206 128
rect 42518 116 42524 128
rect 26200 88 42524 116
rect 26200 76 26206 88
rect 42518 76 42524 88
rect 42576 76 42582 128
<< via1 >>
rect 14096 10888 14148 10940
rect 30104 10888 30156 10940
rect 11152 10820 11204 10872
rect 37004 10820 37056 10872
rect 4436 10752 4488 10804
rect 26884 10752 26936 10804
rect 5080 10684 5132 10736
rect 34060 10684 34112 10736
rect 6368 10616 6420 10668
rect 37096 10616 37148 10668
rect 8668 10548 8720 10600
rect 19156 10548 19208 10600
rect 30748 10480 30800 10532
rect 9220 10412 9272 10464
rect 11520 10412 11572 10464
rect 16856 10412 16908 10464
rect 21916 10412 21968 10464
rect 26700 10412 26752 10464
rect 8116 10344 8168 10396
rect 12164 10344 12216 10396
rect 14372 10344 14424 10396
rect 19616 10344 19668 10396
rect 25136 10344 25188 10396
rect 33232 10412 33284 10464
rect 33876 10412 33928 10464
rect 37280 10412 37332 10464
rect 37740 10412 37792 10464
rect 39764 10412 39816 10464
rect 30012 10344 30064 10396
rect 32588 10344 32640 10396
rect 36912 10344 36964 10396
rect 39212 10344 39264 10396
rect 7840 10276 7892 10328
rect 11796 10276 11848 10328
rect 29184 10276 29236 10328
rect 31852 10276 31904 10328
rect 36636 10276 36688 10328
rect 39028 10276 39080 10328
rect 7288 10208 7340 10260
rect 10968 10208 11020 10260
rect 11060 10208 11112 10260
rect 12624 10208 12676 10260
rect 13268 10208 13320 10260
rect 16212 10208 16264 10260
rect 29736 10208 29788 10260
rect 31576 10208 31628 10260
rect 32772 10208 32824 10260
rect 36912 10208 36964 10260
rect 37464 10208 37516 10260
rect 39488 10208 39540 10260
rect 7196 10140 7248 10192
rect 10416 10140 10468 10192
rect 22192 10140 22244 10192
rect 35348 10140 35400 10192
rect 36084 10140 36136 10192
rect 37832 10140 37884 10192
rect 7748 10072 7800 10124
rect 10692 10072 10744 10124
rect 13544 10072 13596 10124
rect 15108 10072 15160 10124
rect 19432 10072 19484 10124
rect 6644 10004 6696 10056
rect 10140 10004 10192 10056
rect 10232 10004 10284 10056
rect 14004 10004 14056 10056
rect 8300 9936 8352 9988
rect 9864 9936 9916 9988
rect 9956 9936 10008 9988
rect 13728 9936 13780 9988
rect 6460 9868 6512 9920
rect 8760 9868 8812 9920
rect 9128 9868 9180 9920
rect 11060 9868 11112 9920
rect 11336 9868 11388 9920
rect 15476 9936 15528 9988
rect 19340 10004 19392 10056
rect 21364 10004 21416 10056
rect 24676 10072 24728 10124
rect 30472 10072 30524 10124
rect 31392 10072 31444 10124
rect 34888 10072 34940 10124
rect 35532 10072 35584 10124
rect 38200 10072 38252 10124
rect 38292 10072 38344 10124
rect 40040 10072 40092 10124
rect 23204 10004 23256 10056
rect 28908 10004 28960 10056
rect 30012 10004 30064 10056
rect 30840 10004 30892 10056
rect 34796 10004 34848 10056
rect 36360 10004 36412 10056
rect 38660 10004 38712 10056
rect 38844 10004 38896 10056
rect 41052 10004 41104 10056
rect 14464 9868 14516 9920
rect 16488 9868 16540 9920
rect 5816 9800 5868 9852
rect 9036 9800 9088 9852
rect 9772 9800 9824 9852
rect 12072 9800 12124 9852
rect 13360 9800 13412 9852
rect 14280 9800 14332 9852
rect 15108 9800 15160 9852
rect 16764 9800 16816 9852
rect 25136 9936 25188 9988
rect 17132 9868 17184 9920
rect 28448 9936 28500 9988
rect 28632 9936 28684 9988
rect 29644 9936 29696 9988
rect 31116 9936 31168 9988
rect 32128 9936 32180 9988
rect 35808 9936 35860 9988
rect 37556 9936 37608 9988
rect 38568 9936 38620 9988
rect 40684 9936 40736 9988
rect 25320 9868 25372 9920
rect 27160 9868 27212 9920
rect 33324 9868 33376 9920
rect 34612 9868 34664 9920
rect 34980 9868 35032 9920
rect 36636 9868 36688 9920
rect 38016 9868 38068 9920
rect 39948 9868 40000 9920
rect 21272 9800 21324 9852
rect 21364 9800 21416 9852
rect 22928 9800 22980 9852
rect 24768 9800 24820 9852
rect 25964 9800 26016 9852
rect 27252 9800 27304 9852
rect 27896 9800 27948 9852
rect 28356 9800 28408 9852
rect 29276 9800 29328 9852
rect 29460 9800 29512 9852
rect 31484 9800 31536 9852
rect 34336 9800 34388 9852
rect 35256 9800 35308 9852
rect 35348 9800 35400 9852
rect 42524 10344 42576 10396
rect 4160 9732 4212 9784
rect 7104 9732 7156 9784
rect 7472 9732 7524 9784
rect 9312 9732 9364 9784
rect 9496 9732 9548 9784
rect 13452 9732 13504 9784
rect 13636 9732 13688 9784
rect 14556 9732 14608 9784
rect 16304 9732 16356 9784
rect 17592 9732 17644 9784
rect 17684 9732 17736 9784
rect 19524 9732 19576 9784
rect 19616 9732 19668 9784
rect 6736 9664 6788 9716
rect 7380 9664 7432 9716
rect 8576 9664 8628 9716
rect 11244 9664 11296 9716
rect 13176 9664 13228 9716
rect 13820 9664 13872 9716
rect 16028 9664 16080 9716
rect 17316 9664 17368 9716
rect 19156 9664 19208 9716
rect 20628 9664 20680 9716
rect 21180 9664 21232 9716
rect 22100 9664 22152 9716
rect 23388 9664 23440 9716
rect 23664 9664 23716 9716
rect 23940 9664 23992 9716
rect 25504 9664 25556 9716
rect 25596 9664 25648 9716
rect 26516 9664 26568 9716
rect 26976 9732 27028 9784
rect 27988 9732 28040 9784
rect 28080 9732 28132 9784
rect 29092 9732 29144 9784
rect 39120 9732 39172 9784
rect 41696 9732 41748 9784
rect 5908 9596 5960 9648
rect 15844 9596 15896 9648
rect 16488 9596 16540 9648
rect 27528 9664 27580 9716
rect 29184 9664 29236 9716
rect 32312 9664 32364 9716
rect 32496 9664 32548 9716
rect 33692 9664 33744 9716
rect 34152 9664 34204 9716
rect 35624 9664 35676 9716
rect 37188 9664 37240 9716
rect 39304 9664 39356 9716
rect 39396 9664 39448 9716
rect 40316 9664 40368 9716
rect 5264 9528 5316 9580
rect 8484 9528 8536 9580
rect 15752 9528 15804 9580
rect 28632 9596 28684 9648
rect 31668 9596 31720 9648
rect 35440 9596 35492 9648
rect 39856 9596 39908 9648
rect 4528 9460 4580 9512
rect 13728 9460 13780 9512
rect 16396 9460 16448 9512
rect 26792 9460 26844 9512
rect 29736 9528 29788 9580
rect 31208 9460 31260 9512
rect 7012 9392 7064 9444
rect 23296 9392 23348 9444
rect 7288 9324 7340 9376
rect 17960 9324 18012 9376
rect 21272 9324 21324 9376
rect 27436 9392 27488 9444
rect 31392 9392 31444 9444
rect 32588 9392 32640 9444
rect 23848 9324 23900 9376
rect 43628 9324 43680 9376
rect 4344 9256 4396 9308
rect 15568 9256 15620 9308
rect 18144 9256 18196 9308
rect 40500 9256 40552 9308
rect 4712 9188 4764 9240
rect 6920 9188 6972 9240
rect 11888 9188 11940 9240
rect 34152 9188 34204 9240
rect 5632 9120 5684 9172
rect 3516 9052 3568 9104
rect 5724 9052 5776 9104
rect 6184 9052 6236 9104
rect 10968 9052 11020 9104
rect 11612 9052 11664 9104
rect 16212 9120 16264 9172
rect 35900 9120 35952 9172
rect 7104 8984 7156 9036
rect 18512 9052 18564 9104
rect 19616 9052 19668 9104
rect 6092 8916 6144 8968
rect 11152 8916 11204 8968
rect 4896 8848 4948 8900
rect 8208 8848 8260 8900
rect 19432 8984 19484 9036
rect 13912 8916 13964 8968
rect 20536 8916 20588 8968
rect 26792 9052 26844 9104
rect 29000 9052 29052 9104
rect 30656 9052 30708 9104
rect 35808 9052 35860 9104
rect 26884 8984 26936 9036
rect 41144 8984 41196 9036
rect 29828 8916 29880 8968
rect 31668 8916 31720 8968
rect 32128 8916 32180 8968
rect 39580 8916 39632 8968
rect 42616 8916 42668 8968
rect 17500 8848 17552 8900
rect 21916 8848 21968 8900
rect 23664 8848 23716 8900
rect 24124 8848 24176 8900
rect 34244 8848 34296 8900
rect 35716 8848 35768 8900
rect 42984 8848 43036 8900
rect 3240 8780 3292 8832
rect 4804 8780 4856 8832
rect 8484 8780 8536 8832
rect 8668 8780 8720 8832
rect 9864 8780 9916 8832
rect 11336 8780 11388 8832
rect 12532 8780 12584 8832
rect 14096 8780 14148 8832
rect 15292 8780 15344 8832
rect 19524 8780 19576 8832
rect 22744 8780 22796 8832
rect 28816 8780 28868 8832
rect 30472 8780 30524 8832
rect 42708 8780 42760 8832
rect 2658 8678 2710 8730
rect 2722 8678 2774 8730
rect 2786 8678 2838 8730
rect 2850 8678 2902 8730
rect 2914 8678 2966 8730
rect 2978 8678 3030 8730
rect 8658 8678 8710 8730
rect 8722 8678 8774 8730
rect 8786 8678 8838 8730
rect 8850 8678 8902 8730
rect 8914 8678 8966 8730
rect 8978 8678 9030 8730
rect 14658 8678 14710 8730
rect 14722 8678 14774 8730
rect 14786 8678 14838 8730
rect 14850 8678 14902 8730
rect 14914 8678 14966 8730
rect 14978 8678 15030 8730
rect 20658 8678 20710 8730
rect 20722 8678 20774 8730
rect 20786 8678 20838 8730
rect 20850 8678 20902 8730
rect 20914 8678 20966 8730
rect 20978 8678 21030 8730
rect 26658 8678 26710 8730
rect 26722 8678 26774 8730
rect 26786 8678 26838 8730
rect 26850 8678 26902 8730
rect 26914 8678 26966 8730
rect 26978 8678 27030 8730
rect 32658 8678 32710 8730
rect 32722 8678 32774 8730
rect 32786 8678 32838 8730
rect 32850 8678 32902 8730
rect 32914 8678 32966 8730
rect 32978 8678 33030 8730
rect 38658 8678 38710 8730
rect 38722 8678 38774 8730
rect 38786 8678 38838 8730
rect 38850 8678 38902 8730
rect 38914 8678 38966 8730
rect 38978 8678 39030 8730
rect 6276 8576 6328 8628
rect 6644 8576 6696 8628
rect 6000 8508 6052 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5632 8440 5684 8492
rect 6092 8440 6144 8492
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 14372 8576 14424 8628
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 15108 8576 15160 8628
rect 15384 8576 15436 8628
rect 16028 8619 16080 8628
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 16304 8619 16356 8628
rect 16304 8585 16313 8619
rect 16313 8585 16347 8619
rect 16347 8585 16356 8619
rect 16304 8576 16356 8585
rect 16764 8576 16816 8628
rect 17592 8576 17644 8628
rect 17868 8576 17920 8628
rect 18420 8576 18472 8628
rect 19432 8576 19484 8628
rect 24124 8576 24176 8628
rect 24860 8576 24912 8628
rect 7104 8508 7156 8560
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7564 8440 7616 8492
rect 3332 8372 3384 8424
rect 3516 8304 3568 8356
rect 4160 8279 4212 8288
rect 4160 8245 4169 8279
rect 4169 8245 4203 8279
rect 4203 8245 4212 8279
rect 4160 8236 4212 8245
rect 5540 8304 5592 8356
rect 5816 8304 5868 8356
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 6092 8236 6144 8288
rect 6828 8236 6880 8288
rect 7196 8304 7248 8356
rect 7380 8304 7432 8356
rect 7656 8304 7708 8356
rect 7840 8372 7892 8424
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8300 8372 8352 8424
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 10784 8508 10836 8560
rect 13728 8508 13780 8560
rect 9312 8440 9364 8449
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11152 8440 11204 8492
rect 10600 8372 10652 8424
rect 8116 8304 8168 8356
rect 9128 8304 9180 8356
rect 9496 8304 9548 8356
rect 9956 8347 10008 8356
rect 9956 8313 9965 8347
rect 9965 8313 9999 8347
rect 9999 8313 10008 8347
rect 9956 8304 10008 8313
rect 10232 8347 10284 8356
rect 10232 8313 10241 8347
rect 10241 8313 10275 8347
rect 10275 8313 10284 8347
rect 10232 8304 10284 8313
rect 10876 8372 10928 8424
rect 11428 8372 11480 8424
rect 11060 8304 11112 8356
rect 8852 8236 8904 8288
rect 11152 8236 11204 8288
rect 11336 8236 11388 8288
rect 13452 8440 13504 8492
rect 14372 8440 14424 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 18604 8508 18656 8560
rect 12808 8304 12860 8356
rect 12716 8236 12768 8288
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 17592 8440 17644 8492
rect 17868 8440 17920 8492
rect 18144 8483 18196 8492
rect 18144 8449 18153 8483
rect 18153 8449 18187 8483
rect 18187 8449 18196 8483
rect 18144 8440 18196 8449
rect 19432 8440 19484 8492
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 20076 8440 20128 8492
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 14648 8304 14700 8356
rect 15292 8304 15344 8356
rect 17040 8304 17092 8356
rect 17776 8304 17828 8356
rect 18788 8304 18840 8356
rect 19248 8304 19300 8356
rect 13728 8236 13780 8288
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 14464 8236 14516 8288
rect 17592 8236 17644 8288
rect 18328 8236 18380 8288
rect 18880 8236 18932 8288
rect 20720 8372 20772 8424
rect 21732 8372 21784 8424
rect 19616 8304 19668 8356
rect 23112 8508 23164 8560
rect 24032 8508 24084 8560
rect 24768 8508 24820 8560
rect 26240 8508 26292 8560
rect 22836 8440 22888 8492
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 24308 8440 24360 8492
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 25504 8483 25556 8492
rect 25504 8449 25513 8483
rect 25513 8449 25547 8483
rect 25547 8449 25556 8483
rect 25504 8440 25556 8449
rect 25964 8440 26016 8492
rect 27344 8576 27396 8628
rect 29000 8551 29052 8560
rect 29000 8517 29009 8551
rect 29009 8517 29043 8551
rect 29043 8517 29052 8551
rect 29000 8508 29052 8517
rect 29184 8551 29236 8560
rect 29184 8517 29193 8551
rect 29193 8517 29227 8551
rect 29227 8517 29236 8551
rect 29184 8508 29236 8517
rect 28264 8440 28316 8492
rect 22652 8372 22704 8424
rect 24400 8415 24452 8424
rect 24400 8381 24409 8415
rect 24409 8381 24443 8415
rect 24443 8381 24452 8415
rect 24400 8372 24452 8381
rect 25228 8372 25280 8424
rect 27344 8372 27396 8424
rect 27712 8372 27764 8424
rect 29000 8372 29052 8424
rect 29920 8440 29972 8492
rect 30104 8440 30156 8492
rect 23112 8304 23164 8356
rect 23204 8304 23256 8356
rect 19708 8236 19760 8288
rect 22008 8236 22060 8288
rect 22836 8236 22888 8288
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 26884 8304 26936 8356
rect 27252 8236 27304 8288
rect 29552 8304 29604 8356
rect 30748 8440 30800 8492
rect 32036 8508 32088 8560
rect 33140 8508 33192 8560
rect 31852 8440 31904 8492
rect 33324 8440 33376 8492
rect 33600 8508 33652 8560
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 34796 8440 34848 8492
rect 34888 8440 34940 8492
rect 35900 8483 35952 8492
rect 35900 8449 35909 8483
rect 35909 8449 35943 8483
rect 35943 8449 35952 8483
rect 35900 8440 35952 8449
rect 36820 8483 36872 8492
rect 36820 8449 36829 8483
rect 36829 8449 36863 8483
rect 36863 8449 36872 8483
rect 36820 8440 36872 8449
rect 36912 8483 36964 8492
rect 36912 8449 36921 8483
rect 36921 8449 36955 8483
rect 36955 8449 36964 8483
rect 36912 8440 36964 8449
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 38476 8483 38528 8492
rect 38476 8449 38485 8483
rect 38485 8449 38519 8483
rect 38519 8449 38528 8483
rect 38476 8440 38528 8449
rect 40224 8508 40276 8560
rect 39396 8440 39448 8492
rect 39580 8483 39632 8492
rect 39580 8449 39589 8483
rect 39589 8449 39623 8483
rect 39623 8449 39632 8483
rect 39580 8440 39632 8449
rect 41788 8508 41840 8560
rect 32956 8372 33008 8424
rect 33968 8372 34020 8424
rect 34980 8415 35032 8424
rect 34980 8381 34989 8415
rect 34989 8381 35023 8415
rect 35023 8381 35032 8415
rect 34980 8372 35032 8381
rect 35072 8372 35124 8424
rect 33784 8304 33836 8356
rect 36636 8347 36688 8356
rect 36636 8313 36645 8347
rect 36645 8313 36679 8347
rect 36679 8313 36688 8347
rect 36636 8304 36688 8313
rect 38200 8304 38252 8356
rect 38660 8347 38712 8356
rect 38660 8313 38669 8347
rect 38669 8313 38703 8347
rect 38703 8313 38712 8347
rect 38660 8304 38712 8313
rect 39120 8347 39172 8356
rect 39120 8313 39129 8347
rect 39129 8313 39163 8347
rect 39163 8313 39172 8347
rect 39120 8304 39172 8313
rect 39304 8304 39356 8356
rect 39948 8347 40000 8356
rect 39948 8313 39957 8347
rect 39957 8313 39991 8347
rect 39991 8313 40000 8347
rect 39948 8304 40000 8313
rect 40040 8304 40092 8356
rect 41420 8440 41472 8492
rect 41604 8483 41656 8492
rect 41604 8449 41613 8483
rect 41613 8449 41647 8483
rect 41647 8449 41656 8483
rect 41604 8440 41656 8449
rect 42800 8576 42852 8628
rect 43444 8619 43496 8628
rect 43444 8585 43453 8619
rect 43453 8585 43487 8619
rect 43487 8585 43496 8619
rect 43444 8576 43496 8585
rect 42708 8440 42760 8492
rect 42984 8440 43036 8492
rect 41512 8372 41564 8424
rect 41328 8304 41380 8356
rect 41696 8304 41748 8356
rect 43076 8347 43128 8356
rect 43076 8313 43085 8347
rect 43085 8313 43119 8347
rect 43119 8313 43128 8347
rect 43076 8304 43128 8313
rect 30656 8236 30708 8288
rect 30748 8279 30800 8288
rect 30748 8245 30757 8279
rect 30757 8245 30791 8279
rect 30791 8245 30800 8279
rect 30748 8236 30800 8245
rect 30840 8236 30892 8288
rect 31760 8279 31812 8288
rect 31760 8245 31769 8279
rect 31769 8245 31803 8279
rect 31803 8245 31812 8279
rect 31760 8236 31812 8245
rect 33048 8236 33100 8288
rect 36912 8236 36964 8288
rect 40684 8279 40736 8288
rect 40684 8245 40693 8279
rect 40693 8245 40727 8279
rect 40727 8245 40736 8279
rect 40684 8236 40736 8245
rect 41052 8279 41104 8288
rect 41052 8245 41061 8279
rect 41061 8245 41095 8279
rect 41095 8245 41104 8279
rect 41052 8236 41104 8245
rect 41144 8236 41196 8288
rect 42432 8236 42484 8288
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 13918 8134 13970 8186
rect 13982 8134 14034 8186
rect 14046 8134 14098 8186
rect 14110 8134 14162 8186
rect 14174 8134 14226 8186
rect 14238 8134 14290 8186
rect 19918 8134 19970 8186
rect 19982 8134 20034 8186
rect 20046 8134 20098 8186
rect 20110 8134 20162 8186
rect 20174 8134 20226 8186
rect 20238 8134 20290 8186
rect 25918 8134 25970 8186
rect 25982 8134 26034 8186
rect 26046 8134 26098 8186
rect 26110 8134 26162 8186
rect 26174 8134 26226 8186
rect 26238 8134 26290 8186
rect 31918 8134 31970 8186
rect 31982 8134 32034 8186
rect 32046 8134 32098 8186
rect 32110 8134 32162 8186
rect 32174 8134 32226 8186
rect 32238 8134 32290 8186
rect 37918 8134 37970 8186
rect 37982 8134 38034 8186
rect 38046 8134 38098 8186
rect 38110 8134 38162 8186
rect 38174 8134 38226 8186
rect 38238 8134 38290 8186
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 5448 8032 5500 8084
rect 6092 8075 6144 8084
rect 6092 8041 6101 8075
rect 6101 8041 6135 8075
rect 6135 8041 6144 8075
rect 6092 8032 6144 8041
rect 6460 8075 6512 8084
rect 6460 8041 6469 8075
rect 6469 8041 6503 8075
rect 6503 8041 6512 8075
rect 6460 8032 6512 8041
rect 4068 7964 4120 8016
rect 5632 7964 5684 8016
rect 5724 7964 5776 8016
rect 7748 8032 7800 8084
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 8760 8032 8812 8084
rect 10324 8032 10376 8084
rect 10508 8032 10560 8084
rect 8852 7964 8904 8016
rect 3792 7896 3844 7948
rect 3884 7896 3936 7948
rect 1492 7871 1544 7880
rect 1492 7837 1501 7871
rect 1501 7837 1535 7871
rect 1535 7837 1544 7871
rect 1492 7828 1544 7837
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2320 7828 2372 7880
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 6092 7896 6144 7948
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 4344 7828 4396 7880
rect 4712 7828 4764 7880
rect 6368 7896 6420 7948
rect 1676 7760 1728 7812
rect 2412 7803 2464 7812
rect 2412 7769 2421 7803
rect 2421 7769 2455 7803
rect 2455 7769 2464 7803
rect 2412 7760 2464 7769
rect 3332 7760 3384 7812
rect 3424 7803 3476 7812
rect 3424 7769 3433 7803
rect 3433 7769 3467 7803
rect 3467 7769 3476 7803
rect 3424 7760 3476 7769
rect 5448 7760 5500 7812
rect 8944 7939 8996 7948
rect 6552 7828 6604 7880
rect 7012 7871 7064 7880
rect 7012 7837 7042 7871
rect 7042 7837 7064 7871
rect 7012 7828 7064 7837
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 14464 7896 14516 7948
rect 8484 7828 8536 7880
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 9128 7828 9180 7880
rect 5172 7692 5224 7744
rect 5264 7692 5316 7744
rect 7656 7760 7708 7812
rect 6276 7692 6328 7744
rect 6460 7692 6512 7744
rect 7012 7692 7064 7744
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8300 7692 8352 7744
rect 8576 7692 8628 7744
rect 10140 7692 10192 7744
rect 12072 7760 12124 7812
rect 12256 7871 12308 7880
rect 12256 7837 12290 7871
rect 12290 7837 12308 7871
rect 12256 7828 12308 7837
rect 12624 7828 12676 7880
rect 12808 7692 12860 7744
rect 13268 7760 13320 7812
rect 14096 7828 14148 7880
rect 14832 7871 14884 7880
rect 14832 7837 14841 7871
rect 14841 7837 14875 7871
rect 14875 7837 14884 7871
rect 14832 7828 14884 7837
rect 15108 7871 15160 7880
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 15660 8032 15712 8084
rect 17408 8032 17460 8084
rect 18420 8032 18472 8084
rect 18696 8032 18748 8084
rect 18972 8032 19024 8084
rect 19524 8032 19576 8084
rect 21916 8032 21968 8084
rect 22560 8032 22612 8084
rect 16764 7964 16816 8016
rect 17868 8007 17920 8016
rect 17868 7973 17877 8007
rect 17877 7973 17911 8007
rect 17911 7973 17920 8007
rect 17868 7964 17920 7973
rect 15384 7896 15436 7948
rect 22192 8007 22244 8016
rect 22192 7973 22201 8007
rect 22201 7973 22235 8007
rect 22235 7973 22244 8007
rect 22192 7964 22244 7973
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 15844 7871 15896 7880
rect 15844 7837 15874 7871
rect 15874 7837 15896 7871
rect 15844 7828 15896 7837
rect 13452 7692 13504 7744
rect 13912 7692 13964 7744
rect 18604 7896 18656 7948
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17408 7828 17460 7880
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 18972 7828 19024 7880
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 19432 7896 19484 7948
rect 19524 7896 19576 7948
rect 19708 7828 19760 7880
rect 21088 7896 21140 7948
rect 21180 7828 21232 7880
rect 21640 7828 21692 7880
rect 21916 7871 21968 7880
rect 21916 7837 21925 7871
rect 21925 7837 21959 7871
rect 21959 7837 21968 7871
rect 21916 7828 21968 7837
rect 22928 7871 22980 7880
rect 22928 7837 22937 7871
rect 22937 7837 22971 7871
rect 22971 7837 22980 7871
rect 22928 7828 22980 7837
rect 23204 7871 23256 7880
rect 23204 7837 23213 7871
rect 23213 7837 23247 7871
rect 23247 7837 23256 7871
rect 23204 7828 23256 7837
rect 23480 7828 23532 7880
rect 18420 7760 18472 7812
rect 24492 7896 24544 7948
rect 25412 7964 25464 8016
rect 26792 7896 26844 7948
rect 29920 8032 29972 8084
rect 32588 8032 32640 8084
rect 34336 8075 34388 8084
rect 34336 8041 34345 8075
rect 34345 8041 34379 8075
rect 34379 8041 34388 8075
rect 34336 8032 34388 8041
rect 34520 8032 34572 8084
rect 30748 7964 30800 8016
rect 25044 7871 25096 7880
rect 25044 7837 25053 7871
rect 25053 7837 25087 7871
rect 25087 7837 25096 7871
rect 25044 7828 25096 7837
rect 25412 7828 25464 7880
rect 25964 7871 26016 7880
rect 25964 7837 25973 7871
rect 25973 7837 26007 7871
rect 26007 7837 26016 7871
rect 25964 7828 26016 7837
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 26240 7828 26292 7837
rect 27620 7828 27672 7880
rect 27712 7828 27764 7880
rect 28172 7871 28224 7880
rect 28172 7837 28181 7871
rect 28181 7837 28215 7871
rect 28215 7837 28224 7871
rect 28172 7828 28224 7837
rect 24216 7760 24268 7812
rect 24584 7760 24636 7812
rect 29184 7803 29236 7812
rect 29184 7769 29193 7803
rect 29193 7769 29227 7803
rect 29227 7769 29236 7803
rect 29184 7760 29236 7769
rect 17408 7692 17460 7744
rect 17592 7692 17644 7744
rect 18696 7692 18748 7744
rect 19800 7692 19852 7744
rect 19984 7692 20036 7744
rect 20444 7692 20496 7744
rect 27068 7692 27120 7744
rect 29000 7692 29052 7744
rect 29368 7692 29420 7744
rect 29460 7692 29512 7744
rect 30932 7939 30984 7948
rect 30932 7905 30941 7939
rect 30941 7905 30975 7939
rect 30975 7905 30984 7939
rect 30932 7896 30984 7905
rect 34704 7964 34756 8016
rect 32956 7939 33008 7948
rect 32956 7905 32965 7939
rect 32965 7905 32999 7939
rect 32999 7905 33008 7939
rect 32956 7896 33008 7905
rect 37464 8032 37516 8084
rect 37556 8075 37608 8084
rect 37556 8041 37565 8075
rect 37565 8041 37599 8075
rect 37599 8041 37608 8075
rect 37556 8032 37608 8041
rect 37832 8032 37884 8084
rect 39212 8032 39264 8084
rect 39764 8032 39816 8084
rect 40132 8032 40184 8084
rect 41512 8075 41564 8084
rect 41512 8041 41521 8075
rect 41521 8041 41555 8075
rect 41555 8041 41564 8075
rect 41512 8032 41564 8041
rect 43168 8032 43220 8084
rect 37188 7964 37240 8016
rect 39488 7964 39540 8016
rect 41328 7964 41380 8016
rect 41696 7964 41748 8016
rect 30196 7871 30248 7880
rect 30196 7837 30205 7871
rect 30205 7837 30239 7871
rect 30239 7837 30248 7871
rect 30196 7828 30248 7837
rect 31024 7871 31076 7880
rect 31024 7837 31058 7871
rect 31058 7837 31076 7871
rect 31024 7828 31076 7837
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 33048 7871 33100 7880
rect 33048 7837 33057 7871
rect 33057 7837 33091 7871
rect 33091 7837 33100 7871
rect 33048 7828 33100 7837
rect 33324 7871 33376 7880
rect 33324 7837 33333 7871
rect 33333 7837 33367 7871
rect 33367 7837 33376 7871
rect 33324 7828 33376 7837
rect 33416 7828 33468 7880
rect 43352 7964 43404 8016
rect 34796 7828 34848 7880
rect 35164 7828 35216 7880
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 35716 7871 35768 7880
rect 35716 7837 35725 7871
rect 35725 7837 35759 7871
rect 35759 7837 35768 7871
rect 35716 7828 35768 7837
rect 36452 7871 36504 7880
rect 36452 7837 36461 7871
rect 36461 7837 36495 7871
rect 36495 7837 36504 7871
rect 36452 7828 36504 7837
rect 36544 7871 36596 7880
rect 36544 7837 36578 7871
rect 36578 7837 36596 7871
rect 36544 7828 36596 7837
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 37832 7828 37884 7880
rect 32036 7760 32088 7812
rect 32128 7760 32180 7812
rect 35440 7760 35492 7812
rect 32312 7692 32364 7744
rect 32680 7692 32732 7744
rect 33324 7692 33376 7744
rect 33876 7692 33928 7744
rect 34152 7692 34204 7744
rect 36452 7692 36504 7744
rect 39120 7828 39172 7880
rect 39304 7760 39356 7812
rect 39212 7692 39264 7744
rect 43536 7896 43588 7948
rect 39672 7828 39724 7880
rect 40132 7871 40184 7880
rect 40132 7837 40141 7871
rect 40141 7837 40175 7871
rect 40175 7837 40184 7871
rect 40132 7828 40184 7837
rect 41512 7828 41564 7880
rect 40408 7760 40460 7812
rect 41880 7828 41932 7880
rect 42156 7871 42208 7880
rect 42156 7837 42165 7871
rect 42165 7837 42199 7871
rect 42199 7837 42208 7871
rect 42156 7828 42208 7837
rect 42524 7871 42576 7880
rect 42524 7837 42533 7871
rect 42533 7837 42567 7871
rect 42567 7837 42576 7871
rect 42524 7828 42576 7837
rect 42984 7828 43036 7880
rect 42800 7760 42852 7812
rect 42156 7692 42208 7744
rect 43076 7735 43128 7744
rect 43076 7701 43085 7735
rect 43085 7701 43119 7735
rect 43119 7701 43128 7735
rect 43076 7692 43128 7701
rect 43444 7735 43496 7744
rect 43444 7701 43453 7735
rect 43453 7701 43487 7735
rect 43487 7701 43496 7735
rect 43444 7692 43496 7701
rect 2658 7590 2710 7642
rect 2722 7590 2774 7642
rect 2786 7590 2838 7642
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 8658 7590 8710 7642
rect 8722 7590 8774 7642
rect 8786 7590 8838 7642
rect 8850 7590 8902 7642
rect 8914 7590 8966 7642
rect 8978 7590 9030 7642
rect 14658 7590 14710 7642
rect 14722 7590 14774 7642
rect 14786 7590 14838 7642
rect 14850 7590 14902 7642
rect 14914 7590 14966 7642
rect 14978 7590 15030 7642
rect 20658 7590 20710 7642
rect 20722 7590 20774 7642
rect 20786 7590 20838 7642
rect 20850 7590 20902 7642
rect 20914 7590 20966 7642
rect 20978 7590 21030 7642
rect 26658 7590 26710 7642
rect 26722 7590 26774 7642
rect 26786 7590 26838 7642
rect 26850 7590 26902 7642
rect 26914 7590 26966 7642
rect 26978 7590 27030 7642
rect 32658 7590 32710 7642
rect 32722 7590 32774 7642
rect 32786 7590 32838 7642
rect 32850 7590 32902 7642
rect 32914 7590 32966 7642
rect 32978 7590 33030 7642
rect 38658 7590 38710 7642
rect 38722 7590 38774 7642
rect 38786 7590 38838 7642
rect 38850 7590 38902 7642
rect 38914 7590 38966 7642
rect 38978 7590 39030 7642
rect 2044 7488 2096 7540
rect 3056 7420 3108 7472
rect 3148 7463 3200 7472
rect 3148 7429 3157 7463
rect 3157 7429 3191 7463
rect 3191 7429 3200 7463
rect 3148 7420 3200 7429
rect 6736 7531 6788 7540
rect 6736 7497 6745 7531
rect 6745 7497 6779 7531
rect 6779 7497 6788 7531
rect 6736 7488 6788 7497
rect 7840 7488 7892 7540
rect 8208 7488 8260 7540
rect 9312 7488 9364 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 12808 7488 12860 7540
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 3240 7352 3292 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 1768 7284 1820 7336
rect 1308 7216 1360 7268
rect 5356 7352 5408 7404
rect 4160 7284 4212 7336
rect 5724 7352 5776 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 5540 7284 5592 7336
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6460 7284 6512 7336
rect 7012 7352 7064 7404
rect 7196 7352 7248 7404
rect 7472 7352 7524 7404
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 5080 7148 5132 7200
rect 7288 7216 7340 7268
rect 7748 7284 7800 7336
rect 9128 7352 9180 7404
rect 9312 7352 9364 7404
rect 9588 7352 9640 7404
rect 9680 7352 9732 7404
rect 8300 7284 8352 7336
rect 9220 7284 9272 7336
rect 10232 7352 10284 7404
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 11060 7352 11112 7404
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 10692 7284 10744 7336
rect 6828 7148 6880 7200
rect 9680 7148 9732 7200
rect 9772 7148 9824 7200
rect 10048 7148 10100 7200
rect 11980 7352 12032 7404
rect 12808 7284 12860 7336
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 14096 7420 14148 7472
rect 15660 7420 15712 7472
rect 14924 7352 14976 7404
rect 15936 7488 15988 7540
rect 17316 7488 17368 7540
rect 18420 7488 18472 7540
rect 18696 7488 18748 7540
rect 19708 7531 19760 7540
rect 19708 7497 19717 7531
rect 19717 7497 19751 7531
rect 19751 7497 19760 7531
rect 19708 7488 19760 7497
rect 15844 7420 15896 7472
rect 16396 7352 16448 7404
rect 16580 7352 16632 7404
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 17960 7352 18012 7404
rect 13544 7148 13596 7200
rect 13728 7148 13780 7200
rect 15752 7284 15804 7336
rect 17776 7327 17828 7336
rect 17776 7293 17785 7327
rect 17785 7293 17819 7327
rect 17819 7293 17828 7327
rect 17776 7284 17828 7293
rect 19800 7420 19852 7472
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 20444 7352 20496 7404
rect 24124 7488 24176 7540
rect 24400 7488 24452 7540
rect 26240 7488 26292 7540
rect 22652 7420 22704 7472
rect 23204 7420 23256 7472
rect 15844 7148 15896 7200
rect 16672 7216 16724 7268
rect 20996 7284 21048 7336
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 19708 7148 19760 7200
rect 20444 7148 20496 7200
rect 20536 7148 20588 7200
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 22008 7284 22060 7336
rect 23572 7395 23624 7404
rect 23572 7361 23581 7395
rect 23581 7361 23615 7395
rect 23615 7361 23624 7395
rect 23572 7352 23624 7361
rect 24032 7395 24084 7404
rect 24032 7361 24066 7395
rect 24066 7361 24084 7395
rect 24032 7352 24084 7361
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24492 7420 24544 7472
rect 26424 7420 26476 7472
rect 27068 7488 27120 7540
rect 27252 7420 27304 7472
rect 27988 7420 28040 7472
rect 26332 7352 26384 7404
rect 22744 7284 22796 7336
rect 22376 7216 22428 7268
rect 23848 7216 23900 7268
rect 23940 7148 23992 7200
rect 24216 7148 24268 7200
rect 29552 7395 29604 7404
rect 29552 7361 29561 7395
rect 29561 7361 29595 7395
rect 29595 7361 29604 7395
rect 29552 7352 29604 7361
rect 30380 7395 30432 7404
rect 30380 7361 30389 7395
rect 30389 7361 30423 7395
rect 30423 7361 30432 7395
rect 30380 7352 30432 7361
rect 25320 7148 25372 7200
rect 25504 7148 25556 7200
rect 27620 7284 27672 7336
rect 28356 7327 28408 7336
rect 28356 7293 28365 7327
rect 28365 7293 28399 7327
rect 28399 7293 28408 7327
rect 28356 7284 28408 7293
rect 28540 7327 28592 7336
rect 28540 7293 28549 7327
rect 28549 7293 28583 7327
rect 28583 7293 28592 7327
rect 28540 7284 28592 7293
rect 29000 7327 29052 7336
rect 29000 7293 29009 7327
rect 29009 7293 29043 7327
rect 29043 7293 29052 7327
rect 29000 7284 29052 7293
rect 26516 7216 26568 7268
rect 29920 7284 29972 7336
rect 31024 7352 31076 7404
rect 26608 7148 26660 7200
rect 27620 7148 27672 7200
rect 27988 7191 28040 7200
rect 27988 7157 27997 7191
rect 27997 7157 28031 7191
rect 28031 7157 28040 7191
rect 27988 7148 28040 7157
rect 28172 7148 28224 7200
rect 29000 7148 29052 7200
rect 30748 7284 30800 7336
rect 31944 7488 31996 7540
rect 32036 7488 32088 7540
rect 31484 7395 31536 7404
rect 31484 7361 31493 7395
rect 31493 7361 31527 7395
rect 31527 7361 31536 7395
rect 31484 7352 31536 7361
rect 31576 7395 31628 7404
rect 31576 7361 31585 7395
rect 31585 7361 31619 7395
rect 31619 7361 31628 7395
rect 31576 7352 31628 7361
rect 31668 7352 31720 7404
rect 33048 7420 33100 7472
rect 32772 7352 32824 7404
rect 33324 7488 33376 7540
rect 35532 7488 35584 7540
rect 36728 7488 36780 7540
rect 37004 7488 37056 7540
rect 39304 7488 39356 7540
rect 30104 7216 30156 7268
rect 33048 7284 33100 7336
rect 30564 7148 30616 7200
rect 30932 7148 30984 7200
rect 32128 7148 32180 7200
rect 35256 7352 35308 7404
rect 33876 7327 33928 7336
rect 33876 7293 33885 7327
rect 33885 7293 33919 7327
rect 33919 7293 33928 7327
rect 33876 7284 33928 7293
rect 34152 7327 34204 7336
rect 34152 7293 34161 7327
rect 34161 7293 34195 7327
rect 34195 7293 34204 7327
rect 34152 7284 34204 7293
rect 34244 7327 34296 7336
rect 34244 7293 34278 7327
rect 34278 7293 34296 7327
rect 34244 7284 34296 7293
rect 34428 7327 34480 7336
rect 34428 7293 34437 7327
rect 34437 7293 34471 7327
rect 34471 7293 34480 7327
rect 34428 7284 34480 7293
rect 36268 7352 36320 7404
rect 38752 7352 38804 7404
rect 39304 7395 39356 7404
rect 39304 7361 39313 7395
rect 39313 7361 39347 7395
rect 39347 7361 39356 7395
rect 39304 7352 39356 7361
rect 39488 7352 39540 7404
rect 37280 7327 37332 7336
rect 37280 7293 37289 7327
rect 37289 7293 37323 7327
rect 37323 7293 37332 7327
rect 37280 7284 37332 7293
rect 38384 7327 38436 7336
rect 38384 7293 38393 7327
rect 38393 7293 38427 7327
rect 38427 7293 38436 7327
rect 38384 7284 38436 7293
rect 34888 7216 34940 7268
rect 36360 7216 36412 7268
rect 34428 7148 34480 7200
rect 35440 7148 35492 7200
rect 38660 7216 38712 7268
rect 39028 7259 39080 7268
rect 39028 7225 39037 7259
rect 39037 7225 39071 7259
rect 39071 7225 39080 7259
rect 39028 7216 39080 7225
rect 40316 7488 40368 7540
rect 40684 7531 40736 7540
rect 40684 7497 40693 7531
rect 40693 7497 40727 7531
rect 40727 7497 40736 7531
rect 40684 7488 40736 7497
rect 41788 7488 41840 7540
rect 42892 7488 42944 7540
rect 43260 7488 43312 7540
rect 42248 7395 42300 7404
rect 42248 7361 42257 7395
rect 42257 7361 42291 7395
rect 42291 7361 42300 7395
rect 42248 7352 42300 7361
rect 42432 7352 42484 7404
rect 42892 7395 42944 7404
rect 42892 7361 42901 7395
rect 42901 7361 42935 7395
rect 42935 7361 42944 7395
rect 42892 7352 42944 7361
rect 42340 7284 42392 7336
rect 41972 7216 42024 7268
rect 42064 7216 42116 7268
rect 43444 7191 43496 7200
rect 43444 7157 43453 7191
rect 43453 7157 43487 7191
rect 43487 7157 43496 7191
rect 43444 7148 43496 7157
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 13918 7046 13970 7098
rect 13982 7046 14034 7098
rect 14046 7046 14098 7098
rect 14110 7046 14162 7098
rect 14174 7046 14226 7098
rect 14238 7046 14290 7098
rect 19918 7046 19970 7098
rect 19982 7046 20034 7098
rect 20046 7046 20098 7098
rect 20110 7046 20162 7098
rect 20174 7046 20226 7098
rect 20238 7046 20290 7098
rect 25918 7046 25970 7098
rect 25982 7046 26034 7098
rect 26046 7046 26098 7098
rect 26110 7046 26162 7098
rect 26174 7046 26226 7098
rect 26238 7046 26290 7098
rect 31918 7046 31970 7098
rect 31982 7046 32034 7098
rect 32046 7046 32098 7098
rect 32110 7046 32162 7098
rect 32174 7046 32226 7098
rect 32238 7046 32290 7098
rect 37918 7046 37970 7098
rect 37982 7046 38034 7098
rect 38046 7046 38098 7098
rect 38110 7046 38162 7098
rect 38174 7046 38226 7098
rect 38238 7046 38290 7098
rect 6000 6944 6052 6996
rect 7840 6944 7892 6996
rect 10232 6944 10284 6996
rect 3976 6919 4028 6928
rect 3976 6885 3985 6919
rect 3985 6885 4019 6919
rect 4019 6885 4028 6919
rect 3976 6876 4028 6885
rect 4896 6876 4948 6928
rect 5080 6919 5132 6928
rect 5080 6885 5089 6919
rect 5089 6885 5123 6919
rect 5123 6885 5132 6919
rect 5080 6876 5132 6885
rect 10416 6944 10468 6996
rect 12624 6944 12676 6996
rect 13452 6987 13504 6996
rect 13452 6953 13461 6987
rect 13461 6953 13495 6987
rect 13495 6953 13504 6987
rect 13452 6944 13504 6953
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 4344 6808 4396 6860
rect 5172 6808 5224 6860
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 5540 6808 5592 6860
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 7288 6808 7340 6860
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 3056 6740 3108 6792
rect 3240 6740 3292 6792
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 2228 6672 2280 6724
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 4068 6672 4120 6724
rect 6828 6740 6880 6792
rect 8116 6740 8168 6792
rect 9312 6808 9364 6860
rect 12164 6876 12216 6928
rect 12716 6876 12768 6928
rect 19340 6944 19392 6996
rect 19432 6944 19484 6996
rect 27988 6944 28040 6996
rect 28356 6944 28408 6996
rect 30932 6944 30984 6996
rect 31024 6944 31076 6996
rect 32036 6944 32088 6996
rect 32220 6944 32272 6996
rect 32588 6944 32640 6996
rect 18512 6876 18564 6928
rect 19064 6876 19116 6928
rect 10232 6851 10284 6860
rect 10232 6817 10241 6851
rect 10241 6817 10275 6851
rect 10275 6817 10284 6851
rect 10232 6808 10284 6817
rect 10324 6808 10376 6860
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10508 6740 10560 6792
rect 10784 6740 10836 6792
rect 11152 6740 11204 6792
rect 11520 6740 11572 6792
rect 14188 6808 14240 6860
rect 14280 6740 14332 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 17684 6851 17736 6860
rect 17684 6817 17693 6851
rect 17693 6817 17727 6851
rect 17727 6817 17736 6851
rect 17684 6808 17736 6817
rect 14924 6783 14976 6792
rect 14924 6749 14933 6783
rect 14933 6749 14967 6783
rect 14967 6749 14976 6783
rect 14924 6740 14976 6749
rect 8300 6672 8352 6724
rect 6368 6604 6420 6656
rect 6460 6604 6512 6656
rect 7288 6604 7340 6656
rect 8208 6604 8260 6656
rect 9128 6604 9180 6656
rect 11060 6672 11112 6724
rect 16856 6740 16908 6792
rect 17316 6740 17368 6792
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 17960 6740 18012 6792
rect 18328 6672 18380 6724
rect 10232 6604 10284 6656
rect 12072 6604 12124 6656
rect 14740 6604 14792 6656
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 17316 6604 17368 6656
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 20996 6808 21048 6860
rect 19156 6740 19208 6792
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 19984 6740 20036 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 21364 6740 21416 6792
rect 22468 6851 22520 6860
rect 22468 6817 22477 6851
rect 22477 6817 22511 6851
rect 22511 6817 22520 6851
rect 22468 6808 22520 6817
rect 23112 6808 23164 6860
rect 24216 6808 24268 6860
rect 26240 6808 26292 6860
rect 27528 6851 27580 6860
rect 27528 6817 27537 6851
rect 27537 6817 27571 6851
rect 27571 6817 27580 6851
rect 27528 6808 27580 6817
rect 28632 6919 28684 6928
rect 28632 6885 28641 6919
rect 28641 6885 28675 6919
rect 28675 6885 28684 6919
rect 28632 6876 28684 6885
rect 29000 6876 29052 6928
rect 29368 6808 29420 6860
rect 31576 6876 31628 6928
rect 33048 6944 33100 6996
rect 33416 6944 33468 6996
rect 34244 6944 34296 6996
rect 34152 6876 34204 6928
rect 36544 6944 36596 6996
rect 37004 6944 37056 6996
rect 37464 6944 37516 6996
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 22744 6783 22796 6792
rect 22744 6749 22753 6783
rect 22753 6749 22787 6783
rect 22787 6749 22796 6783
rect 22744 6740 22796 6749
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 25504 6783 25556 6792
rect 25504 6749 25513 6783
rect 25513 6749 25547 6783
rect 25547 6749 25556 6783
rect 25504 6740 25556 6749
rect 25596 6740 25648 6792
rect 26424 6783 26476 6792
rect 26424 6749 26433 6783
rect 26433 6749 26467 6783
rect 26467 6749 26476 6783
rect 26424 6740 26476 6749
rect 26516 6783 26568 6792
rect 26516 6749 26550 6783
rect 26550 6749 26568 6783
rect 26516 6740 26568 6749
rect 26700 6783 26752 6792
rect 26700 6749 26709 6783
rect 26709 6749 26743 6783
rect 26743 6749 26752 6783
rect 26700 6740 26752 6749
rect 28080 6740 28132 6792
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 19340 6604 19392 6656
rect 23020 6672 23072 6724
rect 23112 6672 23164 6724
rect 19892 6604 19944 6656
rect 20168 6604 20220 6656
rect 20444 6604 20496 6656
rect 20536 6604 20588 6656
rect 21732 6604 21784 6656
rect 23204 6604 23256 6656
rect 23480 6647 23532 6656
rect 23480 6613 23489 6647
rect 23489 6613 23523 6647
rect 23523 6613 23532 6647
rect 23480 6604 23532 6613
rect 23664 6672 23716 6724
rect 23940 6604 23992 6656
rect 24952 6604 25004 6656
rect 26424 6604 26476 6656
rect 27804 6604 27856 6656
rect 29276 6740 29328 6792
rect 29644 6740 29696 6792
rect 30012 6783 30064 6792
rect 30012 6749 30021 6783
rect 30021 6749 30055 6783
rect 30055 6749 30064 6783
rect 30012 6740 30064 6749
rect 31392 6808 31444 6860
rect 30288 6740 30340 6792
rect 30380 6740 30432 6792
rect 30564 6783 30616 6792
rect 30564 6749 30573 6783
rect 30573 6749 30607 6783
rect 30607 6749 30616 6783
rect 30564 6740 30616 6749
rect 30840 6740 30892 6792
rect 30932 6783 30984 6792
rect 30932 6749 30941 6783
rect 30941 6749 30975 6783
rect 30975 6749 30984 6783
rect 30932 6740 30984 6749
rect 31300 6740 31352 6792
rect 32588 6851 32640 6860
rect 32588 6817 32597 6851
rect 32597 6817 32631 6851
rect 32631 6817 32640 6851
rect 32588 6808 32640 6817
rect 33692 6851 33744 6860
rect 33692 6817 33701 6851
rect 33701 6817 33735 6851
rect 33735 6817 33744 6851
rect 33692 6808 33744 6817
rect 29000 6672 29052 6724
rect 29184 6604 29236 6656
rect 29276 6604 29328 6656
rect 29552 6647 29604 6656
rect 29552 6613 29561 6647
rect 29561 6613 29595 6647
rect 29595 6613 29604 6647
rect 29552 6604 29604 6613
rect 31392 6672 31444 6724
rect 32312 6740 32364 6792
rect 32496 6783 32548 6792
rect 32496 6749 32505 6783
rect 32505 6749 32539 6783
rect 32539 6749 32548 6783
rect 32496 6740 32548 6749
rect 33232 6740 33284 6792
rect 34612 6808 34664 6860
rect 37556 6876 37608 6928
rect 36084 6851 36136 6860
rect 36084 6817 36093 6851
rect 36093 6817 36127 6851
rect 36127 6817 36136 6851
rect 36084 6808 36136 6817
rect 36544 6851 36596 6860
rect 36544 6817 36553 6851
rect 36553 6817 36587 6851
rect 36587 6817 36596 6851
rect 36544 6808 36596 6817
rect 36636 6808 36688 6860
rect 37004 6808 37056 6860
rect 37280 6808 37332 6860
rect 38568 6944 38620 6996
rect 39028 6944 39080 6996
rect 39212 6944 39264 6996
rect 41144 6944 41196 6996
rect 35808 6799 35860 6808
rect 35808 6765 35817 6799
rect 35817 6765 35851 6799
rect 35851 6765 35860 6799
rect 35808 6756 35860 6765
rect 37096 6783 37148 6792
rect 37096 6749 37105 6783
rect 37105 6749 37139 6783
rect 37139 6749 37148 6783
rect 37096 6740 37148 6749
rect 37740 6740 37792 6792
rect 38752 6808 38804 6860
rect 38568 6740 38620 6792
rect 30564 6604 30616 6656
rect 31484 6604 31536 6656
rect 33692 6672 33744 6724
rect 35072 6672 35124 6724
rect 35348 6672 35400 6724
rect 32312 6647 32364 6656
rect 32312 6613 32321 6647
rect 32321 6613 32355 6647
rect 32355 6613 32364 6647
rect 32312 6604 32364 6613
rect 32496 6604 32548 6656
rect 32680 6604 32732 6656
rect 33232 6604 33284 6656
rect 33508 6604 33560 6656
rect 34520 6604 34572 6656
rect 35256 6604 35308 6656
rect 35624 6647 35676 6656
rect 35624 6613 35633 6647
rect 35633 6613 35667 6647
rect 35667 6613 35676 6647
rect 35624 6604 35676 6613
rect 37648 6604 37700 6656
rect 38752 6604 38804 6656
rect 39856 6876 39908 6928
rect 42064 6944 42116 6996
rect 42340 6987 42392 6996
rect 42340 6953 42349 6987
rect 42349 6953 42383 6987
rect 42383 6953 42392 6987
rect 42340 6944 42392 6953
rect 39764 6808 39816 6860
rect 41880 6808 41932 6860
rect 41696 6740 41748 6792
rect 42708 6783 42760 6792
rect 42708 6749 42717 6783
rect 42717 6749 42751 6783
rect 42751 6749 42760 6783
rect 42708 6740 42760 6749
rect 40132 6604 40184 6656
rect 42984 6672 43036 6724
rect 43076 6715 43128 6724
rect 43076 6681 43085 6715
rect 43085 6681 43119 6715
rect 43119 6681 43128 6715
rect 43076 6672 43128 6681
rect 42800 6604 42852 6656
rect 42892 6647 42944 6656
rect 42892 6613 42901 6647
rect 42901 6613 42935 6647
rect 42935 6613 42944 6647
rect 42892 6604 42944 6613
rect 43444 6647 43496 6656
rect 43444 6613 43453 6647
rect 43453 6613 43487 6647
rect 43487 6613 43496 6647
rect 43444 6604 43496 6613
rect 2658 6502 2710 6554
rect 2722 6502 2774 6554
rect 2786 6502 2838 6554
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 8658 6502 8710 6554
rect 8722 6502 8774 6554
rect 8786 6502 8838 6554
rect 8850 6502 8902 6554
rect 8914 6502 8966 6554
rect 8978 6502 9030 6554
rect 14658 6502 14710 6554
rect 14722 6502 14774 6554
rect 14786 6502 14838 6554
rect 14850 6502 14902 6554
rect 14914 6502 14966 6554
rect 14978 6502 15030 6554
rect 20658 6502 20710 6554
rect 20722 6502 20774 6554
rect 20786 6502 20838 6554
rect 20850 6502 20902 6554
rect 20914 6502 20966 6554
rect 20978 6502 21030 6554
rect 26658 6502 26710 6554
rect 26722 6502 26774 6554
rect 26786 6502 26838 6554
rect 26850 6502 26902 6554
rect 26914 6502 26966 6554
rect 26978 6502 27030 6554
rect 32658 6502 32710 6554
rect 32722 6502 32774 6554
rect 32786 6502 32838 6554
rect 32850 6502 32902 6554
rect 32914 6502 32966 6554
rect 32978 6502 33030 6554
rect 38658 6502 38710 6554
rect 38722 6502 38774 6554
rect 38786 6502 38838 6554
rect 38850 6502 38902 6554
rect 38914 6502 38966 6554
rect 38978 6502 39030 6554
rect 2780 6400 2832 6452
rect 3424 6400 3476 6452
rect 3608 6400 3660 6452
rect 5816 6400 5868 6452
rect 5908 6400 5960 6452
rect 6644 6400 6696 6452
rect 6460 6332 6512 6384
rect 1676 6264 1728 6316
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 2964 6264 3016 6316
rect 2412 6196 2464 6248
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 3516 6239 3568 6282
rect 3516 6230 3525 6239
rect 3525 6230 3559 6239
rect 3559 6230 3568 6239
rect 3608 6307 3660 6316
rect 3608 6273 3642 6307
rect 3642 6273 3660 6307
rect 3608 6264 3660 6273
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 5724 6264 5776 6316
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 8760 6400 8812 6452
rect 9128 6400 9180 6452
rect 9220 6400 9272 6452
rect 9588 6400 9640 6452
rect 9956 6400 10008 6452
rect 10048 6400 10100 6452
rect 10508 6400 10560 6452
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 13636 6400 13688 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 10232 6332 10284 6384
rect 18880 6400 18932 6452
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 14280 6375 14332 6384
rect 14280 6341 14289 6375
rect 14289 6341 14323 6375
rect 14323 6341 14332 6375
rect 14280 6332 14332 6341
rect 14924 6332 14976 6384
rect 17040 6332 17092 6384
rect 17316 6332 17368 6384
rect 17684 6332 17736 6384
rect 17776 6332 17828 6384
rect 18052 6332 18104 6384
rect 18788 6375 18840 6384
rect 18788 6341 18797 6375
rect 18797 6341 18831 6375
rect 18831 6341 18840 6375
rect 18788 6332 18840 6341
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 5816 6196 5868 6248
rect 3056 6128 3108 6180
rect 4528 6128 4580 6180
rect 3332 6060 3384 6112
rect 6368 6060 6420 6112
rect 7840 6060 7892 6112
rect 8208 6239 8260 6248
rect 8208 6205 8217 6239
rect 8217 6205 8251 6239
rect 8251 6205 8260 6239
rect 8208 6196 8260 6205
rect 8300 6196 8352 6248
rect 8852 6239 8904 6248
rect 8852 6205 8861 6239
rect 8861 6205 8895 6239
rect 8895 6205 8904 6239
rect 8852 6196 8904 6205
rect 10692 6264 10744 6316
rect 11244 6264 11296 6316
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 13544 6264 13596 6316
rect 13820 6264 13872 6316
rect 14188 6264 14240 6316
rect 17592 6307 17644 6316
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 20352 6400 20404 6452
rect 20444 6400 20496 6452
rect 23664 6400 23716 6452
rect 23756 6443 23808 6452
rect 23756 6409 23765 6443
rect 23765 6409 23799 6443
rect 23799 6409 23808 6443
rect 23756 6400 23808 6409
rect 19524 6332 19576 6384
rect 19984 6332 20036 6384
rect 22928 6332 22980 6384
rect 24860 6332 24912 6384
rect 25044 6400 25096 6452
rect 26516 6400 26568 6452
rect 29920 6400 29972 6452
rect 31392 6400 31444 6452
rect 10048 6196 10100 6248
rect 11520 6196 11572 6248
rect 16948 6196 17000 6248
rect 8944 6060 8996 6112
rect 9220 6060 9272 6112
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 9864 6060 9916 6112
rect 11520 6060 11572 6112
rect 11796 6060 11848 6112
rect 12624 6060 12676 6112
rect 17316 6060 17368 6112
rect 17408 6060 17460 6112
rect 19616 6264 19668 6316
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 19800 6307 19852 6316
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 20720 6307 20772 6316
rect 20720 6273 20729 6307
rect 20729 6273 20763 6307
rect 20763 6273 20772 6307
rect 20720 6264 20772 6273
rect 21916 6264 21968 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 23480 6307 23532 6316
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 23756 6264 23808 6316
rect 23940 6307 23992 6316
rect 23940 6273 23949 6307
rect 23949 6273 23983 6307
rect 23983 6273 23992 6307
rect 23940 6264 23992 6273
rect 24124 6307 24176 6316
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 18328 6196 18380 6248
rect 18788 6128 18840 6180
rect 19156 6196 19208 6248
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 20352 6196 20404 6248
rect 20904 6196 20956 6248
rect 21180 6196 21232 6248
rect 21640 6196 21692 6248
rect 22744 6196 22796 6248
rect 24676 6264 24728 6316
rect 27160 6332 27212 6384
rect 27528 6332 27580 6384
rect 26424 6264 26476 6316
rect 27436 6264 27488 6316
rect 27620 6264 27672 6316
rect 27988 6307 28040 6316
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 28172 6307 28224 6316
rect 28172 6273 28181 6307
rect 28181 6273 28215 6307
rect 28215 6273 28224 6307
rect 28172 6264 28224 6273
rect 28356 6307 28408 6316
rect 28356 6273 28365 6307
rect 28365 6273 28399 6307
rect 28399 6273 28408 6307
rect 28356 6264 28408 6273
rect 29368 6307 29420 6316
rect 29368 6273 29377 6307
rect 29377 6273 29411 6307
rect 29411 6273 29420 6307
rect 29368 6264 29420 6273
rect 24400 6196 24452 6248
rect 25136 6239 25188 6248
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 18696 6060 18748 6112
rect 19616 6060 19668 6112
rect 19984 6060 20036 6112
rect 20720 6060 20772 6112
rect 22192 6128 22244 6180
rect 23664 6128 23716 6180
rect 26976 6196 27028 6248
rect 30748 6332 30800 6384
rect 31576 6332 31628 6384
rect 30288 6264 30340 6316
rect 30656 6264 30708 6316
rect 31300 6264 31352 6316
rect 31668 6264 31720 6316
rect 31760 6307 31812 6316
rect 31760 6273 31769 6307
rect 31769 6273 31803 6307
rect 31803 6273 31812 6307
rect 31760 6264 31812 6273
rect 31852 6264 31904 6316
rect 32772 6332 32824 6384
rect 37096 6400 37148 6452
rect 37188 6400 37240 6452
rect 39764 6400 39816 6452
rect 40500 6443 40552 6452
rect 40500 6409 40509 6443
rect 40509 6409 40543 6443
rect 40543 6409 40552 6443
rect 40500 6400 40552 6409
rect 42616 6443 42668 6452
rect 42616 6409 42625 6443
rect 42625 6409 42659 6443
rect 42659 6409 42668 6443
rect 42616 6400 42668 6409
rect 43444 6443 43496 6452
rect 43444 6409 43453 6443
rect 43453 6409 43487 6443
rect 43487 6409 43496 6443
rect 43444 6400 43496 6409
rect 21640 6103 21692 6112
rect 21640 6069 21649 6103
rect 21649 6069 21683 6103
rect 21683 6069 21692 6103
rect 21640 6060 21692 6069
rect 21916 6060 21968 6112
rect 22928 6060 22980 6112
rect 23020 6060 23072 6112
rect 26332 6060 26384 6112
rect 26700 6103 26752 6112
rect 26700 6069 26709 6103
rect 26709 6069 26743 6103
rect 26743 6069 26752 6103
rect 26700 6060 26752 6069
rect 26792 6060 26844 6112
rect 28356 6128 28408 6180
rect 28816 6171 28868 6180
rect 28816 6137 28825 6171
rect 28825 6137 28859 6171
rect 28859 6137 28868 6171
rect 28816 6128 28868 6137
rect 29920 6128 29972 6180
rect 29368 6060 29420 6112
rect 29736 6060 29788 6112
rect 32036 6196 32088 6248
rect 32588 6264 32640 6316
rect 32864 6307 32916 6316
rect 32864 6273 32873 6307
rect 32873 6273 32907 6307
rect 32907 6273 32916 6307
rect 32864 6264 32916 6273
rect 35072 6264 35124 6316
rect 35624 6264 35676 6316
rect 36084 6264 36136 6316
rect 36452 6264 36504 6316
rect 30840 6128 30892 6180
rect 31576 6128 31628 6180
rect 31300 6060 31352 6112
rect 31392 6103 31444 6112
rect 31392 6069 31401 6103
rect 31401 6069 31435 6103
rect 31435 6069 31444 6103
rect 31392 6060 31444 6069
rect 32220 6128 32272 6180
rect 32956 6196 33008 6248
rect 33508 6239 33560 6248
rect 33508 6205 33517 6239
rect 33517 6205 33551 6239
rect 33551 6205 33560 6239
rect 33508 6196 33560 6205
rect 33416 6128 33468 6180
rect 33876 6239 33928 6248
rect 33876 6205 33910 6239
rect 33910 6205 33928 6239
rect 33876 6196 33928 6205
rect 34060 6239 34112 6248
rect 34060 6205 34069 6239
rect 34069 6205 34103 6239
rect 34103 6205 34112 6239
rect 34060 6196 34112 6205
rect 35900 6239 35952 6248
rect 35900 6205 35909 6239
rect 35909 6205 35943 6239
rect 35943 6205 35952 6239
rect 35900 6196 35952 6205
rect 37740 6307 37792 6316
rect 37740 6273 37749 6307
rect 37749 6273 37783 6307
rect 37783 6273 37792 6307
rect 37740 6264 37792 6273
rect 38384 6264 38436 6316
rect 38660 6264 38712 6316
rect 39580 6307 39632 6316
rect 39580 6273 39614 6307
rect 39614 6273 39632 6307
rect 39580 6264 39632 6273
rect 42800 6307 42852 6316
rect 42800 6273 42809 6307
rect 42809 6273 42843 6307
rect 42843 6273 42852 6307
rect 42800 6264 42852 6273
rect 37188 6196 37240 6248
rect 37464 6239 37516 6248
rect 37464 6205 37473 6239
rect 37473 6205 37507 6239
rect 37507 6205 37516 6239
rect 37464 6196 37516 6205
rect 34612 6128 34664 6180
rect 39304 6196 39356 6248
rect 39764 6239 39816 6248
rect 39764 6205 39773 6239
rect 39773 6205 39807 6239
rect 39807 6205 39816 6239
rect 39764 6196 39816 6205
rect 39948 6196 40000 6248
rect 43352 6264 43404 6316
rect 34520 6060 34572 6112
rect 34888 6060 34940 6112
rect 35532 6060 35584 6112
rect 36268 6060 36320 6112
rect 36636 6060 36688 6112
rect 39212 6171 39264 6180
rect 39212 6137 39221 6171
rect 39221 6137 39255 6171
rect 39255 6137 39264 6171
rect 39212 6128 39264 6137
rect 39764 6060 39816 6112
rect 43076 6103 43128 6112
rect 43076 6069 43085 6103
rect 43085 6069 43119 6103
rect 43119 6069 43128 6103
rect 43076 6060 43128 6069
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 13918 5958 13970 6010
rect 13982 5958 14034 6010
rect 14046 5958 14098 6010
rect 14110 5958 14162 6010
rect 14174 5958 14226 6010
rect 14238 5958 14290 6010
rect 19918 5958 19970 6010
rect 19982 5958 20034 6010
rect 20046 5958 20098 6010
rect 20110 5958 20162 6010
rect 20174 5958 20226 6010
rect 20238 5958 20290 6010
rect 25918 5958 25970 6010
rect 25982 5958 26034 6010
rect 26046 5958 26098 6010
rect 26110 5958 26162 6010
rect 26174 5958 26226 6010
rect 26238 5958 26290 6010
rect 31918 5958 31970 6010
rect 31982 5958 32034 6010
rect 32046 5958 32098 6010
rect 32110 5958 32162 6010
rect 32174 5958 32226 6010
rect 32238 5958 32290 6010
rect 37918 5958 37970 6010
rect 37982 5958 38034 6010
rect 38046 5958 38098 6010
rect 38110 5958 38162 6010
rect 38174 5958 38226 6010
rect 38238 5958 38290 6010
rect 3056 5899 3108 5908
rect 3056 5865 3065 5899
rect 3065 5865 3099 5899
rect 3099 5865 3108 5899
rect 3056 5856 3108 5865
rect 4436 5899 4488 5908
rect 4436 5865 4445 5899
rect 4445 5865 4479 5899
rect 4479 5865 4488 5899
rect 4436 5856 4488 5865
rect 4620 5856 4672 5908
rect 5448 5856 5500 5908
rect 6920 5856 6972 5908
rect 3424 5831 3476 5840
rect 3424 5797 3433 5831
rect 3433 5797 3467 5831
rect 3467 5797 3476 5831
rect 3424 5788 3476 5797
rect 5356 5788 5408 5840
rect 1768 5720 1820 5772
rect 3240 5720 3292 5772
rect 4528 5720 4580 5772
rect 4620 5763 4672 5772
rect 4620 5729 4629 5763
rect 4629 5729 4663 5763
rect 4663 5729 4672 5763
rect 4620 5720 4672 5729
rect 5816 5720 5868 5772
rect 6368 5831 6420 5840
rect 6368 5797 6377 5831
rect 6377 5797 6411 5831
rect 6411 5797 6420 5831
rect 6368 5788 6420 5797
rect 6000 5720 6052 5772
rect 6736 5720 6788 5772
rect 7564 5856 7616 5908
rect 8760 5856 8812 5908
rect 11980 5856 12032 5908
rect 12532 5856 12584 5908
rect 13176 5856 13228 5908
rect 13360 5899 13412 5908
rect 13360 5865 13369 5899
rect 13369 5865 13403 5899
rect 13403 5865 13412 5899
rect 13360 5856 13412 5865
rect 13728 5856 13780 5908
rect 14188 5856 14240 5908
rect 14372 5856 14424 5908
rect 15200 5856 15252 5908
rect 7380 5788 7432 5840
rect 7748 5788 7800 5840
rect 8024 5788 8076 5840
rect 8668 5788 8720 5840
rect 10140 5831 10192 5840
rect 10140 5797 10149 5831
rect 10149 5797 10183 5831
rect 10183 5797 10192 5831
rect 10140 5788 10192 5797
rect 12072 5831 12124 5840
rect 12072 5797 12081 5831
rect 12081 5797 12115 5831
rect 12115 5797 12124 5831
rect 12072 5788 12124 5797
rect 1492 5695 1544 5704
rect 1492 5661 1501 5695
rect 1501 5661 1535 5695
rect 1535 5661 1544 5695
rect 1492 5652 1544 5661
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 4252 5652 4304 5704
rect 5540 5652 5592 5704
rect 2504 5584 2556 5636
rect 3424 5584 3476 5636
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 3516 5516 3568 5568
rect 3608 5516 3660 5568
rect 4712 5516 4764 5568
rect 6828 5516 6880 5568
rect 10048 5720 10100 5772
rect 10784 5763 10836 5772
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 11152 5720 11204 5772
rect 7932 5652 7984 5704
rect 9772 5695 9824 5704
rect 9772 5661 9790 5695
rect 9790 5661 9824 5695
rect 9772 5652 9824 5661
rect 8576 5627 8628 5636
rect 8576 5593 8585 5627
rect 8585 5593 8619 5627
rect 8619 5593 8628 5627
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 14372 5720 14424 5772
rect 15292 5788 15344 5840
rect 15384 5720 15436 5772
rect 16396 5788 16448 5840
rect 17408 5788 17460 5840
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 13452 5652 13504 5704
rect 8576 5584 8628 5593
rect 8392 5516 8444 5568
rect 9496 5516 9548 5568
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 13360 5584 13412 5636
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 14924 5652 14976 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 15936 5695 15988 5704
rect 15936 5661 15954 5695
rect 15954 5661 15988 5695
rect 15936 5652 15988 5661
rect 17592 5652 17644 5704
rect 17776 5652 17828 5704
rect 18604 5856 18656 5908
rect 19064 5856 19116 5908
rect 19248 5899 19300 5908
rect 19248 5865 19257 5899
rect 19257 5865 19291 5899
rect 19291 5865 19300 5899
rect 19248 5856 19300 5865
rect 19616 5856 19668 5908
rect 19984 5856 20036 5908
rect 20260 5856 20312 5908
rect 20720 5856 20772 5908
rect 20904 5856 20956 5908
rect 21548 5856 21600 5908
rect 21640 5856 21692 5908
rect 23940 5899 23992 5908
rect 23940 5865 23949 5899
rect 23949 5865 23983 5899
rect 23983 5865 23992 5899
rect 23940 5856 23992 5865
rect 24124 5856 24176 5908
rect 20352 5788 20404 5840
rect 20444 5831 20496 5840
rect 20444 5797 20453 5831
rect 20453 5797 20487 5831
rect 20487 5797 20496 5831
rect 20444 5788 20496 5797
rect 19340 5652 19392 5704
rect 19616 5652 19668 5704
rect 19800 5695 19852 5704
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 24584 5788 24636 5840
rect 19984 5720 20036 5729
rect 25688 5720 25740 5772
rect 29184 5856 29236 5908
rect 30196 5856 30248 5908
rect 30288 5856 30340 5908
rect 31024 5856 31076 5908
rect 32956 5856 33008 5908
rect 34060 5856 34112 5908
rect 34336 5899 34388 5908
rect 34336 5865 34345 5899
rect 34345 5865 34379 5899
rect 34379 5865 34388 5899
rect 34336 5856 34388 5865
rect 34704 5899 34756 5908
rect 34704 5865 34713 5899
rect 34713 5865 34747 5899
rect 34747 5865 34756 5899
rect 34704 5856 34756 5865
rect 26608 5788 26660 5840
rect 27804 5788 27856 5840
rect 29920 5788 29972 5840
rect 31300 5788 31352 5840
rect 36544 5856 36596 5908
rect 37372 5899 37424 5908
rect 37372 5865 37381 5899
rect 37381 5865 37415 5899
rect 37415 5865 37424 5899
rect 37372 5856 37424 5865
rect 37464 5856 37516 5908
rect 37648 5788 37700 5840
rect 39212 5899 39264 5908
rect 39212 5865 39221 5899
rect 39221 5865 39255 5899
rect 39255 5865 39264 5899
rect 39212 5856 39264 5865
rect 42892 5788 42944 5840
rect 43444 5831 43496 5840
rect 43444 5797 43453 5831
rect 43453 5797 43487 5831
rect 43487 5797 43496 5831
rect 43444 5788 43496 5797
rect 26240 5763 26292 5772
rect 26240 5729 26249 5763
rect 26249 5729 26283 5763
rect 26283 5729 26292 5763
rect 26240 5720 26292 5729
rect 26332 5720 26384 5772
rect 18880 5627 18932 5636
rect 18880 5593 18889 5627
rect 18889 5593 18923 5627
rect 18923 5593 18932 5627
rect 18880 5584 18932 5593
rect 18972 5584 19024 5636
rect 15476 5516 15528 5568
rect 15660 5516 15712 5568
rect 16488 5516 16540 5568
rect 18788 5516 18840 5568
rect 19156 5584 19208 5636
rect 19340 5516 19392 5568
rect 19708 5516 19760 5568
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 20904 5652 20956 5704
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 21548 5584 21600 5636
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 24768 5652 24820 5704
rect 23848 5584 23900 5636
rect 25596 5652 25648 5704
rect 25964 5652 26016 5704
rect 26994 5695 27046 5704
rect 26994 5661 27003 5695
rect 27003 5661 27037 5695
rect 27037 5661 27046 5695
rect 26994 5652 27046 5661
rect 27252 5695 27304 5704
rect 27252 5661 27261 5695
rect 27261 5661 27295 5695
rect 27295 5661 27304 5695
rect 27252 5652 27304 5661
rect 27896 5720 27948 5772
rect 28172 5720 28224 5772
rect 28356 5652 28408 5704
rect 29736 5695 29788 5704
rect 29736 5661 29745 5695
rect 29745 5661 29779 5695
rect 29779 5661 29788 5695
rect 29736 5652 29788 5661
rect 30748 5763 30800 5772
rect 30748 5729 30757 5763
rect 30757 5729 30791 5763
rect 30791 5729 30800 5763
rect 30748 5720 30800 5729
rect 31484 5720 31536 5772
rect 32680 5763 32732 5772
rect 32680 5729 32689 5763
rect 32689 5729 32723 5763
rect 32723 5729 32732 5763
rect 32680 5720 32732 5729
rect 36452 5720 36504 5772
rect 30932 5695 30984 5704
rect 30932 5661 30941 5695
rect 30941 5661 30975 5695
rect 30975 5661 30984 5695
rect 30932 5652 30984 5661
rect 31668 5695 31720 5704
rect 31668 5661 31677 5695
rect 31677 5661 31711 5695
rect 31711 5661 31720 5695
rect 31668 5652 31720 5661
rect 31760 5695 31812 5704
rect 31760 5661 31794 5695
rect 31794 5661 31812 5695
rect 31760 5652 31812 5661
rect 33048 5652 33100 5704
rect 34520 5695 34572 5704
rect 34520 5661 34529 5695
rect 34529 5661 34563 5695
rect 34563 5661 34572 5695
rect 34520 5652 34572 5661
rect 35440 5695 35492 5704
rect 35440 5661 35449 5695
rect 35449 5661 35483 5695
rect 35483 5661 35492 5695
rect 35440 5652 35492 5661
rect 21640 5516 21692 5568
rect 22008 5516 22060 5568
rect 24860 5516 24912 5568
rect 25044 5516 25096 5568
rect 26240 5584 26292 5636
rect 27988 5584 28040 5636
rect 29368 5584 29420 5636
rect 25596 5516 25648 5568
rect 27804 5516 27856 5568
rect 28264 5516 28316 5568
rect 29184 5516 29236 5568
rect 30748 5516 30800 5568
rect 31392 5516 31444 5568
rect 31944 5516 31996 5568
rect 32772 5516 32824 5568
rect 35992 5652 36044 5704
rect 37556 5695 37608 5704
rect 37556 5661 37565 5695
rect 37565 5661 37599 5695
rect 37599 5661 37608 5695
rect 37556 5652 37608 5661
rect 38200 5763 38252 5772
rect 38200 5729 38209 5763
rect 38209 5729 38243 5763
rect 38243 5729 38252 5763
rect 38200 5720 38252 5729
rect 37464 5584 37516 5636
rect 37740 5584 37792 5636
rect 39212 5652 39264 5704
rect 40224 5652 40276 5704
rect 41880 5652 41932 5704
rect 43536 5720 43588 5772
rect 38200 5584 38252 5636
rect 39672 5584 39724 5636
rect 36084 5516 36136 5568
rect 39304 5516 39356 5568
rect 42984 5516 43036 5568
rect 43076 5559 43128 5568
rect 43076 5525 43085 5559
rect 43085 5525 43119 5559
rect 43119 5525 43128 5559
rect 43076 5516 43128 5525
rect 2658 5414 2710 5466
rect 2722 5414 2774 5466
rect 2786 5414 2838 5466
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 8658 5414 8710 5466
rect 8722 5414 8774 5466
rect 8786 5414 8838 5466
rect 8850 5414 8902 5466
rect 8914 5414 8966 5466
rect 8978 5414 9030 5466
rect 14658 5414 14710 5466
rect 14722 5414 14774 5466
rect 14786 5414 14838 5466
rect 14850 5414 14902 5466
rect 14914 5414 14966 5466
rect 14978 5414 15030 5466
rect 20658 5414 20710 5466
rect 20722 5414 20774 5466
rect 20786 5414 20838 5466
rect 20850 5414 20902 5466
rect 20914 5414 20966 5466
rect 20978 5414 21030 5466
rect 26658 5414 26710 5466
rect 26722 5414 26774 5466
rect 26786 5414 26838 5466
rect 26850 5414 26902 5466
rect 26914 5414 26966 5466
rect 26978 5414 27030 5466
rect 32658 5414 32710 5466
rect 32722 5414 32774 5466
rect 32786 5414 32838 5466
rect 32850 5414 32902 5466
rect 32914 5414 32966 5466
rect 32978 5414 33030 5466
rect 38658 5414 38710 5466
rect 38722 5414 38774 5466
rect 38786 5414 38838 5466
rect 38850 5414 38902 5466
rect 38914 5414 38966 5466
rect 38978 5414 39030 5466
rect 2780 5312 2832 5364
rect 1584 5176 1636 5228
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2504 5176 2556 5228
rect 4804 5312 4856 5364
rect 4528 5244 4580 5296
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3884 5176 3936 5228
rect 4988 5176 5040 5228
rect 5172 5176 5224 5228
rect 6460 5244 6512 5296
rect 7104 5312 7156 5364
rect 7656 5312 7708 5364
rect 2688 5151 2740 5160
rect 2688 5117 2697 5151
rect 2697 5117 2731 5151
rect 2731 5117 2740 5151
rect 2688 5108 2740 5117
rect 3056 5108 3108 5160
rect 3148 5040 3200 5092
rect 3424 5083 3476 5092
rect 3424 5049 3433 5083
rect 3433 5049 3467 5083
rect 3467 5049 3476 5083
rect 3424 5040 3476 5049
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 6460 4972 6512 5024
rect 7104 5176 7156 5228
rect 8668 5312 8720 5364
rect 9956 5312 10008 5364
rect 10324 5312 10376 5364
rect 10784 5244 10836 5296
rect 11520 5312 11572 5364
rect 11612 5244 11664 5296
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 11060 5176 11112 5228
rect 12716 5312 12768 5364
rect 12992 5312 13044 5364
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 13636 5176 13688 5228
rect 13912 5176 13964 5228
rect 17224 5312 17276 5364
rect 17592 5312 17644 5364
rect 14188 5287 14240 5296
rect 14188 5253 14197 5287
rect 14197 5253 14231 5287
rect 14231 5253 14240 5287
rect 14188 5244 14240 5253
rect 16488 5244 16540 5296
rect 15016 5176 15068 5228
rect 15844 5219 15896 5228
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 16856 5176 16908 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 19248 5312 19300 5364
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 8300 5108 8352 5160
rect 9312 5108 9364 5160
rect 8576 5083 8628 5092
rect 8576 5049 8585 5083
rect 8585 5049 8619 5083
rect 8619 5049 8628 5083
rect 8576 5040 8628 5049
rect 10324 5040 10376 5092
rect 10784 4972 10836 5024
rect 11796 5108 11848 5160
rect 13360 5108 13412 5160
rect 11888 5040 11940 5092
rect 14464 5108 14516 5160
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 15200 5108 15252 5160
rect 15384 5108 15436 5160
rect 15660 5108 15712 5160
rect 16028 5108 16080 5160
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 18972 5176 19024 5228
rect 19432 5244 19484 5296
rect 19800 5244 19852 5296
rect 19984 5244 20036 5296
rect 22100 5312 22152 5364
rect 22192 5312 22244 5364
rect 23296 5312 23348 5364
rect 23940 5312 23992 5364
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 25504 5312 25556 5364
rect 30472 5312 30524 5364
rect 31208 5312 31260 5364
rect 31760 5355 31812 5364
rect 31760 5321 31769 5355
rect 31769 5321 31803 5355
rect 31803 5321 31812 5355
rect 31760 5312 31812 5321
rect 13728 5040 13780 5092
rect 13452 4972 13504 5024
rect 13912 4972 13964 5024
rect 14740 5040 14792 5092
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 19156 5108 19208 5160
rect 19708 5176 19760 5228
rect 15200 4972 15252 5024
rect 16212 4972 16264 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 18696 4972 18748 5024
rect 18788 4972 18840 5024
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 20076 5108 20128 5160
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 25780 5244 25832 5296
rect 25964 5287 26016 5296
rect 25964 5253 25973 5287
rect 25973 5253 26007 5287
rect 26007 5253 26016 5287
rect 25964 5244 26016 5253
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 20904 5108 20956 5160
rect 21180 5108 21232 5160
rect 21824 5108 21876 5160
rect 22468 5108 22520 5160
rect 19708 5040 19760 5092
rect 20536 5040 20588 5092
rect 21456 5040 21508 5092
rect 21548 4972 21600 5024
rect 22192 5040 22244 5092
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 23940 5219 23992 5228
rect 23940 5185 23974 5219
rect 23974 5185 23992 5219
rect 23940 5176 23992 5185
rect 24124 5219 24176 5228
rect 24124 5185 24133 5219
rect 24133 5185 24167 5219
rect 24167 5185 24176 5219
rect 24124 5176 24176 5185
rect 26608 5176 26660 5228
rect 26976 5176 27028 5228
rect 22744 5108 22796 5160
rect 23296 5108 23348 5160
rect 24492 5108 24544 5160
rect 25596 5108 25648 5160
rect 25872 5108 25924 5160
rect 27344 5176 27396 5228
rect 28264 5219 28316 5228
rect 28264 5185 28273 5219
rect 28273 5185 28307 5219
rect 28307 5185 28316 5219
rect 28264 5176 28316 5185
rect 30564 5244 30616 5296
rect 35624 5312 35676 5364
rect 32036 5244 32088 5296
rect 35716 5244 35768 5296
rect 43168 5312 43220 5364
rect 43444 5355 43496 5364
rect 43444 5321 43453 5355
rect 43453 5321 43487 5355
rect 43487 5321 43496 5355
rect 43444 5312 43496 5321
rect 36636 5244 36688 5296
rect 42708 5244 42760 5296
rect 21916 4972 21968 5024
rect 23296 4972 23348 5024
rect 23664 5040 23716 5092
rect 25228 5040 25280 5092
rect 24032 4972 24084 5024
rect 25320 5015 25372 5024
rect 25320 4981 25329 5015
rect 25329 4981 25363 5015
rect 25363 4981 25372 5015
rect 25320 4972 25372 4981
rect 26424 4972 26476 5024
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 27528 4972 27580 5024
rect 27896 4972 27948 5024
rect 28632 5108 28684 5160
rect 28908 5108 28960 5160
rect 29736 5219 29788 5228
rect 29736 5185 29745 5219
rect 29745 5185 29779 5219
rect 29779 5185 29788 5219
rect 29736 5176 29788 5185
rect 30012 5219 30064 5228
rect 30012 5185 30021 5219
rect 30021 5185 30055 5219
rect 30055 5185 30064 5219
rect 30012 5176 30064 5185
rect 31944 5219 31996 5228
rect 31944 5185 31953 5219
rect 31953 5185 31987 5219
rect 31987 5185 31996 5219
rect 31944 5176 31996 5185
rect 32404 5219 32456 5228
rect 32404 5185 32413 5219
rect 32413 5185 32447 5219
rect 32447 5185 32456 5219
rect 32404 5176 32456 5185
rect 33324 5176 33376 5228
rect 33692 5219 33744 5228
rect 33692 5185 33701 5219
rect 33701 5185 33735 5219
rect 33735 5185 33744 5219
rect 33692 5176 33744 5185
rect 34612 5219 34664 5228
rect 34612 5185 34621 5219
rect 34621 5185 34655 5219
rect 34655 5185 34664 5219
rect 34612 5176 34664 5185
rect 34888 5219 34940 5228
rect 34888 5185 34897 5219
rect 34897 5185 34931 5219
rect 34931 5185 34940 5219
rect 34888 5176 34940 5185
rect 36084 5219 36136 5228
rect 36084 5185 36093 5219
rect 36093 5185 36127 5219
rect 36127 5185 36136 5219
rect 36084 5176 36136 5185
rect 36452 5176 36504 5228
rect 37464 5176 37516 5228
rect 39212 5219 39264 5228
rect 39212 5185 39221 5219
rect 39221 5185 39255 5219
rect 39255 5185 39264 5219
rect 39212 5176 39264 5185
rect 42892 5219 42944 5228
rect 42892 5185 42901 5219
rect 42901 5185 42935 5219
rect 42935 5185 42944 5219
rect 42892 5176 42944 5185
rect 43260 5219 43312 5228
rect 43260 5185 43269 5219
rect 43269 5185 43303 5219
rect 43303 5185 43312 5219
rect 43260 5176 43312 5185
rect 30564 5108 30616 5160
rect 31576 5108 31628 5160
rect 28540 5040 28592 5092
rect 29460 5083 29512 5092
rect 29460 5049 29469 5083
rect 29469 5049 29503 5083
rect 29503 5049 29512 5083
rect 29460 5040 29512 5049
rect 30932 5040 30984 5092
rect 31300 5040 31352 5092
rect 34428 5108 34480 5160
rect 28080 5015 28132 5024
rect 28080 4981 28089 5015
rect 28089 4981 28123 5015
rect 28123 4981 28132 5015
rect 28080 4972 28132 4981
rect 28172 4972 28224 5024
rect 29184 4972 29236 5024
rect 31484 4972 31536 5024
rect 33048 4972 33100 5024
rect 33692 4972 33744 5024
rect 34704 4972 34756 5024
rect 35256 4972 35308 5024
rect 37188 5108 37240 5160
rect 36912 5040 36964 5092
rect 38476 5083 38528 5092
rect 38476 5049 38485 5083
rect 38485 5049 38519 5083
rect 38519 5049 38528 5083
rect 38476 5040 38528 5049
rect 36820 4972 36872 5024
rect 37372 4972 37424 5024
rect 38660 4972 38712 5024
rect 43076 5015 43128 5024
rect 43076 4981 43085 5015
rect 43085 4981 43119 5015
rect 43119 4981 43128 5015
rect 43076 4972 43128 4981
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 13918 4870 13970 4922
rect 13982 4870 14034 4922
rect 14046 4870 14098 4922
rect 14110 4870 14162 4922
rect 14174 4870 14226 4922
rect 14238 4870 14290 4922
rect 19918 4870 19970 4922
rect 19982 4870 20034 4922
rect 20046 4870 20098 4922
rect 20110 4870 20162 4922
rect 20174 4870 20226 4922
rect 20238 4870 20290 4922
rect 25918 4870 25970 4922
rect 25982 4870 26034 4922
rect 26046 4870 26098 4922
rect 26110 4870 26162 4922
rect 26174 4870 26226 4922
rect 26238 4870 26290 4922
rect 31918 4870 31970 4922
rect 31982 4870 32034 4922
rect 32046 4870 32098 4922
rect 32110 4870 32162 4922
rect 32174 4870 32226 4922
rect 32238 4870 32290 4922
rect 37918 4870 37970 4922
rect 37982 4870 38034 4922
rect 38046 4870 38098 4922
rect 38110 4870 38162 4922
rect 38174 4870 38226 4922
rect 38238 4870 38290 4922
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 3700 4768 3752 4820
rect 3332 4632 3384 4684
rect 3608 4632 3660 4684
rect 4804 4632 4856 4684
rect 5540 4632 5592 4684
rect 1400 4564 1452 4616
rect 1676 4564 1728 4616
rect 2596 4564 2648 4616
rect 2780 4564 2832 4616
rect 3056 4564 3108 4616
rect 2044 4539 2096 4548
rect 2044 4505 2053 4539
rect 2053 4505 2087 4539
rect 2087 4505 2096 4539
rect 2044 4496 2096 4505
rect 3148 4496 3200 4548
rect 5816 4632 5868 4684
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 2504 4428 2556 4480
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 6276 4607 6328 4616
rect 6276 4573 6310 4607
rect 6310 4573 6328 4607
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 7564 4632 7616 4684
rect 8576 4768 8628 4820
rect 9128 4768 9180 4820
rect 9312 4768 9364 4820
rect 9036 4700 9088 4752
rect 12716 4768 12768 4820
rect 12992 4768 13044 4820
rect 14372 4768 14424 4820
rect 11796 4700 11848 4752
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 10324 4632 10376 4684
rect 6276 4564 6328 4573
rect 5356 4496 5408 4548
rect 7196 4496 7248 4548
rect 7748 4496 7800 4548
rect 9680 4607 9732 4616
rect 9680 4573 9686 4607
rect 9686 4573 9720 4607
rect 9720 4573 9732 4607
rect 9680 4564 9732 4573
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 11428 4564 11480 4616
rect 6736 4428 6788 4480
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 11152 4496 11204 4548
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12808 4632 12860 4684
rect 14740 4768 14792 4820
rect 14832 4768 14884 4820
rect 15108 4768 15160 4820
rect 15384 4700 15436 4752
rect 15568 4700 15620 4752
rect 16396 4632 16448 4684
rect 16856 4768 16908 4820
rect 17316 4768 17368 4820
rect 17500 4811 17552 4820
rect 17500 4777 17509 4811
rect 17509 4777 17543 4811
rect 17543 4777 17552 4811
rect 17500 4768 17552 4777
rect 18052 4768 18104 4820
rect 18328 4768 18380 4820
rect 19156 4768 19208 4820
rect 17592 4700 17644 4752
rect 18420 4700 18472 4752
rect 19248 4743 19300 4752
rect 19248 4709 19257 4743
rect 19257 4709 19291 4743
rect 19291 4709 19300 4743
rect 19248 4700 19300 4709
rect 18604 4632 18656 4684
rect 18788 4675 18840 4684
rect 18788 4641 18797 4675
rect 18797 4641 18831 4675
rect 18831 4641 18840 4675
rect 18788 4632 18840 4641
rect 12624 4564 12676 4616
rect 14096 4564 14148 4616
rect 14372 4564 14424 4616
rect 14924 4564 14976 4616
rect 15292 4564 15344 4616
rect 15568 4564 15620 4616
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 16212 4564 16264 4616
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 19064 4564 19116 4616
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 11060 4428 11112 4480
rect 18788 4496 18840 4548
rect 20904 4768 20956 4820
rect 22008 4768 22060 4820
rect 22100 4768 22152 4820
rect 22284 4768 22336 4820
rect 20260 4632 20312 4684
rect 20536 4675 20588 4684
rect 20536 4641 20545 4675
rect 20545 4641 20579 4675
rect 20579 4641 20588 4675
rect 20536 4632 20588 4641
rect 21548 4700 21600 4752
rect 21732 4700 21784 4752
rect 26056 4768 26108 4820
rect 26424 4768 26476 4820
rect 26976 4768 27028 4820
rect 27804 4768 27856 4820
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 21640 4632 21692 4684
rect 23204 4675 23256 4684
rect 23204 4641 23222 4675
rect 23222 4641 23256 4675
rect 23204 4632 23256 4641
rect 23296 4675 23348 4684
rect 23296 4641 23305 4675
rect 23305 4641 23339 4675
rect 23339 4641 23348 4675
rect 23296 4632 23348 4641
rect 26424 4664 26476 4673
rect 26424 4630 26433 4664
rect 26433 4630 26467 4664
rect 26467 4630 26476 4664
rect 26424 4621 26476 4630
rect 27896 4632 27948 4684
rect 19892 4607 19944 4616
rect 19892 4573 19901 4607
rect 19901 4573 19935 4607
rect 19935 4573 19944 4607
rect 19892 4564 19944 4573
rect 20904 4607 20956 4616
rect 20904 4573 20938 4607
rect 20938 4573 20956 4607
rect 20904 4564 20956 4573
rect 21088 4607 21140 4616
rect 21088 4573 21097 4607
rect 21097 4573 21131 4607
rect 21131 4573 21140 4607
rect 21088 4564 21140 4573
rect 22192 4564 22244 4616
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 13360 4428 13412 4480
rect 13728 4428 13780 4480
rect 14556 4428 14608 4480
rect 15476 4428 15528 4480
rect 19064 4428 19116 4480
rect 21824 4539 21876 4548
rect 21824 4505 21833 4539
rect 21833 4505 21867 4539
rect 21867 4505 21876 4539
rect 21824 4496 21876 4505
rect 24768 4564 24820 4616
rect 25228 4564 25280 4616
rect 25412 4564 25464 4616
rect 25964 4564 26016 4616
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 26332 4564 26384 4573
rect 26700 4607 26752 4616
rect 26700 4573 26709 4607
rect 26709 4573 26743 4607
rect 26743 4573 26752 4607
rect 26700 4564 26752 4573
rect 27436 4564 27488 4616
rect 27620 4564 27672 4616
rect 30012 4768 30064 4820
rect 29736 4700 29788 4752
rect 30564 4768 30616 4820
rect 31392 4768 31444 4820
rect 32588 4768 32640 4820
rect 28264 4675 28316 4684
rect 28264 4641 28273 4675
rect 28273 4641 28307 4675
rect 28307 4641 28316 4675
rect 28264 4632 28316 4641
rect 28908 4632 28960 4684
rect 28540 4607 28592 4616
rect 28540 4573 28549 4607
rect 28549 4573 28583 4607
rect 28583 4573 28592 4607
rect 28540 4564 28592 4573
rect 28632 4564 28684 4616
rect 30656 4632 30708 4684
rect 31760 4632 31812 4684
rect 32404 4675 32456 4684
rect 32404 4641 32413 4675
rect 32413 4641 32447 4675
rect 32447 4641 32456 4675
rect 32404 4632 32456 4641
rect 33324 4811 33376 4820
rect 33324 4777 33333 4811
rect 33333 4777 33367 4811
rect 33367 4777 33376 4811
rect 33324 4768 33376 4777
rect 34060 4768 34112 4820
rect 36636 4768 36688 4820
rect 35072 4743 35124 4752
rect 35072 4709 35081 4743
rect 35081 4709 35115 4743
rect 35115 4709 35124 4743
rect 35072 4700 35124 4709
rect 36544 4700 36596 4752
rect 39764 4768 39816 4820
rect 42892 4768 42944 4820
rect 36820 4743 36872 4752
rect 36820 4709 36829 4743
rect 36829 4709 36863 4743
rect 36863 4709 36872 4743
rect 36820 4700 36872 4709
rect 43444 4743 43496 4752
rect 43444 4709 43453 4743
rect 43453 4709 43487 4743
rect 43487 4709 43496 4743
rect 43444 4700 43496 4709
rect 37372 4675 37424 4684
rect 37372 4641 37381 4675
rect 37381 4641 37415 4675
rect 37415 4641 37424 4675
rect 37372 4632 37424 4641
rect 37556 4632 37608 4684
rect 22100 4428 22152 4480
rect 22376 4471 22428 4480
rect 22376 4437 22385 4471
rect 22385 4437 22419 4471
rect 22419 4437 22428 4471
rect 22376 4428 22428 4437
rect 22928 4428 22980 4480
rect 28908 4496 28960 4548
rect 25228 4471 25280 4480
rect 25228 4437 25237 4471
rect 25237 4437 25271 4471
rect 25271 4437 25280 4471
rect 25228 4428 25280 4437
rect 25596 4428 25648 4480
rect 25964 4428 26016 4480
rect 26424 4471 26476 4480
rect 26424 4437 26433 4471
rect 26433 4437 26467 4471
rect 26467 4437 26476 4471
rect 26424 4428 26476 4437
rect 26700 4428 26752 4480
rect 30748 4607 30800 4616
rect 30748 4573 30757 4607
rect 30757 4573 30791 4607
rect 30791 4573 30800 4607
rect 30748 4564 30800 4573
rect 31484 4607 31536 4616
rect 31484 4573 31493 4607
rect 31493 4573 31527 4607
rect 31527 4573 31536 4607
rect 31484 4564 31536 4573
rect 32588 4564 32640 4616
rect 32680 4607 32732 4616
rect 32680 4573 32689 4607
rect 32689 4573 32723 4607
rect 32723 4573 32732 4607
rect 32680 4564 32732 4573
rect 34152 4564 34204 4616
rect 36084 4564 36136 4616
rect 31300 4496 31352 4548
rect 30472 4428 30524 4480
rect 30656 4428 30708 4480
rect 34244 4539 34296 4548
rect 34244 4505 34253 4539
rect 34253 4505 34287 4539
rect 34287 4505 34296 4539
rect 34244 4496 34296 4505
rect 32956 4428 33008 4480
rect 33508 4428 33560 4480
rect 36360 4607 36412 4616
rect 36360 4573 36369 4607
rect 36369 4573 36403 4607
rect 36403 4573 36412 4607
rect 36360 4564 36412 4573
rect 37096 4607 37148 4616
rect 37096 4573 37105 4607
rect 37105 4573 37139 4607
rect 37139 4573 37148 4607
rect 37096 4564 37148 4573
rect 38384 4632 38436 4684
rect 38660 4564 38712 4616
rect 42800 4564 42852 4616
rect 43168 4564 43220 4616
rect 36636 4428 36688 4480
rect 37280 4428 37332 4480
rect 43076 4471 43128 4480
rect 43076 4437 43085 4471
rect 43085 4437 43119 4471
rect 43119 4437 43128 4471
rect 43076 4428 43128 4437
rect 2658 4326 2710 4378
rect 2722 4326 2774 4378
rect 2786 4326 2838 4378
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 8658 4326 8710 4378
rect 8722 4326 8774 4378
rect 8786 4326 8838 4378
rect 8850 4326 8902 4378
rect 8914 4326 8966 4378
rect 8978 4326 9030 4378
rect 14658 4326 14710 4378
rect 14722 4326 14774 4378
rect 14786 4326 14838 4378
rect 14850 4326 14902 4378
rect 14914 4326 14966 4378
rect 14978 4326 15030 4378
rect 20658 4326 20710 4378
rect 20722 4326 20774 4378
rect 20786 4326 20838 4378
rect 20850 4326 20902 4378
rect 20914 4326 20966 4378
rect 20978 4326 21030 4378
rect 26658 4326 26710 4378
rect 26722 4326 26774 4378
rect 26786 4326 26838 4378
rect 26850 4326 26902 4378
rect 26914 4326 26966 4378
rect 26978 4326 27030 4378
rect 32658 4326 32710 4378
rect 32722 4326 32774 4378
rect 32786 4326 32838 4378
rect 32850 4326 32902 4378
rect 32914 4326 32966 4378
rect 32978 4326 33030 4378
rect 38658 4326 38710 4378
rect 38722 4326 38774 4378
rect 38786 4326 38838 4378
rect 38850 4326 38902 4378
rect 38914 4326 38966 4378
rect 38978 4326 39030 4378
rect 2412 4224 2464 4276
rect 3148 4224 3200 4276
rect 1492 4199 1544 4208
rect 1492 4165 1501 4199
rect 1501 4165 1535 4199
rect 1535 4165 1544 4199
rect 1492 4156 1544 4165
rect 1860 4199 1912 4208
rect 1860 4165 1869 4199
rect 1869 4165 1903 4199
rect 1903 4165 1912 4199
rect 1860 4156 1912 4165
rect 2228 4199 2280 4208
rect 2228 4165 2237 4199
rect 2237 4165 2271 4199
rect 2271 4165 2280 4199
rect 2228 4156 2280 4165
rect 3056 4156 3108 4208
rect 5172 4224 5224 4276
rect 5356 4224 5408 4276
rect 5908 4224 5960 4276
rect 6644 4224 6696 4276
rect 8392 4224 8444 4276
rect 1492 4020 1544 4072
rect 3332 4088 3384 4140
rect 4436 4156 4488 4208
rect 4896 4156 4948 4208
rect 4620 4088 4672 4140
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 7288 4088 7340 4140
rect 13268 4224 13320 4276
rect 13912 4224 13964 4276
rect 16672 4224 16724 4276
rect 18696 4224 18748 4276
rect 19064 4224 19116 4276
rect 19248 4224 19300 4276
rect 10876 4156 10928 4208
rect 21824 4224 21876 4276
rect 22376 4224 22428 4276
rect 22468 4224 22520 4276
rect 25136 4224 25188 4276
rect 25228 4224 25280 4276
rect 26332 4224 26384 4276
rect 27068 4224 27120 4276
rect 28172 4224 28224 4276
rect 9772 4088 9824 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 3056 3952 3108 4004
rect 4436 3995 4488 4004
rect 4436 3961 4445 3995
rect 4445 3961 4479 3995
rect 4479 3961 4488 3995
rect 4436 3952 4488 3961
rect 1768 3884 1820 3936
rect 2596 3884 2648 3936
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 3884 3884 3936 3936
rect 5448 4020 5500 4072
rect 7748 4020 7800 4072
rect 8576 4020 8628 4072
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 8944 4020 8996 4072
rect 9404 4020 9456 4072
rect 10048 4020 10100 4072
rect 11152 4088 11204 4140
rect 11796 4088 11848 4140
rect 25320 4156 25372 4208
rect 13084 4088 13136 4140
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 15660 4088 15712 4140
rect 16856 4131 16908 4140
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18972 4088 19024 4140
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 12164 3952 12216 4004
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 10968 3884 11020 3936
rect 11520 3884 11572 3936
rect 11888 3884 11940 3936
rect 11980 3884 12032 3936
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 13268 3952 13320 4004
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14464 4020 14516 4072
rect 16764 4020 16816 4072
rect 14740 3952 14792 4004
rect 15568 3884 15620 3936
rect 16488 3952 16540 4004
rect 17684 4063 17736 4072
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 23020 4088 23072 4140
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 17684 4029 17718 4063
rect 17718 4029 17736 4063
rect 17684 4020 17736 4029
rect 18512 3884 18564 3936
rect 20536 4020 20588 4072
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 20904 4020 20956 4072
rect 20996 4063 21048 4072
rect 20996 4029 21005 4063
rect 21005 4029 21039 4063
rect 21039 4029 21048 4063
rect 20996 4020 21048 4029
rect 21640 4020 21692 4072
rect 22192 4020 22244 4072
rect 22836 4020 22888 4072
rect 23204 4020 23256 4072
rect 23664 4020 23716 4072
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 24308 4020 24360 4072
rect 20444 3995 20496 4004
rect 20444 3961 20453 3995
rect 20453 3961 20487 3995
rect 20487 3961 20496 3995
rect 20444 3952 20496 3961
rect 21456 3952 21508 4004
rect 23480 3952 23532 4004
rect 24676 4020 24728 4072
rect 25412 4131 25464 4140
rect 25412 4097 25421 4131
rect 25421 4097 25455 4131
rect 25455 4097 25464 4131
rect 25412 4088 25464 4097
rect 25872 4156 25924 4208
rect 25964 4088 26016 4140
rect 26056 4088 26108 4140
rect 28448 4156 28500 4208
rect 28264 4131 28316 4140
rect 28264 4097 28273 4131
rect 28273 4097 28307 4131
rect 28307 4097 28316 4131
rect 28264 4088 28316 4097
rect 29460 4224 29512 4276
rect 29828 4224 29880 4276
rect 31484 4224 31536 4276
rect 32772 4224 32824 4276
rect 33140 4224 33192 4276
rect 28724 4156 28776 4208
rect 31668 4156 31720 4208
rect 30472 4088 30524 4140
rect 30656 4131 30708 4140
rect 30656 4097 30665 4131
rect 30665 4097 30699 4131
rect 30699 4097 30708 4131
rect 30656 4088 30708 4097
rect 31024 4088 31076 4140
rect 32220 4088 32272 4140
rect 32588 4131 32640 4140
rect 32588 4097 32597 4131
rect 32597 4097 32631 4131
rect 32631 4097 32640 4131
rect 32588 4088 32640 4097
rect 33416 4131 33468 4140
rect 33416 4097 33450 4131
rect 33450 4097 33468 4131
rect 34244 4267 34296 4276
rect 34244 4233 34253 4267
rect 34253 4233 34287 4267
rect 34287 4233 34296 4267
rect 34244 4224 34296 4233
rect 34520 4224 34572 4276
rect 39764 4224 39816 4276
rect 36176 4156 36228 4208
rect 39488 4156 39540 4208
rect 39580 4156 39632 4208
rect 42156 4156 42208 4208
rect 33416 4088 33468 4097
rect 25596 3995 25648 4004
rect 25596 3961 25605 3995
rect 25605 3961 25639 3995
rect 25639 3961 25648 3995
rect 25596 3952 25648 3961
rect 27528 4020 27580 4072
rect 27804 4020 27856 4072
rect 26792 3952 26844 4004
rect 27988 3952 28040 4004
rect 23020 3884 23072 3936
rect 26240 3884 26292 3936
rect 27344 3884 27396 3936
rect 27436 3884 27488 3936
rect 32220 3952 32272 4004
rect 32588 3952 32640 4004
rect 33048 4063 33100 4072
rect 33048 4029 33057 4063
rect 33057 4029 33091 4063
rect 33091 4029 33100 4063
rect 33048 4020 33100 4029
rect 33140 4020 33192 4072
rect 33600 4063 33652 4072
rect 33600 4029 33609 4063
rect 33609 4029 33643 4063
rect 33643 4029 33652 4063
rect 33600 4020 33652 4029
rect 34336 4063 34388 4072
rect 34336 4029 34345 4063
rect 34345 4029 34379 4063
rect 34379 4029 34388 4063
rect 34336 4020 34388 4029
rect 35348 4131 35400 4140
rect 35348 4097 35382 4131
rect 35382 4097 35400 4131
rect 35348 4088 35400 4097
rect 37188 4088 37240 4140
rect 38752 4088 38804 4140
rect 42064 4088 42116 4140
rect 42616 4131 42668 4140
rect 42616 4097 42625 4131
rect 42625 4097 42659 4131
rect 42659 4097 42668 4131
rect 42616 4088 42668 4097
rect 30472 3884 30524 3936
rect 35532 4063 35584 4072
rect 35532 4029 35541 4063
rect 35541 4029 35575 4063
rect 35575 4029 35584 4063
rect 35532 4020 35584 4029
rect 36084 4020 36136 4072
rect 36268 4020 36320 4072
rect 39212 4020 39264 4072
rect 39488 4020 39540 4072
rect 42984 4088 43036 4140
rect 34980 3995 35032 4004
rect 34980 3961 34989 3995
rect 34989 3961 35023 3995
rect 35023 3961 35032 3995
rect 34980 3952 35032 3961
rect 36728 3995 36780 4004
rect 36728 3961 36737 3995
rect 36737 3961 36771 3995
rect 36771 3961 36780 3995
rect 36728 3952 36780 3961
rect 34796 3884 34848 3936
rect 41972 3952 42024 4004
rect 43444 3995 43496 4004
rect 43444 3961 43453 3995
rect 43453 3961 43487 3995
rect 43487 3961 43496 3995
rect 43444 3952 43496 3961
rect 37832 3884 37884 3936
rect 38752 3884 38804 3936
rect 41788 3884 41840 3936
rect 43076 3927 43128 3936
rect 43076 3893 43085 3927
rect 43085 3893 43119 3927
rect 43119 3893 43128 3927
rect 43076 3884 43128 3893
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 13918 3782 13970 3834
rect 13982 3782 14034 3834
rect 14046 3782 14098 3834
rect 14110 3782 14162 3834
rect 14174 3782 14226 3834
rect 14238 3782 14290 3834
rect 19918 3782 19970 3834
rect 19982 3782 20034 3834
rect 20046 3782 20098 3834
rect 20110 3782 20162 3834
rect 20174 3782 20226 3834
rect 20238 3782 20290 3834
rect 25918 3782 25970 3834
rect 25982 3782 26034 3834
rect 26046 3782 26098 3834
rect 26110 3782 26162 3834
rect 26174 3782 26226 3834
rect 26238 3782 26290 3834
rect 31918 3782 31970 3834
rect 31982 3782 32034 3834
rect 32046 3782 32098 3834
rect 32110 3782 32162 3834
rect 32174 3782 32226 3834
rect 32238 3782 32290 3834
rect 37918 3782 37970 3834
rect 37982 3782 38034 3834
rect 38046 3782 38098 3834
rect 38110 3782 38162 3834
rect 38174 3782 38226 3834
rect 38238 3782 38290 3834
rect 1768 3680 1820 3732
rect 2964 3680 3016 3732
rect 3056 3680 3108 3732
rect 6644 3680 6696 3732
rect 7472 3680 7524 3732
rect 3700 3612 3752 3664
rect 4068 3612 4120 3664
rect 4436 3612 4488 3664
rect 4620 3544 4672 3596
rect 4712 3544 4764 3596
rect 7380 3544 7432 3596
rect 1400 3476 1452 3528
rect 2688 3476 2740 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 9864 3680 9916 3732
rect 10416 3612 10468 3664
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 12808 3680 12860 3732
rect 13728 3680 13780 3732
rect 13820 3680 13872 3732
rect 7840 3544 7892 3596
rect 8300 3544 8352 3596
rect 8576 3544 8628 3596
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 7932 3476 7984 3528
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 2228 3451 2280 3460
rect 2228 3417 2237 3451
rect 2237 3417 2271 3451
rect 2271 3417 2280 3451
rect 2228 3408 2280 3417
rect 2412 3408 2464 3460
rect 3976 3408 4028 3460
rect 9772 3544 9824 3596
rect 15108 3612 15160 3664
rect 17868 3680 17920 3732
rect 17960 3680 18012 3732
rect 17500 3612 17552 3664
rect 18328 3680 18380 3732
rect 19248 3612 19300 3664
rect 19340 3655 19392 3664
rect 19340 3621 19349 3655
rect 19349 3621 19383 3655
rect 19383 3621 19392 3655
rect 19340 3612 19392 3621
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 1676 3340 1728 3392
rect 8024 3340 8076 3392
rect 9496 3408 9548 3460
rect 8852 3340 8904 3392
rect 9680 3340 9732 3392
rect 11612 3587 11664 3596
rect 11612 3553 11621 3587
rect 11621 3553 11655 3587
rect 11655 3553 11664 3587
rect 11612 3544 11664 3553
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 10876 3476 10928 3528
rect 13268 3476 13320 3528
rect 13636 3476 13688 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 11336 3340 11388 3392
rect 12532 3340 12584 3392
rect 12716 3340 12768 3392
rect 14464 3408 14516 3460
rect 15108 3408 15160 3460
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 19432 3544 19484 3596
rect 20904 3680 20956 3732
rect 24308 3680 24360 3732
rect 25136 3680 25188 3732
rect 20996 3612 21048 3664
rect 21364 3544 21416 3596
rect 15660 3476 15712 3528
rect 17224 3476 17276 3528
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 17684 3476 17736 3528
rect 18144 3476 18196 3528
rect 19340 3476 19392 3528
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 20536 3476 20588 3528
rect 21824 3519 21876 3528
rect 21824 3485 21833 3519
rect 21833 3485 21867 3519
rect 21867 3485 21876 3519
rect 21824 3476 21876 3485
rect 19800 3408 19852 3460
rect 20904 3408 20956 3460
rect 21180 3408 21232 3460
rect 23480 3612 23532 3664
rect 25044 3612 25096 3664
rect 26332 3680 26384 3732
rect 22652 3587 22704 3596
rect 22652 3553 22661 3587
rect 22661 3553 22695 3587
rect 22695 3553 22704 3587
rect 22652 3544 22704 3553
rect 25688 3587 25740 3596
rect 25688 3553 25697 3587
rect 25697 3553 25731 3587
rect 25731 3553 25740 3587
rect 25688 3544 25740 3553
rect 25872 3587 25924 3596
rect 25872 3553 25881 3587
rect 25881 3553 25915 3587
rect 25915 3553 25924 3587
rect 25872 3544 25924 3553
rect 26332 3587 26384 3596
rect 26332 3553 26341 3587
rect 26341 3553 26375 3587
rect 26375 3553 26384 3587
rect 26332 3544 26384 3553
rect 26608 3587 26660 3596
rect 26608 3553 26617 3587
rect 26617 3553 26651 3587
rect 26651 3553 26660 3587
rect 26608 3544 26660 3553
rect 26792 3544 26844 3596
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 26884 3544 26936 3553
rect 27068 3544 27120 3596
rect 12992 3340 13044 3392
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 13544 3383 13596 3392
rect 13544 3349 13553 3383
rect 13553 3349 13587 3383
rect 13587 3349 13596 3383
rect 13544 3340 13596 3349
rect 13636 3340 13688 3392
rect 14004 3340 14056 3392
rect 14188 3340 14240 3392
rect 15660 3340 15712 3392
rect 16764 3340 16816 3392
rect 17868 3340 17920 3392
rect 18144 3340 18196 3392
rect 20444 3340 20496 3392
rect 21456 3340 21508 3392
rect 22008 3383 22060 3392
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 23848 3476 23900 3528
rect 25228 3476 25280 3528
rect 28264 3680 28316 3732
rect 28264 3587 28316 3596
rect 28264 3553 28273 3587
rect 28273 3553 28307 3587
rect 28307 3553 28316 3587
rect 28264 3544 28316 3553
rect 30564 3723 30616 3732
rect 30564 3689 30573 3723
rect 30573 3689 30607 3723
rect 30607 3689 30616 3723
rect 30564 3680 30616 3689
rect 31116 3680 31168 3732
rect 30748 3612 30800 3664
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 33600 3680 33652 3732
rect 34980 3680 35032 3732
rect 35532 3680 35584 3732
rect 41512 3680 41564 3732
rect 38476 3612 38528 3664
rect 38752 3612 38804 3664
rect 41420 3612 41472 3664
rect 43444 3655 43496 3664
rect 43444 3621 43453 3655
rect 43453 3621 43487 3655
rect 43487 3621 43496 3655
rect 43444 3612 43496 3621
rect 28448 3476 28500 3528
rect 28632 3476 28684 3528
rect 29460 3476 29512 3528
rect 25044 3340 25096 3392
rect 29736 3408 29788 3460
rect 31852 3519 31904 3528
rect 31852 3485 31861 3519
rect 31861 3485 31895 3519
rect 31895 3485 31904 3519
rect 31852 3476 31904 3485
rect 32956 3519 33008 3528
rect 32956 3485 32965 3519
rect 32965 3485 32999 3519
rect 32999 3485 33008 3519
rect 32956 3476 33008 3485
rect 35072 3544 35124 3596
rect 30104 3408 30156 3460
rect 27160 3340 27212 3392
rect 27344 3340 27396 3392
rect 28540 3340 28592 3392
rect 32312 3408 32364 3460
rect 34888 3519 34940 3528
rect 34888 3485 34897 3519
rect 34897 3485 34931 3519
rect 34931 3485 34940 3519
rect 34888 3476 34940 3485
rect 30472 3340 30524 3392
rect 33416 3408 33468 3460
rect 33876 3408 33928 3460
rect 36268 3587 36320 3596
rect 36268 3553 36277 3587
rect 36277 3553 36311 3587
rect 36311 3553 36320 3587
rect 36268 3544 36320 3553
rect 35900 3476 35952 3528
rect 36544 3476 36596 3528
rect 37648 3476 37700 3528
rect 38292 3476 38344 3528
rect 36360 3408 36412 3460
rect 37740 3408 37792 3460
rect 38752 3451 38804 3460
rect 38752 3417 38761 3451
rect 38761 3417 38795 3451
rect 38795 3417 38804 3451
rect 38752 3408 38804 3417
rect 33048 3340 33100 3392
rect 34704 3383 34756 3392
rect 34704 3349 34713 3383
rect 34713 3349 34747 3383
rect 34747 3349 34756 3383
rect 34704 3340 34756 3349
rect 35164 3340 35216 3392
rect 39304 3476 39356 3528
rect 39212 3408 39264 3460
rect 41972 3408 42024 3460
rect 42524 3519 42576 3528
rect 42524 3485 42533 3519
rect 42533 3485 42567 3519
rect 42567 3485 42576 3519
rect 42524 3476 42576 3485
rect 42708 3408 42760 3460
rect 43260 3519 43312 3528
rect 43260 3485 43269 3519
rect 43269 3485 43303 3519
rect 43303 3485 43312 3519
rect 43260 3476 43312 3485
rect 43076 3383 43128 3392
rect 43076 3349 43085 3383
rect 43085 3349 43119 3383
rect 43119 3349 43128 3383
rect 43076 3340 43128 3349
rect 43260 3340 43312 3392
rect 2658 3238 2710 3290
rect 2722 3238 2774 3290
rect 2786 3238 2838 3290
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 8658 3238 8710 3290
rect 8722 3238 8774 3290
rect 8786 3238 8838 3290
rect 8850 3238 8902 3290
rect 8914 3238 8966 3290
rect 8978 3238 9030 3290
rect 14658 3238 14710 3290
rect 14722 3238 14774 3290
rect 14786 3238 14838 3290
rect 14850 3238 14902 3290
rect 14914 3238 14966 3290
rect 14978 3238 15030 3290
rect 20658 3238 20710 3290
rect 20722 3238 20774 3290
rect 20786 3238 20838 3290
rect 20850 3238 20902 3290
rect 20914 3238 20966 3290
rect 20978 3238 21030 3290
rect 26658 3238 26710 3290
rect 26722 3238 26774 3290
rect 26786 3238 26838 3290
rect 26850 3238 26902 3290
rect 26914 3238 26966 3290
rect 26978 3238 27030 3290
rect 32658 3238 32710 3290
rect 32722 3238 32774 3290
rect 32786 3238 32838 3290
rect 32850 3238 32902 3290
rect 32914 3238 32966 3290
rect 32978 3238 33030 3290
rect 38658 3238 38710 3290
rect 38722 3238 38774 3290
rect 38786 3238 38838 3290
rect 38850 3238 38902 3290
rect 38914 3238 38966 3290
rect 38978 3238 39030 3290
rect 6184 3136 6236 3188
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 7748 3136 7800 3188
rect 2780 3111 2832 3120
rect 2780 3077 2789 3111
rect 2789 3077 2823 3111
rect 2823 3077 2832 3111
rect 2780 3068 2832 3077
rect 3056 3068 3108 3120
rect 8024 3068 8076 3120
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 5172 3000 5224 3052
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 4712 2932 4764 2984
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 7840 2932 7892 2984
rect 8300 2932 8352 2984
rect 8668 2932 8720 2984
rect 8944 2975 8996 2984
rect 8944 2941 8978 2975
rect 8978 2941 8996 2975
rect 8944 2932 8996 2941
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 9128 2932 9180 2941
rect 2504 2907 2556 2916
rect 2504 2873 2513 2907
rect 2513 2873 2547 2907
rect 2547 2873 2556 2907
rect 2504 2864 2556 2873
rect 7840 2796 7892 2848
rect 8576 2907 8628 2916
rect 8576 2873 8585 2907
rect 8585 2873 8619 2907
rect 8619 2873 8628 2907
rect 8576 2864 8628 2873
rect 10508 3000 10560 3052
rect 10784 3068 10836 3120
rect 10692 3000 10744 3052
rect 14280 3136 14332 3188
rect 15936 3136 15988 3188
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 16856 3179 16908 3188
rect 16856 3145 16865 3179
rect 16865 3145 16899 3179
rect 16899 3145 16908 3179
rect 16856 3136 16908 3145
rect 17224 3179 17276 3188
rect 17224 3145 17233 3179
rect 17233 3145 17267 3179
rect 17267 3145 17276 3179
rect 17224 3136 17276 3145
rect 19524 3136 19576 3188
rect 19800 3136 19852 3188
rect 13636 3068 13688 3120
rect 10048 2932 10100 2984
rect 10324 2975 10376 2984
rect 10324 2941 10333 2975
rect 10333 2941 10367 2975
rect 10367 2941 10376 2975
rect 10324 2932 10376 2941
rect 11520 2975 11572 2984
rect 11520 2941 11529 2975
rect 11529 2941 11563 2975
rect 11563 2941 11572 2975
rect 11520 2932 11572 2941
rect 12624 3000 12676 3052
rect 13360 3000 13412 3052
rect 13820 3068 13872 3120
rect 14464 3068 14516 3120
rect 22652 3068 22704 3120
rect 14004 3000 14056 3052
rect 10140 2796 10192 2848
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 14556 2839 14608 2848
rect 14556 2805 14565 2839
rect 14565 2805 14599 2839
rect 14599 2805 14608 2839
rect 14556 2796 14608 2805
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 16764 3043 16816 3052
rect 16764 3009 16773 3043
rect 16773 3009 16807 3043
rect 16807 3009 16816 3043
rect 16764 3000 16816 3009
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 18328 3043 18380 3052
rect 18328 3009 18346 3043
rect 18346 3009 18380 3043
rect 18328 3000 18380 3009
rect 19156 3043 19208 3052
rect 19156 3009 19165 3043
rect 19165 3009 19199 3043
rect 19199 3009 19208 3043
rect 19156 3000 19208 3009
rect 20444 3043 20496 3052
rect 20444 3009 20478 3043
rect 20478 3009 20496 3043
rect 20444 3000 20496 3009
rect 21916 3043 21968 3052
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 21916 3000 21968 3009
rect 22928 3043 22980 3052
rect 22928 3009 22937 3043
rect 22937 3009 22971 3043
rect 22971 3009 22980 3043
rect 22928 3000 22980 3009
rect 23572 3000 23624 3052
rect 24124 3043 24176 3052
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 24952 3043 25004 3052
rect 24952 3009 24961 3043
rect 24961 3009 24995 3043
rect 24995 3009 25004 3043
rect 24952 3000 25004 3009
rect 26424 3136 26476 3188
rect 27160 3136 27212 3188
rect 28816 3136 28868 3188
rect 30288 3179 30340 3188
rect 30288 3145 30297 3179
rect 30297 3145 30331 3179
rect 30331 3145 30340 3179
rect 30288 3136 30340 3145
rect 32496 3136 32548 3188
rect 34888 3136 34940 3188
rect 36360 3136 36412 3188
rect 38476 3136 38528 3188
rect 25872 3068 25924 3120
rect 17592 2932 17644 2984
rect 17960 2932 18012 2984
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 18696 2907 18748 2916
rect 18696 2873 18705 2907
rect 18705 2873 18739 2907
rect 18739 2873 18748 2907
rect 18696 2864 18748 2873
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 19800 2932 19852 2984
rect 20352 2975 20404 2984
rect 20352 2941 20361 2975
rect 20361 2941 20395 2975
rect 20395 2941 20404 2975
rect 20352 2932 20404 2941
rect 21364 2932 21416 2984
rect 27344 3043 27396 3052
rect 27344 3009 27353 3043
rect 27353 3009 27387 3043
rect 27387 3009 27396 3043
rect 27344 3000 27396 3009
rect 29460 3068 29512 3120
rect 31852 3068 31904 3120
rect 39120 3136 39172 3188
rect 40408 3179 40460 3188
rect 40408 3145 40417 3179
rect 40417 3145 40451 3179
rect 40451 3145 40460 3179
rect 40408 3136 40460 3145
rect 41144 3179 41196 3188
rect 41144 3145 41153 3179
rect 41153 3145 41187 3179
rect 41187 3145 41196 3179
rect 41144 3136 41196 3145
rect 41604 3179 41656 3188
rect 41604 3145 41613 3179
rect 41613 3145 41647 3179
rect 41647 3145 41656 3179
rect 41604 3136 41656 3145
rect 41880 3136 41932 3188
rect 41972 3136 42024 3188
rect 39396 3068 39448 3120
rect 27620 3000 27672 3052
rect 28540 3043 28592 3052
rect 28540 3009 28574 3043
rect 28574 3009 28592 3043
rect 28540 3000 28592 3009
rect 30104 3043 30156 3052
rect 30104 3009 30113 3043
rect 30113 3009 30147 3043
rect 30147 3009 30156 3043
rect 30104 3000 30156 3009
rect 30472 3043 30524 3052
rect 30472 3009 30481 3043
rect 30481 3009 30515 3043
rect 30515 3009 30524 3043
rect 30472 3000 30524 3009
rect 30748 3043 30800 3052
rect 30748 3009 30757 3043
rect 30757 3009 30791 3043
rect 30791 3009 30800 3043
rect 30748 3000 30800 3009
rect 32404 3043 32456 3052
rect 32404 3009 32413 3043
rect 32413 3009 32447 3043
rect 32447 3009 32456 3043
rect 32404 3000 32456 3009
rect 32588 3043 32640 3052
rect 32588 3009 32597 3043
rect 32597 3009 32631 3043
rect 32631 3009 32640 3043
rect 32588 3000 32640 3009
rect 33324 3043 33376 3052
rect 33324 3009 33333 3043
rect 33333 3009 33367 3043
rect 33367 3009 33376 3043
rect 33324 3000 33376 3009
rect 33600 3043 33652 3052
rect 33600 3009 33609 3043
rect 33609 3009 33643 3043
rect 33643 3009 33652 3043
rect 33600 3000 33652 3009
rect 34244 3000 34296 3052
rect 34428 3000 34480 3052
rect 35256 3043 35308 3052
rect 35256 3009 35265 3043
rect 35265 3009 35299 3043
rect 35299 3009 35308 3043
rect 35256 3000 35308 3009
rect 38384 3043 38436 3052
rect 38384 3009 38393 3043
rect 38393 3009 38427 3043
rect 38427 3009 38436 3043
rect 38384 3000 38436 3009
rect 39120 3000 39172 3052
rect 26424 2932 26476 2984
rect 28448 2975 28500 2984
rect 19616 2864 19668 2916
rect 19800 2796 19852 2848
rect 22284 2864 22336 2916
rect 20352 2796 20404 2848
rect 21088 2796 21140 2848
rect 21456 2796 21508 2848
rect 23572 2796 23624 2848
rect 24860 2907 24912 2916
rect 24860 2873 24869 2907
rect 24869 2873 24903 2907
rect 24903 2873 24912 2907
rect 24860 2864 24912 2873
rect 26516 2864 26568 2916
rect 27160 2907 27212 2916
rect 27160 2873 27169 2907
rect 27169 2873 27203 2907
rect 27203 2873 27212 2907
rect 27160 2864 27212 2873
rect 28448 2941 28457 2975
rect 28457 2941 28491 2975
rect 28491 2941 28500 2975
rect 28448 2932 28500 2941
rect 28724 2975 28776 2984
rect 28724 2941 28733 2975
rect 28733 2941 28767 2975
rect 28767 2941 28776 2975
rect 28724 2932 28776 2941
rect 33048 2975 33100 2984
rect 33048 2941 33057 2975
rect 33057 2941 33091 2975
rect 33091 2941 33100 2975
rect 33048 2932 33100 2941
rect 33416 2975 33468 2984
rect 33416 2941 33450 2975
rect 33450 2941 33468 2975
rect 33416 2932 33468 2941
rect 35348 2975 35400 2984
rect 35348 2941 35382 2975
rect 35382 2941 35400 2975
rect 35348 2932 35400 2941
rect 35532 2975 35584 2984
rect 35532 2941 35541 2975
rect 35541 2941 35575 2975
rect 35575 2941 35584 2975
rect 35532 2932 35584 2941
rect 37188 2932 37240 2984
rect 40592 3043 40644 3052
rect 40592 3009 40601 3043
rect 40601 3009 40635 3043
rect 40635 3009 40644 3043
rect 40592 3000 40644 3009
rect 41328 3043 41380 3052
rect 41328 3009 41337 3043
rect 41337 3009 41371 3043
rect 41371 3009 41380 3043
rect 41328 3000 41380 3009
rect 41420 3043 41472 3052
rect 41420 3009 41429 3043
rect 41429 3009 41463 3043
rect 41463 3009 41472 3043
rect 41420 3000 41472 3009
rect 41972 3043 42024 3052
rect 41972 3009 41981 3043
rect 41981 3009 42015 3043
rect 42015 3009 42024 3043
rect 41972 3000 42024 3009
rect 42248 3043 42300 3052
rect 42248 3009 42257 3043
rect 42257 3009 42291 3043
rect 42291 3009 42300 3043
rect 42248 3000 42300 3009
rect 43444 3179 43496 3188
rect 43444 3145 43453 3179
rect 43453 3145 43487 3179
rect 43487 3145 43496 3179
rect 43444 3136 43496 3145
rect 39396 2932 39448 2984
rect 28172 2907 28224 2916
rect 28172 2873 28181 2907
rect 28181 2873 28215 2907
rect 28215 2873 28224 2907
rect 28172 2864 28224 2873
rect 27712 2796 27764 2848
rect 29184 2796 29236 2848
rect 29460 2839 29512 2848
rect 29460 2805 29469 2839
rect 29469 2805 29503 2839
rect 29503 2805 29512 2839
rect 29460 2796 29512 2805
rect 29736 2796 29788 2848
rect 33968 2796 34020 2848
rect 34152 2796 34204 2848
rect 34704 2864 34756 2916
rect 37004 2864 37056 2916
rect 40960 2864 41012 2916
rect 42892 2864 42944 2916
rect 38292 2796 38344 2848
rect 38568 2796 38620 2848
rect 43076 2839 43128 2848
rect 43076 2805 43085 2839
rect 43085 2805 43119 2839
rect 43119 2805 43128 2839
rect 43076 2796 43128 2805
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 13918 2694 13970 2746
rect 13982 2694 14034 2746
rect 14046 2694 14098 2746
rect 14110 2694 14162 2746
rect 14174 2694 14226 2746
rect 14238 2694 14290 2746
rect 19918 2694 19970 2746
rect 19982 2694 20034 2746
rect 20046 2694 20098 2746
rect 20110 2694 20162 2746
rect 20174 2694 20226 2746
rect 20238 2694 20290 2746
rect 25918 2694 25970 2746
rect 25982 2694 26034 2746
rect 26046 2694 26098 2746
rect 26110 2694 26162 2746
rect 26174 2694 26226 2746
rect 26238 2694 26290 2746
rect 31918 2694 31970 2746
rect 31982 2694 32034 2746
rect 32046 2694 32098 2746
rect 32110 2694 32162 2746
rect 32174 2694 32226 2746
rect 32238 2694 32290 2746
rect 37918 2694 37970 2746
rect 37982 2694 38034 2746
rect 38046 2694 38098 2746
rect 38110 2694 38162 2746
rect 38174 2694 38226 2746
rect 38238 2694 38290 2746
rect 7196 2592 7248 2644
rect 5908 2524 5960 2576
rect 8576 2592 8628 2644
rect 9312 2592 9364 2644
rect 9864 2592 9916 2644
rect 10324 2592 10376 2644
rect 9128 2524 9180 2576
rect 1308 2456 1360 2508
rect 3240 2456 3292 2508
rect 5724 2456 5776 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 1768 2388 1820 2440
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 3332 2363 3384 2372
rect 3332 2329 3341 2363
rect 3341 2329 3375 2363
rect 3375 2329 3384 2363
rect 3332 2320 3384 2329
rect 5724 2363 5776 2372
rect 5724 2329 5733 2363
rect 5733 2329 5767 2363
rect 5767 2329 5776 2363
rect 5724 2320 5776 2329
rect 7380 2456 7432 2508
rect 12716 2592 12768 2644
rect 12624 2524 12676 2576
rect 14096 2524 14148 2576
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7380 2320 7432 2372
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 9772 2388 9824 2440
rect 9404 2320 9456 2372
rect 10048 2397 10057 2430
rect 10057 2397 10091 2430
rect 10091 2397 10100 2430
rect 10048 2378 10100 2397
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 12440 2388 12492 2440
rect 11612 2320 11664 2372
rect 3516 2252 3568 2304
rect 4528 2252 4580 2304
rect 6920 2252 6972 2304
rect 7288 2252 7340 2304
rect 12716 2320 12768 2372
rect 14556 2388 14608 2440
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 12900 2252 12952 2304
rect 13544 2295 13596 2304
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 14372 2363 14424 2372
rect 14372 2329 14381 2363
rect 14381 2329 14415 2363
rect 14415 2329 14424 2363
rect 14372 2320 14424 2329
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 18696 2592 18748 2644
rect 18788 2592 18840 2644
rect 20352 2592 20404 2644
rect 21272 2592 21324 2644
rect 21364 2635 21416 2644
rect 21364 2601 21373 2635
rect 21373 2601 21407 2635
rect 21407 2601 21416 2635
rect 21364 2592 21416 2601
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 17500 2320 17552 2372
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 20352 2320 20404 2372
rect 20536 2388 20588 2440
rect 24032 2592 24084 2644
rect 22376 2499 22428 2508
rect 22376 2465 22385 2499
rect 22385 2465 22419 2499
rect 22419 2465 22428 2499
rect 22376 2456 22428 2465
rect 24952 2499 25004 2508
rect 24952 2465 24961 2499
rect 24961 2465 24995 2499
rect 24995 2465 25004 2499
rect 24952 2456 25004 2465
rect 14464 2252 14516 2304
rect 15292 2252 15344 2304
rect 16580 2252 16632 2304
rect 17684 2252 17736 2304
rect 18052 2252 18104 2304
rect 22468 2320 22520 2372
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 26332 2592 26384 2644
rect 28172 2635 28224 2644
rect 28172 2601 28181 2635
rect 28181 2601 28215 2635
rect 28215 2601 28224 2635
rect 28172 2592 28224 2601
rect 28724 2592 28776 2644
rect 28816 2592 28868 2644
rect 30104 2592 30156 2644
rect 25780 2456 25832 2508
rect 27068 2499 27120 2508
rect 27068 2465 27077 2499
rect 27077 2465 27111 2499
rect 27111 2465 27120 2499
rect 27068 2456 27120 2465
rect 29184 2499 29236 2508
rect 29184 2465 29193 2499
rect 29193 2465 29227 2499
rect 29227 2465 29236 2499
rect 30380 2499 30432 2508
rect 29184 2456 29236 2465
rect 30380 2465 30389 2499
rect 30389 2465 30423 2499
rect 30423 2465 30432 2499
rect 30380 2456 30432 2465
rect 28816 2388 28868 2440
rect 28908 2431 28960 2440
rect 28908 2397 28917 2431
rect 28917 2397 28951 2431
rect 28951 2397 28960 2431
rect 28908 2388 28960 2397
rect 22928 2320 22980 2372
rect 26424 2320 26476 2372
rect 22560 2252 22612 2304
rect 22652 2252 22704 2304
rect 31668 2592 31720 2644
rect 33508 2592 33560 2644
rect 34704 2635 34756 2644
rect 34704 2601 34713 2635
rect 34713 2601 34747 2635
rect 34747 2601 34756 2635
rect 34704 2592 34756 2601
rect 35624 2592 35676 2644
rect 42800 2524 42852 2576
rect 43444 2567 43496 2576
rect 43444 2533 43453 2567
rect 43453 2533 43487 2567
rect 43487 2533 43496 2567
rect 43444 2524 43496 2533
rect 31116 2456 31168 2508
rect 32128 2499 32180 2508
rect 32128 2465 32137 2499
rect 32137 2465 32171 2499
rect 32171 2465 32180 2499
rect 32128 2456 32180 2465
rect 33784 2456 33836 2508
rect 39304 2456 39356 2508
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 34428 2388 34480 2440
rect 35348 2388 35400 2440
rect 35440 2431 35492 2440
rect 35440 2397 35449 2431
rect 35449 2397 35483 2431
rect 35483 2397 35492 2431
rect 35440 2388 35492 2397
rect 35992 2388 36044 2440
rect 36544 2431 36596 2440
rect 36544 2397 36553 2431
rect 36553 2397 36587 2431
rect 36587 2397 36596 2431
rect 36544 2388 36596 2397
rect 32128 2252 32180 2304
rect 36912 2320 36964 2372
rect 33968 2295 34020 2304
rect 33968 2261 33977 2295
rect 33977 2261 34011 2295
rect 34011 2261 34020 2295
rect 33968 2252 34020 2261
rect 39488 2252 39540 2304
rect 42892 2252 42944 2304
rect 43076 2295 43128 2304
rect 43076 2261 43085 2295
rect 43085 2261 43119 2295
rect 43119 2261 43128 2295
rect 43076 2252 43128 2261
rect 2658 2150 2710 2202
rect 2722 2150 2774 2202
rect 2786 2150 2838 2202
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 8658 2150 8710 2202
rect 8722 2150 8774 2202
rect 8786 2150 8838 2202
rect 8850 2150 8902 2202
rect 8914 2150 8966 2202
rect 8978 2150 9030 2202
rect 14658 2150 14710 2202
rect 14722 2150 14774 2202
rect 14786 2150 14838 2202
rect 14850 2150 14902 2202
rect 14914 2150 14966 2202
rect 14978 2150 15030 2202
rect 20658 2150 20710 2202
rect 20722 2150 20774 2202
rect 20786 2150 20838 2202
rect 20850 2150 20902 2202
rect 20914 2150 20966 2202
rect 20978 2150 21030 2202
rect 26658 2150 26710 2202
rect 26722 2150 26774 2202
rect 26786 2150 26838 2202
rect 26850 2150 26902 2202
rect 26914 2150 26966 2202
rect 26978 2150 27030 2202
rect 32658 2150 32710 2202
rect 32722 2150 32774 2202
rect 32786 2150 32838 2202
rect 32850 2150 32902 2202
rect 32914 2150 32966 2202
rect 32978 2150 33030 2202
rect 38658 2150 38710 2202
rect 38722 2150 38774 2202
rect 38786 2150 38838 2202
rect 38850 2150 38902 2202
rect 38914 2150 38966 2202
rect 38978 2150 39030 2202
rect 9864 2048 9916 2100
rect 13176 2048 13228 2100
rect 17500 2048 17552 2100
rect 19156 2048 19208 2100
rect 19432 2048 19484 2100
rect 30012 2048 30064 2100
rect 32772 2048 32824 2100
rect 35808 2048 35860 2100
rect 4804 1980 4856 2032
rect 11336 1980 11388 2032
rect 15660 1980 15712 2032
rect 4068 1912 4120 1964
rect 11152 1912 11204 1964
rect 9772 1844 9824 1896
rect 10600 1844 10652 1896
rect 5172 1776 5224 1828
rect 13544 1912 13596 1964
rect 15476 1912 15528 1964
rect 21088 1912 21140 1964
rect 11796 1844 11848 1896
rect 19984 1844 20036 1896
rect 13084 1776 13136 1828
rect 24400 1844 24452 1896
rect 29000 1980 29052 2032
rect 29092 1912 29144 1964
rect 33048 1980 33100 2032
rect 36912 1980 36964 2032
rect 20168 1776 20220 1828
rect 24584 1776 24636 1828
rect 37832 1912 37884 1964
rect 6552 1708 6604 1760
rect 13452 1708 13504 1760
rect 17040 1708 17092 1760
rect 32312 1708 32364 1760
rect 39396 1776 39448 1828
rect 9404 1640 9456 1692
rect 17592 1640 17644 1692
rect 17776 1640 17828 1692
rect 22652 1640 22704 1692
rect 25044 1640 25096 1692
rect 35716 1640 35768 1692
rect 35900 1708 35952 1760
rect 39672 1708 39724 1760
rect 37096 1640 37148 1692
rect 40040 1640 40092 1692
rect 41972 1640 42024 1692
rect 5540 1572 5592 1624
rect 1676 1504 1728 1556
rect 12348 1504 12400 1556
rect 14464 1572 14516 1624
rect 17408 1572 17460 1624
rect 22008 1572 22060 1624
rect 16212 1504 16264 1556
rect 10600 1436 10652 1488
rect 25228 1504 25280 1556
rect 32036 1504 32088 1556
rect 34060 1504 34112 1556
rect 19616 1436 19668 1488
rect 22100 1436 22152 1488
rect 34428 1436 34480 1488
rect 4988 1300 5040 1352
rect 9956 1300 10008 1352
rect 11704 1300 11756 1352
rect 4436 1232 4488 1284
rect 15108 1232 15160 1284
rect 28356 1368 28408 1420
rect 39120 1504 39172 1556
rect 37280 1436 37332 1488
rect 42248 1436 42300 1488
rect 20076 1232 20128 1284
rect 21916 1232 21968 1284
rect 22008 1232 22060 1284
rect 28080 1232 28132 1284
rect 11704 1164 11756 1216
rect 12808 1164 12860 1216
rect 19156 1164 19208 1216
rect 23756 1164 23808 1216
rect 4620 1096 4672 1148
rect 23480 1096 23532 1148
rect 8484 1028 8536 1080
rect 15476 1028 15528 1080
rect 15568 1028 15620 1080
rect 30840 1096 30892 1148
rect 33324 1232 33376 1284
rect 34428 1300 34480 1352
rect 40592 1368 40644 1420
rect 40408 1300 40460 1352
rect 41420 1300 41472 1352
rect 39212 1232 39264 1284
rect 43260 1232 43312 1284
rect 38016 1164 38068 1216
rect 42156 1164 42208 1216
rect 35900 1096 35952 1148
rect 36820 1096 36872 1148
rect 39580 1096 39632 1148
rect 23664 1028 23716 1080
rect 29000 1028 29052 1080
rect 29644 1028 29696 1080
rect 38384 1028 38436 1080
rect 6276 960 6328 1012
rect 27436 960 27488 1012
rect 11520 892 11572 944
rect 29552 892 29604 944
rect 13728 824 13780 876
rect 26240 824 26292 876
rect 6092 756 6144 808
rect 39304 756 39356 808
rect 1584 688 1636 740
rect 37464 688 37516 740
rect 2504 620 2556 672
rect 36452 620 36504 672
rect 10784 552 10836 604
rect 21824 552 21876 604
rect 23480 552 23532 604
rect 33140 552 33192 604
rect 3792 484 3844 536
rect 14464 484 14516 536
rect 16672 484 16724 536
rect 22008 484 22060 536
rect 35716 484 35768 536
rect 42616 484 42668 536
rect 4896 416 4948 468
rect 19064 416 19116 468
rect 7104 348 7156 400
rect 15568 348 15620 400
rect 30932 348 30984 400
rect 42064 348 42116 400
rect 28540 280 28592 332
rect 40040 280 40092 332
rect 24952 212 25004 264
rect 37280 212 37332 264
rect 27344 144 27396 196
rect 41328 144 41380 196
rect 15200 76 15252 128
rect 21180 76 21232 128
rect 26148 76 26200 128
rect 42524 76 42576 128
<< metal2 >>
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 3422 9888 3478 9897
rect 3422 9823 3478 9832
rect 3054 9616 3110 9625
rect 3054 9551 3110 9560
rect 1398 9344 1454 9353
rect 1398 9279 1454 9288
rect 1412 8498 1440 9279
rect 2318 8800 2374 8809
rect 2318 8735 2374 8744
rect 1674 8528 1730 8537
rect 1400 8492 1452 8498
rect 1674 8463 1730 8472
rect 1400 8434 1452 8440
rect 1490 7984 1546 7993
rect 1490 7919 1546 7928
rect 1504 7886 1532 7919
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1688 7818 1716 8463
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 2332 7886 2360 8735
rect 2656 8732 3032 8741
rect 2712 8730 2736 8732
rect 2792 8730 2816 8732
rect 2872 8730 2896 8732
rect 2952 8730 2976 8732
rect 2712 8678 2722 8730
rect 2966 8678 2976 8730
rect 2712 8676 2736 8678
rect 2792 8676 2816 8678
rect 2872 8676 2896 8678
rect 2952 8676 2976 8678
rect 2656 8667 3032 8676
rect 3068 8514 3096 9551
rect 3330 9480 3386 9489
rect 3330 9415 3386 9424
rect 3146 9072 3202 9081
rect 3146 9007 3202 9016
rect 2976 8486 3096 8514
rect 2976 7886 3004 8486
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 3068 8090 3096 8191
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2320 7880 2372 7886
rect 2964 7880 3016 7886
rect 2320 7822 2372 7828
rect 2410 7848 2466 7857
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 2056 7546 2084 7822
rect 2964 7822 3016 7828
rect 2410 7783 2412 7792
rect 2464 7783 2466 7792
rect 2412 7754 2464 7760
rect 2656 7644 3032 7653
rect 2712 7642 2736 7644
rect 2792 7642 2816 7644
rect 2872 7642 2896 7644
rect 2952 7642 2976 7644
rect 2712 7590 2722 7642
rect 2966 7590 2976 7642
rect 2712 7588 2736 7590
rect 2792 7588 2816 7590
rect 2872 7588 2896 7590
rect 2952 7588 2976 7590
rect 2656 7579 3032 7588
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 3068 7478 3096 7919
rect 3160 7478 3188 9007
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8498 3280 8774
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3344 8430 3372 9415
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3436 7818 3464 9823
rect 4160 9784 4212 9790
rect 4160 9726 4212 9732
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3528 8362 3556 9046
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3238 7576 3294 7585
rect 3238 7511 3294 7520
rect 3056 7472 3108 7478
rect 2318 7440 2374 7449
rect 2962 7440 3018 7449
rect 2318 7375 2374 7384
rect 2412 7404 2464 7410
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1308 7268 1360 7274
rect 1308 7210 1360 7216
rect 1320 2514 1348 7210
rect 1412 7177 1440 7278
rect 1398 7168 1454 7177
rect 1398 7103 1454 7112
rect 1398 6896 1454 6905
rect 1398 6831 1400 6840
rect 1452 6831 1454 6840
rect 1400 6802 1452 6808
rect 1490 6624 1546 6633
rect 1490 6559 1546 6568
rect 1398 6080 1454 6089
rect 1398 6015 1454 6024
rect 1412 4622 1440 6015
rect 1504 5710 1532 6559
rect 1780 6322 1808 7278
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 2332 6798 2360 7375
rect 3056 7414 3108 7420
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3252 7410 3280 7511
rect 2962 7375 3018 7384
rect 3240 7404 3292 7410
rect 2412 7346 2464 7352
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1688 5896 1716 6258
rect 2240 6236 2268 6666
rect 2318 6352 2374 6361
rect 2424 6338 2452 7346
rect 2976 7324 3004 7375
rect 3240 7346 3292 7352
rect 2976 7296 3188 7324
rect 3344 7313 3372 7754
rect 3056 6792 3108 6798
rect 3160 6780 3188 7296
rect 3330 7304 3386 7313
rect 3330 7239 3386 7248
rect 3422 6896 3478 6905
rect 3422 6831 3478 6840
rect 3240 6792 3292 6798
rect 3160 6752 3240 6780
rect 3056 6734 3108 6740
rect 3240 6734 3292 6740
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6361 2544 6598
rect 2656 6556 3032 6565
rect 2712 6554 2736 6556
rect 2792 6554 2816 6556
rect 2872 6554 2896 6556
rect 2952 6554 2976 6556
rect 2712 6502 2722 6554
rect 2966 6502 2976 6554
rect 2712 6500 2736 6502
rect 2792 6500 2816 6502
rect 2872 6500 2896 6502
rect 2952 6500 2976 6502
rect 2656 6491 3032 6500
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2374 6310 2452 6338
rect 2502 6352 2558 6361
rect 2318 6287 2374 6296
rect 2502 6287 2558 6296
rect 2792 6254 2820 6394
rect 3068 6338 3096 6734
rect 3330 6488 3386 6497
rect 3436 6458 3464 6831
rect 3620 6458 3648 8434
rect 4172 8294 4200 9726
rect 4344 9308 4396 9314
rect 4344 9250 4396 9256
rect 4356 8498 4384 9250
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3804 8078 4292 8106
rect 3804 7954 3832 8078
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3790 6488 3846 6497
rect 3330 6423 3386 6432
rect 3424 6452 3476 6458
rect 2976 6322 3280 6338
rect 2964 6316 3280 6322
rect 3016 6310 3280 6316
rect 2964 6258 3016 6264
rect 2412 6248 2464 6254
rect 2240 6208 2360 6236
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 1688 5868 1808 5896
rect 1674 5808 1730 5817
rect 1780 5778 1808 5868
rect 1674 5743 1730 5752
rect 1768 5772 1820 5778
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1490 4992 1546 5001
rect 1490 4927 1546 4936
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1412 3534 1440 4383
rect 1504 4214 1532 4927
rect 1492 4208 1544 4214
rect 1492 4150 1544 4156
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3913 1532 4014
rect 1490 3904 1546 3913
rect 1490 3839 1546 3848
rect 1596 3641 1624 5170
rect 1688 4622 1716 5743
rect 1768 5714 1820 5720
rect 1780 5137 1808 5714
rect 2332 5710 2360 6208
rect 2412 6190 2464 6196
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2424 5386 2452 6190
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2516 5545 2544 5578
rect 2792 5556 2820 6190
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3068 5914 3096 6122
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3252 5778 3280 6310
rect 3344 6118 3372 6423
rect 3424 6394 3476 6400
rect 3608 6452 3660 6458
rect 3790 6423 3846 6432
rect 3608 6394 3660 6400
rect 3804 6322 3832 6423
rect 3608 6316 3660 6322
rect 3516 6282 3568 6288
rect 3608 6258 3660 6264
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3422 6216 3478 6225
rect 3516 6224 3568 6230
rect 3422 6151 3478 6160
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3436 5846 3464 6151
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3238 5672 3294 5681
rect 3528 5658 3556 6224
rect 3620 6089 3648 6258
rect 3606 6080 3662 6089
rect 3606 6015 3662 6024
rect 3896 5760 3924 7890
rect 4080 7449 4108 7958
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4066 7440 4122 7449
rect 4066 7375 4122 7384
rect 4172 7342 4200 7822
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3988 6769 4016 6870
rect 3974 6760 4030 6769
rect 3974 6695 4030 6704
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3974 6080 4030 6089
rect 3974 6015 4030 6024
rect 3804 5732 3924 5760
rect 3238 5607 3294 5616
rect 3424 5636 3476 5642
rect 2502 5536 2558 5545
rect 2792 5528 3096 5556
rect 2502 5471 2558 5480
rect 2656 5468 3032 5477
rect 2712 5466 2736 5468
rect 2792 5466 2816 5468
rect 2872 5466 2896 5468
rect 2952 5466 2976 5468
rect 2712 5414 2722 5466
rect 2966 5414 2976 5466
rect 2712 5412 2736 5414
rect 2792 5412 2816 5414
rect 2872 5412 2896 5414
rect 2952 5412 2976 5414
rect 2656 5403 3032 5412
rect 2424 5358 2544 5386
rect 2516 5234 2544 5358
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 1766 5128 1822 5137
rect 1766 5063 1822 5072
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 1858 4720 1914 4729
rect 1858 4655 1914 4664
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1872 4214 1900 4655
rect 2042 4584 2098 4593
rect 2042 4519 2044 4528
rect 2096 4519 2098 4528
rect 2044 4490 2096 4496
rect 2424 4282 2452 5170
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2596 4616 2648 4622
rect 2700 4604 2728 5102
rect 2792 4622 2820 5306
rect 3068 5166 3096 5528
rect 3146 5536 3202 5545
rect 3146 5471 3202 5480
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3160 5098 3188 5471
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 2648 4576 2728 4604
rect 2780 4616 2832 4622
rect 2596 4558 2648 4564
rect 2780 4558 2832 4564
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1860 4208 1912 4214
rect 2228 4208 2280 4214
rect 1860 4150 1912 4156
rect 2226 4176 2228 4185
rect 2280 4176 2282 4185
rect 2226 4111 2282 4120
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3738 1808 3878
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 2516 3641 2544 4422
rect 2656 4380 3032 4389
rect 2712 4378 2736 4380
rect 2792 4378 2816 4380
rect 2872 4378 2896 4380
rect 2952 4378 2976 4380
rect 2712 4326 2722 4378
rect 2966 4326 2976 4378
rect 2712 4324 2736 4326
rect 2792 4324 2816 4326
rect 2872 4324 2896 4326
rect 2952 4324 2976 4326
rect 2656 4315 3032 4324
rect 3068 4214 3096 4558
rect 3148 4548 3200 4554
rect 3148 4490 3200 4496
rect 3160 4282 3188 4490
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 2502 3632 2558 3641
rect 2502 3567 2558 3576
rect 1400 3528 1452 3534
rect 2608 3482 2636 3878
rect 2700 3534 2728 3878
rect 3068 3738 3096 3946
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 1400 3470 1452 3476
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2516 3454 2636 3482
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1676 3392 1728 3398
rect 1872 3369 1900 3402
rect 1676 3334 1728 3340
rect 1858 3360 1914 3369
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2553 1440 2926
rect 1398 2544 1454 2553
rect 1308 2508 1360 2514
rect 1398 2479 1454 2488
rect 1308 2450 1360 2456
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 2281 1440 2382
rect 1398 2272 1454 2281
rect 1398 2207 1454 2216
rect 1596 746 1624 3334
rect 1688 1562 1716 3334
rect 1858 3295 1914 3304
rect 2240 3233 2268 3402
rect 2226 3224 2282 3233
rect 2226 3159 2282 3168
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 1780 2009 1808 2382
rect 1766 2000 1822 2009
rect 1766 1935 1822 1944
rect 2332 1578 2360 2994
rect 1676 1556 1728 1562
rect 1676 1498 1728 1504
rect 2148 1550 2360 1578
rect 2148 800 2176 1550
rect 2424 1465 2452 3402
rect 2516 3040 2544 3454
rect 2976 3448 3004 3674
rect 2976 3420 3096 3448
rect 2656 3292 3032 3301
rect 2712 3290 2736 3292
rect 2792 3290 2816 3292
rect 2872 3290 2896 3292
rect 2952 3290 2976 3292
rect 2712 3238 2722 3290
rect 2966 3238 2976 3290
rect 2712 3236 2736 3238
rect 2792 3236 2816 3238
rect 2872 3236 2896 3238
rect 2952 3236 2976 3238
rect 2656 3227 3032 3236
rect 3068 3126 3096 3420
rect 2780 3120 2832 3126
rect 2778 3088 2780 3097
rect 3056 3120 3108 3126
rect 2832 3088 2834 3097
rect 2516 3012 2636 3040
rect 3056 3062 3108 3068
rect 2778 3023 2834 3032
rect 2502 2952 2558 2961
rect 2502 2887 2504 2896
rect 2556 2887 2558 2896
rect 2504 2858 2556 2864
rect 2608 2292 2636 3012
rect 3252 2514 3280 5607
rect 3528 5630 3740 5658
rect 3424 5578 3476 5584
rect 3436 5273 3464 5578
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3422 5264 3478 5273
rect 3422 5199 3478 5208
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 4826 3464 5034
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3344 4146 3372 4626
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3528 3097 3556 5510
rect 3620 4690 3648 5510
rect 3712 5409 3740 5630
rect 3698 5400 3754 5409
rect 3698 5335 3754 5344
rect 3712 5234 3740 5335
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3712 3670 3740 4762
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3514 3088 3570 3097
rect 3514 3023 3570 3032
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 2516 2264 2636 2292
rect 2410 1456 2466 1465
rect 2410 1391 2466 1400
rect 1584 740 1636 746
rect 1584 682 1636 688
rect 2134 0 2190 800
rect 2516 678 2544 2264
rect 2656 2204 3032 2213
rect 2712 2202 2736 2204
rect 2792 2202 2816 2204
rect 2872 2202 2896 2204
rect 2952 2202 2976 2204
rect 2712 2150 2722 2202
rect 2966 2150 2976 2202
rect 2712 2148 2736 2150
rect 2792 2148 2816 2150
rect 2872 2148 2896 2150
rect 2952 2148 2976 2150
rect 2656 2139 3032 2148
rect 3344 1737 3372 2314
rect 3516 2304 3568 2310
rect 3436 2264 3516 2292
rect 3330 1728 3386 1737
rect 3330 1663 3386 1672
rect 3436 1170 3464 2264
rect 3516 2246 3568 2252
rect 3344 1142 3464 1170
rect 3344 800 3372 1142
rect 2504 672 2556 678
rect 2504 614 2556 620
rect 3330 0 3386 800
rect 3804 542 3832 5732
rect 3884 5228 3936 5234
rect 3988 5216 4016 6015
rect 3936 5188 4016 5216
rect 3884 5170 3936 5176
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 1193 3924 3878
rect 4080 3670 4108 6666
rect 4172 5545 4200 7278
rect 4264 5710 4292 8078
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7721 4384 7822
rect 4342 7712 4398 7721
rect 4342 7647 4398 7656
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4158 5536 4214 5545
rect 4158 5471 4214 5480
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3882 1184 3938 1193
rect 3882 1119 3938 1128
rect 3988 921 4016 3402
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 1970 4108 2382
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4356 1329 4384 6802
rect 4448 5914 4476 10746
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 4540 6186 4568 9454
rect 4712 9240 4764 9246
rect 4712 9182 4764 9188
rect 4724 8498 4752 9182
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4632 5914 4660 6734
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4618 5808 4674 5817
rect 4528 5772 4580 5778
rect 4618 5743 4620 5752
rect 4528 5714 4580 5720
rect 4672 5743 4674 5752
rect 4620 5714 4672 5720
rect 4540 5302 4568 5714
rect 4724 5574 4752 7822
rect 4816 5681 4844 8774
rect 4908 8294 4936 8842
rect 5092 8498 5120 10678
rect 5170 10450 5226 11250
rect 5446 10450 5502 11250
rect 5722 10450 5778 11250
rect 5998 10450 6054 11250
rect 6274 10450 6330 11250
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4986 8392 5042 8401
rect 4986 8327 5042 8336
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4802 5672 4858 5681
rect 4802 5607 4858 5616
rect 4712 5568 4764 5574
rect 4908 5556 4936 6870
rect 4712 5510 4764 5516
rect 4816 5528 4936 5556
rect 4816 5370 4844 5528
rect 4804 5364 4856 5370
rect 5000 5352 5028 8327
rect 5078 8120 5134 8129
rect 5078 8055 5134 8064
rect 5092 7290 5120 8055
rect 5184 7750 5212 10450
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 8294 5304 9522
rect 5354 8392 5410 8401
rect 5354 8327 5410 8336
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5172 7744 5224 7750
rect 5264 7744 5316 7750
rect 5172 7686 5224 7692
rect 5262 7712 5264 7721
rect 5368 7732 5396 8327
rect 5460 8090 5488 10450
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5644 8498 5672 9114
rect 5736 9110 5764 10450
rect 5816 9852 5868 9858
rect 5816 9794 5868 9800
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5828 8362 5856 9794
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5446 7984 5502 7993
rect 5446 7919 5502 7928
rect 5460 7818 5488 7919
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5316 7712 5396 7732
rect 5318 7704 5396 7712
rect 5262 7647 5318 7656
rect 5460 7562 5488 7754
rect 5368 7534 5488 7562
rect 5368 7410 5396 7534
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5552 7342 5580 8298
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5540 7336 5592 7342
rect 5092 7262 5212 7290
rect 5540 7278 5592 7284
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6934 5120 7142
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5184 6866 5212 7262
rect 5538 6896 5594 6905
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5356 6860 5408 6866
rect 5644 6866 5672 7958
rect 5736 7410 5764 7958
rect 5814 7712 5870 7721
rect 5814 7647 5870 7656
rect 5828 7410 5856 7647
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5538 6831 5540 6840
rect 5356 6802 5408 6808
rect 5592 6831 5594 6840
rect 5632 6860 5684 6866
rect 5540 6802 5592 6808
rect 5632 6802 5684 6808
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5184 5817 5212 6258
rect 5368 6089 5396 6802
rect 5736 6322 5764 7346
rect 5920 6458 5948 9590
rect 6012 8566 6040 10450
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6104 8498 6132 8910
rect 6196 8498 6224 9046
rect 6288 8634 6316 10450
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 8090 6132 8230
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6380 7954 6408 10610
rect 6550 10450 6606 11250
rect 6826 10450 6882 11250
rect 7102 10450 7158 11250
rect 7378 10450 7434 11250
rect 7654 10450 7710 11250
rect 7930 10450 7986 11250
rect 8206 10450 8262 11250
rect 8482 10450 8538 11250
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 8090 6500 9862
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6564 7970 6592 10450
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 8634 6684 9998
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6368 7948 6420 7954
rect 6564 7942 6684 7970
rect 6368 7890 6420 7896
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5828 6338 5856 6394
rect 5724 6316 5776 6322
rect 5828 6310 5948 6338
rect 5724 6258 5776 6264
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5354 6080 5410 6089
rect 5354 6015 5410 6024
rect 5368 5846 5396 6015
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5356 5840 5408 5846
rect 5170 5808 5226 5817
rect 5356 5782 5408 5788
rect 5170 5743 5226 5752
rect 5262 5672 5318 5681
rect 5262 5607 5318 5616
rect 4804 5306 4856 5312
rect 4908 5324 5028 5352
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 4010 4476 4150
rect 4632 4146 4660 4966
rect 4816 4690 4844 5306
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4342 1320 4398 1329
rect 4448 1290 4476 3606
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4342 1255 4398 1264
rect 4436 1284 4488 1290
rect 4436 1226 4488 1232
rect 3974 912 4030 921
rect 3974 847 4030 856
rect 4540 800 4568 2246
rect 4632 1154 4660 3538
rect 4724 2990 4752 3538
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4816 2038 4844 4422
rect 4908 4214 4936 5324
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4804 2032 4856 2038
rect 4804 1974 4856 1980
rect 4620 1148 4672 1154
rect 4620 1090 4672 1096
rect 3792 536 3844 542
rect 3792 478 3844 484
rect 4526 0 4582 800
rect 4908 474 4936 2382
rect 5000 1358 5028 5170
rect 5080 4480 5132 4486
rect 5078 4448 5080 4457
rect 5132 4448 5134 4457
rect 5078 4383 5134 4392
rect 5184 4282 5212 5170
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5092 3534 5120 4082
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5184 3058 5212 4218
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5276 2938 5304 5607
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4282 5396 4490
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4078 5488 5850
rect 5828 5778 5856 6190
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5540 5704 5592 5710
rect 5538 5672 5540 5681
rect 5592 5672 5594 5681
rect 5538 5607 5594 5616
rect 5722 5128 5778 5137
rect 5722 5063 5778 5072
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5184 2910 5304 2938
rect 5184 1834 5212 2910
rect 5172 1828 5224 1834
rect 5172 1770 5224 1776
rect 5552 1630 5580 4626
rect 5736 2514 5764 5063
rect 5920 4808 5948 6310
rect 6012 5778 6040 6938
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5920 4780 6040 4808
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5828 3369 5856 4626
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 5814 3360 5870 3369
rect 5814 3295 5870 3304
rect 5920 2582 5948 4218
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5540 1624 5592 1630
rect 5540 1566 5592 1572
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5736 800 5764 2314
rect 6012 1465 6040 4780
rect 5998 1456 6054 1465
rect 5998 1391 6054 1400
rect 6104 814 6132 7890
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6276 7744 6328 7750
rect 6182 7712 6238 7721
rect 6276 7686 6328 7692
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6182 7647 6238 7656
rect 6196 7410 6224 7647
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6288 5273 6316 7686
rect 6472 7342 6500 7686
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6662 6500 6734
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6380 6322 6408 6598
rect 6472 6390 6500 6598
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5846 6408 6054
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6472 5302 6500 6326
rect 6460 5296 6512 5302
rect 6274 5264 6330 5273
rect 6274 5199 6330 5208
rect 6380 5256 6460 5284
rect 6182 4720 6238 4729
rect 6182 4655 6238 4664
rect 6196 3194 6224 4655
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6288 4457 6316 4558
rect 6274 4448 6330 4457
rect 6274 4383 6330 4392
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6184 2440 6236 2446
rect 6182 2408 6184 2417
rect 6236 2408 6238 2417
rect 6182 2343 6238 2352
rect 6288 1018 6316 4383
rect 6380 2990 6408 5256
rect 6460 5238 6512 5244
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4690 6500 4966
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6564 1766 6592 7822
rect 6656 6458 6684 7942
rect 6748 7546 6776 9658
rect 6840 8294 6868 10450
rect 7116 9790 7144 10450
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7196 10192 7248 10198
rect 7196 10134 7248 10140
rect 7104 9784 7156 9790
rect 7104 9726 7156 9732
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6920 9240 6972 9246
rect 6920 9182 6972 9188
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6798 6868 7142
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6734 6488 6790 6497
rect 6644 6452 6696 6458
rect 6734 6423 6790 6432
rect 6644 6394 6696 6400
rect 6748 6338 6776 6423
rect 6656 6310 6776 6338
rect 6656 5710 6684 6310
rect 6932 5914 6960 9182
rect 7024 8129 7052 9386
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7116 8673 7144 8978
rect 7102 8664 7158 8673
rect 7102 8599 7158 8608
rect 7104 8560 7156 8566
rect 7104 8502 7156 8508
rect 7010 8120 7066 8129
rect 7010 8055 7066 8064
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7750 7052 7822
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6734 5808 6790 5817
rect 6734 5743 6736 5752
rect 6788 5743 6790 5752
rect 6736 5714 6788 5720
rect 6644 5704 6696 5710
rect 6920 5704 6972 5710
rect 6644 5646 6696 5652
rect 6840 5664 6920 5692
rect 6656 5409 6684 5646
rect 6840 5574 6868 5664
rect 6920 5646 6972 5652
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6642 5400 6698 5409
rect 6642 5335 6698 5344
rect 6656 4282 6684 5335
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6656 2446 6684 3674
rect 6748 3516 6776 4422
rect 6828 3528 6880 3534
rect 6748 3496 6828 3516
rect 6880 3496 6882 3505
rect 6748 3488 6826 3496
rect 6826 3431 6882 3440
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 6276 1012 6328 1018
rect 6276 954 6328 960
rect 6092 808 6144 814
rect 4896 468 4948 474
rect 4896 410 4948 416
rect 5722 0 5778 800
rect 6932 800 6960 2246
rect 6092 750 6144 756
rect 6918 0 6974 800
rect 7024 785 7052 7346
rect 7116 5370 7144 8502
rect 7208 8362 7236 10134
rect 7300 9466 7328 10202
rect 7392 9722 7420 10450
rect 7472 9784 7524 9790
rect 7472 9726 7524 9732
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7300 9438 7420 9466
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8498 7328 9318
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7392 8362 7420 9438
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7484 7868 7512 9726
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7300 7840 7512 7868
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7116 4826 7144 5170
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7208 4706 7236 7346
rect 7300 7274 7328 7840
rect 7378 7712 7434 7721
rect 7378 7647 7434 7656
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7300 6662 7328 6802
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7392 5846 7420 7647
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7116 4678 7236 4706
rect 7010 776 7066 785
rect 7010 711 7066 720
rect 7116 406 7144 4678
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7208 2650 7236 4490
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7300 2310 7328 4082
rect 7484 3738 7512 7346
rect 7576 5914 7604 8434
rect 7668 8362 7696 10450
rect 7840 10328 7892 10334
rect 7840 10270 7892 10276
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7654 8256 7710 8265
rect 7654 8191 7710 8200
rect 7668 7818 7696 8191
rect 7760 8090 7788 10066
rect 7852 8430 7880 10270
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7944 8276 7972 10450
rect 8116 10396 8168 10402
rect 8116 10338 8168 10344
rect 8022 9072 8078 9081
rect 8022 9007 8078 9016
rect 8036 8498 8064 9007
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8128 8362 8156 10338
rect 8220 8906 8248 10450
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8312 8430 8340 9930
rect 8496 9586 8524 10450
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8390 8936 8446 8945
rect 8390 8871 8446 8880
rect 8404 8498 8432 8871
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 7852 8248 7972 8276
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7748 7744 7800 7750
rect 7746 7712 7748 7721
rect 7800 7712 7802 7721
rect 7746 7647 7802 7656
rect 7852 7546 7880 8248
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 8496 7970 8524 8774
rect 8588 8090 8616 9658
rect 8680 8838 8708 10542
rect 8758 10450 8814 11250
rect 9034 10450 9090 11250
rect 9220 10464 9272 10470
rect 8772 9926 8800 10450
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 9048 9858 9076 10450
rect 9310 10450 9366 11250
rect 9586 10450 9642 11250
rect 9862 10450 9918 11250
rect 10138 10450 10194 11250
rect 10414 10450 10470 11250
rect 10690 10450 10746 11250
rect 10966 10450 11022 11250
rect 11152 10872 11204 10878
rect 11152 10814 11204 10820
rect 9220 10406 9272 10412
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9852 9088 9858
rect 9036 9794 9088 9800
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8656 8732 9032 8741
rect 8712 8730 8736 8732
rect 8792 8730 8816 8732
rect 8872 8730 8896 8732
rect 8952 8730 8976 8732
rect 8712 8678 8722 8730
rect 8966 8678 8976 8730
rect 8712 8676 8736 8678
rect 8792 8676 8816 8678
rect 8872 8676 8896 8678
rect 8952 8676 8976 8678
rect 8656 8667 9032 8676
rect 9140 8362 9168 9862
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8666 8120 8722 8129
rect 8576 8084 8628 8090
rect 8666 8055 8722 8064
rect 8760 8084 8812 8090
rect 8576 8026 8628 8032
rect 8220 7942 8524 7970
rect 8220 7546 8248 7942
rect 8484 7880 8536 7886
rect 8390 7848 8446 7857
rect 8680 7857 8708 8055
rect 8760 8026 8812 8032
rect 8772 7886 8800 8026
rect 8864 8022 8892 8230
rect 9232 8072 9260 10406
rect 9324 9790 9352 10450
rect 9312 9784 9364 9790
rect 9312 9726 9364 9732
rect 9496 9784 9548 9790
rect 9496 9726 9548 9732
rect 9310 9616 9366 9625
rect 9310 9551 9366 9560
rect 9324 8498 9352 9551
rect 9402 9208 9458 9217
rect 9402 9143 9458 9152
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9232 8044 9352 8072
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8944 7948 8996 7954
rect 9048 7942 9260 7970
rect 9048 7936 9076 7942
rect 8996 7908 9076 7936
rect 8944 7890 8996 7896
rect 8760 7880 8812 7886
rect 8484 7822 8536 7828
rect 8666 7848 8722 7857
rect 8390 7783 8446 7792
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7760 6984 7788 7278
rect 7852 7002 7880 7346
rect 8312 7342 8340 7686
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 8404 7041 8432 7783
rect 8390 7032 8446 7041
rect 7668 6956 7788 6984
rect 7840 6996 7892 7002
rect 7668 6440 7696 6956
rect 8390 6967 8446 6976
rect 7840 6938 7892 6944
rect 7748 6860 7800 6866
rect 7800 6820 7880 6848
rect 7748 6802 7800 6808
rect 7668 6412 7788 6440
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7668 5370 7696 6258
rect 7760 5846 7788 6412
rect 7852 6202 7880 6820
rect 8116 6792 8168 6798
rect 7944 6752 8116 6780
rect 7944 6497 7972 6752
rect 8116 6734 8168 6740
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 7930 6488 7986 6497
rect 7930 6423 7986 6432
rect 7944 6322 7972 6423
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 8220 6254 8248 6598
rect 8312 6254 8340 6666
rect 8208 6248 8260 6254
rect 7852 6174 7972 6202
rect 8208 6190 8260 6196
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 7840 6112 7892 6118
rect 7944 6100 7972 6174
rect 7944 6072 8432 6100
rect 7840 6054 7892 6060
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7852 5692 7880 6054
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 7932 5704 7984 5710
rect 7852 5664 7932 5692
rect 7932 5646 7984 5652
rect 8036 5545 8064 5782
rect 8404 5574 8432 6072
rect 8392 5568 8444 5574
rect 8022 5536 8078 5545
rect 8392 5510 8444 5516
rect 8022 5471 8078 5480
rect 8298 5400 8354 5409
rect 7656 5364 7708 5370
rect 8298 5335 8354 5344
rect 7656 5306 7708 5312
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7930 5264 7986 5273
rect 7930 5199 7986 5208
rect 7562 5128 7618 5137
rect 7562 5063 7618 5072
rect 7576 4690 7604 5063
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7392 3194 7420 3538
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7576 2774 7604 4422
rect 7484 2746 7604 2774
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7392 2378 7420 2450
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7484 649 7512 2746
rect 7668 1057 7696 5199
rect 7944 5166 7972 5199
rect 8312 5166 8340 5335
rect 7932 5160 7984 5166
rect 7746 5128 7802 5137
rect 7932 5102 7984 5108
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 7746 5063 7802 5072
rect 7760 4554 7788 5063
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 8404 4282 8432 5510
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8390 4176 8446 4185
rect 8390 4111 8446 4120
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7838 4040 7894 4049
rect 7760 3534 7788 4014
rect 7838 3975 7894 3984
rect 7852 3602 7880 3975
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7760 2446 7788 3130
rect 7852 2990 7880 3538
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7840 2984 7892 2990
rect 7944 2961 7972 3470
rect 8024 3392 8076 3398
rect 8312 3369 8340 3538
rect 8024 3334 8076 3340
rect 8298 3360 8354 3369
rect 8036 3126 8064 3334
rect 8298 3295 8354 3304
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8300 2984 8352 2990
rect 7840 2926 7892 2932
rect 7930 2952 7986 2961
rect 8404 2972 8432 4111
rect 8352 2944 8432 2972
rect 8300 2926 8352 2932
rect 7930 2887 7986 2896
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7654 1048 7710 1057
rect 7654 983 7710 992
rect 7852 762 7880 2790
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 8496 1086 8524 7822
rect 8760 7822 8812 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8666 7783 8722 7792
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8588 5642 8616 7686
rect 8656 7644 9032 7653
rect 8712 7642 8736 7644
rect 8792 7642 8816 7644
rect 8872 7642 8896 7644
rect 8952 7642 8976 7644
rect 8712 7590 8722 7642
rect 8966 7590 8976 7642
rect 8712 7588 8736 7590
rect 8792 7588 8816 7590
rect 8872 7588 8896 7590
rect 8952 7588 8976 7590
rect 8656 7579 9032 7588
rect 9140 7410 9168 7822
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9232 7342 9260 7942
rect 9324 7546 9352 8044
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9324 6984 9352 7346
rect 9232 6956 9352 6984
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 8656 6556 9032 6565
rect 8712 6554 8736 6556
rect 8792 6554 8816 6556
rect 8872 6554 8896 6556
rect 8952 6554 8976 6556
rect 8712 6502 8722 6554
rect 8966 6502 8976 6554
rect 8712 6500 8736 6502
rect 8792 6500 8816 6502
rect 8872 6500 8896 6502
rect 8952 6500 8976 6502
rect 8656 6491 9032 6500
rect 9140 6458 9168 6598
rect 9232 6458 9260 6956
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9324 6497 9352 6802
rect 9310 6488 9366 6497
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9220 6452 9272 6458
rect 9310 6423 9366 6432
rect 9220 6394 9272 6400
rect 8666 6080 8722 6089
rect 8666 6015 8722 6024
rect 8680 5846 8708 6015
rect 8772 5914 8800 6394
rect 9416 6338 9444 9143
rect 9508 8362 9536 9726
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9600 7410 9628 10450
rect 9876 9994 9904 10450
rect 10152 10062 10180 10450
rect 10428 10198 10456 10450
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10704 10130 10732 10450
rect 10980 10266 11008 10450
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9772 9852 9824 9858
rect 9772 9794 9824 9800
rect 9784 7546 9812 9794
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 7290 9720 7346
rect 9600 7262 9720 7290
rect 9600 6458 9628 7262
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9692 6798 9720 7142
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 8864 6310 9444 6338
rect 8864 6254 8892 6310
rect 9784 6304 9812 7142
rect 9692 6276 9812 6304
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 9140 6174 9352 6202
rect 8944 6112 8996 6118
rect 9140 6100 9168 6174
rect 8996 6072 9168 6100
rect 9220 6112 9272 6118
rect 8944 6054 8996 6060
rect 9220 6054 9272 6060
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8656 5468 9032 5477
rect 8712 5466 8736 5468
rect 8792 5466 8816 5468
rect 8872 5466 8896 5468
rect 8952 5466 8976 5468
rect 8712 5414 8722 5466
rect 8966 5414 8976 5466
rect 8712 5412 8736 5414
rect 8792 5412 8816 5414
rect 8872 5412 8896 5414
rect 8952 5412 8976 5414
rect 8656 5403 9032 5412
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8588 4826 8616 5034
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8680 4468 8708 5306
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9034 4856 9090 4865
rect 9140 4826 9168 5170
rect 9034 4791 9090 4800
rect 9128 4820 9180 4826
rect 9048 4758 9076 4791
rect 9128 4762 9180 4768
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8588 4440 8708 4468
rect 8588 4078 8616 4440
rect 8656 4380 9032 4389
rect 8712 4378 8736 4380
rect 8792 4378 8816 4380
rect 8872 4378 8896 4380
rect 8952 4378 8976 4380
rect 8712 4326 8722 4378
rect 8966 4326 8976 4378
rect 8712 4324 8736 4326
rect 8792 4324 8816 4326
rect 8872 4324 8896 4326
rect 8952 4324 8976 4326
rect 8656 4315 9032 4324
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8588 3074 8616 3538
rect 8864 3398 8892 4014
rect 8956 3777 8984 4014
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 8956 3602 8984 3703
rect 9126 3632 9182 3641
rect 8944 3596 8996 3602
rect 9126 3567 9182 3576
rect 8944 3538 8996 3544
rect 8852 3392 8904 3398
rect 9140 3369 9168 3567
rect 8852 3334 8904 3340
rect 9126 3360 9182 3369
rect 8656 3292 9032 3301
rect 9126 3295 9182 3304
rect 8712 3290 8736 3292
rect 8792 3290 8816 3292
rect 8872 3290 8896 3292
rect 8952 3290 8976 3292
rect 8712 3238 8722 3290
rect 8966 3238 8976 3290
rect 8712 3236 8736 3238
rect 8792 3236 8816 3238
rect 8872 3236 8896 3238
rect 8952 3236 8976 3238
rect 8656 3227 9032 3236
rect 9126 3224 9182 3233
rect 8956 3168 9126 3176
rect 8956 3159 9182 3168
rect 8956 3148 9168 3159
rect 8588 3046 8708 3074
rect 8680 2990 8708 3046
rect 8956 2990 8984 3148
rect 8668 2984 8720 2990
rect 8666 2952 8668 2961
rect 8944 2984 8996 2990
rect 8720 2952 8722 2961
rect 8576 2916 8628 2922
rect 8944 2926 8996 2932
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 8666 2887 8722 2896
rect 8576 2858 8628 2864
rect 8588 2650 8616 2858
rect 8956 2825 8984 2926
rect 8942 2816 8998 2825
rect 8942 2751 8998 2760
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 9140 2582 9168 2926
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 8656 2204 9032 2213
rect 8712 2202 8736 2204
rect 8792 2202 8816 2204
rect 8872 2202 8896 2204
rect 8952 2202 8976 2204
rect 8712 2150 8722 2202
rect 8966 2150 8976 2202
rect 8712 2148 8736 2150
rect 8792 2148 8816 2150
rect 8872 2148 8896 2150
rect 8952 2148 8976 2150
rect 8656 2139 9032 2148
rect 9232 1601 9260 6054
rect 9324 5166 9352 6174
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9324 4826 9352 5102
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9402 4312 9458 4321
rect 9402 4247 9458 4256
rect 9416 4078 9444 4247
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9324 2650 9352 3946
rect 9508 3924 9536 5510
rect 9416 3896 9536 3924
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9416 2378 9444 3896
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9416 1698 9444 2314
rect 9508 2009 9536 3402
rect 9600 2281 9628 6054
rect 9692 5137 9720 6276
rect 9876 6202 9904 8774
rect 9968 8362 9996 9930
rect 10046 9888 10102 9897
rect 10046 9823 10102 9832
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 10060 7206 10088 9823
rect 10244 8362 10272 9998
rect 11072 9926 11100 10202
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10322 9344 10378 9353
rect 10322 9279 10378 9288
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10336 8090 10364 9279
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10784 8560 10836 8566
rect 10414 8528 10470 8537
rect 10784 8502 10836 8508
rect 10414 8463 10416 8472
rect 10468 8463 10470 8472
rect 10416 8434 10468 8440
rect 10600 8424 10652 8430
rect 10506 8392 10562 8401
rect 10600 8366 10652 8372
rect 10506 8327 10562 8336
rect 10520 8090 10548 8327
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9956 6792 10008 6798
rect 10008 6752 10088 6780
rect 9956 6734 10008 6740
rect 10060 6633 10088 6752
rect 10046 6624 10102 6633
rect 10046 6559 10102 6568
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9784 6174 9904 6202
rect 9784 5953 9812 6174
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9770 5944 9826 5953
rect 9770 5879 9826 5888
rect 9876 5817 9904 6054
rect 9862 5808 9918 5817
rect 9862 5743 9918 5752
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5409 9812 5646
rect 9770 5400 9826 5409
rect 9968 5370 9996 6394
rect 10060 6254 10088 6394
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 10046 5944 10102 5953
rect 10046 5879 10102 5888
rect 10060 5778 10088 5879
rect 10152 5846 10180 7686
rect 10230 7576 10286 7585
rect 10230 7511 10286 7520
rect 10244 7410 10272 7511
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 6996 10284 7002
rect 10336 6984 10364 7346
rect 10284 6956 10364 6984
rect 10416 6996 10468 7002
rect 10232 6938 10284 6944
rect 10416 6938 10468 6944
rect 10428 6905 10456 6938
rect 10414 6896 10470 6905
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10324 6860 10376 6866
rect 10414 6831 10470 6840
rect 10324 6802 10376 6808
rect 10244 6662 10272 6802
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9770 5335 9826 5344
rect 9956 5364 10008 5370
rect 9678 5128 9734 5137
rect 9678 5063 9734 5072
rect 9692 4622 9720 5063
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9784 4146 9812 5335
rect 9956 5306 10008 5312
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 9968 4690 9996 4791
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9954 4448 10010 4457
rect 9954 4383 10010 4392
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9770 3904 9826 3913
rect 9770 3839 9826 3848
rect 9784 3602 9812 3839
rect 9876 3738 9904 4082
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9862 3632 9918 3641
rect 9772 3596 9824 3602
rect 9862 3567 9918 3576
rect 9772 3538 9824 3544
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9586 2272 9642 2281
rect 9586 2207 9642 2216
rect 9494 2000 9550 2009
rect 9494 1935 9550 1944
rect 9404 1692 9456 1698
rect 9404 1634 9456 1640
rect 9218 1592 9274 1601
rect 9218 1527 9274 1536
rect 8484 1080 8536 1086
rect 8484 1022 8536 1028
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 9324 870 9444 898
rect 9324 800 9352 870
rect 7852 734 8064 762
rect 7470 640 7526 649
rect 7470 575 7526 584
rect 7104 400 7156 406
rect 7104 342 7156 348
rect 8114 0 8170 800
rect 9310 0 9366 800
rect 9416 762 9444 870
rect 9692 762 9720 3334
rect 9876 3097 9904 3567
rect 9862 3088 9918 3097
rect 9862 3023 9918 3032
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9784 1902 9812 2382
rect 9876 2106 9904 2586
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9968 1358 9996 4383
rect 10060 4078 10088 5714
rect 10244 5234 10272 6326
rect 10336 5370 10364 6802
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 6458 10548 6734
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10506 5672 10562 5681
rect 10506 5607 10562 5616
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10336 5234 10364 5306
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10322 5128 10378 5137
rect 10322 5063 10324 5072
rect 10376 5063 10378 5072
rect 10324 5034 10376 5040
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10060 2436 10088 2926
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10048 2430 10100 2436
rect 10048 2372 10100 2378
rect 9956 1352 10008 1358
rect 9956 1294 10008 1300
rect 9416 734 9720 762
rect 10152 762 10180 2790
rect 10244 1204 10272 4422
rect 10336 2990 10364 4626
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10428 3777 10456 4558
rect 10414 3768 10470 3777
rect 10414 3703 10470 3712
rect 10428 3670 10456 3703
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10520 3058 10548 5607
rect 10612 3942 10640 8366
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 6322 10732 7278
rect 10796 6798 10824 8502
rect 10876 8424 10928 8430
rect 10874 8392 10876 8401
rect 10928 8392 10930 8401
rect 10874 8327 10930 8336
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10888 6089 10916 6831
rect 10874 6080 10930 6089
rect 10874 6015 10930 6024
rect 10782 5808 10838 5817
rect 10782 5743 10784 5752
rect 10836 5743 10838 5752
rect 10784 5714 10836 5720
rect 10796 5302 10824 5714
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10784 5296 10836 5302
rect 10690 5264 10746 5273
rect 10784 5238 10836 5244
rect 10690 5199 10746 5208
rect 10704 4729 10732 5199
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10690 4720 10746 4729
rect 10690 4655 10746 4664
rect 10704 4622 10732 4655
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10796 4146 10824 4966
rect 10888 4214 10916 5510
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10980 3942 11008 9046
rect 11164 8974 11192 10814
rect 11242 10450 11298 11250
rect 11518 10464 11574 11250
rect 11518 10450 11520 10464
rect 11256 9722 11284 10450
rect 11572 10450 11574 10464
rect 11794 10450 11850 11250
rect 12070 10450 12126 11250
rect 12346 10554 12402 11250
rect 12176 10526 12402 10554
rect 11520 10406 11572 10412
rect 11808 10334 11836 10450
rect 11796 10328 11848 10334
rect 11796 10270 11848 10276
rect 11702 10024 11758 10033
rect 11702 9959 11758 9968
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11348 8838 11376 9862
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 7546 11100 8298
rect 11164 8294 11192 8434
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11348 7410 11376 8230
rect 11440 7585 11468 8366
rect 11426 7576 11482 7585
rect 11426 7511 11482 7520
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11072 6730 11100 7346
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11164 5778 11192 6734
rect 11334 6624 11390 6633
rect 11334 6559 11390 6568
rect 11242 6488 11298 6497
rect 11242 6423 11298 6432
rect 11256 6322 11284 6423
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11256 6089 11284 6258
rect 11242 6080 11298 6089
rect 11242 6015 11298 6024
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 5137 11100 5170
rect 11058 5128 11114 5137
rect 11058 5063 11114 5072
rect 11072 4486 11100 5063
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11164 4146 11192 4490
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 10600 3936 10652 3942
rect 10968 3936 11020 3942
rect 10600 3878 10652 3884
rect 10874 3904 10930 3913
rect 10968 3878 11020 3884
rect 10874 3839 10930 3848
rect 10888 3534 10916 3839
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10796 3126 10824 3470
rect 11348 3398 11376 6559
rect 11440 4622 11468 7511
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11532 6254 11560 6734
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11532 6118 11560 6190
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11532 5370 11560 5646
rect 11624 5409 11652 9046
rect 11610 5400 11666 5409
rect 11520 5364 11572 5370
rect 11610 5335 11666 5344
rect 11520 5306 11572 5312
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11532 3738 11560 3878
rect 11624 3777 11652 5238
rect 11610 3768 11666 3777
rect 11520 3732 11572 3738
rect 11610 3703 11666 3712
rect 11520 3674 11572 3680
rect 11624 3602 11652 3703
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10324 2984 10376 2990
rect 10704 2961 10732 2994
rect 10324 2926 10376 2932
rect 10690 2952 10746 2961
rect 10336 2650 10364 2926
rect 10690 2887 10746 2896
rect 10796 2774 10824 3062
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 10796 2746 10916 2774
rect 10324 2644 10376 2650
rect 10888 2632 10916 2746
rect 10324 2586 10376 2592
rect 10796 2604 10916 2632
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10612 1902 10640 2382
rect 10600 1896 10652 1902
rect 10600 1838 10652 1844
rect 10612 1494 10640 1838
rect 10600 1488 10652 1494
rect 10600 1430 10652 1436
rect 10244 1176 10732 1204
rect 10428 870 10548 898
rect 10428 762 10456 870
rect 10520 800 10548 870
rect 10152 734 10456 762
rect 10506 0 10562 800
rect 10704 490 10732 1176
rect 10796 610 10824 2604
rect 11334 2136 11390 2145
rect 11334 2071 11390 2080
rect 11348 2038 11376 2071
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11164 1873 11192 1906
rect 11150 1864 11206 1873
rect 11150 1799 11206 1808
rect 11532 950 11560 2926
rect 11624 2378 11652 3538
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11716 1358 11744 9959
rect 12084 9858 12112 10450
rect 12176 10402 12204 10526
rect 12346 10450 12402 10526
rect 12622 10450 12678 11250
rect 12898 10450 12954 11250
rect 13174 10450 13230 11250
rect 13450 10450 13506 11250
rect 13726 10450 13782 11250
rect 14002 10450 14058 11250
rect 14096 10940 14148 10946
rect 14096 10882 14148 10888
rect 12164 10396 12216 10402
rect 12164 10338 12216 10344
rect 12636 10266 12664 10450
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12072 9852 12124 9858
rect 12072 9794 12124 9800
rect 11888 9240 11940 9246
rect 11888 9182 11940 9188
rect 11794 7440 11850 7449
rect 11794 7375 11850 7384
rect 11808 6118 11836 7375
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11796 5704 11848 5710
rect 11900 5692 11928 9182
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12254 8392 12310 8401
rect 12254 8327 12310 8336
rect 12268 7886 12296 8327
rect 12256 7880 12308 7886
rect 12070 7848 12126 7857
rect 12256 7822 12308 7828
rect 12070 7783 12072 7792
rect 12124 7783 12126 7792
rect 12072 7754 12124 7760
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 6458 12020 7346
rect 12254 7304 12310 7313
rect 12254 7239 12310 7248
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11848 5664 11928 5692
rect 11796 5646 11848 5652
rect 11808 5166 11836 5646
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11808 4758 11836 5102
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11808 1902 11836 4082
rect 11900 3942 11928 5034
rect 11992 3942 12020 5850
rect 12084 5846 12112 6598
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12070 5536 12126 5545
rect 12070 5471 12126 5480
rect 12084 4729 12112 5471
rect 12070 4720 12126 4729
rect 12070 4655 12126 4664
rect 12084 4622 12112 4655
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12176 4010 12204 6870
rect 12164 4004 12216 4010
rect 12164 3946 12216 3952
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 12268 3233 12296 7239
rect 12544 6633 12572 8774
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 8288 12768 8294
rect 12820 8265 12848 8298
rect 12716 8230 12768 8236
rect 12806 8256 12862 8265
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7002 12664 7822
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12530 6624 12586 6633
rect 12530 6559 12586 6568
rect 12636 6474 12664 6938
rect 12728 6934 12756 8230
rect 12806 8191 12862 8200
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7546 12848 7686
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12636 6446 12756 6474
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12544 5658 12572 5850
rect 12452 5630 12572 5658
rect 12346 4992 12402 5001
rect 12346 4927 12402 4936
rect 12254 3224 12310 3233
rect 12254 3159 12310 3168
rect 11796 1896 11848 1902
rect 11796 1838 11848 1844
rect 12360 1562 12388 4927
rect 12452 4321 12480 5630
rect 12530 5264 12586 5273
rect 12530 5199 12586 5208
rect 12438 4312 12494 4321
rect 12438 4247 12494 4256
rect 12544 3584 12572 5199
rect 12636 4622 12664 6054
rect 12728 5778 12756 6446
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5370 12756 5714
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12728 4826 12756 5170
rect 12820 5080 12848 7278
rect 12912 5352 12940 10450
rect 13188 9722 13216 10450
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13280 7818 13308 10202
rect 13360 9852 13412 9858
rect 13360 9794 13412 9800
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 13082 7032 13138 7041
rect 13280 7018 13308 7239
rect 13082 6967 13138 6976
rect 13188 6990 13308 7018
rect 13096 5930 13124 6967
rect 13004 5902 13124 5930
rect 13188 5914 13216 6990
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13176 5908 13228 5914
rect 13004 5681 13032 5902
rect 13176 5850 13228 5856
rect 13084 5704 13136 5710
rect 12990 5672 13046 5681
rect 13084 5646 13136 5652
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12990 5607 13046 5616
rect 12992 5364 13044 5370
rect 12912 5324 12992 5352
rect 12992 5306 13044 5312
rect 13096 5216 13124 5646
rect 13004 5188 13124 5216
rect 12820 5052 12940 5080
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12820 3738 12848 4626
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12452 3556 12756 3584
rect 12452 2446 12480 3556
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 2564 12572 3334
rect 12636 3058 12664 3431
rect 12728 3398 12756 3556
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12728 2650 12756 2926
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12624 2576 12676 2582
rect 12544 2536 12624 2564
rect 12624 2518 12676 2524
rect 12440 2440 12492 2446
rect 12912 2428 12940 5052
rect 13004 4826 13032 5188
rect 13082 5128 13138 5137
rect 13082 5063 13138 5072
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13096 4457 13124 5063
rect 13082 4448 13138 4457
rect 13082 4383 13138 4392
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13004 2553 13032 3334
rect 13096 3097 13124 4082
rect 13082 3088 13138 3097
rect 13082 3023 13138 3032
rect 12990 2544 13046 2553
rect 12990 2479 13046 2488
rect 12912 2400 13032 2428
rect 12440 2382 12492 2388
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 12728 2145 12756 2314
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12714 2136 12770 2145
rect 12714 2071 12770 2080
rect 12348 1556 12400 1562
rect 12348 1498 12400 1504
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 12820 1222 12848 2246
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 12808 1216 12860 1222
rect 12808 1158 12860 1164
rect 11520 944 11572 950
rect 11520 886 11572 892
rect 11716 800 11744 1158
rect 12912 800 12940 2246
rect 13004 1737 13032 2400
rect 13096 1834 13124 3023
rect 13188 2106 13216 5646
rect 13280 4282 13308 6258
rect 13372 5914 13400 9794
rect 13464 9790 13492 10450
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13452 9784 13504 9790
rect 13452 9726 13504 9732
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13464 7993 13492 8434
rect 13450 7984 13506 7993
rect 13450 7919 13506 7928
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7002 13492 7686
rect 13556 7206 13584 10066
rect 13740 9994 13768 10450
rect 14016 10062 14044 10450
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13636 9784 13688 9790
rect 13636 9726 13688 9732
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13648 6458 13676 9726
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 8566 13768 9454
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 7410 13768 8230
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 7206 13768 7346
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13450 6080 13506 6089
rect 13450 6015 13506 6024
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13464 5710 13492 6015
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13372 5409 13400 5578
rect 13358 5400 13414 5409
rect 13358 5335 13414 5344
rect 13372 5166 13400 5335
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13372 4078 13400 4422
rect 13360 4072 13412 4078
rect 13266 4040 13322 4049
rect 13360 4014 13412 4020
rect 13266 3975 13268 3984
rect 13320 3975 13322 3984
rect 13268 3946 13320 3952
rect 13358 3904 13414 3913
rect 13358 3839 13414 3848
rect 13266 3768 13322 3777
rect 13266 3703 13322 3712
rect 13280 3534 13308 3703
rect 13268 3528 13320 3534
rect 13372 3505 13400 3839
rect 13464 3516 13492 4966
rect 13556 3652 13584 6258
rect 13740 5914 13768 7142
rect 13832 6458 13860 9658
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8294 13952 8910
rect 14108 8838 14136 10882
rect 14278 10450 14334 11250
rect 14554 10450 14610 11250
rect 14830 10450 14886 11250
rect 15106 10450 15162 11250
rect 15382 10450 15438 11250
rect 15658 10450 15714 11250
rect 15934 10450 15990 11250
rect 16210 10450 16266 11250
rect 16486 10450 16542 11250
rect 16762 10450 16818 11250
rect 16856 10464 16908 10470
rect 14292 9858 14320 10450
rect 14372 10396 14424 10402
rect 14372 10338 14424 10344
rect 14280 9852 14332 9858
rect 14280 9794 14332 9800
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14384 8634 14412 10338
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 8634 14504 9862
rect 14568 9790 14596 10450
rect 14556 9784 14608 9790
rect 14556 9726 14608 9732
rect 14844 8922 14872 10450
rect 15120 10130 15148 10450
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15108 9852 15160 9858
rect 15108 9794 15160 9800
rect 14568 8894 14872 8922
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13916 8188 14292 8197
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14156 8188
rect 14212 8186 14236 8188
rect 13972 8134 13982 8186
rect 14226 8134 14236 8186
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14156 8134
rect 14212 8132 14236 8134
rect 13916 8123 14292 8132
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13924 7585 13952 7686
rect 13910 7576 13966 7585
rect 13910 7511 13966 7520
rect 14108 7478 14136 7822
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 13916 7100 14292 7109
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14156 7100
rect 14212 7098 14236 7100
rect 13972 7046 13982 7098
rect 14226 7046 14236 7098
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14156 7046
rect 14212 7044 14236 7046
rect 13916 7035 14292 7044
rect 14186 6896 14242 6905
rect 14186 6831 14188 6840
rect 14240 6831 14242 6840
rect 14188 6802 14240 6808
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14200 6322 14228 6802
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6390 14320 6734
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13648 4865 13676 5170
rect 13740 5098 13768 5578
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13634 4856 13690 4865
rect 13634 4791 13690 4800
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13648 3913 13676 4082
rect 13634 3904 13690 3913
rect 13634 3839 13690 3848
rect 13740 3738 13768 4422
rect 13832 3738 13860 6258
rect 13916 6012 14292 6021
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14156 6012
rect 14212 6010 14236 6012
rect 13972 5958 13982 6010
rect 14226 5958 14236 6010
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14156 5958
rect 14212 5956 14236 5958
rect 13916 5947 14292 5956
rect 14384 5914 14412 8434
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7954 14504 8230
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14568 7018 14596 8894
rect 14656 8732 15032 8741
rect 14712 8730 14736 8732
rect 14792 8730 14816 8732
rect 14872 8730 14896 8732
rect 14952 8730 14976 8732
rect 14712 8678 14722 8730
rect 14966 8678 14976 8730
rect 14712 8676 14736 8678
rect 14792 8676 14816 8678
rect 14872 8676 14896 8678
rect 14952 8676 14976 8678
rect 14656 8667 15032 8676
rect 15120 8634 15148 9794
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 14660 8362 14688 8434
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14832 7880 14884 7886
rect 14830 7848 14832 7857
rect 14884 7848 14886 7857
rect 14830 7783 14886 7792
rect 15028 7732 15056 8434
rect 15304 8362 15332 8774
rect 15396 8634 15424 10450
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15384 7948 15436 7954
rect 15384 7890 15436 7896
rect 15108 7880 15160 7886
rect 15160 7840 15240 7868
rect 15108 7822 15160 7828
rect 15028 7704 15148 7732
rect 14656 7644 15032 7653
rect 14712 7642 14736 7644
rect 14792 7642 14816 7644
rect 14872 7642 14896 7644
rect 14952 7642 14976 7644
rect 14712 7590 14722 7642
rect 14966 7590 14976 7642
rect 14712 7588 14736 7590
rect 14792 7588 14816 7590
rect 14872 7588 14896 7590
rect 14952 7588 14976 7590
rect 14656 7579 15032 7588
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14568 6990 14780 7018
rect 14462 6896 14518 6905
rect 14462 6831 14518 6840
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14200 5302 14228 5850
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13924 5030 13952 5170
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13916 4924 14292 4933
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14156 4924
rect 14212 4922 14236 4924
rect 13972 4870 13982 4922
rect 14226 4870 14236 4922
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14156 4870
rect 14212 4868 14236 4870
rect 13916 4859 14292 4868
rect 14384 4826 14412 5714
rect 14476 5409 14504 6831
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14568 5953 14596 6734
rect 14752 6662 14780 6990
rect 14936 6798 14964 7346
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14656 6556 15032 6565
rect 14712 6554 14736 6556
rect 14792 6554 14816 6556
rect 14872 6554 14896 6556
rect 14952 6554 14976 6556
rect 14712 6502 14722 6554
rect 14966 6502 14976 6554
rect 14712 6500 14736 6502
rect 14792 6500 14816 6502
rect 14872 6500 14896 6502
rect 14952 6500 14976 6502
rect 14656 6491 15032 6500
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14646 6080 14702 6089
rect 14646 6015 14702 6024
rect 14554 5944 14610 5953
rect 14554 5879 14610 5888
rect 14660 5556 14688 6015
rect 14936 5710 14964 6326
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14568 5528 14688 5556
rect 14462 5400 14518 5409
rect 14462 5335 14518 5344
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14096 4616 14148 4622
rect 14094 4584 14096 4593
rect 14372 4616 14424 4622
rect 14148 4584 14150 4593
rect 14094 4519 14150 4528
rect 14278 4584 14334 4593
rect 14372 4558 14424 4564
rect 14278 4519 14334 4528
rect 14002 4448 14058 4457
rect 14002 4383 14058 4392
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13924 4185 13952 4218
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13912 4072 13964 4078
rect 14016 4060 14044 4383
rect 14292 4321 14320 4519
rect 14278 4312 14334 4321
rect 14278 4247 14334 4256
rect 14384 4162 14412 4558
rect 14476 4264 14504 5102
rect 14568 4604 14596 5528
rect 14656 5468 15032 5477
rect 14712 5466 14736 5468
rect 14792 5466 14816 5468
rect 14872 5466 14896 5468
rect 14952 5466 14976 5468
rect 14712 5414 14722 5466
rect 14966 5414 14976 5466
rect 14712 5412 14736 5414
rect 14792 5412 14816 5414
rect 14872 5412 14896 5414
rect 14952 5412 14976 5414
rect 14656 5403 15032 5412
rect 14830 5264 14886 5273
rect 14830 5199 14886 5208
rect 15016 5228 15068 5234
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4706 14688 5102
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4826 14780 5034
rect 14844 5001 14872 5199
rect 15016 5170 15068 5176
rect 14830 4992 14886 5001
rect 14830 4927 14886 4936
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14844 4706 14872 4762
rect 14660 4678 14872 4706
rect 14924 4616 14976 4622
rect 14568 4576 14924 4604
rect 14568 4486 14596 4576
rect 14924 4558 14976 4564
rect 14556 4480 14608 4486
rect 15028 4468 15056 5170
rect 15120 4826 15148 7704
rect 15212 6089 15240 7840
rect 15396 7313 15424 7890
rect 15488 7886 15516 9930
rect 15568 9308 15620 9314
rect 15568 9250 15620 9256
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15382 7304 15438 7313
rect 15382 7239 15438 7248
rect 15198 6080 15254 6089
rect 15198 6015 15254 6024
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15212 5166 15240 5850
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15028 4440 15148 4468
rect 14556 4422 14608 4428
rect 14656 4380 15032 4389
rect 14712 4378 14736 4380
rect 14792 4378 14816 4380
rect 14872 4378 14896 4380
rect 14952 4378 14976 4380
rect 14712 4326 14722 4378
rect 14966 4326 14976 4378
rect 14712 4324 14736 4326
rect 14792 4324 14816 4326
rect 14872 4324 14896 4326
rect 14952 4324 14976 4326
rect 14656 4315 15032 4324
rect 14476 4236 14780 4264
rect 14384 4134 14688 4162
rect 13964 4032 14044 4060
rect 14464 4072 14516 4078
rect 13912 4014 13964 4020
rect 14660 4049 14688 4134
rect 14464 4014 14516 4020
rect 14646 4040 14702 4049
rect 13916 3836 14292 3845
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14156 3836
rect 14212 3834 14236 3836
rect 13972 3782 13982 3834
rect 14226 3782 14236 3834
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14156 3782
rect 14212 3780 14236 3782
rect 13916 3771 14292 3780
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13556 3624 13676 3652
rect 13648 3618 13676 3624
rect 13648 3590 13768 3618
rect 13636 3528 13688 3534
rect 13268 3470 13320 3476
rect 13358 3496 13414 3505
rect 13280 3097 13308 3470
rect 13464 3488 13636 3516
rect 13636 3470 13688 3476
rect 13358 3431 13414 3440
rect 13360 3392 13412 3398
rect 13544 3392 13596 3398
rect 13360 3334 13412 3340
rect 13464 3352 13544 3380
rect 13266 3088 13322 3097
rect 13372 3058 13400 3334
rect 13266 3023 13322 3032
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13084 1828 13136 1834
rect 13084 1770 13136 1776
rect 13464 1766 13492 3352
rect 13544 3334 13596 3340
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3126 13676 3334
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 1970 13584 2246
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 13452 1760 13504 1766
rect 12990 1728 13046 1737
rect 13452 1702 13504 1708
rect 12990 1663 13046 1672
rect 13740 882 13768 3590
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14004 3392 14056 3398
rect 13818 3360 13874 3369
rect 14004 3334 14056 3340
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 13818 3295 13874 3304
rect 13832 3126 13860 3295
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 14016 3058 14044 3334
rect 14200 3233 14228 3334
rect 14186 3224 14242 3233
rect 14292 3194 14320 3470
rect 14476 3466 14504 4014
rect 14752 4010 14780 4236
rect 14646 3975 14702 3984
rect 14740 4004 14792 4010
rect 14660 3534 14688 3975
rect 14740 3946 14792 3952
rect 15120 3670 15148 4440
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 14656 3292 15032 3301
rect 14712 3290 14736 3292
rect 14792 3290 14816 3292
rect 14872 3290 14896 3292
rect 14952 3290 14976 3292
rect 14712 3238 14722 3290
rect 14966 3238 14976 3290
rect 14712 3236 14736 3238
rect 14792 3236 14816 3238
rect 14872 3236 14896 3238
rect 14952 3236 14976 3238
rect 14656 3227 15032 3236
rect 14186 3159 14242 3168
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14464 3120 14516 3126
rect 14278 3088 14334 3097
rect 14004 3052 14056 3058
rect 14462 3088 14464 3097
rect 14516 3088 14518 3097
rect 14334 3046 14412 3074
rect 14278 3023 14334 3032
rect 14004 2994 14056 3000
rect 14384 2825 14412 3046
rect 14462 3023 14518 3032
rect 14370 2816 14426 2825
rect 13916 2748 14292 2757
rect 14370 2751 14426 2760
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14156 2748
rect 14212 2746 14236 2748
rect 13972 2694 13982 2746
rect 14226 2694 14236 2746
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14156 2694
rect 14212 2692 14236 2694
rect 13916 2683 14292 2692
rect 14370 2680 14426 2689
rect 14370 2615 14426 2624
rect 14096 2576 14148 2582
rect 14384 2530 14412 2615
rect 14096 2518 14148 2524
rect 13728 876 13780 882
rect 13728 818 13780 824
rect 14108 800 14136 2518
rect 14200 2502 14412 2530
rect 14200 2417 14228 2502
rect 14186 2408 14242 2417
rect 14186 2343 14242 2352
rect 14370 2408 14426 2417
rect 14370 2343 14372 2352
rect 14424 2343 14426 2352
rect 14372 2314 14424 2320
rect 14476 2310 14504 3023
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14568 2446 14596 2790
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14464 2304 14516 2310
rect 14370 2272 14426 2281
rect 14464 2246 14516 2252
rect 14370 2207 14426 2216
rect 14384 1329 14412 2207
rect 14656 2204 15032 2213
rect 14712 2202 14736 2204
rect 14792 2202 14816 2204
rect 14872 2202 14896 2204
rect 14952 2202 14976 2204
rect 14712 2150 14722 2202
rect 14966 2150 14976 2202
rect 14712 2148 14736 2150
rect 14792 2148 14816 2150
rect 14872 2148 14896 2150
rect 14952 2148 14976 2150
rect 14656 2139 15032 2148
rect 14464 1624 14516 1630
rect 14464 1566 14516 1572
rect 14370 1320 14426 1329
rect 14370 1255 14426 1264
rect 10784 604 10836 610
rect 10784 546 10836 552
rect 10782 504 10838 513
rect 10704 462 10782 490
rect 10782 439 10838 448
rect 11702 0 11758 800
rect 12898 0 12954 800
rect 14094 0 14150 800
rect 14476 542 14504 1566
rect 15120 1290 15148 3402
rect 15108 1284 15160 1290
rect 15108 1226 15160 1232
rect 14464 536 14516 542
rect 14464 478 14516 484
rect 15212 134 15240 4966
rect 15304 4622 15332 5782
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15396 5166 15424 5714
rect 15476 5568 15528 5574
rect 15580 5545 15608 9250
rect 15672 8090 15700 10450
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 8498 15792 9522
rect 15856 8498 15884 9590
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 7478 15884 7822
rect 15948 7546 15976 10450
rect 16224 10266 16252 10450
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16500 9926 16528 10450
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16776 9858 16804 10450
rect 17038 10450 17094 11250
rect 17314 10450 17370 11250
rect 17590 10450 17646 11250
rect 17866 10450 17922 11250
rect 18142 10450 18198 11250
rect 18418 10450 18474 11250
rect 18694 10450 18750 11250
rect 18970 10450 19026 11250
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 16856 10406 16908 10412
rect 16764 9852 16816 9858
rect 16764 9794 16816 9800
rect 16304 9784 16356 9790
rect 16304 9726 16356 9732
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16040 8634 16068 9658
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16118 8392 16174 8401
rect 16118 8327 16174 8336
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15660 7472 15712 7478
rect 15844 7472 15896 7478
rect 15712 7420 15792 7426
rect 15660 7414 15792 7420
rect 15844 7414 15896 7420
rect 15672 7398 15792 7414
rect 15764 7342 15792 7398
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15672 5574 15700 6598
rect 15764 5710 15792 6598
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15660 5568 15712 5574
rect 15476 5510 15528 5516
rect 15566 5536 15622 5545
rect 15488 5386 15516 5510
rect 15660 5510 15712 5516
rect 15750 5536 15806 5545
rect 15566 5471 15622 5480
rect 15750 5471 15806 5480
rect 15488 5358 15700 5386
rect 15566 5264 15622 5273
rect 15566 5199 15622 5208
rect 15384 5160 15436 5166
rect 15436 5120 15516 5148
rect 15384 5102 15436 5108
rect 15382 4856 15438 4865
rect 15382 4791 15438 4800
rect 15396 4758 15424 4791
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15488 4486 15516 5120
rect 15580 4758 15608 5199
rect 15672 5166 15700 5358
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15580 3942 15608 4558
rect 15672 4146 15700 4558
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15488 3058 15516 3538
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15672 3398 15700 3470
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15764 3058 15792 5471
rect 15856 5234 15884 7142
rect 16132 5794 16160 8327
rect 16224 6905 16252 9114
rect 16316 8634 16344 9726
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16408 7698 16436 9454
rect 16500 8498 16528 9590
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16776 8022 16804 8570
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16578 7848 16634 7857
rect 16578 7783 16634 7792
rect 16316 7670 16436 7698
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 15948 5766 16160 5794
rect 15948 5710 15976 5766
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15934 5400 15990 5409
rect 15934 5335 15990 5344
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15948 3194 15976 5335
rect 16040 5166 16068 5766
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4622 16252 4966
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16316 4434 16344 7670
rect 16592 7528 16620 7783
rect 16408 7500 16620 7528
rect 16408 7410 16436 7500
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16672 7404 16724 7410
rect 16724 7364 16804 7392
rect 16672 7346 16724 7352
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16408 4690 16436 5782
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16500 5302 16528 5510
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16224 4406 16344 4434
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 800 15332 2246
rect 15672 2038 15700 2382
rect 15660 2032 15712 2038
rect 15660 1974 15712 1980
rect 15476 1964 15528 1970
rect 15476 1906 15528 1912
rect 15488 1086 15516 1906
rect 16224 1562 16252 4406
rect 16302 4312 16358 4321
rect 16302 4247 16358 4256
rect 16316 2689 16344 4247
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16500 3194 16528 3946
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16592 2774 16620 7346
rect 16776 7313 16804 7364
rect 16762 7304 16818 7313
rect 16672 7268 16724 7274
rect 16762 7239 16818 7248
rect 16672 7210 16724 7216
rect 16684 4282 16712 7210
rect 16868 6882 16896 10406
rect 17052 8362 17080 10450
rect 17132 9920 17184 9926
rect 17130 9888 17132 9897
rect 17184 9888 17186 9897
rect 17130 9823 17186 9832
rect 17328 9722 17356 10450
rect 17604 9790 17632 10450
rect 17880 9874 17908 10450
rect 17788 9846 17908 9874
rect 17592 9784 17644 9790
rect 17592 9726 17644 9732
rect 17684 9784 17736 9790
rect 17684 9726 17736 9732
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8498 17540 8842
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17604 8498 17632 8570
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17420 7886 17448 8026
rect 17604 7886 17632 8230
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17038 7712 17094 7721
rect 17038 7647 17094 7656
rect 16946 7440 17002 7449
rect 16946 7375 16948 7384
rect 17000 7375 17002 7384
rect 16948 7346 17000 7352
rect 16776 6854 16896 6882
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16776 4078 16804 6854
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 5234 16896 6734
rect 17052 6390 17080 7647
rect 17328 7546 17356 7822
rect 17604 7750 17632 7822
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17420 6798 17448 7686
rect 17696 6866 17724 9726
rect 17788 8362 17816 9846
rect 18156 9738 18184 10450
rect 17880 9710 18184 9738
rect 17880 8634 17908 9710
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9081 18000 9318
rect 18144 9308 18196 9314
rect 18144 9250 18196 9256
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 18156 8498 18184 9250
rect 18432 8634 18460 10450
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17880 8022 17908 8434
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18050 8120 18106 8129
rect 18050 8055 18106 8064
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17788 6798 17816 7278
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17328 6662 17356 6734
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17682 6624 17738 6633
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 17130 6352 17186 6361
rect 17130 6287 17186 6296
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16960 5234 16988 6190
rect 17038 5944 17094 5953
rect 17038 5879 17094 5888
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16868 4826 16896 5170
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16854 4448 16910 4457
rect 16854 4383 16910 4392
rect 16868 4146 16896 4383
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16776 3058 16804 3334
rect 16854 3224 16910 3233
rect 16854 3159 16856 3168
rect 16908 3159 16910 3168
rect 16856 3130 16908 3136
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16592 2746 16712 2774
rect 16302 2680 16358 2689
rect 16302 2615 16358 2624
rect 16580 2304 16632 2310
rect 16580 2246 16632 2252
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 16592 1170 16620 2246
rect 16500 1142 16620 1170
rect 15476 1080 15528 1086
rect 15476 1022 15528 1028
rect 15568 1080 15620 1086
rect 15568 1022 15620 1028
rect 15200 128 15252 134
rect 15200 70 15252 76
rect 15290 0 15346 800
rect 15580 406 15608 1022
rect 16500 800 16528 1142
rect 15568 400 15620 406
rect 15568 342 15620 348
rect 16486 0 16542 800
rect 16684 542 16712 2746
rect 17052 1766 17080 5879
rect 17144 5273 17172 6287
rect 17236 5370 17264 6598
rect 17682 6559 17738 6568
rect 17696 6390 17724 6559
rect 17788 6390 17816 6734
rect 17316 6384 17368 6390
rect 17684 6384 17736 6390
rect 17316 6326 17368 6332
rect 17590 6352 17646 6361
rect 17328 6118 17356 6326
rect 17684 6326 17736 6332
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17590 6287 17592 6296
rect 17644 6287 17646 6296
rect 17592 6258 17644 6264
rect 17498 6216 17554 6225
rect 17498 6151 17554 6160
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17314 5944 17370 5953
rect 17314 5879 17370 5888
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17130 5264 17186 5273
rect 17328 5250 17356 5879
rect 17420 5846 17448 6054
rect 17408 5840 17460 5846
rect 17408 5782 17460 5788
rect 17130 5199 17186 5208
rect 17236 5222 17356 5250
rect 17236 3534 17264 5222
rect 17512 4978 17540 6151
rect 17604 5710 17632 6258
rect 17682 5944 17738 5953
rect 17682 5879 17738 5888
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17420 4950 17540 4978
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17328 3913 17356 4762
rect 17314 3904 17370 3913
rect 17314 3839 17370 3848
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17222 3224 17278 3233
rect 17222 3159 17224 3168
rect 17276 3159 17278 3168
rect 17224 3130 17276 3136
rect 17040 1760 17092 1766
rect 17040 1702 17092 1708
rect 17420 1630 17448 4950
rect 17498 4856 17554 4865
rect 17498 4791 17500 4800
rect 17552 4791 17554 4800
rect 17500 4762 17552 4768
rect 17604 4758 17632 5306
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17696 4622 17724 5879
rect 17776 5704 17828 5710
rect 17880 5692 17908 7783
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17972 6798 18000 7346
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18064 6474 18092 8055
rect 18340 7886 18368 8230
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18340 7721 18368 7822
rect 18432 7818 18460 8026
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18326 7712 18382 7721
rect 18326 7647 18382 7656
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18328 6724 18380 6730
rect 18328 6666 18380 6672
rect 17828 5664 17908 5692
rect 17972 6446 18092 6474
rect 17776 5646 17828 5652
rect 17972 5556 18000 6446
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17880 5528 18000 5556
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17684 4616 17736 4622
rect 17788 4593 17816 4966
rect 17684 4558 17736 4564
rect 17774 4584 17830 4593
rect 17696 4078 17724 4558
rect 17774 4519 17830 4528
rect 17774 4312 17830 4321
rect 17880 4298 17908 5528
rect 18064 5386 18092 6326
rect 18340 6254 18368 6666
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18432 5624 18460 7482
rect 18524 6934 18552 9046
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18616 7954 18644 8502
rect 18708 8090 18736 10450
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18708 7546 18736 7686
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18800 6390 18828 8298
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18892 7313 18920 8230
rect 18984 8090 19012 10450
rect 19168 10305 19196 10542
rect 19246 10450 19302 11250
rect 19522 10450 19578 11250
rect 19798 10450 19854 11250
rect 20074 10450 20130 11250
rect 20350 10450 20406 11250
rect 20626 10450 20682 11250
rect 20902 10450 20958 11250
rect 21178 10450 21234 11250
rect 21454 10554 21510 11250
rect 21730 10554 21786 11250
rect 21454 10526 21680 10554
rect 21454 10450 21510 10526
rect 19154 10296 19210 10305
rect 19154 10231 19210 10240
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18878 7304 18934 7313
rect 18878 7239 18934 7248
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6458 18920 6598
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18984 6236 19012 7822
rect 19076 7041 19104 7822
rect 19062 7032 19118 7041
rect 19062 6967 19118 6976
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 19076 6338 19104 6870
rect 19168 6798 19196 9658
rect 19260 8362 19288 10450
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19260 6905 19288 7346
rect 19352 7002 19380 9998
rect 19444 9042 19472 10066
rect 19536 9790 19564 10450
rect 19616 10396 19668 10402
rect 19616 10338 19668 10344
rect 19628 9790 19656 10338
rect 19524 9784 19576 9790
rect 19524 9726 19576 9732
rect 19616 9784 19668 9790
rect 19616 9726 19668 9732
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19444 8498 19472 8570
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19536 8090 19564 8774
rect 19628 8498 19656 9046
rect 19812 8809 19840 10450
rect 19798 8800 19854 8809
rect 19798 8735 19854 8744
rect 20088 8498 20116 10450
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19444 7002 19472 7890
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19536 6905 19564 7890
rect 19246 6896 19302 6905
rect 19246 6831 19302 6840
rect 19522 6896 19578 6905
rect 19522 6831 19578 6840
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19260 6458 19288 6831
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19076 6310 19288 6338
rect 18892 6225 19012 6236
rect 18694 6216 18750 6225
rect 18878 6216 19012 6225
rect 18694 6151 18750 6160
rect 18788 6180 18840 6186
rect 18708 6118 18736 6151
rect 18934 6208 19012 6216
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 18878 6151 18934 6160
rect 18788 6122 18840 6128
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18696 6112 18748 6118
rect 18800 6089 18828 6122
rect 18696 6054 18748 6060
rect 18786 6080 18842 6089
rect 18616 5914 18644 6054
rect 18970 6080 19026 6089
rect 18786 6015 18842 6024
rect 18892 6038 18970 6066
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18892 5642 18920 6038
rect 18970 6015 19026 6024
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18880 5636 18932 5642
rect 18432 5596 18736 5624
rect 18708 5545 18736 5596
rect 18880 5578 18932 5584
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18788 5568 18840 5574
rect 18142 5536 18198 5545
rect 18142 5471 18198 5480
rect 18510 5536 18566 5545
rect 18694 5536 18750 5545
rect 18566 5494 18644 5522
rect 18510 5471 18566 5480
rect 17972 5358 18092 5386
rect 17972 4706 18000 5358
rect 18156 4842 18184 5471
rect 18616 5234 18644 5494
rect 18788 5510 18840 5516
rect 18694 5471 18750 5480
rect 18512 5228 18564 5234
rect 18432 5188 18512 5216
rect 18064 4826 18184 4842
rect 18052 4820 18184 4826
rect 18104 4814 18184 4820
rect 18326 4856 18382 4865
rect 18326 4791 18328 4800
rect 18052 4762 18104 4768
rect 18380 4791 18382 4800
rect 18328 4762 18380 4768
rect 18432 4758 18460 5188
rect 18512 5170 18564 5176
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18800 5030 18828 5510
rect 18984 5234 19012 5578
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19076 5166 19104 5850
rect 19168 5642 19196 6190
rect 19260 5914 19288 6310
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19352 5710 19380 6598
rect 19536 6497 19564 6831
rect 19522 6488 19578 6497
rect 19522 6423 19578 6432
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19156 5636 19208 5642
rect 19536 5624 19564 6326
rect 19628 6322 19656 8298
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19720 8129 19748 8230
rect 19916 8188 20292 8197
rect 19972 8186 19996 8188
rect 20052 8186 20076 8188
rect 20132 8186 20156 8188
rect 20212 8186 20236 8188
rect 19972 8134 19982 8186
rect 20226 8134 20236 8186
rect 19972 8132 19996 8134
rect 20052 8132 20076 8134
rect 20132 8132 20156 8134
rect 20212 8132 20236 8134
rect 19706 8120 19762 8129
rect 19916 8123 20292 8132
rect 19706 8055 19762 8064
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7546 19748 7822
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19812 7478 19840 7686
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19708 7200 19760 7206
rect 19996 7188 20024 7686
rect 19708 7142 19760 7148
rect 19812 7160 20024 7188
rect 19720 6322 19748 7142
rect 19812 6322 19840 7160
rect 19916 7100 20292 7109
rect 19972 7098 19996 7100
rect 20052 7098 20076 7100
rect 20132 7098 20156 7100
rect 20212 7098 20236 7100
rect 19972 7046 19982 7098
rect 20226 7046 20236 7098
rect 19972 7044 19996 7046
rect 20052 7044 20076 7046
rect 20132 7044 20156 7046
rect 20212 7044 20236 7046
rect 19916 7035 20292 7044
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 19904 6662 19932 6734
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19996 6390 20024 6734
rect 20180 6662 20208 6734
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20364 6458 20392 10450
rect 20640 9722 20668 10450
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20916 9194 20944 10450
rect 21192 9722 21220 10450
rect 21546 10296 21602 10305
rect 21546 10231 21602 10240
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21376 9858 21404 9998
rect 21560 9897 21588 10231
rect 21546 9888 21602 9897
rect 21272 9852 21324 9858
rect 21272 9794 21324 9800
rect 21364 9852 21416 9858
rect 21546 9823 21602 9832
rect 21364 9794 21416 9800
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21284 9382 21312 9794
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 20916 9166 21128 9194
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20442 8664 20498 8673
rect 20442 8599 20498 8608
rect 20456 8265 20484 8599
rect 20442 8256 20498 8265
rect 20442 8191 20498 8200
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 7410 20484 7686
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20548 7206 20576 8910
rect 20656 8732 21032 8741
rect 20712 8730 20736 8732
rect 20792 8730 20816 8732
rect 20872 8730 20896 8732
rect 20952 8730 20976 8732
rect 20712 8678 20722 8730
rect 20966 8678 20976 8730
rect 20712 8676 20736 8678
rect 20792 8676 20816 8678
rect 20872 8676 20896 8678
rect 20952 8676 20976 8678
rect 20656 8667 21032 8676
rect 20720 8424 20772 8430
rect 20718 8392 20720 8401
rect 20772 8392 20774 8401
rect 20718 8327 20774 8336
rect 21100 7954 21128 9166
rect 21652 8498 21680 10526
rect 21730 10526 21864 10554
rect 21730 10450 21786 10526
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 21180 7880 21232 7886
rect 21640 7880 21692 7886
rect 21232 7840 21312 7868
rect 21180 7822 21232 7828
rect 20656 7644 21032 7653
rect 20712 7642 20736 7644
rect 20792 7642 20816 7644
rect 20872 7642 20896 7644
rect 20952 7642 20976 7644
rect 20712 7590 20722 7642
rect 20966 7590 20976 7642
rect 20712 7588 20736 7590
rect 20792 7588 20816 7590
rect 20872 7588 20896 7590
rect 20952 7588 20976 7590
rect 20656 7579 21032 7588
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20626 7168 20682 7177
rect 20456 6866 20484 7142
rect 20626 7103 20682 7112
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20640 6746 20668 7103
rect 21008 6866 21036 7278
rect 20996 6860 21048 6866
rect 21048 6820 21128 6848
rect 20996 6802 21048 6808
rect 20456 6718 20668 6746
rect 20456 6662 20484 6718
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 19984 6384 20036 6390
rect 20456 6338 20484 6394
rect 19984 6326 20036 6332
rect 19616 6316 19668 6322
rect 19616 6258 19668 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 20364 6310 20484 6338
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19706 6080 19762 6089
rect 19628 5953 19656 6054
rect 19812 6066 19840 6258
rect 20364 6254 20392 6310
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 19996 6118 20024 6190
rect 19762 6038 19840 6066
rect 19984 6112 20036 6118
rect 20548 6066 20576 6598
rect 20656 6556 21032 6565
rect 20712 6554 20736 6556
rect 20792 6554 20816 6556
rect 20872 6554 20896 6556
rect 20952 6554 20976 6556
rect 20712 6502 20722 6554
rect 20966 6502 20976 6554
rect 20712 6500 20736 6502
rect 20792 6500 20816 6502
rect 20872 6500 20896 6502
rect 20952 6500 20976 6502
rect 20656 6491 21032 6500
rect 21100 6440 21128 6820
rect 20732 6412 21128 6440
rect 20732 6322 20760 6412
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 19984 6054 20036 6060
rect 19706 6015 19762 6024
rect 19614 5944 19670 5953
rect 19614 5879 19616 5888
rect 19668 5879 19670 5888
rect 19616 5850 19668 5856
rect 19812 5710 19840 6038
rect 20364 6038 20576 6066
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 19916 6012 20292 6021
rect 19972 6010 19996 6012
rect 20052 6010 20076 6012
rect 20132 6010 20156 6012
rect 20212 6010 20236 6012
rect 19972 5958 19982 6010
rect 20226 5958 20236 6010
rect 19972 5956 19996 5958
rect 20052 5956 20076 5958
rect 20132 5956 20156 5958
rect 20212 5956 20236 5958
rect 19916 5947 20292 5956
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 19996 5778 20024 5850
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19616 5704 19668 5710
rect 19156 5578 19208 5584
rect 19444 5596 19564 5624
rect 19614 5672 19616 5681
rect 19800 5704 19852 5710
rect 19668 5672 19670 5681
rect 19800 5646 19852 5652
rect 19614 5607 19670 5616
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19444 5522 19472 5596
rect 19708 5568 19760 5574
rect 19352 5409 19380 5510
rect 19444 5494 19564 5522
rect 19708 5510 19760 5516
rect 19338 5400 19394 5409
rect 19248 5364 19300 5370
rect 19338 5335 19394 5344
rect 19248 5306 19300 5312
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19156 5160 19208 5166
rect 19156 5102 19208 5108
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18510 4856 18566 4865
rect 18510 4791 18566 4800
rect 18420 4752 18472 4758
rect 17972 4678 18092 4706
rect 18420 4694 18472 4700
rect 17830 4270 17908 4298
rect 17774 4247 17830 4256
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17684 4072 17736 4078
rect 17512 4032 17684 4060
rect 17512 3670 17540 4032
rect 17684 4014 17736 4020
rect 17880 3738 17908 4082
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17512 2836 17540 3470
rect 17592 2984 17644 2990
rect 17696 2938 17724 3470
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17644 2932 17724 2938
rect 17592 2926 17724 2932
rect 17604 2910 17724 2926
rect 17512 2808 17632 2836
rect 17604 2446 17632 2808
rect 17696 2774 17724 2910
rect 17880 2825 17908 3334
rect 17972 2990 18000 3674
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17866 2816 17922 2825
rect 17696 2746 17816 2774
rect 17866 2751 17922 2760
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 17512 2106 17540 2314
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 17604 1698 17632 2382
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17592 1692 17644 1698
rect 17592 1634 17644 1640
rect 17408 1624 17460 1630
rect 17408 1566 17460 1572
rect 17696 800 17724 2246
rect 17788 1698 17816 2746
rect 17880 2446 17908 2751
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18064 2310 18092 4678
rect 18234 4584 18290 4593
rect 18234 4519 18290 4528
rect 18142 3768 18198 3777
rect 18142 3703 18198 3712
rect 18156 3534 18184 3703
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18156 3058 18184 3334
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18248 1873 18276 4519
rect 18524 3942 18552 4791
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18616 4457 18644 4626
rect 18602 4448 18658 4457
rect 18602 4383 18658 4392
rect 18708 4282 18736 4966
rect 18800 4690 18828 4966
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18800 4554 18828 4626
rect 19076 4622 19104 5102
rect 19168 4826 19196 5102
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19260 4758 19288 5306
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19444 4865 19472 5238
rect 19536 5216 19564 5494
rect 19720 5234 19748 5510
rect 19798 5400 19854 5409
rect 19798 5335 19854 5344
rect 19812 5302 19840 5335
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19984 5296 20036 5302
rect 20272 5284 20300 5850
rect 20364 5846 20392 6038
rect 20732 5914 20760 6054
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20444 5840 20496 5846
rect 20496 5800 20576 5828
rect 20444 5782 20496 5788
rect 20548 5658 20576 5800
rect 20036 5256 20300 5284
rect 20456 5630 20576 5658
rect 20720 5704 20772 5710
rect 20824 5692 20852 6412
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 20916 5953 20944 6190
rect 20902 5944 20958 5953
rect 20902 5879 20904 5888
rect 20956 5879 20958 5888
rect 20904 5850 20956 5856
rect 20916 5710 20944 5850
rect 20772 5664 20852 5692
rect 20904 5704 20956 5710
rect 20720 5646 20772 5652
rect 20904 5646 20956 5652
rect 20996 5704 21048 5710
rect 21048 5664 21128 5692
rect 20996 5646 21048 5652
rect 19984 5238 20036 5244
rect 19708 5228 19760 5234
rect 19536 5188 19656 5216
rect 19430 4856 19486 4865
rect 19430 4791 19486 4800
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 19064 4480 19116 4486
rect 18970 4448 19026 4457
rect 19064 4422 19116 4428
rect 18970 4383 19026 4392
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18878 4176 18934 4185
rect 18984 4146 19012 4383
rect 19076 4282 19104 4422
rect 19338 4312 19394 4321
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19248 4276 19300 4282
rect 19338 4247 19394 4256
rect 19248 4218 19300 4224
rect 18878 4111 18934 4120
rect 18972 4140 19024 4146
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18340 3058 18368 3674
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18420 2984 18472 2990
rect 18418 2952 18420 2961
rect 18472 2952 18474 2961
rect 18418 2887 18474 2896
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18708 2650 18736 2858
rect 18786 2680 18842 2689
rect 18696 2644 18748 2650
rect 18786 2615 18788 2624
rect 18696 2586 18748 2592
rect 18840 2615 18842 2624
rect 18788 2586 18840 2592
rect 18234 1864 18290 1873
rect 18234 1799 18290 1808
rect 17776 1692 17828 1698
rect 17776 1634 17828 1640
rect 18892 800 18920 4111
rect 18972 4082 19024 4088
rect 19260 3670 19288 4218
rect 19352 3670 19380 4247
rect 19430 3904 19486 3913
rect 19430 3839 19486 3848
rect 19248 3664 19300 3670
rect 19062 3632 19118 3641
rect 19248 3606 19300 3612
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19444 3602 19472 3839
rect 19062 3567 19118 3576
rect 19432 3596 19484 3602
rect 16672 536 16724 542
rect 16672 478 16724 484
rect 17682 0 17738 800
rect 18878 0 18934 800
rect 19076 474 19104 3567
rect 19432 3538 19484 3544
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19154 3224 19210 3233
rect 19154 3159 19210 3168
rect 19168 3058 19196 3159
rect 19352 3074 19380 3470
rect 19536 3194 19564 3470
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19156 3052 19208 3058
rect 19352 3046 19564 3074
rect 19156 2994 19208 3000
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 2106 19472 2926
rect 19536 2446 19564 3046
rect 19628 2922 19656 5188
rect 19708 5170 19760 5176
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 20076 5160 20128 5166
rect 20128 5120 20392 5148
rect 20076 5102 20128 5108
rect 19708 5092 19760 5098
rect 19708 5034 19760 5040
rect 19720 5001 19748 5034
rect 19706 4992 19762 5001
rect 19706 4927 19762 4936
rect 19812 4604 19840 5102
rect 19916 4924 20292 4933
rect 19972 4922 19996 4924
rect 20052 4922 20076 4924
rect 20132 4922 20156 4924
rect 20212 4922 20236 4924
rect 19972 4870 19982 4922
rect 20226 4870 20236 4922
rect 19972 4868 19996 4870
rect 20052 4868 20076 4870
rect 20132 4868 20156 4870
rect 20212 4868 20236 4870
rect 19916 4859 20292 4868
rect 20260 4684 20312 4690
rect 20364 4672 20392 5120
rect 20312 4644 20392 4672
rect 20456 4672 20484 5630
rect 20656 5468 21032 5477
rect 20712 5466 20736 5468
rect 20792 5466 20816 5468
rect 20872 5466 20896 5468
rect 20952 5466 20976 5468
rect 20712 5414 20722 5466
rect 20966 5414 20976 5466
rect 20712 5412 20736 5414
rect 20792 5412 20816 5414
rect 20872 5412 20896 5414
rect 20952 5412 20976 5414
rect 20656 5403 21032 5412
rect 20720 5160 20772 5166
rect 20626 5128 20682 5137
rect 20548 5098 20626 5114
rect 20536 5092 20626 5098
rect 20588 5086 20626 5092
rect 20904 5160 20956 5166
rect 20772 5120 20852 5148
rect 20720 5102 20772 5108
rect 20626 5063 20682 5072
rect 20536 5034 20588 5040
rect 20626 4992 20682 5001
rect 20626 4927 20682 4936
rect 20536 4684 20588 4690
rect 20456 4644 20536 4672
rect 20260 4626 20312 4632
rect 19892 4616 19944 4622
rect 19812 4576 19892 4604
rect 19892 4558 19944 4564
rect 19904 4185 19932 4558
rect 19890 4176 19946 4185
rect 19890 4111 19946 4120
rect 20456 4010 20484 4644
rect 20640 4672 20668 4927
rect 20824 4690 20852 5120
rect 20904 5102 20956 5108
rect 20916 4826 20944 5102
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20588 4644 20668 4672
rect 20812 4684 20864 4690
rect 20536 4626 20588 4632
rect 20812 4626 20864 4632
rect 20916 4622 20944 4762
rect 21100 4622 21128 5664
rect 21192 5166 21220 6190
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 20656 4380 21032 4389
rect 20712 4378 20736 4380
rect 20792 4378 20816 4380
rect 20872 4378 20896 4380
rect 20952 4378 20976 4380
rect 20712 4326 20722 4378
rect 20966 4326 20976 4378
rect 20712 4324 20736 4326
rect 20792 4324 20816 4326
rect 20872 4324 20896 4326
rect 20952 4324 20976 4326
rect 20656 4315 21032 4324
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20996 4072 21048 4078
rect 21100 4060 21128 4558
rect 21178 4312 21234 4321
rect 21178 4247 21234 4256
rect 21048 4032 21128 4060
rect 20996 4014 21048 4020
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20548 3913 20576 4014
rect 20534 3904 20590 3913
rect 19916 3836 20292 3845
rect 20534 3839 20590 3848
rect 19972 3834 19996 3836
rect 20052 3834 20076 3836
rect 20132 3834 20156 3836
rect 20212 3834 20236 3836
rect 19972 3782 19982 3834
rect 20226 3782 20236 3834
rect 19972 3780 19996 3782
rect 20052 3780 20076 3782
rect 20132 3780 20156 3782
rect 20212 3780 20236 3782
rect 19916 3771 20292 3780
rect 20732 3584 20760 4014
rect 20916 3738 20944 4014
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 21008 3670 21036 4014
rect 20996 3664 21048 3670
rect 20996 3606 21048 3612
rect 20732 3556 20944 3584
rect 19892 3528 19944 3534
rect 19890 3496 19892 3505
rect 20536 3528 20588 3534
rect 19944 3496 19946 3505
rect 19800 3460 19852 3466
rect 20536 3470 20588 3476
rect 19890 3431 19946 3440
rect 19800 3402 19852 3408
rect 19812 3194 19840 3402
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 20456 3058 20484 3334
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 20352 2984 20404 2990
rect 20404 2932 20484 2938
rect 20352 2926 20484 2932
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19168 1222 19196 2042
rect 19628 1494 19656 2858
rect 19812 2854 19840 2926
rect 20364 2910 20484 2926
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 20352 2848 20404 2854
rect 20456 2825 20484 2910
rect 20352 2790 20404 2796
rect 20442 2816 20498 2825
rect 19916 2748 20292 2757
rect 19972 2746 19996 2748
rect 20052 2746 20076 2748
rect 20132 2746 20156 2748
rect 20212 2746 20236 2748
rect 19972 2694 19982 2746
rect 20226 2694 20236 2746
rect 19972 2692 19996 2694
rect 20052 2692 20076 2694
rect 20132 2692 20156 2694
rect 20212 2692 20236 2694
rect 19916 2683 20292 2692
rect 20364 2650 20392 2790
rect 20442 2751 20498 2760
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20364 2378 20392 2450
rect 20548 2446 20576 3470
rect 20916 3466 20944 3556
rect 21192 3466 21220 4247
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 20656 3292 21032 3301
rect 20712 3290 20736 3292
rect 20792 3290 20816 3292
rect 20872 3290 20896 3292
rect 20952 3290 20976 3292
rect 20712 3238 20722 3290
rect 20966 3238 20976 3290
rect 20712 3236 20736 3238
rect 20792 3236 20816 3238
rect 20872 3236 20896 3238
rect 20952 3236 20976 3238
rect 20656 3227 21032 3236
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 20656 2204 21032 2213
rect 20712 2202 20736 2204
rect 20792 2202 20816 2204
rect 20872 2202 20896 2204
rect 20952 2202 20976 2204
rect 20712 2150 20722 2202
rect 20966 2150 20976 2202
rect 20712 2148 20736 2150
rect 20792 2148 20816 2150
rect 20872 2148 20896 2150
rect 20952 2148 20976 2150
rect 20656 2139 21032 2148
rect 21100 1970 21128 2790
rect 21284 2689 21312 7840
rect 21640 7822 21692 7828
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21560 7041 21588 7278
rect 21546 7032 21602 7041
rect 21546 6967 21602 6976
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21376 3992 21404 6734
rect 21546 6624 21602 6633
rect 21546 6559 21602 6568
rect 21454 6352 21510 6361
rect 21454 6287 21510 6296
rect 21468 6089 21496 6287
rect 21454 6080 21510 6089
rect 21454 6015 21510 6024
rect 21560 5914 21588 6559
rect 21652 6254 21680 7822
rect 21744 6662 21772 8366
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21836 6304 21864 10526
rect 21916 10464 21968 10470
rect 22006 10450 22062 11250
rect 22282 10450 22338 11250
rect 22558 10450 22614 11250
rect 22834 10450 22890 11250
rect 23110 10450 23166 11250
rect 23386 10554 23442 11250
rect 23386 10526 23612 10554
rect 23386 10450 23442 10526
rect 21916 10406 21968 10412
rect 21928 8906 21956 10406
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21914 8664 21970 8673
rect 21914 8599 21970 8608
rect 21928 8090 21956 8599
rect 22020 8498 22048 10450
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 22008 8288 22060 8294
rect 22006 8256 22008 8265
rect 22060 8256 22062 8265
rect 22006 8191 22062 8200
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21914 7984 21970 7993
rect 21914 7919 21970 7928
rect 21928 7886 21956 7919
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21928 7041 21956 7822
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21914 7032 21970 7041
rect 21914 6967 21970 6976
rect 21914 6896 21970 6905
rect 22020 6882 22048 7278
rect 21970 6854 22048 6882
rect 21914 6831 21970 6840
rect 21928 6798 21956 6831
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22112 6322 22140 9658
rect 22204 8673 22232 10134
rect 22190 8664 22246 8673
rect 22190 8599 22246 8608
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 21916 6316 21968 6322
rect 21836 6276 21916 6304
rect 21916 6258 21968 6264
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 21640 6248 21692 6254
rect 21692 6208 21772 6236
rect 21640 6190 21692 6196
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21652 5914 21680 6054
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21744 5794 21772 6208
rect 22204 6186 22232 7958
rect 22296 7392 22324 10450
rect 22572 8090 22600 10450
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22664 7970 22692 8366
rect 22572 7942 22692 7970
rect 22376 7404 22428 7410
rect 22296 7364 22376 7392
rect 22376 7346 22428 7352
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22388 6497 22416 7210
rect 22466 6896 22522 6905
rect 22466 6831 22468 6840
rect 22520 6831 22522 6840
rect 22468 6802 22520 6808
rect 22374 6488 22430 6497
rect 22374 6423 22430 6432
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 21652 5766 21772 5794
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21468 4593 21496 5034
rect 21560 5030 21588 5578
rect 21652 5574 21680 5766
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21822 5264 21878 5273
rect 21822 5199 21878 5208
rect 21836 5166 21864 5199
rect 21824 5160 21876 5166
rect 21824 5102 21876 5108
rect 21928 5030 21956 6054
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 22098 5536 22154 5545
rect 22020 5234 22048 5510
rect 22098 5471 22154 5480
rect 22112 5370 22140 5471
rect 22204 5370 22232 5646
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 21548 5024 21600 5030
rect 21916 5024 21968 5030
rect 21548 4966 21600 4972
rect 21730 4992 21786 5001
rect 21916 4966 21968 4972
rect 22006 4992 22062 5001
rect 21730 4927 21786 4936
rect 22006 4927 22062 4936
rect 21744 4758 21772 4927
rect 22020 4826 22048 4927
rect 22112 4826 22140 5170
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22192 5092 22244 5098
rect 22192 5034 22244 5040
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 21548 4752 21600 4758
rect 21548 4694 21600 4700
rect 21732 4752 21784 4758
rect 21732 4694 21784 4700
rect 21454 4584 21510 4593
rect 21454 4519 21510 4528
rect 21560 4321 21588 4694
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21546 4312 21602 4321
rect 21546 4247 21602 4256
rect 21652 4078 21680 4626
rect 22204 4622 22232 5034
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21824 4548 21876 4554
rect 21824 4490 21876 4496
rect 21836 4282 21864 4490
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 22112 4146 22140 4422
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22204 4078 22232 4558
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 21456 4004 21508 4010
rect 21376 3964 21456 3992
rect 21376 3602 21404 3964
rect 21456 3946 21508 3952
rect 22098 3632 22154 3641
rect 21364 3596 21416 3602
rect 22098 3567 22154 3576
rect 21364 3538 21416 3544
rect 21824 3528 21876 3534
rect 21454 3496 21510 3505
rect 21824 3470 21876 3476
rect 21454 3431 21510 3440
rect 21468 3398 21496 3431
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21270 2680 21326 2689
rect 21376 2650 21404 2926
rect 21468 2854 21496 3334
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21270 2615 21272 2624
rect 21324 2615 21326 2624
rect 21364 2644 21416 2650
rect 21272 2586 21324 2592
rect 21364 2586 21416 2592
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 19984 1896 20036 1902
rect 20036 1844 20116 1850
rect 19984 1838 20116 1844
rect 19996 1822 20116 1838
rect 20088 1816 20116 1822
rect 20168 1828 20220 1834
rect 20088 1788 20168 1816
rect 20168 1770 20220 1776
rect 19616 1488 19668 1494
rect 19616 1430 19668 1436
rect 20076 1284 20128 1290
rect 20076 1226 20128 1232
rect 19156 1216 19208 1222
rect 19156 1158 19208 1164
rect 20088 800 20116 1226
rect 21192 836 21312 864
rect 19064 468 19116 474
rect 19064 410 19116 416
rect 20074 0 20130 800
rect 21192 134 21220 836
rect 21284 800 21312 836
rect 21180 128 21232 134
rect 21180 70 21232 76
rect 21270 0 21326 800
rect 21836 610 21864 3470
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 21928 1290 21956 2994
rect 22020 1630 22048 3334
rect 22008 1624 22060 1630
rect 22008 1566 22060 1572
rect 22112 1494 22140 3567
rect 22190 2952 22246 2961
rect 22296 2922 22324 4762
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22388 4282 22416 4422
rect 22480 4282 22508 5102
rect 22572 4321 22600 7942
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22558 4312 22614 4321
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22468 4276 22520 4282
rect 22558 4247 22614 4256
rect 22468 4218 22520 4224
rect 22664 3602 22692 7414
rect 22756 7342 22784 8774
rect 22848 8498 22876 10450
rect 22928 9852 22980 9858
rect 22928 9794 22980 9800
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22756 7177 22784 7278
rect 22742 7168 22798 7177
rect 22742 7103 22798 7112
rect 22742 7032 22798 7041
rect 22742 6967 22798 6976
rect 22756 6798 22784 6967
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 22756 5166 22784 6190
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22848 4078 22876 8230
rect 22940 7886 22968 9794
rect 23124 8566 23152 10450
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23216 8362 23244 9998
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 23112 8356 23164 8362
rect 23112 8298 23164 8304
rect 23204 8356 23256 8362
rect 23204 8298 23256 8304
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22940 6390 22968 7822
rect 23124 6866 23152 8298
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23216 7478 23244 7822
rect 23204 7472 23256 7478
rect 23308 7449 23336 9386
rect 23400 8498 23428 9658
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23204 7414 23256 7420
rect 23294 7440 23350 7449
rect 23294 7375 23350 7384
rect 23386 6896 23442 6905
rect 23112 6860 23164 6866
rect 23386 6831 23442 6840
rect 23112 6802 23164 6808
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 23032 6118 23060 6666
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22940 5234 22968 6054
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22940 4486 22968 5170
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 23020 4140 23072 4146
rect 23124 4128 23152 6666
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23216 5352 23244 6598
rect 23296 5364 23348 5370
rect 23216 5324 23296 5352
rect 23216 4690 23244 5324
rect 23296 5306 23348 5312
rect 23400 5284 23428 6831
rect 23492 6746 23520 7822
rect 23584 7410 23612 10526
rect 23662 10450 23718 11250
rect 23938 10450 23994 11250
rect 24214 10450 24270 11250
rect 24490 10450 24546 11250
rect 24766 10450 24822 11250
rect 25042 10554 25098 11250
rect 24872 10526 25098 10554
rect 23676 9722 23704 10450
rect 23952 9722 23980 10450
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23676 8498 23704 8842
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23754 8256 23810 8265
rect 23754 8191 23810 8200
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23492 6718 23612 6746
rect 23480 6656 23532 6662
rect 23480 6598 23532 6604
rect 23492 6322 23520 6598
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23400 5256 23520 5284
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 23308 5030 23336 5102
rect 23296 5024 23348 5030
rect 23296 4966 23348 4972
rect 23308 4690 23336 4966
rect 23492 4808 23520 5256
rect 23584 5001 23612 6718
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23676 6458 23704 6666
rect 23768 6458 23796 8191
rect 23860 7274 23888 9318
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 24136 8634 24164 8842
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 24044 7410 24072 8502
rect 24228 7818 24256 10450
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24136 7410 24164 7482
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 23940 7200 23992 7206
rect 23940 7142 23992 7148
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 23952 6662 23980 7142
rect 24228 6866 24256 7142
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 23664 6180 23716 6186
rect 23664 6122 23716 6128
rect 23676 5098 23704 6122
rect 23768 5710 23796 6258
rect 23952 5914 23980 6258
rect 24136 5914 24164 6258
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23860 5545 23888 5578
rect 23846 5536 23902 5545
rect 23846 5471 23902 5480
rect 23846 5400 23902 5409
rect 23846 5335 23902 5344
rect 23940 5364 23992 5370
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23570 4992 23626 5001
rect 23570 4927 23626 4936
rect 23492 4780 23612 4808
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23072 4100 23152 4128
rect 23020 4082 23072 4088
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 23032 3942 23060 4082
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23020 3936 23072 3942
rect 23216 3913 23244 4014
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23020 3878 23072 3884
rect 23202 3904 23258 3913
rect 23202 3839 23258 3848
rect 23216 3641 23244 3839
rect 23492 3670 23520 3946
rect 23480 3664 23532 3670
rect 23202 3632 23258 3641
rect 22652 3596 22704 3602
rect 23480 3606 23532 3612
rect 23202 3567 23258 3576
rect 22652 3538 22704 3544
rect 22664 3126 22692 3538
rect 22652 3120 22704 3126
rect 22572 3080 22652 3108
rect 22190 2887 22246 2896
rect 22284 2916 22336 2922
rect 22204 1873 22232 2887
rect 22284 2858 22336 2864
rect 22376 2508 22428 2514
rect 22572 2496 22600 3080
rect 22652 3062 22704 3068
rect 23584 3058 23612 4780
rect 23676 4078 23704 5034
rect 23754 4584 23810 4593
rect 23754 4519 23810 4528
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 22428 2468 22600 2496
rect 22376 2450 22428 2456
rect 22940 2394 22968 2994
rect 23584 2854 23612 2994
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 22572 2378 22968 2394
rect 22468 2372 22520 2378
rect 22468 2314 22520 2320
rect 22572 2372 22980 2378
rect 22572 2366 22928 2372
rect 22190 1864 22246 1873
rect 22190 1799 22246 1808
rect 22100 1488 22152 1494
rect 22100 1430 22152 1436
rect 21916 1284 21968 1290
rect 21916 1226 21968 1232
rect 22008 1284 22060 1290
rect 22008 1226 22060 1232
rect 21824 604 21876 610
rect 21824 546 21876 552
rect 22020 542 22048 1226
rect 22480 800 22508 2314
rect 22572 2310 22600 2366
rect 22928 2314 22980 2320
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 22664 1698 22692 2246
rect 22652 1692 22704 1698
rect 22652 1634 22704 1640
rect 23768 1222 23796 4519
rect 23860 4078 23888 5335
rect 23940 5306 23992 5312
rect 23952 5234 23980 5306
rect 24122 5264 24178 5273
rect 23940 5228 23992 5234
rect 24122 5199 24124 5208
rect 23940 5170 23992 5176
rect 24176 5199 24178 5208
rect 24124 5170 24176 5176
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24044 4622 24072 4966
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 24044 4457 24072 4558
rect 24030 4448 24086 4457
rect 24030 4383 24086 4392
rect 24136 4146 24164 5170
rect 24124 4140 24176 4146
rect 24044 4100 24124 4128
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23860 3534 23888 4014
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 24044 2650 24072 4100
rect 24124 4082 24176 4088
rect 24320 4078 24348 8434
rect 24400 8424 24452 8430
rect 24400 8366 24452 8372
rect 24412 7546 24440 8366
rect 24504 7954 24532 10450
rect 24674 10160 24730 10169
rect 24674 10095 24676 10104
rect 24728 10095 24730 10104
rect 24676 10066 24728 10072
rect 24780 9858 24808 10450
rect 24768 9852 24820 9858
rect 24768 9794 24820 9800
rect 24872 9704 24900 10526
rect 25042 10450 25098 10526
rect 25318 10450 25374 11250
rect 25594 10450 25650 11250
rect 25870 10554 25926 11250
rect 25870 10526 26096 10554
rect 25870 10450 25926 10526
rect 25136 10396 25188 10402
rect 25136 10338 25188 10344
rect 25148 9994 25176 10338
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25332 9926 25360 10450
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25608 9722 25636 10450
rect 25964 9852 26016 9858
rect 25964 9794 26016 9800
rect 24780 9676 24900 9704
rect 25504 9716 25556 9722
rect 24780 8566 24808 9676
rect 25504 9658 25556 9664
rect 25596 9716 25648 9722
rect 25596 9658 25648 9664
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24492 7948 24544 7954
rect 24492 7890 24544 7896
rect 24584 7812 24636 7818
rect 24584 7754 24636 7760
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24412 6254 24440 7482
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 24400 6248 24452 6254
rect 24400 6190 24452 6196
rect 24504 6100 24532 7414
rect 24412 6072 24532 6100
rect 24308 4072 24360 4078
rect 24308 4014 24360 4020
rect 24320 3738 24348 4014
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24122 3088 24178 3097
rect 24122 3023 24124 3032
rect 24176 3023 24178 3032
rect 24124 2994 24176 3000
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24412 1902 24440 6072
rect 24596 5846 24624 7754
rect 24688 6798 24716 8434
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24872 6633 24900 8570
rect 25516 8498 25544 9658
rect 25976 8498 26004 9794
rect 26068 9704 26096 10526
rect 26146 10450 26202 11250
rect 26422 10450 26478 11250
rect 26698 10464 26754 11250
rect 26884 10804 26936 10810
rect 26884 10746 26936 10752
rect 26698 10450 26700 10464
rect 26160 9874 26188 10450
rect 26160 9846 26372 9874
rect 26068 9676 26280 9704
rect 26252 8566 26280 9676
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 25504 8492 25556 8498
rect 25504 8434 25556 8440
rect 25964 8492 26016 8498
rect 25964 8434 26016 8440
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24952 6656 25004 6662
rect 24858 6624 24914 6633
rect 24952 6598 25004 6604
rect 24858 6559 24914 6568
rect 24964 6497 24992 6598
rect 24950 6488 25006 6497
rect 25056 6458 25084 7822
rect 25134 6488 25190 6497
rect 24950 6423 25006 6432
rect 25044 6452 25096 6458
rect 25134 6423 25190 6432
rect 25044 6394 25096 6400
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 24584 5840 24636 5846
rect 24584 5782 24636 5788
rect 24490 5536 24546 5545
rect 24490 5471 24546 5480
rect 24504 5166 24532 5471
rect 24596 5273 24624 5782
rect 24582 5264 24638 5273
rect 24582 5199 24638 5208
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 24582 4176 24638 4185
rect 24582 4111 24638 4120
rect 24400 1896 24452 1902
rect 24400 1838 24452 1844
rect 24596 1834 24624 4111
rect 24688 4078 24716 6258
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 5370 24808 5646
rect 24872 5574 24900 6326
rect 25148 6254 25176 6423
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24780 3641 24808 4558
rect 24766 3632 24822 3641
rect 24766 3567 24822 3576
rect 24872 2922 24900 5510
rect 25056 3670 25084 5510
rect 25148 4865 25176 6190
rect 25240 5409 25268 8366
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25424 8022 25452 8230
rect 25916 8188 26292 8197
rect 25972 8186 25996 8188
rect 26052 8186 26076 8188
rect 26132 8186 26156 8188
rect 26212 8186 26236 8188
rect 25972 8134 25982 8186
rect 26226 8134 26236 8186
rect 25972 8132 25996 8134
rect 26052 8132 26076 8134
rect 26132 8132 26156 8134
rect 26212 8132 26236 8134
rect 25916 8123 26292 8132
rect 25412 8016 25464 8022
rect 25412 7958 25464 7964
rect 25412 7880 25464 7886
rect 25964 7880 26016 7886
rect 25464 7840 25544 7868
rect 25412 7822 25464 7828
rect 25516 7206 25544 7840
rect 25964 7822 26016 7828
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 25976 7721 26004 7822
rect 25962 7712 26018 7721
rect 25962 7647 26018 7656
rect 26252 7546 26280 7822
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26344 7410 26372 9846
rect 26436 7478 26464 10450
rect 26752 10450 26754 10464
rect 26700 10406 26752 10412
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 26528 7970 26556 9658
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 26804 9110 26832 9454
rect 26792 9104 26844 9110
rect 26792 9046 26844 9052
rect 26896 9042 26924 10746
rect 26974 10450 27030 11250
rect 27250 10450 27306 11250
rect 27526 10450 27582 11250
rect 27802 10450 27858 11250
rect 28078 10450 28134 11250
rect 28354 10450 28410 11250
rect 28630 10450 28686 11250
rect 28906 10450 28962 11250
rect 29182 10450 29238 11250
rect 29458 10450 29514 11250
rect 29734 10450 29790 11250
rect 30010 10450 30066 11250
rect 30104 10940 30156 10946
rect 30104 10882 30156 10888
rect 26988 9790 27016 10450
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 26976 9784 27028 9790
rect 26976 9726 27028 9732
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26656 8732 27032 8741
rect 26712 8730 26736 8732
rect 26792 8730 26816 8732
rect 26872 8730 26896 8732
rect 26952 8730 26976 8732
rect 26712 8678 26722 8730
rect 26966 8678 26976 8730
rect 26712 8676 26736 8678
rect 26792 8676 26816 8678
rect 26872 8676 26896 8678
rect 26952 8676 26976 8678
rect 26656 8667 27032 8676
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 26528 7954 26832 7970
rect 26528 7948 26844 7954
rect 26528 7942 26792 7948
rect 26792 7890 26844 7896
rect 26896 7857 26924 8298
rect 26882 7848 26938 7857
rect 26882 7783 26938 7792
rect 27068 7744 27120 7750
rect 27068 7686 27120 7692
rect 26656 7644 27032 7653
rect 26712 7642 26736 7644
rect 26792 7642 26816 7644
rect 26872 7642 26896 7644
rect 26952 7642 26976 7644
rect 26712 7590 26722 7642
rect 26966 7590 26976 7642
rect 26712 7588 26736 7590
rect 26792 7588 26816 7590
rect 26872 7588 26896 7590
rect 26952 7588 26976 7590
rect 26656 7579 27032 7588
rect 27080 7546 27108 7686
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 26424 7472 26476 7478
rect 26424 7414 26476 7420
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26516 7268 26568 7274
rect 26516 7210 26568 7216
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25332 5556 25360 7142
rect 25516 6798 25544 7142
rect 25916 7100 26292 7109
rect 25972 7098 25996 7100
rect 26052 7098 26076 7100
rect 26132 7098 26156 7100
rect 26212 7098 26236 7100
rect 25972 7046 25982 7098
rect 26226 7046 26236 7098
rect 25972 7044 25996 7046
rect 26052 7044 26076 7046
rect 26132 7044 26156 7046
rect 26212 7044 26236 7046
rect 25916 7035 26292 7044
rect 26528 7018 26556 7210
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 26436 6990 26556 7018
rect 26146 6896 26202 6905
rect 26202 6866 26280 6882
rect 26202 6860 26292 6866
rect 26202 6854 26240 6860
rect 26146 6831 26202 6840
rect 26240 6802 26292 6808
rect 26436 6798 26464 6990
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26516 6792 26568 6798
rect 26620 6780 26648 7142
rect 26700 6792 26752 6798
rect 26620 6752 26700 6780
rect 26516 6734 26568 6740
rect 26700 6734 26752 6740
rect 25608 5710 25636 6734
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26436 6322 26464 6598
rect 26528 6458 26556 6734
rect 26656 6556 27032 6565
rect 26712 6554 26736 6556
rect 26792 6554 26816 6556
rect 26872 6554 26896 6556
rect 26952 6554 26976 6556
rect 26712 6502 26722 6554
rect 26966 6502 26976 6554
rect 26712 6500 26736 6502
rect 26792 6500 26816 6502
rect 26872 6500 26896 6502
rect 26952 6500 26976 6502
rect 26656 6491 27032 6500
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 27172 6390 27200 9862
rect 27264 9858 27292 10450
rect 27252 9852 27304 9858
rect 27252 9794 27304 9800
rect 27342 9752 27398 9761
rect 27540 9722 27568 10450
rect 27342 9687 27398 9696
rect 27528 9716 27580 9722
rect 27356 8634 27384 9687
rect 27528 9658 27580 9664
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 27264 7721 27292 8230
rect 27356 7732 27384 8366
rect 27448 7857 27476 9386
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27724 7886 27752 8366
rect 27620 7880 27672 7886
rect 27434 7848 27490 7857
rect 27620 7822 27672 7828
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27434 7783 27490 7792
rect 27250 7712 27306 7721
rect 27356 7704 27476 7732
rect 27250 7647 27306 7656
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 27160 6384 27212 6390
rect 27160 6326 27212 6332
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 26792 6112 26844 6118
rect 26792 6054 26844 6060
rect 25916 6012 26292 6021
rect 25972 6010 25996 6012
rect 26052 6010 26076 6012
rect 26132 6010 26156 6012
rect 26212 6010 26236 6012
rect 25972 5958 25982 6010
rect 26226 5958 26236 6010
rect 25972 5956 25996 5958
rect 26052 5956 26076 5958
rect 26132 5956 26156 5958
rect 26212 5956 26236 5958
rect 25916 5947 26292 5956
rect 26344 5896 26372 6054
rect 26712 5953 26740 6054
rect 26160 5868 26372 5896
rect 26698 5944 26754 5953
rect 26698 5879 26754 5888
rect 25688 5772 25740 5778
rect 25688 5714 25740 5720
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25596 5568 25648 5574
rect 25332 5528 25596 5556
rect 25596 5510 25648 5516
rect 25226 5400 25282 5409
rect 25226 5335 25282 5344
rect 25504 5364 25556 5370
rect 25504 5306 25556 5312
rect 25228 5092 25280 5098
rect 25228 5034 25280 5040
rect 25134 4856 25190 4865
rect 25134 4791 25190 4800
rect 25240 4622 25268 5034
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25228 4480 25280 4486
rect 25228 4422 25280 4428
rect 25240 4282 25268 4422
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25148 3738 25176 4218
rect 25332 4214 25360 4966
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25320 4208 25372 4214
rect 25320 4150 25372 4156
rect 25424 4146 25452 4558
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25516 4026 25544 5306
rect 25596 5160 25648 5166
rect 25596 5102 25648 5108
rect 25608 4486 25636 5102
rect 25596 4480 25648 4486
rect 25596 4422 25648 4428
rect 25424 3998 25544 4026
rect 25596 4004 25648 4010
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25044 3664 25096 3670
rect 25044 3606 25096 3612
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 24952 3052 25004 3058
rect 24952 2994 25004 3000
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24964 2514 24992 2994
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 24584 1828 24636 1834
rect 24584 1770 24636 1776
rect 25056 1698 25084 3334
rect 25240 2446 25268 3470
rect 25424 2825 25452 3998
rect 25596 3946 25648 3952
rect 25608 3777 25636 3946
rect 25594 3768 25650 3777
rect 25594 3703 25650 3712
rect 25700 3602 25728 5714
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 25870 5536 25926 5545
rect 25976 5522 26004 5646
rect 26054 5536 26110 5545
rect 25976 5494 26054 5522
rect 25870 5471 25926 5480
rect 26054 5471 26110 5480
rect 25780 5296 25832 5302
rect 25780 5238 25832 5244
rect 25792 3924 25820 5238
rect 25884 5166 25912 5471
rect 25962 5400 26018 5409
rect 25962 5335 26018 5344
rect 25976 5302 26004 5335
rect 25964 5296 26016 5302
rect 25964 5238 26016 5244
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 26160 5012 26188 5868
rect 26608 5840 26660 5846
rect 26606 5808 26608 5817
rect 26660 5808 26662 5817
rect 26240 5772 26292 5778
rect 26240 5714 26292 5720
rect 26332 5772 26384 5778
rect 26606 5743 26662 5752
rect 26332 5714 26384 5720
rect 26252 5642 26280 5714
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 26344 5556 26372 5714
rect 26804 5556 26832 6054
rect 26988 5794 27016 6190
rect 27264 6089 27292 7414
rect 27342 6760 27398 6769
rect 27342 6695 27398 6704
rect 27250 6080 27306 6089
rect 27250 6015 27306 6024
rect 26988 5766 27200 5794
rect 26994 5704 27046 5710
rect 26344 5528 26832 5556
rect 26896 5664 26994 5692
rect 26896 5556 26924 5664
rect 27172 5692 27200 5766
rect 27252 5704 27304 5710
rect 27172 5664 27252 5692
rect 26994 5646 27046 5652
rect 27252 5646 27304 5652
rect 26896 5528 27108 5556
rect 27080 5522 27108 5528
rect 27080 5494 27200 5522
rect 26656 5468 27032 5477
rect 26712 5466 26736 5468
rect 26792 5466 26816 5468
rect 26872 5466 26896 5468
rect 26952 5466 26976 5468
rect 26712 5414 26722 5466
rect 26966 5414 26976 5466
rect 26712 5412 26736 5414
rect 26792 5412 26816 5414
rect 26872 5412 26896 5414
rect 26952 5412 26976 5414
rect 26514 5400 26570 5409
rect 26656 5403 27032 5412
rect 26570 5344 27108 5352
rect 26514 5335 27108 5344
rect 26528 5324 27108 5335
rect 26698 5264 26754 5273
rect 26608 5228 26660 5234
rect 26698 5199 26754 5208
rect 26974 5264 27030 5273
rect 26974 5199 26976 5208
rect 26608 5170 26660 5176
rect 26424 5024 26476 5030
rect 26160 4984 26372 5012
rect 25916 4924 26292 4933
rect 25972 4922 25996 4924
rect 26052 4922 26076 4924
rect 26132 4922 26156 4924
rect 26212 4922 26236 4924
rect 25972 4870 25982 4922
rect 26226 4870 26236 4922
rect 25972 4868 25996 4870
rect 26052 4868 26076 4870
rect 26132 4868 26156 4870
rect 26212 4868 26236 4870
rect 25916 4859 26292 4868
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 25962 4720 26018 4729
rect 25962 4655 26018 4664
rect 25976 4622 26004 4655
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25964 4480 26016 4486
rect 25964 4422 26016 4428
rect 25870 4312 25926 4321
rect 25870 4247 25926 4256
rect 25884 4214 25912 4247
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25976 4146 26004 4422
rect 26068 4146 26096 4762
rect 26344 4622 26372 4984
rect 26424 4966 26476 4972
rect 26436 4826 26464 4966
rect 26620 4865 26648 5170
rect 26606 4856 26662 4865
rect 26424 4820 26476 4826
rect 26606 4791 26662 4800
rect 26424 4762 26476 4768
rect 26436 4679 26464 4762
rect 26424 4673 26476 4679
rect 26332 4616 26384 4622
rect 26712 4622 26740 5199
rect 27028 5199 27030 5208
rect 26976 5170 27028 5176
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26988 4826 27016 4966
rect 26976 4820 27028 4826
rect 26976 4762 27028 4768
rect 26424 4615 26476 4621
rect 26700 4616 26752 4622
rect 26332 4558 26384 4564
rect 26700 4558 26752 4564
rect 26424 4480 26476 4486
rect 26344 4440 26424 4468
rect 26344 4282 26372 4440
rect 26700 4480 26752 4486
rect 26424 4422 26476 4428
rect 26574 4440 26700 4468
rect 26574 4298 26602 4440
rect 26700 4422 26752 4428
rect 26656 4380 27032 4389
rect 26712 4378 26736 4380
rect 26792 4378 26816 4380
rect 26872 4378 26896 4380
rect 26952 4378 26976 4380
rect 26712 4326 26722 4378
rect 26966 4326 26976 4378
rect 26712 4324 26736 4326
rect 26792 4324 26816 4326
rect 26872 4324 26896 4326
rect 26952 4324 26976 4326
rect 26656 4315 27032 4324
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 26528 4270 26602 4298
rect 27080 4282 27108 5324
rect 27068 4276 27120 4282
rect 26528 4162 26556 4270
rect 27068 4218 27120 4224
rect 25964 4140 26016 4146
rect 25964 4082 26016 4088
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26252 4134 26556 4162
rect 25976 4026 26004 4082
rect 26252 4026 26280 4134
rect 25976 3998 26280 4026
rect 26330 4040 26386 4049
rect 26330 3975 26386 3984
rect 26514 4040 26570 4049
rect 26514 3975 26570 3984
rect 26792 4004 26844 4010
rect 26240 3936 26292 3942
rect 25792 3896 26240 3924
rect 26240 3878 26292 3884
rect 25916 3836 26292 3845
rect 25972 3834 25996 3836
rect 26052 3834 26076 3836
rect 26132 3834 26156 3836
rect 26212 3834 26236 3836
rect 25972 3782 25982 3834
rect 26226 3782 26236 3834
rect 25972 3780 25996 3782
rect 26052 3780 26076 3782
rect 26132 3780 26156 3782
rect 26212 3780 26236 3782
rect 25916 3771 26292 3780
rect 26344 3738 26372 3975
rect 26422 3768 26478 3777
rect 26332 3732 26384 3738
rect 26422 3703 26478 3712
rect 26332 3674 26384 3680
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 26332 3596 26384 3602
rect 26332 3538 26384 3544
rect 25884 3126 25912 3538
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 25410 2816 25466 2825
rect 25410 2751 25466 2760
rect 25916 2748 26292 2757
rect 25972 2746 25996 2748
rect 26052 2746 26076 2748
rect 26132 2746 26156 2748
rect 26212 2746 26236 2748
rect 25972 2694 25982 2746
rect 26226 2694 26236 2746
rect 25972 2692 25996 2694
rect 26052 2692 26076 2694
rect 26132 2692 26156 2694
rect 26212 2692 26236 2694
rect 25778 2680 25834 2689
rect 25916 2683 26292 2692
rect 26344 2650 26372 3538
rect 26436 3194 26464 3703
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 25778 2615 25834 2624
rect 26332 2644 26384 2650
rect 25792 2514 25820 2615
rect 26332 2586 26384 2592
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25044 1692 25096 1698
rect 25044 1634 25096 1640
rect 25240 1562 25268 2382
rect 26436 2378 26464 2926
rect 26528 2922 26556 3975
rect 26792 3946 26844 3952
rect 26606 3904 26662 3913
rect 26606 3839 26662 3848
rect 26620 3602 26648 3839
rect 26804 3602 26832 3946
rect 27172 3913 27200 5494
rect 27356 5234 27384 6695
rect 27448 6497 27476 7704
rect 27632 7342 27660 7822
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27526 6896 27582 6905
rect 27526 6831 27528 6840
rect 27580 6831 27582 6840
rect 27528 6802 27580 6808
rect 27434 6488 27490 6497
rect 27632 6474 27660 7142
rect 27434 6423 27490 6432
rect 27540 6446 27660 6474
rect 27540 6390 27568 6446
rect 27528 6384 27580 6390
rect 27528 6326 27580 6332
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27448 5760 27476 6258
rect 27448 5732 27568 5760
rect 27434 5672 27490 5681
rect 27434 5607 27490 5616
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27342 4856 27398 4865
rect 27342 4791 27398 4800
rect 27356 3942 27384 4791
rect 27448 4622 27476 5607
rect 27540 5030 27568 5732
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27632 4729 27660 6258
rect 27618 4720 27674 4729
rect 27618 4655 27674 4664
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27528 4072 27580 4078
rect 27632 4060 27660 4558
rect 27580 4032 27660 4060
rect 27528 4014 27580 4020
rect 27344 3936 27396 3942
rect 27158 3904 27214 3913
rect 27344 3878 27396 3884
rect 27436 3936 27488 3942
rect 27436 3878 27488 3884
rect 27158 3839 27214 3848
rect 26882 3768 26938 3777
rect 26882 3703 26938 3712
rect 26896 3602 26924 3703
rect 26608 3596 26660 3602
rect 26608 3538 26660 3544
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 26656 3292 27032 3301
rect 26712 3290 26736 3292
rect 26792 3290 26816 3292
rect 26872 3290 26896 3292
rect 26952 3290 26976 3292
rect 26712 3238 26722 3290
rect 26966 3238 26976 3290
rect 26712 3236 26736 3238
rect 26792 3236 26816 3238
rect 26872 3236 26896 3238
rect 26952 3236 26976 3238
rect 26656 3227 27032 3236
rect 26516 2916 26568 2922
rect 26516 2858 26568 2864
rect 27080 2514 27108 3538
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 27344 3392 27396 3398
rect 27344 3334 27396 3340
rect 27172 3194 27200 3334
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27356 3058 27384 3334
rect 27344 3052 27396 3058
rect 27344 2994 27396 3000
rect 27158 2952 27214 2961
rect 27158 2887 27160 2896
rect 27212 2887 27214 2896
rect 27160 2858 27212 2864
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 26656 2204 27032 2213
rect 26712 2202 26736 2204
rect 26792 2202 26816 2204
rect 26872 2202 26896 2204
rect 26952 2202 26976 2204
rect 26712 2150 26722 2202
rect 26966 2150 26976 2202
rect 26712 2148 26736 2150
rect 26792 2148 26816 2150
rect 26872 2148 26896 2150
rect 26952 2148 26976 2150
rect 26656 2139 27032 2148
rect 26238 1864 26294 1873
rect 26238 1799 26294 1808
rect 25228 1556 25280 1562
rect 25228 1498 25280 1504
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 23480 1148 23532 1154
rect 23480 1090 23532 1096
rect 22008 536 22060 542
rect 22008 478 22060 484
rect 22466 0 22522 800
rect 23492 610 23520 1090
rect 23664 1080 23716 1086
rect 23664 1022 23716 1028
rect 23676 800 23704 1022
rect 24872 870 24992 898
rect 24872 800 24900 870
rect 23480 604 23532 610
rect 23480 546 23532 552
rect 23662 0 23718 800
rect 24858 0 24914 800
rect 24964 270 24992 870
rect 26068 870 26188 898
rect 26252 882 26280 1799
rect 27448 1018 27476 3878
rect 27540 3040 27568 4014
rect 27620 3052 27672 3058
rect 27540 3012 27620 3040
rect 27620 2994 27672 3000
rect 27724 2854 27752 7822
rect 27816 6662 27844 10450
rect 27896 9852 27948 9858
rect 27896 9794 27948 9800
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27804 5840 27856 5846
rect 27804 5782 27856 5788
rect 27816 5574 27844 5782
rect 27908 5778 27936 9794
rect 28092 9790 28120 10450
rect 28368 9858 28396 10450
rect 28644 9994 28672 10450
rect 28920 10062 28948 10450
rect 29196 10334 29224 10450
rect 29184 10328 29236 10334
rect 29184 10270 29236 10276
rect 28908 10056 28960 10062
rect 28908 9998 28960 10004
rect 28448 9988 28500 9994
rect 28448 9930 28500 9936
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28356 9852 28408 9858
rect 28356 9794 28408 9800
rect 27988 9784 28040 9790
rect 27988 9726 28040 9732
rect 28080 9784 28132 9790
rect 28080 9726 28132 9732
rect 28000 7478 28028 9726
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28170 8120 28226 8129
rect 28170 8055 28226 8064
rect 28184 7886 28212 8055
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 27988 7472 28040 7478
rect 27988 7414 28040 7420
rect 28184 7206 28212 7822
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28000 7002 28028 7142
rect 28078 7032 28134 7041
rect 27988 6996 28040 7002
rect 28078 6967 28134 6976
rect 27988 6938 28040 6944
rect 28092 6882 28120 6967
rect 28000 6854 28120 6882
rect 28000 6322 28028 6854
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 27896 5772 27948 5778
rect 27896 5714 27948 5720
rect 27988 5636 28040 5642
rect 27988 5578 28040 5584
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 27896 5024 27948 5030
rect 27896 4966 27948 4972
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 27816 4078 27844 4762
rect 27908 4690 27936 4966
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27804 4072 27856 4078
rect 27804 4014 27856 4020
rect 28000 4010 28028 5578
rect 28092 5137 28120 6734
rect 28276 6361 28304 8434
rect 28356 7336 28408 7342
rect 28356 7278 28408 7284
rect 28368 7002 28396 7278
rect 28356 6996 28408 7002
rect 28356 6938 28408 6944
rect 28262 6352 28318 6361
rect 28172 6316 28224 6322
rect 28368 6322 28396 6938
rect 28262 6287 28318 6296
rect 28356 6316 28408 6322
rect 28172 6258 28224 6264
rect 28356 6258 28408 6264
rect 28184 5778 28212 6258
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 28368 5817 28396 6122
rect 28354 5808 28410 5817
rect 28172 5772 28224 5778
rect 28354 5743 28410 5752
rect 28172 5714 28224 5720
rect 28368 5710 28396 5743
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 28170 5400 28226 5409
rect 28170 5335 28226 5344
rect 28078 5128 28134 5137
rect 28078 5063 28134 5072
rect 28184 5030 28212 5335
rect 28276 5234 28304 5510
rect 28264 5228 28316 5234
rect 28264 5170 28316 5176
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 27988 4004 28040 4010
rect 27988 3946 28040 3952
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 28092 1290 28120 4966
rect 28262 4720 28318 4729
rect 28262 4655 28264 4664
rect 28316 4655 28318 4664
rect 28264 4626 28316 4632
rect 28172 4276 28224 4282
rect 28172 4218 28224 4224
rect 28184 3641 28212 4218
rect 28276 4146 28304 4626
rect 28460 4214 28488 9930
rect 29472 9858 29500 10450
rect 29748 10266 29776 10450
rect 30024 10402 30052 10450
rect 30012 10396 30064 10402
rect 30012 10338 30064 10344
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 29644 9988 29696 9994
rect 29644 9930 29696 9936
rect 29276 9852 29328 9858
rect 29276 9794 29328 9800
rect 29460 9852 29512 9858
rect 29460 9794 29512 9800
rect 29092 9784 29144 9790
rect 29092 9726 29144 9732
rect 28632 9648 28684 9654
rect 28632 9590 28684 9596
rect 28540 7336 28592 7342
rect 28540 7278 28592 7284
rect 28552 5098 28580 7278
rect 28644 6934 28672 9590
rect 28722 9480 28778 9489
rect 28722 9415 28778 9424
rect 28632 6928 28684 6934
rect 28632 6870 28684 6876
rect 28630 6624 28686 6633
rect 28630 6559 28686 6568
rect 28644 5166 28672 6559
rect 28736 5409 28764 9415
rect 29000 9104 29052 9110
rect 29000 9046 29052 9052
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 28828 6633 28856 8774
rect 29012 8566 29040 9046
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 29000 8424 29052 8430
rect 29000 8366 29052 8372
rect 29012 7834 29040 8366
rect 28920 7806 29040 7834
rect 28920 7041 28948 7806
rect 29104 7800 29132 9726
rect 29184 9716 29236 9722
rect 29184 9658 29236 9664
rect 29196 8566 29224 9658
rect 29184 8560 29236 8566
rect 29184 8502 29236 8508
rect 29184 7812 29236 7818
rect 29104 7772 29184 7800
rect 29184 7754 29236 7760
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7342 29040 7686
rect 29000 7336 29052 7342
rect 29000 7278 29052 7284
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 28906 7032 28962 7041
rect 28906 6967 28962 6976
rect 29012 6934 29040 7142
rect 29000 6928 29052 6934
rect 29000 6870 29052 6876
rect 29288 6798 29316 9794
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29380 7449 29408 7686
rect 29366 7440 29422 7449
rect 29366 7375 29422 7384
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29000 6724 29052 6730
rect 29000 6666 29052 6672
rect 28814 6624 28870 6633
rect 28814 6559 28870 6568
rect 28906 6216 28962 6225
rect 28816 6180 28868 6186
rect 29012 6202 29040 6666
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 29276 6656 29328 6662
rect 29276 6598 29328 6604
rect 28962 6174 29040 6202
rect 28906 6151 28962 6160
rect 28816 6122 28868 6128
rect 28722 5400 28778 5409
rect 28722 5335 28778 5344
rect 28632 5160 28684 5166
rect 28632 5102 28684 5108
rect 28540 5092 28592 5098
rect 28540 5034 28592 5040
rect 28538 4720 28594 4729
rect 28538 4655 28594 4664
rect 28552 4622 28580 4655
rect 28644 4622 28672 5102
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28448 4208 28500 4214
rect 28552 4185 28580 4558
rect 28724 4208 28776 4214
rect 28448 4150 28500 4156
rect 28538 4176 28594 4185
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 28276 3738 28304 4082
rect 28460 3754 28488 4150
rect 28724 4150 28776 4156
rect 28538 4111 28594 4120
rect 28264 3732 28316 3738
rect 28460 3726 28672 3754
rect 28264 3674 28316 3680
rect 28170 3632 28226 3641
rect 28276 3602 28304 3674
rect 28446 3632 28502 3641
rect 28170 3567 28226 3576
rect 28264 3596 28316 3602
rect 28446 3567 28502 3576
rect 28264 3538 28316 3544
rect 28460 3534 28488 3567
rect 28644 3534 28672 3726
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 28540 3392 28592 3398
rect 28736 3380 28764 4150
rect 28540 3334 28592 3340
rect 28644 3352 28764 3380
rect 28552 3074 28580 3334
rect 28368 3058 28580 3074
rect 28368 3052 28592 3058
rect 28368 3046 28540 3052
rect 28172 2916 28224 2922
rect 28172 2858 28224 2864
rect 28184 2650 28212 2858
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 28368 1426 28396 3046
rect 28540 2994 28592 3000
rect 28448 2984 28500 2990
rect 28644 2938 28672 3352
rect 28828 3194 28856 6122
rect 29196 5914 29224 6598
rect 29184 5908 29236 5914
rect 29184 5850 29236 5856
rect 29182 5808 29238 5817
rect 29182 5743 29238 5752
rect 29196 5574 29224 5743
rect 29288 5624 29316 6598
rect 29380 6322 29408 6802
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 29368 6112 29420 6118
rect 29368 6054 29420 6060
rect 29380 5953 29408 6054
rect 29366 5944 29422 5953
rect 29366 5879 29422 5888
rect 29368 5636 29420 5642
rect 29288 5596 29368 5624
rect 29368 5578 29420 5584
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 28908 5160 28960 5166
rect 29380 5137 29408 5578
rect 29472 5273 29500 7686
rect 29564 7410 29592 8298
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29656 6798 29684 9930
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29552 6656 29604 6662
rect 29552 6598 29604 6604
rect 29458 5264 29514 5273
rect 29458 5199 29514 5208
rect 28908 5102 28960 5108
rect 29366 5128 29422 5137
rect 28920 4690 28948 5102
rect 29366 5063 29422 5072
rect 29460 5092 29512 5098
rect 29460 5034 29512 5040
rect 29184 5024 29236 5030
rect 29184 4966 29236 4972
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28920 4554 28948 4626
rect 29196 4593 29224 4966
rect 29182 4584 29238 4593
rect 28908 4548 28960 4554
rect 29182 4519 29238 4528
rect 28908 4490 28960 4496
rect 29472 4282 29500 5034
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 28906 3768 28962 3777
rect 28906 3703 28962 3712
rect 28816 3188 28868 3194
rect 28816 3130 28868 3136
rect 28500 2932 28672 2938
rect 28448 2926 28672 2932
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 28460 2910 28672 2926
rect 28736 2650 28764 2926
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 28828 2446 28856 2586
rect 28920 2446 28948 3703
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 29472 3126 29500 3470
rect 29460 3120 29512 3126
rect 29460 3062 29512 3068
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29196 2514 29224 2790
rect 29184 2508 29236 2514
rect 29184 2450 29236 2456
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29000 2032 29052 2038
rect 29000 1974 29052 1980
rect 28356 1420 28408 1426
rect 28356 1362 28408 1368
rect 28080 1284 28132 1290
rect 28080 1226 28132 1232
rect 29012 1086 29040 1974
rect 29092 1964 29144 1970
rect 29092 1906 29144 1912
rect 29000 1080 29052 1086
rect 29000 1022 29052 1028
rect 27436 1012 27488 1018
rect 27436 954 27488 960
rect 29104 921 29132 1906
rect 29472 1465 29500 2790
rect 29458 1456 29514 1465
rect 29458 1391 29514 1400
rect 29564 950 29592 6598
rect 29748 6202 29776 9522
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29656 6174 29776 6202
rect 29656 5817 29684 6174
rect 29736 6112 29788 6118
rect 29736 6054 29788 6060
rect 29642 5808 29698 5817
rect 29642 5743 29698 5752
rect 29748 5710 29776 6054
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29736 5228 29788 5234
rect 29736 5170 29788 5176
rect 29748 4758 29776 5170
rect 29736 4752 29788 4758
rect 29736 4694 29788 4700
rect 29840 4282 29868 8910
rect 29920 8492 29972 8498
rect 29920 8434 29972 8440
rect 29932 8090 29960 8434
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29932 7993 29960 8026
rect 29918 7984 29974 7993
rect 29918 7919 29974 7928
rect 29920 7336 29972 7342
rect 29920 7278 29972 7284
rect 29932 6458 29960 7278
rect 30024 6798 30052 9998
rect 30116 8498 30144 10882
rect 30286 10554 30342 11250
rect 30286 10526 30420 10554
rect 30286 10450 30342 10526
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 29920 6452 29972 6458
rect 29920 6394 29972 6400
rect 29920 6180 29972 6186
rect 29920 6122 29972 6128
rect 29932 5846 29960 6122
rect 29920 5840 29972 5846
rect 29920 5782 29972 5788
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 30024 4826 30052 5170
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 30116 4706 30144 7210
rect 30208 5914 30236 7822
rect 30392 7410 30420 10526
rect 30562 10450 30618 11250
rect 30654 10568 30710 10577
rect 30654 10503 30710 10512
rect 30748 10532 30800 10538
rect 30472 10124 30524 10130
rect 30472 10066 30524 10072
rect 30484 8838 30512 10066
rect 30472 8832 30524 8838
rect 30472 8774 30524 8780
rect 30470 7984 30526 7993
rect 30470 7919 30526 7928
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30380 6792 30432 6798
rect 30484 6780 30512 7919
rect 30576 7392 30604 10450
rect 30668 9110 30696 10503
rect 30748 10474 30800 10480
rect 30656 9104 30708 9110
rect 30656 9046 30708 9052
rect 30760 8498 30788 10474
rect 30838 10450 30894 11250
rect 31114 10450 31170 11250
rect 31390 10450 31446 11250
rect 31666 10450 31722 11250
rect 31942 10450 31998 11250
rect 32218 10450 32274 11250
rect 32494 10450 32550 11250
rect 32770 10450 32826 11250
rect 33046 10450 33102 11250
rect 33232 10464 33284 10470
rect 30852 10062 30880 10450
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 31128 9994 31156 10450
rect 31404 10130 31432 10450
rect 31576 10260 31628 10266
rect 31576 10202 31628 10208
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31116 9988 31168 9994
rect 31116 9930 31168 9936
rect 31484 9852 31536 9858
rect 31484 9794 31536 9800
rect 31298 9616 31354 9625
rect 31298 9551 31354 9560
rect 31208 9512 31260 9518
rect 31208 9454 31260 9460
rect 30930 8936 30986 8945
rect 30930 8871 30986 8880
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30944 8378 30972 8871
rect 30668 8350 30972 8378
rect 30668 8294 30696 8350
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 30840 8288 30892 8294
rect 30840 8230 30892 8236
rect 30760 8022 30788 8230
rect 30748 8016 30800 8022
rect 30748 7958 30800 7964
rect 30746 7712 30802 7721
rect 30746 7647 30802 7656
rect 30576 7364 30696 7392
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6798 30604 7142
rect 30432 6752 30512 6780
rect 30564 6792 30616 6798
rect 30380 6734 30432 6740
rect 30564 6734 30616 6740
rect 30300 6322 30328 6734
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30286 5944 30342 5953
rect 30196 5908 30248 5914
rect 30286 5879 30288 5888
rect 30196 5850 30248 5856
rect 30340 5879 30342 5888
rect 30470 5944 30526 5953
rect 30470 5879 30526 5888
rect 30288 5850 30340 5856
rect 30286 5808 30342 5817
rect 30286 5743 30342 5752
rect 30024 4678 30144 4706
rect 29828 4276 29880 4282
rect 29828 4218 29880 4224
rect 29736 3460 29788 3466
rect 29736 3402 29788 3408
rect 29748 2854 29776 3402
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 30024 2106 30052 4678
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 30116 3369 30144 3402
rect 30102 3360 30158 3369
rect 30158 3318 30236 3346
rect 30102 3295 30158 3304
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 30116 2650 30144 2994
rect 30208 2961 30236 3318
rect 30300 3194 30328 5743
rect 30484 5370 30512 5879
rect 30576 5386 30604 6598
rect 30668 6322 30696 7364
rect 30760 7342 30788 7647
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30852 7188 30880 8230
rect 30944 7954 30972 8350
rect 30932 7948 30984 7954
rect 30932 7890 30984 7896
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31036 7410 31064 7822
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 30760 7160 30880 7188
rect 30932 7200 30984 7206
rect 30760 6390 30788 7160
rect 30932 7142 30984 7148
rect 30944 7002 30972 7142
rect 31036 7002 31064 7346
rect 31114 7168 31170 7177
rect 31114 7103 31170 7112
rect 30932 6996 30984 7002
rect 30932 6938 30984 6944
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30932 6792 30984 6798
rect 30932 6734 30984 6740
rect 30748 6384 30800 6390
rect 30748 6326 30800 6332
rect 30656 6316 30708 6322
rect 30656 6258 30708 6264
rect 30852 6186 30880 6734
rect 30944 6361 30972 6734
rect 30930 6352 30986 6361
rect 30930 6287 30986 6296
rect 30840 6180 30892 6186
rect 30840 6122 30892 6128
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 30748 5772 30800 5778
rect 30748 5714 30800 5720
rect 30760 5574 30788 5714
rect 30932 5704 30984 5710
rect 30932 5646 30984 5652
rect 30748 5568 30800 5574
rect 30748 5510 30800 5516
rect 30472 5364 30524 5370
rect 30576 5358 30696 5386
rect 30472 5306 30524 5312
rect 30564 5296 30616 5302
rect 30484 5244 30564 5250
rect 30484 5238 30616 5244
rect 30484 5222 30604 5238
rect 30484 4486 30512 5222
rect 30564 5160 30616 5166
rect 30564 5102 30616 5108
rect 30576 4978 30604 5102
rect 30668 5080 30696 5358
rect 30944 5098 30972 5646
rect 30932 5092 30984 5098
rect 30668 5052 30788 5080
rect 30576 4950 30696 4978
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30484 3942 30512 4082
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30576 3738 30604 4762
rect 30668 4690 30696 4950
rect 30760 4706 30788 5052
rect 30932 5034 30984 5040
rect 30930 4992 30986 5001
rect 30930 4927 30986 4936
rect 30656 4684 30708 4690
rect 30760 4678 30880 4706
rect 30656 4626 30708 4632
rect 30748 4616 30800 4622
rect 30748 4558 30800 4564
rect 30656 4480 30708 4486
rect 30656 4422 30708 4428
rect 30668 4146 30696 4422
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 30564 3732 30616 3738
rect 30564 3674 30616 3680
rect 30760 3670 30788 4558
rect 30748 3664 30800 3670
rect 30748 3606 30800 3612
rect 30472 3392 30524 3398
rect 30472 3334 30524 3340
rect 30288 3188 30340 3194
rect 30288 3130 30340 3136
rect 30484 3058 30512 3334
rect 30746 3088 30802 3097
rect 30472 3052 30524 3058
rect 30746 3023 30748 3032
rect 30472 2994 30524 3000
rect 30800 3023 30802 3032
rect 30748 2994 30800 3000
rect 30194 2952 30250 2961
rect 30194 2887 30250 2896
rect 30484 2774 30512 2994
rect 30392 2746 30512 2774
rect 30104 2644 30156 2650
rect 30104 2586 30156 2592
rect 30392 2514 30420 2746
rect 30380 2508 30432 2514
rect 30380 2450 30432 2456
rect 30012 2100 30064 2106
rect 30012 2042 30064 2048
rect 30852 1154 30880 4678
rect 30944 4185 30972 4927
rect 30930 4176 30986 4185
rect 31036 4146 31064 5850
rect 30930 4111 30986 4120
rect 31024 4140 31076 4146
rect 31024 4082 31076 4088
rect 31128 3738 31156 7103
rect 31220 5370 31248 9454
rect 31312 6798 31340 9551
rect 31392 9444 31444 9450
rect 31392 9386 31444 9392
rect 31404 6866 31432 9386
rect 31496 7410 31524 9794
rect 31588 7410 31616 10202
rect 31680 9654 31708 10450
rect 31852 10328 31904 10334
rect 31852 10270 31904 10276
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 31758 9208 31814 9217
rect 31758 9143 31814 9152
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31680 8106 31708 8910
rect 31772 8294 31800 9143
rect 31864 8498 31892 10270
rect 31956 8548 31984 10450
rect 32128 9988 32180 9994
rect 32232 9976 32260 10450
rect 32232 9948 32444 9976
rect 32128 9930 32180 9936
rect 32140 8974 32168 9930
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 32324 8673 32352 9658
rect 32310 8664 32366 8673
rect 32310 8599 32366 8608
rect 32036 8560 32088 8566
rect 31956 8520 32036 8548
rect 32036 8502 32088 8508
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31916 8188 32292 8197
rect 31972 8186 31996 8188
rect 32052 8186 32076 8188
rect 32132 8186 32156 8188
rect 32212 8186 32236 8188
rect 31972 8134 31982 8186
rect 32226 8134 32236 8186
rect 31972 8132 31996 8134
rect 32052 8132 32076 8134
rect 32132 8132 32156 8134
rect 32212 8132 32236 8134
rect 31916 8123 32292 8132
rect 31680 8078 31800 8106
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31668 7404 31720 7410
rect 31668 7346 31720 7352
rect 31576 6928 31628 6934
rect 31576 6870 31628 6876
rect 31392 6860 31444 6866
rect 31392 6802 31444 6808
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31392 6724 31444 6730
rect 31392 6666 31444 6672
rect 31404 6458 31432 6666
rect 31484 6656 31536 6662
rect 31484 6598 31536 6604
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 31298 6352 31354 6361
rect 31298 6287 31300 6296
rect 31352 6287 31354 6296
rect 31300 6258 31352 6264
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31392 6112 31444 6118
rect 31392 6054 31444 6060
rect 31312 5846 31340 6054
rect 31300 5840 31352 5846
rect 31300 5782 31352 5788
rect 31404 5574 31432 6054
rect 31496 5778 31524 6598
rect 31588 6390 31616 6870
rect 31680 6633 31708 7346
rect 31666 6624 31722 6633
rect 31666 6559 31722 6568
rect 31576 6384 31628 6390
rect 31576 6326 31628 6332
rect 31772 6322 31800 8078
rect 32036 7812 32088 7818
rect 32036 7754 32088 7760
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 32048 7546 32076 7754
rect 31944 7540 31996 7546
rect 31944 7482 31996 7488
rect 32036 7540 32088 7546
rect 32036 7482 32088 7488
rect 31956 7449 31984 7482
rect 31942 7440 31998 7449
rect 31942 7375 31998 7384
rect 32140 7206 32168 7754
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 31916 7100 32292 7109
rect 31972 7098 31996 7100
rect 32052 7098 32076 7100
rect 32132 7098 32156 7100
rect 32212 7098 32236 7100
rect 31972 7046 31982 7098
rect 32226 7046 32236 7098
rect 31972 7044 31996 7046
rect 32052 7044 32076 7046
rect 32132 7044 32156 7046
rect 32212 7044 32236 7046
rect 31916 7035 32292 7044
rect 32036 6996 32088 7002
rect 32036 6938 32088 6944
rect 32220 6996 32272 7002
rect 32220 6938 32272 6944
rect 31850 6624 31906 6633
rect 31850 6559 31906 6568
rect 31864 6322 31892 6559
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31760 6316 31812 6322
rect 31760 6258 31812 6264
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 31576 6180 31628 6186
rect 31576 6122 31628 6128
rect 31484 5772 31536 5778
rect 31484 5714 31536 5720
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 31208 5364 31260 5370
rect 31208 5306 31260 5312
rect 31300 5092 31352 5098
rect 31300 5034 31352 5040
rect 31312 4706 31340 5034
rect 31404 4826 31432 5510
rect 31588 5166 31616 6122
rect 31680 5953 31708 6258
rect 32048 6254 32076 6938
rect 32036 6248 32088 6254
rect 32036 6190 32088 6196
rect 32232 6186 32260 6938
rect 32324 6798 32352 7686
rect 32416 7392 32444 9948
rect 32508 9722 32536 10450
rect 32588 10396 32640 10402
rect 32588 10338 32640 10344
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 32600 9450 32628 10338
rect 32784 10266 32812 10450
rect 32772 10260 32824 10266
rect 32772 10202 32824 10208
rect 33060 9738 33088 10450
rect 33322 10450 33378 11250
rect 33598 10450 33654 11250
rect 33874 10464 33930 11250
rect 34060 10736 34112 10742
rect 34060 10678 34112 10684
rect 33874 10450 33876 10464
rect 33232 10406 33284 10412
rect 33060 9710 33180 9738
rect 32588 9444 32640 9450
rect 32588 9386 32640 9392
rect 32656 8732 33032 8741
rect 32712 8730 32736 8732
rect 32792 8730 32816 8732
rect 32872 8730 32896 8732
rect 32952 8730 32976 8732
rect 32712 8678 32722 8730
rect 32966 8678 32976 8730
rect 32712 8676 32736 8678
rect 32792 8676 32816 8678
rect 32872 8676 32896 8678
rect 32952 8676 32976 8678
rect 32656 8667 33032 8676
rect 33152 8566 33180 9710
rect 33140 8560 33192 8566
rect 33140 8502 33192 8508
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 32968 8129 32996 8366
rect 33048 8288 33100 8294
rect 33100 8248 33180 8276
rect 33048 8230 33100 8236
rect 32954 8120 33010 8129
rect 32588 8084 32640 8090
rect 32954 8055 33010 8064
rect 32588 8026 32640 8032
rect 32600 7460 32628 8026
rect 32968 7954 32996 8055
rect 32956 7948 33008 7954
rect 32956 7890 33008 7896
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 32692 7750 32720 7822
rect 32680 7744 32732 7750
rect 32680 7686 32732 7692
rect 32656 7644 33032 7653
rect 32712 7642 32736 7644
rect 32792 7642 32816 7644
rect 32872 7642 32896 7644
rect 32952 7642 32976 7644
rect 32712 7590 32722 7642
rect 32966 7590 32976 7642
rect 32712 7588 32736 7590
rect 32792 7588 32816 7590
rect 32872 7588 32896 7590
rect 32952 7588 32976 7590
rect 32656 7579 33032 7588
rect 33060 7478 33088 7822
rect 33048 7472 33100 7478
rect 32600 7432 32720 7460
rect 32692 7392 32720 7432
rect 33048 7414 33100 7420
rect 32772 7404 32824 7410
rect 32416 7364 32628 7392
rect 32692 7364 32772 7392
rect 32600 7324 32628 7364
rect 32772 7346 32824 7352
rect 32600 7296 32720 7324
rect 32494 7168 32550 7177
rect 32494 7103 32550 7112
rect 32508 6798 32536 7103
rect 32586 7032 32642 7041
rect 32586 6967 32588 6976
rect 32640 6967 32642 6976
rect 32588 6938 32640 6944
rect 32586 6896 32642 6905
rect 32586 6831 32588 6840
rect 32640 6831 32642 6840
rect 32588 6802 32640 6808
rect 32312 6792 32364 6798
rect 32312 6734 32364 6740
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32312 6656 32364 6662
rect 32312 6598 32364 6604
rect 32496 6656 32548 6662
rect 32496 6598 32548 6604
rect 32220 6180 32272 6186
rect 32220 6122 32272 6128
rect 31916 6012 32292 6021
rect 31972 6010 31996 6012
rect 32052 6010 32076 6012
rect 32132 6010 32156 6012
rect 32212 6010 32236 6012
rect 31972 5958 31982 6010
rect 32226 5958 32236 6010
rect 31972 5956 31996 5958
rect 32052 5956 32076 5958
rect 32132 5956 32156 5958
rect 32212 5956 32236 5958
rect 31666 5944 31722 5953
rect 31916 5947 32292 5956
rect 31666 5879 31722 5888
rect 31680 5710 31708 5879
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 31772 5545 31800 5646
rect 31944 5568 31996 5574
rect 31758 5536 31814 5545
rect 31680 5494 31758 5522
rect 31576 5160 31628 5166
rect 31482 5128 31538 5137
rect 31576 5102 31628 5108
rect 31482 5063 31538 5072
rect 31496 5030 31524 5063
rect 31484 5024 31536 5030
rect 31484 4966 31536 4972
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31312 4678 31524 4706
rect 31496 4622 31524 4678
rect 31484 4616 31536 4622
rect 31298 4584 31354 4593
rect 31484 4558 31536 4564
rect 31298 4519 31300 4528
rect 31352 4519 31354 4528
rect 31300 4490 31352 4496
rect 31496 4282 31524 4558
rect 31484 4276 31536 4282
rect 31484 4218 31536 4224
rect 31116 3732 31168 3738
rect 31116 3674 31168 3680
rect 31128 2514 31156 3674
rect 31588 3602 31616 5102
rect 31680 4214 31708 5494
rect 31944 5510 31996 5516
rect 32034 5536 32090 5545
rect 31758 5471 31814 5480
rect 31758 5400 31814 5409
rect 31758 5335 31760 5344
rect 31812 5335 31814 5344
rect 31760 5306 31812 5312
rect 31956 5234 31984 5510
rect 32034 5471 32090 5480
rect 32048 5302 32076 5471
rect 32036 5296 32088 5302
rect 32036 5238 32088 5244
rect 31944 5228 31996 5234
rect 31944 5170 31996 5176
rect 31916 4924 32292 4933
rect 31972 4922 31996 4924
rect 32052 4922 32076 4924
rect 32132 4922 32156 4924
rect 32212 4922 32236 4924
rect 31972 4870 31982 4922
rect 32226 4870 32236 4922
rect 31972 4868 31996 4870
rect 32052 4868 32076 4870
rect 32132 4868 32156 4870
rect 32212 4868 32236 4870
rect 31916 4859 32292 4868
rect 31760 4684 31812 4690
rect 31760 4626 31812 4632
rect 31668 4208 31720 4214
rect 31668 4150 31720 4156
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31772 2938 31800 4626
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 32232 4010 32260 4082
rect 32220 4004 32272 4010
rect 32220 3946 32272 3952
rect 31916 3836 32292 3845
rect 31972 3834 31996 3836
rect 32052 3834 32076 3836
rect 32132 3834 32156 3836
rect 32212 3834 32236 3836
rect 31972 3782 31982 3834
rect 32226 3782 32236 3834
rect 31972 3780 31996 3782
rect 32052 3780 32076 3782
rect 32132 3780 32156 3782
rect 32212 3780 32236 3782
rect 31916 3771 32292 3780
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 31864 3126 31892 3470
rect 32324 3466 32352 6598
rect 32508 6304 32536 6598
rect 32600 6440 32628 6802
rect 32692 6662 32720 7296
rect 32680 6656 32732 6662
rect 32784 6644 32812 7346
rect 33048 7336 33100 7342
rect 33048 7278 33100 7284
rect 33060 7002 33088 7278
rect 33048 6996 33100 7002
rect 33048 6938 33100 6944
rect 32784 6616 33088 6644
rect 32680 6598 32732 6604
rect 32656 6556 33032 6565
rect 32712 6554 32736 6556
rect 32792 6554 32816 6556
rect 32872 6554 32896 6556
rect 32952 6554 32976 6556
rect 32712 6502 32722 6554
rect 32966 6502 32976 6554
rect 32712 6500 32736 6502
rect 32792 6500 32816 6502
rect 32872 6500 32896 6502
rect 32952 6500 32976 6502
rect 32656 6491 33032 6500
rect 32600 6412 32720 6440
rect 32588 6316 32640 6322
rect 32508 6276 32588 6304
rect 32588 6258 32640 6264
rect 32692 6089 32720 6412
rect 32772 6384 32824 6390
rect 32772 6326 32824 6332
rect 32862 6352 32918 6361
rect 32678 6080 32734 6089
rect 32678 6015 32734 6024
rect 32692 5778 32720 6015
rect 32680 5772 32732 5778
rect 32680 5714 32732 5720
rect 32784 5574 32812 6326
rect 32862 6287 32864 6296
rect 32916 6287 32918 6296
rect 32864 6258 32916 6264
rect 32956 6248 33008 6254
rect 32956 6190 33008 6196
rect 32968 5914 32996 6190
rect 32956 5908 33008 5914
rect 32956 5850 33008 5856
rect 33060 5710 33088 6616
rect 33048 5704 33100 5710
rect 33048 5646 33100 5652
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32656 5468 33032 5477
rect 32712 5466 32736 5468
rect 32792 5466 32816 5468
rect 32872 5466 32896 5468
rect 32952 5466 32976 5468
rect 32712 5414 32722 5466
rect 32966 5414 32976 5466
rect 32712 5412 32736 5414
rect 32792 5412 32816 5414
rect 32872 5412 32896 5414
rect 32952 5412 32976 5414
rect 32656 5403 33032 5412
rect 32404 5228 32456 5234
rect 32404 5170 32456 5176
rect 32416 4865 32444 5170
rect 33048 5024 33100 5030
rect 32494 4992 32550 5001
rect 33048 4966 33100 4972
rect 32494 4927 32550 4936
rect 32402 4856 32458 4865
rect 32402 4791 32458 4800
rect 32404 4684 32456 4690
rect 32508 4672 32536 4927
rect 32588 4820 32640 4826
rect 32588 4762 32640 4768
rect 32456 4644 32536 4672
rect 32404 4626 32456 4632
rect 32600 4622 32628 4762
rect 32954 4720 33010 4729
rect 32954 4655 33010 4664
rect 32588 4616 32640 4622
rect 32588 4558 32640 4564
rect 32680 4616 32732 4622
rect 32732 4576 32812 4604
rect 32680 4558 32732 4564
rect 32784 4468 32812 4576
rect 32968 4486 32996 4655
rect 32600 4440 32812 4468
rect 32956 4480 33008 4486
rect 32600 4264 32628 4440
rect 32956 4422 33008 4428
rect 32656 4380 33032 4389
rect 32712 4378 32736 4380
rect 32792 4378 32816 4380
rect 32872 4378 32896 4380
rect 32952 4378 32976 4380
rect 32712 4326 32722 4378
rect 32966 4326 32976 4378
rect 32712 4324 32736 4326
rect 32792 4324 32816 4326
rect 32872 4324 32896 4326
rect 32952 4324 32976 4326
rect 32656 4315 33032 4324
rect 32508 4236 32628 4264
rect 32772 4276 32824 4282
rect 32312 3460 32364 3466
rect 32312 3402 32364 3408
rect 32402 3224 32458 3233
rect 32508 3194 32536 4236
rect 32772 4218 32824 4224
rect 32586 4176 32642 4185
rect 32586 4111 32588 4120
rect 32640 4111 32642 4120
rect 32588 4082 32640 4088
rect 32588 4004 32640 4010
rect 32588 3946 32640 3952
rect 32600 3777 32628 3946
rect 32784 3913 32812 4218
rect 33060 4078 33088 4966
rect 33152 4282 33180 8248
rect 33244 6798 33272 10406
rect 33336 9926 33364 10450
rect 33506 10024 33562 10033
rect 33506 9959 33562 9968
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 33324 8492 33376 8498
rect 33324 8434 33376 8440
rect 33336 7886 33364 8434
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 33336 7750 33364 7822
rect 33324 7744 33376 7750
rect 33324 7686 33376 7692
rect 33336 7546 33364 7686
rect 33324 7540 33376 7546
rect 33324 7482 33376 7488
rect 33232 6792 33284 6798
rect 33232 6734 33284 6740
rect 33232 6656 33284 6662
rect 33336 6644 33364 7482
rect 33428 7002 33456 7822
rect 33416 6996 33468 7002
rect 33416 6938 33468 6944
rect 33520 6905 33548 9959
rect 33612 8566 33640 10450
rect 33928 10450 33930 10464
rect 33876 10406 33928 10412
rect 33692 9716 33744 9722
rect 33692 9658 33744 9664
rect 33600 8560 33652 8566
rect 33600 8502 33652 8508
rect 33598 7440 33654 7449
rect 33598 7375 33654 7384
rect 33506 6896 33562 6905
rect 33506 6831 33562 6840
rect 33284 6616 33364 6644
rect 33508 6656 33560 6662
rect 33232 6598 33284 6604
rect 33508 6598 33560 6604
rect 33140 4276 33192 4282
rect 33140 4218 33192 4224
rect 33152 4078 33180 4218
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 33244 3924 33272 6598
rect 33520 6254 33548 6598
rect 33508 6248 33560 6254
rect 33508 6190 33560 6196
rect 33416 6180 33468 6186
rect 33416 6122 33468 6128
rect 33324 5228 33376 5234
rect 33324 5170 33376 5176
rect 33336 4826 33364 5170
rect 33324 4820 33376 4826
rect 33324 4762 33376 4768
rect 33428 4706 33456 6122
rect 32770 3904 32826 3913
rect 32770 3839 32826 3848
rect 33152 3896 33272 3924
rect 33336 4678 33456 4706
rect 32586 3768 32642 3777
rect 32586 3703 32642 3712
rect 32402 3159 32458 3168
rect 32496 3188 32548 3194
rect 31852 3120 31904 3126
rect 31852 3062 31904 3068
rect 32310 3088 32366 3097
rect 32416 3058 32444 3159
rect 32496 3130 32548 3136
rect 32600 3058 32628 3703
rect 32954 3632 33010 3641
rect 32954 3567 33010 3576
rect 32968 3534 32996 3567
rect 32956 3528 33008 3534
rect 32956 3470 33008 3476
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32656 3292 33032 3301
rect 32712 3290 32736 3292
rect 32792 3290 32816 3292
rect 32872 3290 32896 3292
rect 32952 3290 32976 3292
rect 32712 3238 32722 3290
rect 32966 3238 32976 3290
rect 32712 3236 32736 3238
rect 32792 3236 32816 3238
rect 32872 3236 32896 3238
rect 32952 3236 32976 3238
rect 32656 3227 33032 3236
rect 32310 3023 32366 3032
rect 32404 3052 32456 3058
rect 31680 2910 31800 2938
rect 31680 2650 31708 2910
rect 31916 2748 32292 2757
rect 31972 2746 31996 2748
rect 32052 2746 32076 2748
rect 32132 2746 32156 2748
rect 32212 2746 32236 2748
rect 31972 2694 31982 2746
rect 32226 2694 32236 2746
rect 31972 2692 31996 2694
rect 32052 2692 32076 2694
rect 32132 2692 32156 2694
rect 32212 2692 32236 2694
rect 31916 2683 32292 2692
rect 31668 2644 31720 2650
rect 31668 2586 31720 2592
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 32128 2508 32180 2514
rect 32128 2450 32180 2456
rect 32140 2310 32168 2450
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 32324 1766 32352 3023
rect 32404 2994 32456 3000
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 33060 2990 33088 3334
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 32656 2204 33032 2213
rect 32712 2202 32736 2204
rect 32792 2202 32816 2204
rect 32872 2202 32896 2204
rect 32952 2202 32976 2204
rect 32712 2150 32722 2202
rect 32966 2150 32976 2202
rect 32712 2148 32736 2150
rect 32792 2148 32816 2150
rect 32872 2148 32896 2150
rect 32952 2148 32976 2150
rect 32656 2139 33032 2148
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 32312 1760 32364 1766
rect 32312 1702 32364 1708
rect 32036 1556 32088 1562
rect 32036 1498 32088 1504
rect 30840 1148 30892 1154
rect 30840 1090 30892 1096
rect 29644 1080 29696 1086
rect 29644 1022 29696 1028
rect 29552 944 29604 950
rect 29090 912 29146 921
rect 26068 800 26096 870
rect 24952 264 25004 270
rect 24952 206 25004 212
rect 26054 0 26110 800
rect 26160 134 26188 870
rect 26240 876 26292 882
rect 26240 818 26292 824
rect 27264 870 27384 898
rect 27264 800 27292 870
rect 26148 128 26200 134
rect 26148 70 26200 76
rect 27250 0 27306 800
rect 27356 202 27384 870
rect 28460 870 28580 898
rect 28460 800 28488 870
rect 27344 196 27396 202
rect 27344 138 27396 144
rect 28446 0 28502 800
rect 28552 338 28580 870
rect 29552 886 29604 892
rect 29090 847 29146 856
rect 29656 800 29684 1022
rect 30852 870 30972 898
rect 30852 800 30880 870
rect 28540 332 28592 338
rect 28540 274 28592 280
rect 29642 0 29698 800
rect 30838 0 30894 800
rect 30944 406 30972 870
rect 32048 800 32076 1498
rect 32784 1329 32812 2042
rect 33048 2032 33100 2038
rect 33048 1974 33100 1980
rect 32770 1320 32826 1329
rect 32770 1255 32826 1264
rect 30932 400 30984 406
rect 30932 342 30984 348
rect 32034 0 32090 800
rect 33060 649 33088 1974
rect 33046 640 33102 649
rect 33152 610 33180 3896
rect 33336 3058 33364 4678
rect 33612 4570 33640 7375
rect 33704 6866 33732 9658
rect 33968 8424 34020 8430
rect 33888 8384 33968 8412
rect 33784 8356 33836 8362
rect 33784 8298 33836 8304
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33692 6724 33744 6730
rect 33692 6666 33744 6672
rect 33704 5234 33732 6666
rect 33692 5228 33744 5234
rect 33692 5170 33744 5176
rect 33692 5024 33744 5030
rect 33692 4966 33744 4972
rect 33428 4542 33640 4570
rect 33428 4185 33456 4542
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33414 4176 33470 4185
rect 33414 4111 33416 4120
rect 33468 4111 33470 4120
rect 33416 4082 33468 4088
rect 33520 3913 33548 4422
rect 33600 4072 33652 4078
rect 33600 4014 33652 4020
rect 33506 3904 33562 3913
rect 33506 3839 33562 3848
rect 33612 3738 33640 4014
rect 33600 3732 33652 3738
rect 33600 3674 33652 3680
rect 33416 3460 33468 3466
rect 33416 3402 33468 3408
rect 33324 3052 33376 3058
rect 33324 2994 33376 3000
rect 33428 2990 33456 3402
rect 33600 3052 33652 3058
rect 33600 2994 33652 3000
rect 33416 2984 33468 2990
rect 33416 2926 33468 2932
rect 33612 2904 33640 2994
rect 33520 2876 33640 2904
rect 33520 2650 33548 2876
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33324 1284 33376 1290
rect 33324 1226 33376 1232
rect 33336 898 33364 1226
rect 33244 870 33364 898
rect 33244 800 33272 870
rect 33046 575 33102 584
rect 33140 604 33192 610
rect 33140 546 33192 552
rect 33230 0 33286 800
rect 33704 785 33732 4966
rect 33796 2514 33824 8298
rect 33888 8265 33916 8384
rect 33968 8366 34020 8372
rect 33874 8256 33930 8265
rect 33874 8191 33930 8200
rect 33876 7744 33928 7750
rect 33876 7686 33928 7692
rect 33888 7342 33916 7686
rect 33876 7336 33928 7342
rect 33876 7278 33928 7284
rect 34072 6780 34100 10678
rect 34150 10450 34206 11250
rect 34426 10450 34482 11250
rect 34702 10450 34758 11250
rect 34978 10450 35034 11250
rect 35254 10450 35310 11250
rect 35530 10450 35586 11250
rect 35806 10450 35862 11250
rect 36082 10450 36138 11250
rect 36358 10450 36414 11250
rect 36634 10450 36690 11250
rect 36910 10450 36966 11250
rect 37004 10872 37056 10878
rect 37004 10814 37056 10820
rect 34164 9722 34192 10450
rect 34336 9852 34388 9858
rect 34336 9794 34388 9800
rect 34152 9716 34204 9722
rect 34152 9658 34204 9664
rect 34152 9240 34204 9246
rect 34152 9182 34204 9188
rect 34164 8498 34192 9182
rect 34244 8900 34296 8906
rect 34244 8842 34296 8848
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 34164 7342 34192 7686
rect 34256 7426 34284 8842
rect 34348 8090 34376 9794
rect 34440 9738 34468 10450
rect 34612 9920 34664 9926
rect 34612 9862 34664 9868
rect 34440 9710 34560 9738
rect 34426 9344 34482 9353
rect 34426 9279 34482 9288
rect 34336 8084 34388 8090
rect 34336 8026 34388 8032
rect 34440 7426 34468 9279
rect 34532 8090 34560 9710
rect 34520 8084 34572 8090
rect 34520 8026 34572 8032
rect 34256 7398 34376 7426
rect 34440 7398 34560 7426
rect 34152 7336 34204 7342
rect 34152 7278 34204 7284
rect 34244 7336 34296 7342
rect 34244 7278 34296 7284
rect 34164 6934 34192 7278
rect 34256 7041 34284 7278
rect 34242 7032 34298 7041
rect 34242 6967 34244 6976
rect 34296 6967 34298 6976
rect 34244 6938 34296 6944
rect 34152 6928 34204 6934
rect 34152 6870 34204 6876
rect 34072 6752 34192 6780
rect 33876 6248 33928 6254
rect 33874 6216 33876 6225
rect 34060 6248 34112 6254
rect 33928 6216 33930 6225
rect 34060 6190 34112 6196
rect 33874 6151 33930 6160
rect 33888 3466 33916 6151
rect 34072 5914 34100 6190
rect 34060 5908 34112 5914
rect 34060 5850 34112 5856
rect 34060 4820 34112 4826
rect 34060 4762 34112 4768
rect 33966 3904 34022 3913
rect 33966 3839 34022 3848
rect 33876 3460 33928 3466
rect 33876 3402 33928 3408
rect 33980 2854 34008 3839
rect 33968 2848 34020 2854
rect 33968 2790 34020 2796
rect 33784 2508 33836 2514
rect 33784 2450 33836 2456
rect 33968 2304 34020 2310
rect 33968 2246 34020 2252
rect 33980 1737 34008 2246
rect 33966 1728 34022 1737
rect 33966 1663 34022 1672
rect 34072 1562 34100 4762
rect 34164 4622 34192 6752
rect 34348 5914 34376 7398
rect 34428 7336 34480 7342
rect 34428 7278 34480 7284
rect 34440 7206 34468 7278
rect 34428 7200 34480 7206
rect 34428 7142 34480 7148
rect 34532 6662 34560 7398
rect 34624 6866 34652 9862
rect 34716 8022 34744 10450
rect 34888 10124 34940 10130
rect 34888 10066 34940 10072
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34808 8498 34836 9998
rect 34900 8498 34928 10066
rect 34992 9926 35020 10450
rect 34980 9920 35032 9926
rect 34980 9862 35032 9868
rect 35268 9858 35296 10450
rect 35438 10432 35494 10441
rect 35438 10367 35494 10376
rect 35348 10192 35400 10198
rect 35348 10134 35400 10140
rect 35360 9858 35388 10134
rect 35256 9852 35308 9858
rect 35256 9794 35308 9800
rect 35348 9852 35400 9858
rect 35348 9794 35400 9800
rect 35452 9654 35480 10367
rect 35544 10130 35572 10450
rect 35714 10296 35770 10305
rect 35714 10231 35770 10240
rect 35532 10124 35584 10130
rect 35532 10066 35584 10072
rect 35624 9716 35676 9722
rect 35624 9658 35676 9664
rect 35440 9648 35492 9654
rect 35440 9590 35492 9596
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 34888 8492 34940 8498
rect 34888 8434 34940 8440
rect 34980 8424 35032 8430
rect 34978 8392 34980 8401
rect 35072 8424 35124 8430
rect 35032 8392 35034 8401
rect 35072 8366 35124 8372
rect 34978 8327 35034 8336
rect 34704 8016 34756 8022
rect 34704 7958 34756 7964
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34612 6180 34664 6186
rect 34612 6122 34664 6128
rect 34520 6112 34572 6118
rect 34520 6054 34572 6060
rect 34336 5908 34388 5914
rect 34336 5850 34388 5856
rect 34532 5710 34560 6054
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34624 5234 34652 6122
rect 34704 5908 34756 5914
rect 34704 5850 34756 5856
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34428 5160 34480 5166
rect 34428 5102 34480 5108
rect 34440 5001 34468 5102
rect 34716 5030 34744 5850
rect 34704 5024 34756 5030
rect 34426 4992 34482 5001
rect 34704 4966 34756 4972
rect 34426 4927 34482 4936
rect 34152 4616 34204 4622
rect 34152 4558 34204 4564
rect 34244 4548 34296 4554
rect 34244 4490 34296 4496
rect 34256 4282 34284 4490
rect 34244 4276 34296 4282
rect 34244 4218 34296 4224
rect 34520 4276 34572 4282
rect 34520 4218 34572 4224
rect 34242 4176 34298 4185
rect 34242 4111 34298 4120
rect 34256 3058 34284 4111
rect 34336 4072 34388 4078
rect 34336 4014 34388 4020
rect 34348 3777 34376 4014
rect 34334 3768 34390 3777
rect 34334 3703 34390 3712
rect 34244 3052 34296 3058
rect 34348 3040 34376 3703
rect 34428 3052 34480 3058
rect 34348 3012 34428 3040
rect 34244 2994 34296 3000
rect 34428 2994 34480 3000
rect 34152 2848 34204 2854
rect 34152 2790 34204 2796
rect 34164 2446 34192 2790
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 34428 2440 34480 2446
rect 34428 2382 34480 2388
rect 34060 1556 34112 1562
rect 34060 1498 34112 1504
rect 34440 1494 34468 2382
rect 34532 2009 34560 4218
rect 34808 3942 34836 7822
rect 34888 7268 34940 7274
rect 34888 7210 34940 7216
rect 34900 6780 34928 7210
rect 34900 6752 35020 6780
rect 34888 6112 34940 6118
rect 34888 6054 34940 6060
rect 34900 5234 34928 6054
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 34992 4468 35020 6752
rect 35084 6730 35112 8366
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35072 6724 35124 6730
rect 35072 6666 35124 6672
rect 35072 6316 35124 6322
rect 35072 6258 35124 6264
rect 35084 5681 35112 6258
rect 35070 5672 35126 5681
rect 35070 5607 35126 5616
rect 35070 4856 35126 4865
rect 35070 4791 35126 4800
rect 35084 4758 35112 4791
rect 35072 4752 35124 4758
rect 35072 4694 35124 4700
rect 34992 4440 35112 4468
rect 34980 4004 35032 4010
rect 34980 3946 35032 3952
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 34992 3738 35020 3946
rect 34980 3732 35032 3738
rect 34980 3674 35032 3680
rect 35084 3602 35112 4440
rect 35072 3596 35124 3602
rect 35072 3538 35124 3544
rect 34888 3528 34940 3534
rect 34888 3470 34940 3476
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34716 3097 34744 3334
rect 34900 3194 34928 3470
rect 35176 3398 35204 7822
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 35268 6769 35296 7346
rect 35254 6760 35310 6769
rect 35360 6730 35388 7822
rect 35440 7812 35492 7818
rect 35440 7754 35492 7760
rect 35452 7206 35480 7754
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 35440 7200 35492 7206
rect 35440 7142 35492 7148
rect 35438 6760 35494 6769
rect 35254 6695 35310 6704
rect 35348 6724 35400 6730
rect 35438 6695 35494 6704
rect 35348 6666 35400 6672
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 35268 5030 35296 6598
rect 35452 5710 35480 6695
rect 35544 6118 35572 7482
rect 35636 6662 35664 9658
rect 35728 8906 35756 10231
rect 35820 9994 35848 10450
rect 36096 10198 36124 10450
rect 36084 10192 36136 10198
rect 36084 10134 36136 10140
rect 36372 10062 36400 10450
rect 36648 10334 36676 10450
rect 36924 10402 36952 10450
rect 36912 10396 36964 10402
rect 36912 10338 36964 10344
rect 36636 10328 36688 10334
rect 36636 10270 36688 10276
rect 36912 10260 36964 10266
rect 36912 10202 36964 10208
rect 36360 10056 36412 10062
rect 36360 9998 36412 10004
rect 35808 9988 35860 9994
rect 35808 9930 35860 9936
rect 36636 9920 36688 9926
rect 36636 9862 36688 9868
rect 35900 9172 35952 9178
rect 35900 9114 35952 9120
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 35716 8900 35768 8906
rect 35716 8842 35768 8848
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35624 6656 35676 6662
rect 35624 6598 35676 6604
rect 35622 6488 35678 6497
rect 35622 6423 35678 6432
rect 35636 6322 35664 6423
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35532 6112 35584 6118
rect 35532 6054 35584 6060
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 35728 5386 35756 7822
rect 35820 7449 35848 9046
rect 35912 8498 35940 9114
rect 36542 8936 36598 8945
rect 36542 8871 36598 8880
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 36556 8242 36584 8871
rect 36648 8362 36676 9862
rect 36924 8498 36952 10202
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36912 8492 36964 8498
rect 36912 8434 36964 8440
rect 36636 8356 36688 8362
rect 36636 8298 36688 8304
rect 36556 8214 36676 8242
rect 36358 8120 36414 8129
rect 36358 8055 36414 8064
rect 35806 7440 35862 7449
rect 36268 7404 36320 7410
rect 35806 7375 35862 7384
rect 36004 7364 36268 7392
rect 35808 6808 35860 6814
rect 35808 6750 35860 6756
rect 35636 5370 35756 5386
rect 35624 5364 35756 5370
rect 35676 5358 35756 5364
rect 35624 5306 35676 5312
rect 35716 5296 35768 5302
rect 35716 5238 35768 5244
rect 35256 5024 35308 5030
rect 35256 4966 35308 4972
rect 35346 4176 35402 4185
rect 35346 4111 35348 4120
rect 35400 4111 35402 4120
rect 35348 4082 35400 4088
rect 35532 4072 35584 4078
rect 35254 4040 35310 4049
rect 35532 4014 35584 4020
rect 35254 3975 35310 3984
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 34888 3188 34940 3194
rect 34888 3130 34940 3136
rect 34702 3088 34758 3097
rect 35268 3058 35296 3975
rect 35544 3738 35572 4014
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35438 3496 35494 3505
rect 35438 3431 35494 3440
rect 34702 3023 34758 3032
rect 35256 3052 35308 3058
rect 35256 2994 35308 3000
rect 35348 2984 35400 2990
rect 35348 2926 35400 2932
rect 34704 2916 34756 2922
rect 34704 2858 34756 2864
rect 34716 2650 34744 2858
rect 34704 2644 34756 2650
rect 34704 2586 34756 2592
rect 35360 2446 35388 2926
rect 35452 2446 35480 3431
rect 35532 2984 35584 2990
rect 35532 2926 35584 2932
rect 35544 2632 35572 2926
rect 35624 2644 35676 2650
rect 35544 2604 35624 2632
rect 35624 2586 35676 2592
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 34518 2000 34574 2009
rect 34518 1935 34574 1944
rect 35728 1698 35756 5238
rect 35820 2106 35848 6750
rect 35900 6248 35952 6254
rect 36004 6236 36032 7364
rect 36268 7346 36320 7352
rect 36082 7304 36138 7313
rect 36372 7274 36400 8055
rect 36452 7880 36504 7886
rect 36452 7822 36504 7828
rect 36544 7880 36596 7886
rect 36544 7822 36596 7828
rect 36464 7750 36492 7822
rect 36452 7744 36504 7750
rect 36452 7686 36504 7692
rect 36082 7239 36138 7248
rect 36360 7268 36412 7274
rect 36096 6866 36124 7239
rect 36360 7210 36412 7216
rect 36556 7002 36584 7822
rect 36544 6996 36596 7002
rect 36544 6938 36596 6944
rect 36648 6866 36676 8214
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36740 7546 36768 7822
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 36084 6860 36136 6866
rect 36084 6802 36136 6808
rect 36544 6860 36596 6866
rect 36544 6802 36596 6808
rect 36636 6860 36688 6866
rect 36636 6802 36688 6808
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 36452 6316 36504 6322
rect 36452 6258 36504 6264
rect 35952 6208 36032 6236
rect 35900 6190 35952 6196
rect 36004 5710 36032 6208
rect 35992 5704 36044 5710
rect 35992 5646 36044 5652
rect 35900 3528 35952 3534
rect 35898 3496 35900 3505
rect 35952 3496 35954 3505
rect 35898 3431 35954 3440
rect 36004 2446 36032 5646
rect 36096 5574 36124 6258
rect 36268 6112 36320 6118
rect 36268 6054 36320 6060
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 36096 5234 36124 5510
rect 36084 5228 36136 5234
rect 36136 5188 36216 5216
rect 36084 5170 36136 5176
rect 36084 4616 36136 4622
rect 36084 4558 36136 4564
rect 36096 4078 36124 4558
rect 36188 4214 36216 5188
rect 36176 4208 36228 4214
rect 36176 4150 36228 4156
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 36188 3584 36216 4150
rect 36280 4078 36308 6054
rect 36464 5778 36492 6258
rect 36556 5914 36584 6802
rect 36648 6118 36676 6802
rect 36832 6202 36860 8434
rect 36912 8288 36964 8294
rect 36912 8230 36964 8236
rect 36740 6174 36860 6202
rect 36636 6112 36688 6118
rect 36636 6054 36688 6060
rect 36544 5908 36596 5914
rect 36544 5850 36596 5856
rect 36452 5772 36504 5778
rect 36452 5714 36504 5720
rect 36464 5234 36492 5714
rect 36636 5296 36688 5302
rect 36636 5238 36688 5244
rect 36452 5228 36504 5234
rect 36452 5170 36504 5176
rect 36358 4720 36414 4729
rect 36358 4655 36414 4664
rect 36372 4622 36400 4655
rect 36360 4616 36412 4622
rect 36360 4558 36412 4564
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 36268 3596 36320 3602
rect 36188 3556 36268 3584
rect 36268 3538 36320 3544
rect 36360 3460 36412 3466
rect 36360 3402 36412 3408
rect 36372 3194 36400 3402
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 35808 2100 35860 2106
rect 35808 2042 35860 2048
rect 35900 1760 35952 1766
rect 35900 1702 35952 1708
rect 35716 1692 35768 1698
rect 35716 1634 35768 1640
rect 34428 1488 34480 1494
rect 34428 1430 34480 1436
rect 34428 1352 34480 1358
rect 34428 1294 34480 1300
rect 34440 800 34468 1294
rect 35912 1154 35940 1702
rect 35900 1148 35952 1154
rect 35900 1090 35952 1096
rect 35636 870 35756 898
rect 35636 800 35664 870
rect 33690 776 33746 785
rect 33690 711 33746 720
rect 34426 0 34482 800
rect 35622 0 35678 800
rect 35728 542 35756 870
rect 36464 678 36492 5170
rect 36648 4826 36676 5238
rect 36636 4820 36688 4826
rect 36636 4762 36688 4768
rect 36544 4752 36596 4758
rect 36544 4694 36596 4700
rect 36634 4720 36690 4729
rect 36556 3618 36584 4694
rect 36634 4655 36690 4664
rect 36648 4486 36676 4655
rect 36636 4480 36688 4486
rect 36636 4422 36688 4428
rect 36740 4010 36768 6174
rect 36924 5098 36952 8230
rect 37016 7546 37044 10814
rect 37096 10668 37148 10674
rect 37096 10610 37148 10616
rect 37108 8004 37136 10610
rect 37186 10450 37242 11250
rect 37280 10464 37332 10470
rect 37200 9722 37228 10450
rect 37462 10450 37518 11250
rect 37738 10464 37794 11250
rect 37738 10450 37740 10464
rect 37280 10406 37332 10412
rect 37188 9716 37240 9722
rect 37188 9658 37240 9664
rect 37292 8498 37320 10406
rect 37476 10266 37504 10450
rect 37792 10450 37794 10464
rect 38014 10450 38070 11250
rect 38290 10450 38346 11250
rect 38566 10450 38622 11250
rect 38842 10450 38898 11250
rect 39118 10450 39174 11250
rect 39394 10450 39450 11250
rect 39670 10554 39726 11250
rect 39670 10526 40172 10554
rect 39670 10450 39726 10526
rect 39764 10464 39816 10470
rect 37740 10406 37792 10412
rect 37464 10260 37516 10266
rect 37464 10202 37516 10208
rect 37832 10192 37884 10198
rect 37832 10134 37884 10140
rect 37556 9988 37608 9994
rect 37556 9930 37608 9936
rect 37370 8528 37426 8537
rect 37280 8492 37332 8498
rect 37370 8463 37426 8472
rect 37280 8434 37332 8440
rect 37188 8016 37240 8022
rect 37108 7976 37188 8004
rect 37188 7958 37240 7964
rect 37004 7540 37056 7546
rect 37004 7482 37056 7488
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 37004 6996 37056 7002
rect 37004 6938 37056 6944
rect 37016 6866 37044 6938
rect 37292 6866 37320 7278
rect 37004 6860 37056 6866
rect 37004 6802 37056 6808
rect 37280 6860 37332 6866
rect 37280 6802 37332 6808
rect 37096 6792 37148 6798
rect 37096 6734 37148 6740
rect 37108 6458 37136 6734
rect 37096 6452 37148 6458
rect 37096 6394 37148 6400
rect 37188 6452 37240 6458
rect 37188 6394 37240 6400
rect 37200 6254 37228 6394
rect 37188 6248 37240 6254
rect 37188 6190 37240 6196
rect 37384 5914 37412 8463
rect 37568 8090 37596 9930
rect 37844 8090 37872 10134
rect 38028 9926 38056 10450
rect 38304 10130 38332 10450
rect 38200 10124 38252 10130
rect 38200 10066 38252 10072
rect 38292 10124 38344 10130
rect 38292 10066 38344 10072
rect 38016 9920 38068 9926
rect 38016 9862 38068 9868
rect 38212 8362 38240 10066
rect 38580 9994 38608 10450
rect 38856 10062 38884 10450
rect 39028 10328 39080 10334
rect 39028 10270 39080 10276
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 38568 9988 38620 9994
rect 38568 9930 38620 9936
rect 38672 8820 38700 9998
rect 39040 9466 39068 10270
rect 39132 9790 39160 10450
rect 39212 10396 39264 10402
rect 39212 10338 39264 10344
rect 39120 9784 39172 9790
rect 39120 9726 39172 9732
rect 39040 9438 39160 9466
rect 38580 8792 38700 8820
rect 38580 8548 38608 8792
rect 38656 8732 39032 8741
rect 38712 8730 38736 8732
rect 38792 8730 38816 8732
rect 38872 8730 38896 8732
rect 38952 8730 38976 8732
rect 38712 8678 38722 8730
rect 38966 8678 38976 8730
rect 38712 8676 38736 8678
rect 38792 8676 38816 8678
rect 38872 8676 38896 8678
rect 38952 8676 38976 8678
rect 38656 8667 39032 8676
rect 38580 8520 38700 8548
rect 38476 8492 38528 8498
rect 38476 8434 38528 8440
rect 38200 8356 38252 8362
rect 38200 8298 38252 8304
rect 37916 8188 38292 8197
rect 37972 8186 37996 8188
rect 38052 8186 38076 8188
rect 38132 8186 38156 8188
rect 38212 8186 38236 8188
rect 37972 8134 37982 8186
rect 38226 8134 38236 8186
rect 37972 8132 37996 8134
rect 38052 8132 38076 8134
rect 38132 8132 38156 8134
rect 38212 8132 38236 8134
rect 37916 8123 38292 8132
rect 37464 8084 37516 8090
rect 37464 8026 37516 8032
rect 37556 8084 37608 8090
rect 37556 8026 37608 8032
rect 37832 8084 37884 8090
rect 37832 8026 37884 8032
rect 37476 7018 37504 8026
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37476 7002 37688 7018
rect 37464 6996 37688 7002
rect 37516 6990 37688 6996
rect 37464 6938 37516 6944
rect 37556 6928 37608 6934
rect 37556 6870 37608 6876
rect 37464 6248 37516 6254
rect 37464 6190 37516 6196
rect 37476 6089 37504 6190
rect 37462 6080 37518 6089
rect 37462 6015 37518 6024
rect 37476 5914 37504 6015
rect 37372 5908 37424 5914
rect 37372 5850 37424 5856
rect 37464 5908 37516 5914
rect 37464 5850 37516 5856
rect 37568 5710 37596 6870
rect 37660 6662 37688 6990
rect 37740 6792 37792 6798
rect 37740 6734 37792 6740
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37752 6497 37780 6734
rect 37738 6488 37794 6497
rect 37738 6423 37794 6432
rect 37740 6316 37792 6322
rect 37740 6258 37792 6264
rect 37648 5840 37700 5846
rect 37648 5782 37700 5788
rect 37556 5704 37608 5710
rect 37556 5646 37608 5652
rect 37464 5636 37516 5642
rect 37464 5578 37516 5584
rect 37476 5234 37504 5578
rect 37464 5228 37516 5234
rect 37464 5170 37516 5176
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 36912 5092 36964 5098
rect 36912 5034 36964 5040
rect 36820 5024 36872 5030
rect 36820 4966 36872 4972
rect 36832 4758 36860 4966
rect 36820 4752 36872 4758
rect 36820 4694 36872 4700
rect 36924 4604 36952 5034
rect 37096 4616 37148 4622
rect 36924 4576 37096 4604
rect 37096 4558 37148 4564
rect 37200 4146 37228 5102
rect 37372 5024 37424 5030
rect 37372 4966 37424 4972
rect 37384 4690 37412 4966
rect 37476 4706 37504 5170
rect 37476 4690 37596 4706
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 37476 4684 37608 4690
rect 37476 4678 37556 4684
rect 37280 4480 37332 4486
rect 37280 4422 37332 4428
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 36728 4004 36780 4010
rect 36728 3946 36780 3952
rect 36556 3590 37136 3618
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 36556 2961 36584 3470
rect 36542 2952 36598 2961
rect 36542 2887 36598 2896
rect 37004 2916 37056 2922
rect 36556 2446 36584 2887
rect 37004 2858 37056 2864
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36912 2372 36964 2378
rect 36912 2314 36964 2320
rect 36924 2038 36952 2314
rect 36912 2032 36964 2038
rect 36912 1974 36964 1980
rect 37016 1193 37044 2858
rect 37108 1698 37136 3590
rect 37188 2984 37240 2990
rect 37188 2926 37240 2932
rect 37096 1692 37148 1698
rect 37096 1634 37148 1640
rect 37002 1184 37058 1193
rect 36820 1148 36872 1154
rect 37002 1119 37058 1128
rect 36820 1090 36872 1096
rect 36832 800 36860 1090
rect 37200 1057 37228 2926
rect 37292 1601 37320 4422
rect 37278 1592 37334 1601
rect 37278 1527 37334 1536
rect 37280 1488 37332 1494
rect 37280 1430 37332 1436
rect 37186 1048 37242 1057
rect 37186 983 37242 992
rect 36452 672 36504 678
rect 36452 614 36504 620
rect 35716 536 35768 542
rect 35716 478 35768 484
rect 36818 0 36874 800
rect 37292 270 37320 1430
rect 37476 746 37504 4678
rect 37556 4626 37608 4632
rect 37660 3534 37688 5782
rect 37752 5642 37780 6258
rect 37740 5636 37792 5642
rect 37740 5578 37792 5584
rect 37844 4026 37872 7822
rect 38384 7336 38436 7342
rect 38384 7278 38436 7284
rect 37916 7100 38292 7109
rect 37972 7098 37996 7100
rect 38052 7098 38076 7100
rect 38132 7098 38156 7100
rect 38212 7098 38236 7100
rect 37972 7046 37982 7098
rect 38226 7046 38236 7098
rect 37972 7044 37996 7046
rect 38052 7044 38076 7046
rect 38132 7044 38156 7046
rect 38212 7044 38236 7046
rect 37916 7035 38292 7044
rect 38396 6322 38424 7278
rect 38384 6316 38436 6322
rect 38384 6258 38436 6264
rect 37916 6012 38292 6021
rect 37972 6010 37996 6012
rect 38052 6010 38076 6012
rect 38132 6010 38156 6012
rect 38212 6010 38236 6012
rect 37972 5958 37982 6010
rect 38226 5958 38236 6010
rect 37972 5956 37996 5958
rect 38052 5956 38076 5958
rect 38132 5956 38156 5958
rect 38212 5956 38236 5958
rect 37916 5947 38292 5956
rect 38200 5772 38252 5778
rect 38200 5714 38252 5720
rect 38212 5642 38240 5714
rect 38200 5636 38252 5642
rect 38200 5578 38252 5584
rect 37916 4924 38292 4933
rect 37972 4922 37996 4924
rect 38052 4922 38076 4924
rect 38132 4922 38156 4924
rect 38212 4922 38236 4924
rect 37972 4870 37982 4922
rect 38226 4870 38236 4922
rect 37972 4868 37996 4870
rect 38052 4868 38076 4870
rect 38132 4868 38156 4870
rect 38212 4868 38236 4870
rect 37916 4859 38292 4868
rect 38396 4808 38424 6258
rect 38488 5250 38516 8434
rect 38672 8362 38700 8520
rect 39132 8362 39160 9438
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 39120 8356 39172 8362
rect 39120 8298 39172 8304
rect 39224 8090 39252 10338
rect 39408 9722 39436 10450
rect 39764 10406 39816 10412
rect 39488 10260 39540 10266
rect 39488 10202 39540 10208
rect 39304 9716 39356 9722
rect 39304 9658 39356 9664
rect 39396 9716 39448 9722
rect 39396 9658 39448 9664
rect 39316 8362 39344 9658
rect 39396 8492 39448 8498
rect 39396 8434 39448 8440
rect 39304 8356 39356 8362
rect 39304 8298 39356 8304
rect 39212 8084 39264 8090
rect 39212 8026 39264 8032
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 38656 7644 39032 7653
rect 38712 7642 38736 7644
rect 38792 7642 38816 7644
rect 38872 7642 38896 7644
rect 38952 7642 38976 7644
rect 38712 7590 38722 7642
rect 38966 7590 38976 7642
rect 38712 7588 38736 7590
rect 38792 7588 38816 7590
rect 38872 7588 38896 7590
rect 38952 7588 38976 7590
rect 38656 7579 39032 7588
rect 38752 7404 38804 7410
rect 38752 7346 38804 7352
rect 38660 7268 38712 7274
rect 38660 7210 38712 7216
rect 38568 6996 38620 7002
rect 38568 6938 38620 6944
rect 38580 6798 38608 6938
rect 38568 6792 38620 6798
rect 38568 6734 38620 6740
rect 38672 6644 38700 7210
rect 38764 6866 38792 7346
rect 39028 7268 39080 7274
rect 39028 7210 39080 7216
rect 39040 7002 39068 7210
rect 39028 6996 39080 7002
rect 39028 6938 39080 6944
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38750 6760 38806 6769
rect 38750 6695 38806 6704
rect 38764 6662 38792 6695
rect 38580 6616 38700 6644
rect 38752 6656 38804 6662
rect 38580 6338 38608 6616
rect 38752 6598 38804 6604
rect 38656 6556 39032 6565
rect 38712 6554 38736 6556
rect 38792 6554 38816 6556
rect 38872 6554 38896 6556
rect 38952 6554 38976 6556
rect 38712 6502 38722 6554
rect 38966 6502 38976 6554
rect 38712 6500 38736 6502
rect 38792 6500 38816 6502
rect 38872 6500 38896 6502
rect 38952 6500 38976 6502
rect 38656 6491 39032 6500
rect 38580 6322 38700 6338
rect 38580 6316 38712 6322
rect 38580 6310 38660 6316
rect 38660 6258 38712 6264
rect 38656 5468 39032 5477
rect 38712 5466 38736 5468
rect 38792 5466 38816 5468
rect 38872 5466 38896 5468
rect 38952 5466 38976 5468
rect 38712 5414 38722 5466
rect 38966 5414 38976 5466
rect 38712 5412 38736 5414
rect 38792 5412 38816 5414
rect 38872 5412 38896 5414
rect 38952 5412 38976 5414
rect 38656 5403 39032 5412
rect 38488 5222 38608 5250
rect 38474 5128 38530 5137
rect 38474 5063 38476 5072
rect 38528 5063 38530 5072
rect 38476 5034 38528 5040
rect 38304 4780 38424 4808
rect 38304 4729 38332 4780
rect 38290 4720 38346 4729
rect 38290 4655 38346 4664
rect 38384 4684 38436 4690
rect 38384 4626 38436 4632
rect 37752 3998 37872 4026
rect 37648 3528 37700 3534
rect 37648 3470 37700 3476
rect 37752 3466 37780 3998
rect 37832 3936 37884 3942
rect 37832 3878 37884 3884
rect 37740 3460 37792 3466
rect 37740 3402 37792 3408
rect 37844 1970 37872 3878
rect 37916 3836 38292 3845
rect 37972 3834 37996 3836
rect 38052 3834 38076 3836
rect 38132 3834 38156 3836
rect 38212 3834 38236 3836
rect 37972 3782 37982 3834
rect 38226 3782 38236 3834
rect 37972 3780 37996 3782
rect 38052 3780 38076 3782
rect 38132 3780 38156 3782
rect 38212 3780 38236 3782
rect 37916 3771 38292 3780
rect 38292 3528 38344 3534
rect 38396 3516 38424 4626
rect 38476 3664 38528 3670
rect 38476 3606 38528 3612
rect 38344 3488 38424 3516
rect 38292 3470 38344 3476
rect 38304 2854 38332 3470
rect 38488 3194 38516 3606
rect 38476 3188 38528 3194
rect 38476 3130 38528 3136
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38292 2848 38344 2854
rect 38292 2790 38344 2796
rect 37916 2748 38292 2757
rect 37972 2746 37996 2748
rect 38052 2746 38076 2748
rect 38132 2746 38156 2748
rect 38212 2746 38236 2748
rect 37972 2694 37982 2746
rect 38226 2694 38236 2746
rect 37972 2692 37996 2694
rect 38052 2692 38076 2694
rect 38132 2692 38156 2694
rect 38212 2692 38236 2694
rect 37916 2683 38292 2692
rect 37832 1964 37884 1970
rect 37832 1906 37884 1912
rect 38016 1216 38068 1222
rect 38016 1158 38068 1164
rect 38028 800 38056 1158
rect 38396 1086 38424 2994
rect 38580 2854 38608 5222
rect 38660 5024 38712 5030
rect 38660 4966 38712 4972
rect 38672 4622 38700 4966
rect 38660 4616 38712 4622
rect 38660 4558 38712 4564
rect 38656 4380 39032 4389
rect 38712 4378 38736 4380
rect 38792 4378 38816 4380
rect 38872 4378 38896 4380
rect 38952 4378 38976 4380
rect 38712 4326 38722 4378
rect 38966 4326 38976 4378
rect 38712 4324 38736 4326
rect 38792 4324 38816 4326
rect 38872 4324 38896 4326
rect 38952 4324 38976 4326
rect 38656 4315 39032 4324
rect 38752 4140 38804 4146
rect 38752 4082 38804 4088
rect 38764 3942 38792 4082
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 38764 3670 38792 3878
rect 38752 3664 38804 3670
rect 38752 3606 38804 3612
rect 38764 3466 38792 3606
rect 38752 3460 38804 3466
rect 38752 3402 38804 3408
rect 38656 3292 39032 3301
rect 38712 3290 38736 3292
rect 38792 3290 38816 3292
rect 38872 3290 38896 3292
rect 38952 3290 38976 3292
rect 38712 3238 38722 3290
rect 38966 3238 38976 3290
rect 38712 3236 38736 3238
rect 38792 3236 38816 3238
rect 38872 3236 38896 3238
rect 38952 3236 38976 3238
rect 38656 3227 39032 3236
rect 39132 3194 39160 7822
rect 39304 7812 39356 7818
rect 39304 7754 39356 7760
rect 39212 7744 39264 7750
rect 39212 7686 39264 7692
rect 39224 7002 39252 7686
rect 39316 7546 39344 7754
rect 39304 7540 39356 7546
rect 39304 7482 39356 7488
rect 39304 7404 39356 7410
rect 39304 7346 39356 7352
rect 39212 6996 39264 7002
rect 39212 6938 39264 6944
rect 39316 6254 39344 7346
rect 39304 6248 39356 6254
rect 39304 6190 39356 6196
rect 39212 6180 39264 6186
rect 39212 6122 39264 6128
rect 39224 5914 39252 6122
rect 39212 5908 39264 5914
rect 39212 5850 39264 5856
rect 39212 5704 39264 5710
rect 39212 5646 39264 5652
rect 39224 5234 39252 5646
rect 39304 5568 39356 5574
rect 39304 5510 39356 5516
rect 39212 5228 39264 5234
rect 39212 5170 39264 5176
rect 39212 4072 39264 4078
rect 39212 4014 39264 4020
rect 39224 3466 39252 4014
rect 39316 3534 39344 5510
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 39212 3460 39264 3466
rect 39212 3402 39264 3408
rect 39120 3188 39172 3194
rect 39120 3130 39172 3136
rect 39408 3126 39436 8434
rect 39500 8022 39528 10202
rect 39580 8968 39632 8974
rect 39580 8910 39632 8916
rect 39592 8498 39620 8910
rect 39580 8492 39632 8498
rect 39580 8434 39632 8440
rect 39776 8090 39804 10406
rect 40040 10124 40092 10130
rect 40040 10066 40092 10072
rect 39948 9920 40000 9926
rect 39948 9862 40000 9868
rect 39856 9648 39908 9654
rect 39856 9590 39908 9596
rect 39764 8084 39816 8090
rect 39764 8026 39816 8032
rect 39488 8016 39540 8022
rect 39488 7958 39540 7964
rect 39672 7880 39724 7886
rect 39672 7822 39724 7828
rect 39488 7404 39540 7410
rect 39540 7364 39620 7392
rect 39488 7346 39540 7352
rect 39592 6769 39620 7364
rect 39578 6760 39634 6769
rect 39578 6695 39634 6704
rect 39592 6322 39620 6695
rect 39580 6316 39632 6322
rect 39580 6258 39632 6264
rect 39684 6202 39712 7822
rect 39868 6934 39896 9590
rect 39960 8362 39988 9862
rect 40052 8362 40080 10066
rect 39948 8356 40000 8362
rect 39948 8298 40000 8304
rect 40040 8356 40092 8362
rect 40040 8298 40092 8304
rect 40144 8090 40172 10526
rect 42524 10396 42576 10402
rect 42524 10338 42576 10344
rect 41052 10056 41104 10062
rect 41052 9998 41104 10004
rect 40684 9988 40736 9994
rect 40684 9930 40736 9936
rect 40316 9716 40368 9722
rect 40316 9658 40368 9664
rect 40224 8560 40276 8566
rect 40224 8502 40276 8508
rect 40132 8084 40184 8090
rect 40132 8026 40184 8032
rect 40132 7880 40184 7886
rect 40132 7822 40184 7828
rect 39856 6928 39908 6934
rect 39856 6870 39908 6876
rect 39764 6860 39816 6866
rect 39764 6802 39816 6808
rect 39776 6458 39804 6802
rect 40144 6662 40172 7822
rect 40132 6656 40184 6662
rect 40132 6598 40184 6604
rect 39764 6452 39816 6458
rect 39764 6394 39816 6400
rect 39500 6174 39712 6202
rect 39764 6248 39816 6254
rect 39764 6190 39816 6196
rect 39948 6248 40000 6254
rect 39948 6190 40000 6196
rect 39500 4214 39528 6174
rect 39776 6118 39804 6190
rect 39764 6112 39816 6118
rect 39764 6054 39816 6060
rect 39672 5636 39724 5642
rect 39672 5578 39724 5584
rect 39488 4208 39540 4214
rect 39488 4150 39540 4156
rect 39580 4208 39632 4214
rect 39580 4150 39632 4156
rect 39488 4072 39540 4078
rect 39488 4014 39540 4020
rect 39396 3120 39448 3126
rect 39396 3062 39448 3068
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 38568 2848 38620 2854
rect 38568 2790 38620 2796
rect 38656 2204 39032 2213
rect 38712 2202 38736 2204
rect 38792 2202 38816 2204
rect 38872 2202 38896 2204
rect 38952 2202 38976 2204
rect 38712 2150 38722 2202
rect 38966 2150 38976 2202
rect 38712 2148 38736 2150
rect 38792 2148 38816 2150
rect 38872 2148 38896 2150
rect 38952 2148 38976 2150
rect 38656 2139 39032 2148
rect 39132 1562 39160 2994
rect 39396 2984 39448 2990
rect 39396 2926 39448 2932
rect 39408 2553 39436 2926
rect 39394 2544 39450 2553
rect 39304 2508 39356 2514
rect 39394 2479 39450 2488
rect 39304 2450 39356 2456
rect 39120 1556 39172 1562
rect 39120 1498 39172 1504
rect 39212 1284 39264 1290
rect 39212 1226 39264 1232
rect 38384 1080 38436 1086
rect 38384 1022 38436 1028
rect 39224 800 39252 1226
rect 39316 814 39344 2450
rect 39500 2394 39528 4014
rect 39408 2366 39528 2394
rect 39408 1834 39436 2366
rect 39488 2304 39540 2310
rect 39488 2246 39540 2252
rect 39396 1828 39448 1834
rect 39396 1770 39448 1776
rect 39304 808 39356 814
rect 37464 740 37516 746
rect 37464 682 37516 688
rect 37280 264 37332 270
rect 37280 206 37332 212
rect 38014 0 38070 800
rect 39210 0 39266 800
rect 39304 750 39356 756
rect 39500 513 39528 2246
rect 39592 1154 39620 4150
rect 39684 1766 39712 5578
rect 39764 4820 39816 4826
rect 39764 4762 39816 4768
rect 39776 4282 39804 4762
rect 39764 4276 39816 4282
rect 39764 4218 39816 4224
rect 39960 2417 39988 6190
rect 40236 5710 40264 8502
rect 40328 7546 40356 9658
rect 40500 9308 40552 9314
rect 40500 9250 40552 9256
rect 40408 7812 40460 7818
rect 40408 7754 40460 7760
rect 40316 7540 40368 7546
rect 40316 7482 40368 7488
rect 40224 5704 40276 5710
rect 40224 5646 40276 5652
rect 40420 3194 40448 7754
rect 40512 6458 40540 9250
rect 40696 8294 40724 9930
rect 41064 8294 41092 9998
rect 41696 9784 41748 9790
rect 41696 9726 41748 9732
rect 41144 9036 41196 9042
rect 41144 8978 41196 8984
rect 41156 8294 41184 8978
rect 41420 8492 41472 8498
rect 41420 8434 41472 8440
rect 41604 8492 41656 8498
rect 41604 8434 41656 8440
rect 41328 8356 41380 8362
rect 41328 8298 41380 8304
rect 40684 8288 40736 8294
rect 40684 8230 40736 8236
rect 41052 8288 41104 8294
rect 41052 8230 41104 8236
rect 41144 8288 41196 8294
rect 41144 8230 41196 8236
rect 41340 8022 41368 8298
rect 41328 8016 41380 8022
rect 41328 7958 41380 7964
rect 40682 7848 40738 7857
rect 40682 7783 40738 7792
rect 40696 7546 40724 7783
rect 40684 7540 40736 7546
rect 40684 7482 40736 7488
rect 41144 6996 41196 7002
rect 41144 6938 41196 6944
rect 40500 6452 40552 6458
rect 40500 6394 40552 6400
rect 40958 3496 41014 3505
rect 40958 3431 41014 3440
rect 40408 3188 40460 3194
rect 40408 3130 40460 3136
rect 40592 3052 40644 3058
rect 40592 2994 40644 3000
rect 39946 2408 40002 2417
rect 39946 2343 40002 2352
rect 39672 1760 39724 1766
rect 39672 1702 39724 1708
rect 40040 1692 40092 1698
rect 40040 1634 40092 1640
rect 39580 1148 39632 1154
rect 39580 1090 39632 1096
rect 39486 504 39542 513
rect 39486 439 39542 448
rect 40052 338 40080 1634
rect 40604 1426 40632 2994
rect 40972 2922 41000 3431
rect 41156 3194 41184 6938
rect 41432 3670 41460 8434
rect 41512 8424 41564 8430
rect 41512 8366 41564 8372
rect 41524 8090 41552 8366
rect 41512 8084 41564 8090
rect 41512 8026 41564 8032
rect 41512 7880 41564 7886
rect 41512 7822 41564 7828
rect 41524 3738 41552 7822
rect 41512 3732 41564 3738
rect 41512 3674 41564 3680
rect 41420 3664 41472 3670
rect 41420 3606 41472 3612
rect 41616 3194 41644 8434
rect 41708 8362 41736 9726
rect 41788 8560 41840 8566
rect 41788 8502 41840 8508
rect 41696 8356 41748 8362
rect 41696 8298 41748 8304
rect 41696 8016 41748 8022
rect 41696 7958 41748 7964
rect 41708 6914 41736 7958
rect 41800 7546 41828 8502
rect 42432 8288 42484 8294
rect 42432 8230 42484 8236
rect 42154 7984 42210 7993
rect 42154 7919 42210 7928
rect 42168 7886 42196 7919
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 42156 7880 42208 7886
rect 42156 7822 42208 7828
rect 41788 7540 41840 7546
rect 41788 7482 41840 7488
rect 41708 6886 41828 6914
rect 41696 6792 41748 6798
rect 41696 6734 41748 6740
rect 41144 3188 41196 3194
rect 41144 3130 41196 3136
rect 41604 3188 41656 3194
rect 41604 3130 41656 3136
rect 41708 3074 41736 6734
rect 41800 3942 41828 6886
rect 41892 6866 41920 7822
rect 42156 7744 42208 7750
rect 42156 7686 42208 7692
rect 41972 7268 42024 7274
rect 41972 7210 42024 7216
rect 42064 7268 42116 7274
rect 42064 7210 42116 7216
rect 41880 6860 41932 6866
rect 41880 6802 41932 6808
rect 41880 5704 41932 5710
rect 41880 5646 41932 5652
rect 41788 3936 41840 3942
rect 41788 3878 41840 3884
rect 41892 3194 41920 5646
rect 41984 4010 42012 7210
rect 42076 7002 42104 7210
rect 42064 6996 42116 7002
rect 42064 6938 42116 6944
rect 42168 4214 42196 7686
rect 42444 7410 42472 8230
rect 42536 7886 42564 10338
rect 43534 9888 43590 9897
rect 43534 9823 43590 9832
rect 43350 9616 43406 9625
rect 43350 9551 43406 9560
rect 43258 9344 43314 9353
rect 43258 9279 43314 9288
rect 43166 9072 43222 9081
rect 43166 9007 43222 9016
rect 42616 8968 42668 8974
rect 42616 8910 42668 8916
rect 42524 7880 42576 7886
rect 42524 7822 42576 7828
rect 42248 7404 42300 7410
rect 42248 7346 42300 7352
rect 42432 7404 42484 7410
rect 42432 7346 42484 7352
rect 42156 4208 42208 4214
rect 42156 4150 42208 4156
rect 42064 4140 42116 4146
rect 42064 4082 42116 4088
rect 41972 4004 42024 4010
rect 41972 3946 42024 3952
rect 41972 3460 42024 3466
rect 41972 3402 42024 3408
rect 41984 3194 42012 3402
rect 41880 3188 41932 3194
rect 41880 3130 41932 3136
rect 41972 3188 42024 3194
rect 41972 3130 42024 3136
rect 41328 3052 41380 3058
rect 41328 2994 41380 3000
rect 41420 3052 41472 3058
rect 41420 2994 41472 3000
rect 41616 3046 41736 3074
rect 41972 3052 42024 3058
rect 40960 2916 41012 2922
rect 40960 2858 41012 2864
rect 40592 1420 40644 1426
rect 40592 1362 40644 1368
rect 40408 1352 40460 1358
rect 40408 1294 40460 1300
rect 40420 800 40448 1294
rect 40040 332 40092 338
rect 40040 274 40092 280
rect 40406 0 40462 800
rect 41340 202 41368 2994
rect 41432 1358 41460 2994
rect 41420 1352 41472 1358
rect 41420 1294 41472 1300
rect 41616 800 41644 3046
rect 41972 2994 42024 3000
rect 41984 1698 42012 2994
rect 41972 1692 42024 1698
rect 41972 1634 42024 1640
rect 41328 196 41380 202
rect 41328 138 41380 144
rect 41602 0 41658 800
rect 42076 406 42104 4082
rect 42260 3210 42288 7346
rect 42340 7336 42392 7342
rect 42340 7278 42392 7284
rect 42352 7002 42380 7278
rect 42340 6996 42392 7002
rect 42340 6938 42392 6944
rect 42628 6458 42656 8910
rect 42984 8900 43036 8906
rect 42984 8842 43036 8848
rect 42708 8832 42760 8838
rect 42708 8774 42760 8780
rect 42798 8800 42854 8809
rect 42720 8498 42748 8774
rect 42798 8735 42854 8744
rect 42812 8634 42840 8735
rect 42800 8628 42852 8634
rect 42800 8570 42852 8576
rect 42996 8498 43024 8842
rect 42708 8492 42760 8498
rect 42708 8434 42760 8440
rect 42984 8492 43036 8498
rect 42984 8434 43036 8440
rect 43076 8356 43128 8362
rect 43076 8298 43128 8304
rect 43088 8265 43116 8298
rect 43074 8256 43130 8265
rect 43074 8191 43130 8200
rect 43180 8090 43208 9007
rect 43168 8084 43220 8090
rect 43168 8026 43220 8032
rect 42890 7984 42946 7993
rect 42890 7919 42946 7928
rect 42800 7812 42852 7818
rect 42800 7754 42852 7760
rect 42708 6792 42760 6798
rect 42708 6734 42760 6740
rect 42616 6452 42668 6458
rect 42616 6394 42668 6400
rect 42720 5817 42748 6734
rect 42812 6662 42840 7754
rect 42904 7546 42932 7919
rect 42984 7880 43036 7886
rect 42984 7822 43036 7828
rect 42892 7540 42944 7546
rect 42892 7482 42944 7488
rect 42890 7440 42946 7449
rect 42890 7375 42892 7384
rect 42944 7375 42946 7384
rect 42892 7346 42944 7352
rect 42996 6730 43024 7822
rect 43076 7744 43128 7750
rect 43076 7686 43128 7692
rect 43088 7449 43116 7686
rect 43272 7546 43300 9279
rect 43364 8022 43392 9551
rect 43444 8628 43496 8634
rect 43444 8570 43496 8576
rect 43456 8537 43484 8570
rect 43442 8528 43498 8537
rect 43442 8463 43498 8472
rect 43352 8016 43404 8022
rect 43352 7958 43404 7964
rect 43548 7954 43576 9823
rect 43628 9376 43680 9382
rect 43628 9318 43680 9324
rect 43536 7948 43588 7954
rect 43536 7890 43588 7896
rect 43444 7744 43496 7750
rect 43442 7712 43444 7721
rect 43496 7712 43498 7721
rect 43442 7647 43498 7656
rect 43260 7540 43312 7546
rect 43260 7482 43312 7488
rect 43074 7440 43130 7449
rect 43074 7375 43130 7384
rect 43444 7200 43496 7206
rect 43442 7168 43444 7177
rect 43496 7168 43498 7177
rect 43442 7103 43498 7112
rect 43640 6914 43668 9318
rect 43442 6896 43498 6905
rect 43442 6831 43498 6840
rect 43548 6886 43668 6914
rect 43074 6760 43130 6769
rect 42984 6724 43036 6730
rect 43074 6695 43076 6704
rect 42984 6666 43036 6672
rect 43128 6695 43130 6704
rect 43076 6666 43128 6672
rect 43456 6662 43484 6831
rect 42800 6656 42852 6662
rect 42892 6656 42944 6662
rect 42800 6598 42852 6604
rect 42890 6624 42892 6633
rect 43444 6656 43496 6662
rect 42944 6624 42946 6633
rect 43444 6598 43496 6604
rect 42890 6559 42946 6568
rect 43444 6452 43496 6458
rect 43444 6394 43496 6400
rect 43456 6361 43484 6394
rect 43442 6352 43498 6361
rect 42800 6316 42852 6322
rect 42800 6258 42852 6264
rect 43352 6316 43404 6322
rect 43442 6287 43498 6296
rect 43352 6258 43404 6264
rect 42706 5808 42762 5817
rect 42706 5743 42762 5752
rect 42812 5692 42840 6258
rect 43076 6112 43128 6118
rect 43074 6080 43076 6089
rect 43128 6080 43130 6089
rect 43074 6015 43130 6024
rect 42892 5840 42944 5846
rect 42892 5782 42944 5788
rect 42720 5664 42840 5692
rect 42720 5302 42748 5664
rect 42904 5386 42932 5782
rect 42984 5568 43036 5574
rect 43076 5568 43128 5574
rect 42984 5510 43036 5516
rect 43074 5536 43076 5545
rect 43128 5536 43130 5545
rect 42812 5358 42932 5386
rect 42708 5296 42760 5302
rect 42708 5238 42760 5244
rect 42812 4622 42840 5358
rect 42892 5228 42944 5234
rect 42892 5170 42944 5176
rect 42904 4826 42932 5170
rect 42892 4820 42944 4826
rect 42892 4762 42944 4768
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 42996 4146 43024 5510
rect 43074 5471 43130 5480
rect 43168 5364 43220 5370
rect 43168 5306 43220 5312
rect 43076 5024 43128 5030
rect 43074 4992 43076 5001
rect 43128 4992 43130 5001
rect 43074 4927 43130 4936
rect 43180 4622 43208 5306
rect 43258 5264 43314 5273
rect 43258 5199 43260 5208
rect 43312 5199 43314 5208
rect 43260 5170 43312 5176
rect 43258 4720 43314 4729
rect 43364 4706 43392 6258
rect 43444 5840 43496 5846
rect 43442 5808 43444 5817
rect 43496 5808 43498 5817
rect 43548 5778 43576 6886
rect 43442 5743 43498 5752
rect 43536 5772 43588 5778
rect 43536 5714 43588 5720
rect 43444 5364 43496 5370
rect 43444 5306 43496 5312
rect 43456 5273 43484 5306
rect 43442 5264 43498 5273
rect 43442 5199 43498 5208
rect 43444 4752 43496 4758
rect 43314 4678 43392 4706
rect 43442 4720 43444 4729
rect 43496 4720 43498 4729
rect 43258 4655 43314 4664
rect 43442 4655 43498 4664
rect 43168 4616 43220 4622
rect 43168 4558 43220 4564
rect 43076 4480 43128 4486
rect 43074 4448 43076 4457
rect 43128 4448 43130 4457
rect 43074 4383 43130 4392
rect 43442 4176 43498 4185
rect 42616 4140 42668 4146
rect 42616 4082 42668 4088
rect 42984 4140 43036 4146
rect 43442 4111 43498 4120
rect 42984 4082 43036 4088
rect 42524 3528 42576 3534
rect 42524 3470 42576 3476
rect 42168 3182 42288 3210
rect 42168 1222 42196 3182
rect 42248 3052 42300 3058
rect 42248 2994 42300 3000
rect 42260 1494 42288 2994
rect 42248 1488 42300 1494
rect 42248 1430 42300 1436
rect 42156 1216 42208 1222
rect 42156 1158 42208 1164
rect 42064 400 42116 406
rect 42064 342 42116 348
rect 42536 134 42564 3470
rect 42628 542 42656 4082
rect 43456 4010 43484 4111
rect 43444 4004 43496 4010
rect 43444 3946 43496 3952
rect 43076 3936 43128 3942
rect 43074 3904 43076 3913
rect 43128 3904 43130 3913
rect 43074 3839 43130 3848
rect 43444 3664 43496 3670
rect 43442 3632 43444 3641
rect 43496 3632 43498 3641
rect 43442 3567 43498 3576
rect 43260 3528 43312 3534
rect 43258 3496 43260 3505
rect 43312 3496 43314 3505
rect 42708 3460 42760 3466
rect 43258 3431 43314 3440
rect 42708 3402 42760 3408
rect 42720 3346 42748 3402
rect 43076 3392 43128 3398
rect 43074 3360 43076 3369
rect 43260 3392 43312 3398
rect 43128 3360 43130 3369
rect 42720 3318 43024 3346
rect 42892 2916 42944 2922
rect 42892 2858 42944 2864
rect 42800 2576 42852 2582
rect 42800 2518 42852 2524
rect 42812 1737 42840 2518
rect 42904 2417 42932 2858
rect 42890 2408 42946 2417
rect 42890 2343 42946 2352
rect 42892 2304 42944 2310
rect 42892 2246 42944 2252
rect 42798 1728 42854 1737
rect 42798 1663 42854 1672
rect 42904 1465 42932 2246
rect 42890 1456 42946 1465
rect 42890 1391 42946 1400
rect 42996 1306 43024 3318
rect 43260 3334 43312 3340
rect 43074 3295 43130 3304
rect 43076 2848 43128 2854
rect 43074 2816 43076 2825
rect 43128 2816 43130 2825
rect 43074 2751 43130 2760
rect 43076 2304 43128 2310
rect 43074 2272 43076 2281
rect 43128 2272 43130 2281
rect 43074 2207 43130 2216
rect 42812 1278 43024 1306
rect 43272 1290 43300 3334
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 43456 3097 43484 3130
rect 43442 3088 43498 3097
rect 43442 3023 43498 3032
rect 43444 2576 43496 2582
rect 43442 2544 43444 2553
rect 43496 2544 43498 2553
rect 43442 2479 43498 2488
rect 43260 1284 43312 1290
rect 42812 800 42840 1278
rect 43260 1226 43312 1232
rect 42616 536 42668 542
rect 42616 478 42668 484
rect 42524 128 42576 134
rect 42524 70 42576 76
rect 42798 0 42854 800
<< via2 >>
rect 3422 9832 3478 9888
rect 3054 9560 3110 9616
rect 1398 9288 1454 9344
rect 2318 8744 2374 8800
rect 1674 8472 1730 8528
rect 1490 7928 1546 7984
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 2656 8730 2712 8732
rect 2736 8730 2792 8732
rect 2816 8730 2872 8732
rect 2896 8730 2952 8732
rect 2976 8730 3032 8732
rect 2656 8678 2658 8730
rect 2658 8678 2710 8730
rect 2710 8678 2712 8730
rect 2736 8678 2774 8730
rect 2774 8678 2786 8730
rect 2786 8678 2792 8730
rect 2816 8678 2838 8730
rect 2838 8678 2850 8730
rect 2850 8678 2872 8730
rect 2896 8678 2902 8730
rect 2902 8678 2914 8730
rect 2914 8678 2952 8730
rect 2976 8678 2978 8730
rect 2978 8678 3030 8730
rect 3030 8678 3032 8730
rect 2656 8676 2712 8678
rect 2736 8676 2792 8678
rect 2816 8676 2872 8678
rect 2896 8676 2952 8678
rect 2976 8676 3032 8678
rect 3330 9424 3386 9480
rect 3146 9016 3202 9072
rect 3054 8200 3110 8256
rect 3054 7928 3110 7984
rect 2410 7812 2466 7848
rect 2410 7792 2412 7812
rect 2412 7792 2464 7812
rect 2464 7792 2466 7812
rect 2656 7642 2712 7644
rect 2736 7642 2792 7644
rect 2816 7642 2872 7644
rect 2896 7642 2952 7644
rect 2976 7642 3032 7644
rect 2656 7590 2658 7642
rect 2658 7590 2710 7642
rect 2710 7590 2712 7642
rect 2736 7590 2774 7642
rect 2774 7590 2786 7642
rect 2786 7590 2792 7642
rect 2816 7590 2838 7642
rect 2838 7590 2850 7642
rect 2850 7590 2872 7642
rect 2896 7590 2902 7642
rect 2902 7590 2914 7642
rect 2914 7590 2952 7642
rect 2976 7590 2978 7642
rect 2978 7590 3030 7642
rect 3030 7590 3032 7642
rect 2656 7588 2712 7590
rect 2736 7588 2792 7590
rect 2816 7588 2872 7590
rect 2896 7588 2952 7590
rect 2976 7588 3032 7590
rect 3238 7520 3294 7576
rect 2318 7384 2374 7440
rect 1398 7112 1454 7168
rect 1398 6860 1454 6896
rect 1398 6840 1400 6860
rect 1400 6840 1452 6860
rect 1452 6840 1454 6860
rect 1490 6568 1546 6624
rect 1398 6024 1454 6080
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 2962 7384 3018 7440
rect 2318 6296 2374 6352
rect 3330 7248 3386 7304
rect 3422 6840 3478 6896
rect 2656 6554 2712 6556
rect 2736 6554 2792 6556
rect 2816 6554 2872 6556
rect 2896 6554 2952 6556
rect 2976 6554 3032 6556
rect 2656 6502 2658 6554
rect 2658 6502 2710 6554
rect 2710 6502 2712 6554
rect 2736 6502 2774 6554
rect 2774 6502 2786 6554
rect 2786 6502 2792 6554
rect 2816 6502 2838 6554
rect 2838 6502 2850 6554
rect 2850 6502 2872 6554
rect 2896 6502 2902 6554
rect 2902 6502 2914 6554
rect 2914 6502 2952 6554
rect 2976 6502 2978 6554
rect 2978 6502 3030 6554
rect 3030 6502 3032 6554
rect 2656 6500 2712 6502
rect 2736 6500 2792 6502
rect 2816 6500 2872 6502
rect 2896 6500 2952 6502
rect 2976 6500 3032 6502
rect 2502 6296 2558 6352
rect 3330 6432 3386 6488
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 1674 5752 1730 5808
rect 1490 4936 1546 4992
rect 1398 4392 1454 4448
rect 1490 3848 1546 3904
rect 3790 6432 3846 6488
rect 3422 6160 3478 6216
rect 3238 5616 3294 5672
rect 3606 6024 3662 6080
rect 4066 7384 4122 7440
rect 3974 6704 4030 6760
rect 3974 6024 4030 6080
rect 2502 5480 2558 5536
rect 2656 5466 2712 5468
rect 2736 5466 2792 5468
rect 2816 5466 2872 5468
rect 2896 5466 2952 5468
rect 2976 5466 3032 5468
rect 2656 5414 2658 5466
rect 2658 5414 2710 5466
rect 2710 5414 2712 5466
rect 2736 5414 2774 5466
rect 2774 5414 2786 5466
rect 2786 5414 2792 5466
rect 2816 5414 2838 5466
rect 2838 5414 2850 5466
rect 2850 5414 2872 5466
rect 2896 5414 2902 5466
rect 2902 5414 2914 5466
rect 2914 5414 2952 5466
rect 2976 5414 2978 5466
rect 2978 5414 3030 5466
rect 3030 5414 3032 5466
rect 2656 5412 2712 5414
rect 2736 5412 2792 5414
rect 2816 5412 2872 5414
rect 2896 5412 2952 5414
rect 2976 5412 3032 5414
rect 1766 5072 1822 5128
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 1858 4664 1914 4720
rect 2042 4548 2098 4584
rect 2042 4528 2044 4548
rect 2044 4528 2096 4548
rect 2096 4528 2098 4548
rect 3146 5480 3202 5536
rect 2226 4156 2228 4176
rect 2228 4156 2280 4176
rect 2280 4156 2282 4176
rect 2226 4120 2282 4156
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 2656 4378 2712 4380
rect 2736 4378 2792 4380
rect 2816 4378 2872 4380
rect 2896 4378 2952 4380
rect 2976 4378 3032 4380
rect 2656 4326 2658 4378
rect 2658 4326 2710 4378
rect 2710 4326 2712 4378
rect 2736 4326 2774 4378
rect 2774 4326 2786 4378
rect 2786 4326 2792 4378
rect 2816 4326 2838 4378
rect 2838 4326 2850 4378
rect 2850 4326 2872 4378
rect 2896 4326 2902 4378
rect 2902 4326 2914 4378
rect 2914 4326 2952 4378
rect 2976 4326 2978 4378
rect 2978 4326 3030 4378
rect 3030 4326 3032 4378
rect 2656 4324 2712 4326
rect 2736 4324 2792 4326
rect 2816 4324 2872 4326
rect 2896 4324 2952 4326
rect 2976 4324 3032 4326
rect 1582 3576 1638 3632
rect 2502 3576 2558 3632
rect 1398 2488 1454 2544
rect 1398 2216 1454 2272
rect 1858 3304 1914 3360
rect 2226 3168 2282 3224
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 1766 1944 1822 2000
rect 2656 3290 2712 3292
rect 2736 3290 2792 3292
rect 2816 3290 2872 3292
rect 2896 3290 2952 3292
rect 2976 3290 3032 3292
rect 2656 3238 2658 3290
rect 2658 3238 2710 3290
rect 2710 3238 2712 3290
rect 2736 3238 2774 3290
rect 2774 3238 2786 3290
rect 2786 3238 2792 3290
rect 2816 3238 2838 3290
rect 2838 3238 2850 3290
rect 2850 3238 2872 3290
rect 2896 3238 2902 3290
rect 2902 3238 2914 3290
rect 2914 3238 2952 3290
rect 2976 3238 2978 3290
rect 2978 3238 3030 3290
rect 3030 3238 3032 3290
rect 2656 3236 2712 3238
rect 2736 3236 2792 3238
rect 2816 3236 2872 3238
rect 2896 3236 2952 3238
rect 2976 3236 3032 3238
rect 2778 3068 2780 3088
rect 2780 3068 2832 3088
rect 2832 3068 2834 3088
rect 2778 3032 2834 3068
rect 2502 2916 2558 2952
rect 2502 2896 2504 2916
rect 2504 2896 2556 2916
rect 2556 2896 2558 2916
rect 3422 5208 3478 5264
rect 3698 5344 3754 5400
rect 3514 3032 3570 3088
rect 2410 1400 2466 1456
rect 2656 2202 2712 2204
rect 2736 2202 2792 2204
rect 2816 2202 2872 2204
rect 2896 2202 2952 2204
rect 2976 2202 3032 2204
rect 2656 2150 2658 2202
rect 2658 2150 2710 2202
rect 2710 2150 2712 2202
rect 2736 2150 2774 2202
rect 2774 2150 2786 2202
rect 2786 2150 2792 2202
rect 2816 2150 2838 2202
rect 2838 2150 2850 2202
rect 2850 2150 2872 2202
rect 2896 2150 2902 2202
rect 2902 2150 2914 2202
rect 2914 2150 2952 2202
rect 2976 2150 2978 2202
rect 2978 2150 3030 2202
rect 3030 2150 3032 2202
rect 2656 2148 2712 2150
rect 2736 2148 2792 2150
rect 2816 2148 2872 2150
rect 2896 2148 2952 2150
rect 2976 2148 3032 2150
rect 3330 1672 3386 1728
rect 4342 7656 4398 7712
rect 4158 5480 4214 5536
rect 3882 1128 3938 1184
rect 4618 5772 4674 5808
rect 4618 5752 4620 5772
rect 4620 5752 4672 5772
rect 4672 5752 4674 5772
rect 4986 8336 5042 8392
rect 4802 5616 4858 5672
rect 5078 8064 5134 8120
rect 5354 8336 5410 8392
rect 5446 7928 5502 7984
rect 5262 7692 5264 7712
rect 5264 7692 5316 7712
rect 5316 7692 5318 7712
rect 5262 7656 5318 7692
rect 5538 6860 5594 6896
rect 5814 7656 5870 7712
rect 5538 6840 5540 6860
rect 5540 6840 5592 6860
rect 5592 6840 5594 6860
rect 5354 6024 5410 6080
rect 5170 5752 5226 5808
rect 5262 5616 5318 5672
rect 4342 1264 4398 1320
rect 3974 856 4030 912
rect 5078 4428 5080 4448
rect 5080 4428 5132 4448
rect 5132 4428 5134 4448
rect 5078 4392 5134 4428
rect 5538 5652 5540 5672
rect 5540 5652 5592 5672
rect 5592 5652 5594 5672
rect 5538 5616 5594 5652
rect 5722 5072 5778 5128
rect 5814 3304 5870 3360
rect 5998 1400 6054 1456
rect 6182 7656 6238 7712
rect 6274 5208 6330 5264
rect 6182 4664 6238 4720
rect 6274 4392 6330 4448
rect 6182 2388 6184 2408
rect 6184 2388 6236 2408
rect 6236 2388 6238 2408
rect 6182 2352 6238 2388
rect 6734 6432 6790 6488
rect 7102 8608 7158 8664
rect 7010 8064 7066 8120
rect 6734 5772 6790 5808
rect 6734 5752 6736 5772
rect 6736 5752 6788 5772
rect 6788 5752 6790 5772
rect 6642 5344 6698 5400
rect 6826 3476 6828 3496
rect 6828 3476 6880 3496
rect 6880 3476 6882 3496
rect 6826 3440 6882 3476
rect 7378 7656 7434 7712
rect 7010 720 7066 776
rect 7654 8200 7710 8256
rect 8022 9016 8078 9072
rect 8390 8880 8446 8936
rect 7746 7692 7748 7712
rect 7748 7692 7800 7712
rect 7800 7692 7802 7712
rect 7746 7656 7802 7692
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 8656 8730 8712 8732
rect 8736 8730 8792 8732
rect 8816 8730 8872 8732
rect 8896 8730 8952 8732
rect 8976 8730 9032 8732
rect 8656 8678 8658 8730
rect 8658 8678 8710 8730
rect 8710 8678 8712 8730
rect 8736 8678 8774 8730
rect 8774 8678 8786 8730
rect 8786 8678 8792 8730
rect 8816 8678 8838 8730
rect 8838 8678 8850 8730
rect 8850 8678 8872 8730
rect 8896 8678 8902 8730
rect 8902 8678 8914 8730
rect 8914 8678 8952 8730
rect 8976 8678 8978 8730
rect 8978 8678 9030 8730
rect 9030 8678 9032 8730
rect 8656 8676 8712 8678
rect 8736 8676 8792 8678
rect 8816 8676 8872 8678
rect 8896 8676 8952 8678
rect 8976 8676 9032 8678
rect 8666 8064 8722 8120
rect 8390 7792 8446 7848
rect 9310 9560 9366 9616
rect 9402 9152 9458 9208
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 8390 6976 8446 7032
rect 7930 6432 7986 6488
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 8022 5480 8078 5536
rect 8298 5344 8354 5400
rect 7654 5208 7710 5264
rect 7930 5208 7986 5264
rect 7562 5072 7618 5128
rect 7746 5072 7802 5128
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 8390 4120 8446 4176
rect 7838 3984 7894 4040
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 8298 3304 8354 3360
rect 7930 2896 7986 2952
rect 7654 992 7710 1048
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 8666 7792 8722 7848
rect 8656 7642 8712 7644
rect 8736 7642 8792 7644
rect 8816 7642 8872 7644
rect 8896 7642 8952 7644
rect 8976 7642 9032 7644
rect 8656 7590 8658 7642
rect 8658 7590 8710 7642
rect 8710 7590 8712 7642
rect 8736 7590 8774 7642
rect 8774 7590 8786 7642
rect 8786 7590 8792 7642
rect 8816 7590 8838 7642
rect 8838 7590 8850 7642
rect 8850 7590 8872 7642
rect 8896 7590 8902 7642
rect 8902 7590 8914 7642
rect 8914 7590 8952 7642
rect 8976 7590 8978 7642
rect 8978 7590 9030 7642
rect 9030 7590 9032 7642
rect 8656 7588 8712 7590
rect 8736 7588 8792 7590
rect 8816 7588 8872 7590
rect 8896 7588 8952 7590
rect 8976 7588 9032 7590
rect 8656 6554 8712 6556
rect 8736 6554 8792 6556
rect 8816 6554 8872 6556
rect 8896 6554 8952 6556
rect 8976 6554 9032 6556
rect 8656 6502 8658 6554
rect 8658 6502 8710 6554
rect 8710 6502 8712 6554
rect 8736 6502 8774 6554
rect 8774 6502 8786 6554
rect 8786 6502 8792 6554
rect 8816 6502 8838 6554
rect 8838 6502 8850 6554
rect 8850 6502 8872 6554
rect 8896 6502 8902 6554
rect 8902 6502 8914 6554
rect 8914 6502 8952 6554
rect 8976 6502 8978 6554
rect 8978 6502 9030 6554
rect 9030 6502 9032 6554
rect 8656 6500 8712 6502
rect 8736 6500 8792 6502
rect 8816 6500 8872 6502
rect 8896 6500 8952 6502
rect 8976 6500 9032 6502
rect 9310 6432 9366 6488
rect 8666 6024 8722 6080
rect 8656 5466 8712 5468
rect 8736 5466 8792 5468
rect 8816 5466 8872 5468
rect 8896 5466 8952 5468
rect 8976 5466 9032 5468
rect 8656 5414 8658 5466
rect 8658 5414 8710 5466
rect 8710 5414 8712 5466
rect 8736 5414 8774 5466
rect 8774 5414 8786 5466
rect 8786 5414 8792 5466
rect 8816 5414 8838 5466
rect 8838 5414 8850 5466
rect 8850 5414 8872 5466
rect 8896 5414 8902 5466
rect 8902 5414 8914 5466
rect 8914 5414 8952 5466
rect 8976 5414 8978 5466
rect 8978 5414 9030 5466
rect 9030 5414 9032 5466
rect 8656 5412 8712 5414
rect 8736 5412 8792 5414
rect 8816 5412 8872 5414
rect 8896 5412 8952 5414
rect 8976 5412 9032 5414
rect 9034 4800 9090 4856
rect 8656 4378 8712 4380
rect 8736 4378 8792 4380
rect 8816 4378 8872 4380
rect 8896 4378 8952 4380
rect 8976 4378 9032 4380
rect 8656 4326 8658 4378
rect 8658 4326 8710 4378
rect 8710 4326 8712 4378
rect 8736 4326 8774 4378
rect 8774 4326 8786 4378
rect 8786 4326 8792 4378
rect 8816 4326 8838 4378
rect 8838 4326 8850 4378
rect 8850 4326 8872 4378
rect 8896 4326 8902 4378
rect 8902 4326 8914 4378
rect 8914 4326 8952 4378
rect 8976 4326 8978 4378
rect 8978 4326 9030 4378
rect 9030 4326 9032 4378
rect 8656 4324 8712 4326
rect 8736 4324 8792 4326
rect 8816 4324 8872 4326
rect 8896 4324 8952 4326
rect 8976 4324 9032 4326
rect 8942 3712 8998 3768
rect 9126 3576 9182 3632
rect 9126 3304 9182 3360
rect 8656 3290 8712 3292
rect 8736 3290 8792 3292
rect 8816 3290 8872 3292
rect 8896 3290 8952 3292
rect 8976 3290 9032 3292
rect 8656 3238 8658 3290
rect 8658 3238 8710 3290
rect 8710 3238 8712 3290
rect 8736 3238 8774 3290
rect 8774 3238 8786 3290
rect 8786 3238 8792 3290
rect 8816 3238 8838 3290
rect 8838 3238 8850 3290
rect 8850 3238 8872 3290
rect 8896 3238 8902 3290
rect 8902 3238 8914 3290
rect 8914 3238 8952 3290
rect 8976 3238 8978 3290
rect 8978 3238 9030 3290
rect 9030 3238 9032 3290
rect 8656 3236 8712 3238
rect 8736 3236 8792 3238
rect 8816 3236 8872 3238
rect 8896 3236 8952 3238
rect 8976 3236 9032 3238
rect 9126 3168 9182 3224
rect 8666 2932 8668 2952
rect 8668 2932 8720 2952
rect 8720 2932 8722 2952
rect 8666 2896 8722 2932
rect 8942 2760 8998 2816
rect 8656 2202 8712 2204
rect 8736 2202 8792 2204
rect 8816 2202 8872 2204
rect 8896 2202 8952 2204
rect 8976 2202 9032 2204
rect 8656 2150 8658 2202
rect 8658 2150 8710 2202
rect 8710 2150 8712 2202
rect 8736 2150 8774 2202
rect 8774 2150 8786 2202
rect 8786 2150 8792 2202
rect 8816 2150 8838 2202
rect 8838 2150 8850 2202
rect 8850 2150 8872 2202
rect 8896 2150 8902 2202
rect 8902 2150 8914 2202
rect 8914 2150 8952 2202
rect 8976 2150 8978 2202
rect 8978 2150 9030 2202
rect 9030 2150 9032 2202
rect 8656 2148 8712 2150
rect 8736 2148 8792 2150
rect 8816 2148 8872 2150
rect 8896 2148 8952 2150
rect 8976 2148 9032 2150
rect 9402 4256 9458 4312
rect 10046 9832 10102 9888
rect 10322 9288 10378 9344
rect 10414 8492 10470 8528
rect 10414 8472 10416 8492
rect 10416 8472 10468 8492
rect 10468 8472 10470 8492
rect 10506 8336 10562 8392
rect 10046 6568 10102 6624
rect 9770 5888 9826 5944
rect 9862 5752 9918 5808
rect 9770 5344 9826 5400
rect 10046 5888 10102 5944
rect 10230 7520 10286 7576
rect 10414 6840 10470 6896
rect 9678 5072 9734 5128
rect 9954 4800 10010 4856
rect 9954 4392 10010 4448
rect 9770 3848 9826 3904
rect 9862 3576 9918 3632
rect 9586 2216 9642 2272
rect 9494 1944 9550 2000
rect 9218 1536 9274 1592
rect 7470 584 7526 640
rect 9862 3032 9918 3088
rect 10506 5616 10562 5672
rect 10322 5092 10378 5128
rect 10322 5072 10324 5092
rect 10324 5072 10376 5092
rect 10376 5072 10378 5092
rect 10414 3712 10470 3768
rect 10874 8372 10876 8392
rect 10876 8372 10928 8392
rect 10928 8372 10930 8392
rect 10874 8336 10930 8372
rect 10874 6840 10930 6896
rect 10874 6024 10930 6080
rect 10782 5772 10838 5808
rect 10782 5752 10784 5772
rect 10784 5752 10836 5772
rect 10836 5752 10838 5772
rect 10690 5208 10746 5264
rect 10690 4664 10746 4720
rect 11702 9968 11758 10024
rect 11426 7520 11482 7576
rect 11334 6568 11390 6624
rect 11242 6432 11298 6488
rect 11242 6024 11298 6080
rect 11058 5072 11114 5128
rect 10874 3848 10930 3904
rect 11610 5344 11666 5400
rect 11610 3712 11666 3768
rect 10690 2896 10746 2952
rect 11334 2080 11390 2136
rect 11150 1808 11206 1864
rect 11794 7384 11850 7440
rect 12254 8336 12310 8392
rect 12070 7812 12126 7848
rect 12070 7792 12072 7812
rect 12072 7792 12124 7812
rect 12124 7792 12126 7812
rect 12254 7248 12310 7304
rect 12070 5480 12126 5536
rect 12070 4664 12126 4720
rect 12530 6568 12586 6624
rect 12806 8200 12862 8256
rect 12346 4936 12402 4992
rect 12254 3168 12310 3224
rect 12530 5208 12586 5264
rect 12438 4256 12494 4312
rect 13266 7248 13322 7304
rect 13082 6976 13138 7032
rect 12990 5616 13046 5672
rect 12622 3440 12678 3496
rect 13082 5072 13138 5128
rect 13082 4392 13138 4448
rect 13082 3032 13138 3088
rect 12990 2488 13046 2544
rect 12714 2080 12770 2136
rect 13450 7928 13506 7984
rect 13450 6024 13506 6080
rect 13358 5344 13414 5400
rect 13266 4004 13322 4040
rect 13266 3984 13268 4004
rect 13268 3984 13320 4004
rect 13320 3984 13322 4004
rect 13358 3848 13414 3904
rect 13266 3712 13322 3768
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 14156 8186 14212 8188
rect 14236 8186 14292 8188
rect 13916 8134 13918 8186
rect 13918 8134 13970 8186
rect 13970 8134 13972 8186
rect 13996 8134 14034 8186
rect 14034 8134 14046 8186
rect 14046 8134 14052 8186
rect 14076 8134 14098 8186
rect 14098 8134 14110 8186
rect 14110 8134 14132 8186
rect 14156 8134 14162 8186
rect 14162 8134 14174 8186
rect 14174 8134 14212 8186
rect 14236 8134 14238 8186
rect 14238 8134 14290 8186
rect 14290 8134 14292 8186
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 14156 8132 14212 8134
rect 14236 8132 14292 8134
rect 13910 7520 13966 7576
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 14156 7098 14212 7100
rect 14236 7098 14292 7100
rect 13916 7046 13918 7098
rect 13918 7046 13970 7098
rect 13970 7046 13972 7098
rect 13996 7046 14034 7098
rect 14034 7046 14046 7098
rect 14046 7046 14052 7098
rect 14076 7046 14098 7098
rect 14098 7046 14110 7098
rect 14110 7046 14132 7098
rect 14156 7046 14162 7098
rect 14162 7046 14174 7098
rect 14174 7046 14212 7098
rect 14236 7046 14238 7098
rect 14238 7046 14290 7098
rect 14290 7046 14292 7098
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 14156 7044 14212 7046
rect 14236 7044 14292 7046
rect 14186 6860 14242 6896
rect 14186 6840 14188 6860
rect 14188 6840 14240 6860
rect 14240 6840 14242 6860
rect 13634 4800 13690 4856
rect 13634 3848 13690 3904
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 14156 6010 14212 6012
rect 14236 6010 14292 6012
rect 13916 5958 13918 6010
rect 13918 5958 13970 6010
rect 13970 5958 13972 6010
rect 13996 5958 14034 6010
rect 14034 5958 14046 6010
rect 14046 5958 14052 6010
rect 14076 5958 14098 6010
rect 14098 5958 14110 6010
rect 14110 5958 14132 6010
rect 14156 5958 14162 6010
rect 14162 5958 14174 6010
rect 14174 5958 14212 6010
rect 14236 5958 14238 6010
rect 14238 5958 14290 6010
rect 14290 5958 14292 6010
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 14156 5956 14212 5958
rect 14236 5956 14292 5958
rect 14656 8730 14712 8732
rect 14736 8730 14792 8732
rect 14816 8730 14872 8732
rect 14896 8730 14952 8732
rect 14976 8730 15032 8732
rect 14656 8678 14658 8730
rect 14658 8678 14710 8730
rect 14710 8678 14712 8730
rect 14736 8678 14774 8730
rect 14774 8678 14786 8730
rect 14786 8678 14792 8730
rect 14816 8678 14838 8730
rect 14838 8678 14850 8730
rect 14850 8678 14872 8730
rect 14896 8678 14902 8730
rect 14902 8678 14914 8730
rect 14914 8678 14952 8730
rect 14976 8678 14978 8730
rect 14978 8678 15030 8730
rect 15030 8678 15032 8730
rect 14656 8676 14712 8678
rect 14736 8676 14792 8678
rect 14816 8676 14872 8678
rect 14896 8676 14952 8678
rect 14976 8676 15032 8678
rect 14830 7828 14832 7848
rect 14832 7828 14884 7848
rect 14884 7828 14886 7848
rect 14830 7792 14886 7828
rect 14656 7642 14712 7644
rect 14736 7642 14792 7644
rect 14816 7642 14872 7644
rect 14896 7642 14952 7644
rect 14976 7642 15032 7644
rect 14656 7590 14658 7642
rect 14658 7590 14710 7642
rect 14710 7590 14712 7642
rect 14736 7590 14774 7642
rect 14774 7590 14786 7642
rect 14786 7590 14792 7642
rect 14816 7590 14838 7642
rect 14838 7590 14850 7642
rect 14850 7590 14872 7642
rect 14896 7590 14902 7642
rect 14902 7590 14914 7642
rect 14914 7590 14952 7642
rect 14976 7590 14978 7642
rect 14978 7590 15030 7642
rect 15030 7590 15032 7642
rect 14656 7588 14712 7590
rect 14736 7588 14792 7590
rect 14816 7588 14872 7590
rect 14896 7588 14952 7590
rect 14976 7588 15032 7590
rect 14462 6840 14518 6896
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 14156 4922 14212 4924
rect 14236 4922 14292 4924
rect 13916 4870 13918 4922
rect 13918 4870 13970 4922
rect 13970 4870 13972 4922
rect 13996 4870 14034 4922
rect 14034 4870 14046 4922
rect 14046 4870 14052 4922
rect 14076 4870 14098 4922
rect 14098 4870 14110 4922
rect 14110 4870 14132 4922
rect 14156 4870 14162 4922
rect 14162 4870 14174 4922
rect 14174 4870 14212 4922
rect 14236 4870 14238 4922
rect 14238 4870 14290 4922
rect 14290 4870 14292 4922
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 14156 4868 14212 4870
rect 14236 4868 14292 4870
rect 14656 6554 14712 6556
rect 14736 6554 14792 6556
rect 14816 6554 14872 6556
rect 14896 6554 14952 6556
rect 14976 6554 15032 6556
rect 14656 6502 14658 6554
rect 14658 6502 14710 6554
rect 14710 6502 14712 6554
rect 14736 6502 14774 6554
rect 14774 6502 14786 6554
rect 14786 6502 14792 6554
rect 14816 6502 14838 6554
rect 14838 6502 14850 6554
rect 14850 6502 14872 6554
rect 14896 6502 14902 6554
rect 14902 6502 14914 6554
rect 14914 6502 14952 6554
rect 14976 6502 14978 6554
rect 14978 6502 15030 6554
rect 15030 6502 15032 6554
rect 14656 6500 14712 6502
rect 14736 6500 14792 6502
rect 14816 6500 14872 6502
rect 14896 6500 14952 6502
rect 14976 6500 15032 6502
rect 14646 6024 14702 6080
rect 14554 5888 14610 5944
rect 14462 5344 14518 5400
rect 14094 4564 14096 4584
rect 14096 4564 14148 4584
rect 14148 4564 14150 4584
rect 14094 4528 14150 4564
rect 14278 4528 14334 4584
rect 14002 4392 14058 4448
rect 13910 4120 13966 4176
rect 14278 4256 14334 4312
rect 14656 5466 14712 5468
rect 14736 5466 14792 5468
rect 14816 5466 14872 5468
rect 14896 5466 14952 5468
rect 14976 5466 15032 5468
rect 14656 5414 14658 5466
rect 14658 5414 14710 5466
rect 14710 5414 14712 5466
rect 14736 5414 14774 5466
rect 14774 5414 14786 5466
rect 14786 5414 14792 5466
rect 14816 5414 14838 5466
rect 14838 5414 14850 5466
rect 14850 5414 14872 5466
rect 14896 5414 14902 5466
rect 14902 5414 14914 5466
rect 14914 5414 14952 5466
rect 14976 5414 14978 5466
rect 14978 5414 15030 5466
rect 15030 5414 15032 5466
rect 14656 5412 14712 5414
rect 14736 5412 14792 5414
rect 14816 5412 14872 5414
rect 14896 5412 14952 5414
rect 14976 5412 15032 5414
rect 14830 5208 14886 5264
rect 14830 4936 14886 4992
rect 15382 7248 15438 7304
rect 15198 6024 15254 6080
rect 14656 4378 14712 4380
rect 14736 4378 14792 4380
rect 14816 4378 14872 4380
rect 14896 4378 14952 4380
rect 14976 4378 15032 4380
rect 14656 4326 14658 4378
rect 14658 4326 14710 4378
rect 14710 4326 14712 4378
rect 14736 4326 14774 4378
rect 14774 4326 14786 4378
rect 14786 4326 14792 4378
rect 14816 4326 14838 4378
rect 14838 4326 14850 4378
rect 14850 4326 14872 4378
rect 14896 4326 14902 4378
rect 14902 4326 14914 4378
rect 14914 4326 14952 4378
rect 14976 4326 14978 4378
rect 14978 4326 15030 4378
rect 15030 4326 15032 4378
rect 14656 4324 14712 4326
rect 14736 4324 14792 4326
rect 14816 4324 14872 4326
rect 14896 4324 14952 4326
rect 14976 4324 15032 4326
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 14156 3834 14212 3836
rect 14236 3834 14292 3836
rect 13916 3782 13918 3834
rect 13918 3782 13970 3834
rect 13970 3782 13972 3834
rect 13996 3782 14034 3834
rect 14034 3782 14046 3834
rect 14046 3782 14052 3834
rect 14076 3782 14098 3834
rect 14098 3782 14110 3834
rect 14110 3782 14132 3834
rect 14156 3782 14162 3834
rect 14162 3782 14174 3834
rect 14174 3782 14212 3834
rect 14236 3782 14238 3834
rect 14238 3782 14290 3834
rect 14290 3782 14292 3834
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 14156 3780 14212 3782
rect 14236 3780 14292 3782
rect 13358 3440 13414 3496
rect 13266 3032 13322 3088
rect 12990 1672 13046 1728
rect 13818 3304 13874 3360
rect 14186 3168 14242 3224
rect 14646 3984 14702 4040
rect 14656 3290 14712 3292
rect 14736 3290 14792 3292
rect 14816 3290 14872 3292
rect 14896 3290 14952 3292
rect 14976 3290 15032 3292
rect 14656 3238 14658 3290
rect 14658 3238 14710 3290
rect 14710 3238 14712 3290
rect 14736 3238 14774 3290
rect 14774 3238 14786 3290
rect 14786 3238 14792 3290
rect 14816 3238 14838 3290
rect 14838 3238 14850 3290
rect 14850 3238 14872 3290
rect 14896 3238 14902 3290
rect 14902 3238 14914 3290
rect 14914 3238 14952 3290
rect 14976 3238 14978 3290
rect 14978 3238 15030 3290
rect 15030 3238 15032 3290
rect 14656 3236 14712 3238
rect 14736 3236 14792 3238
rect 14816 3236 14872 3238
rect 14896 3236 14952 3238
rect 14976 3236 15032 3238
rect 14278 3032 14334 3088
rect 14462 3068 14464 3088
rect 14464 3068 14516 3088
rect 14516 3068 14518 3088
rect 14462 3032 14518 3068
rect 14370 2760 14426 2816
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 14156 2746 14212 2748
rect 14236 2746 14292 2748
rect 13916 2694 13918 2746
rect 13918 2694 13970 2746
rect 13970 2694 13972 2746
rect 13996 2694 14034 2746
rect 14034 2694 14046 2746
rect 14046 2694 14052 2746
rect 14076 2694 14098 2746
rect 14098 2694 14110 2746
rect 14110 2694 14132 2746
rect 14156 2694 14162 2746
rect 14162 2694 14174 2746
rect 14174 2694 14212 2746
rect 14236 2694 14238 2746
rect 14238 2694 14290 2746
rect 14290 2694 14292 2746
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 14156 2692 14212 2694
rect 14236 2692 14292 2694
rect 14370 2624 14426 2680
rect 14186 2352 14242 2408
rect 14370 2372 14426 2408
rect 14370 2352 14372 2372
rect 14372 2352 14424 2372
rect 14424 2352 14426 2372
rect 14370 2216 14426 2272
rect 14656 2202 14712 2204
rect 14736 2202 14792 2204
rect 14816 2202 14872 2204
rect 14896 2202 14952 2204
rect 14976 2202 15032 2204
rect 14656 2150 14658 2202
rect 14658 2150 14710 2202
rect 14710 2150 14712 2202
rect 14736 2150 14774 2202
rect 14774 2150 14786 2202
rect 14786 2150 14792 2202
rect 14816 2150 14838 2202
rect 14838 2150 14850 2202
rect 14850 2150 14872 2202
rect 14896 2150 14902 2202
rect 14902 2150 14914 2202
rect 14914 2150 14952 2202
rect 14976 2150 14978 2202
rect 14978 2150 15030 2202
rect 15030 2150 15032 2202
rect 14656 2148 14712 2150
rect 14736 2148 14792 2150
rect 14816 2148 14872 2150
rect 14896 2148 14952 2150
rect 14976 2148 15032 2150
rect 14370 1264 14426 1320
rect 10782 448 10838 504
rect 16118 8336 16174 8392
rect 15566 5480 15622 5536
rect 15750 5480 15806 5536
rect 15566 5208 15622 5264
rect 15382 4800 15438 4856
rect 16578 7792 16634 7848
rect 16210 6840 16266 6896
rect 15934 5344 15990 5400
rect 16302 4256 16358 4312
rect 16762 7248 16818 7304
rect 17130 9868 17132 9888
rect 17132 9868 17184 9888
rect 17184 9868 17186 9888
rect 17130 9832 17186 9868
rect 17038 7656 17094 7712
rect 16946 7404 17002 7440
rect 16946 7384 16948 7404
rect 16948 7384 17000 7404
rect 17000 7384 17002 7404
rect 17958 9016 18014 9072
rect 18050 8064 18106 8120
rect 17866 7792 17922 7848
rect 17130 6296 17186 6352
rect 17038 5888 17094 5944
rect 16854 4392 16910 4448
rect 16854 3188 16910 3224
rect 16854 3168 16856 3188
rect 16856 3168 16908 3188
rect 16908 3168 16910 3188
rect 16302 2624 16358 2680
rect 17682 6568 17738 6624
rect 17590 6316 17646 6352
rect 17590 6296 17592 6316
rect 17592 6296 17644 6316
rect 17644 6296 17646 6316
rect 17498 6160 17554 6216
rect 17314 5888 17370 5944
rect 17130 5208 17186 5264
rect 17682 5888 17738 5944
rect 17314 3848 17370 3904
rect 17222 3188 17278 3224
rect 17222 3168 17224 3188
rect 17224 3168 17276 3188
rect 17276 3168 17278 3188
rect 17498 4820 17554 4856
rect 17498 4800 17500 4820
rect 17500 4800 17552 4820
rect 17552 4800 17554 4820
rect 18326 7656 18382 7712
rect 17774 4528 17830 4584
rect 17774 4256 17830 4312
rect 19154 10240 19210 10296
rect 18878 7248 18934 7304
rect 19062 6976 19118 7032
rect 19798 8744 19854 8800
rect 19246 6840 19302 6896
rect 19522 6840 19578 6896
rect 18694 6160 18750 6216
rect 18878 6160 18934 6216
rect 18786 6024 18842 6080
rect 18970 6024 19026 6080
rect 18142 5480 18198 5536
rect 18510 5480 18566 5536
rect 18694 5480 18750 5536
rect 18326 4820 18382 4856
rect 18326 4800 18328 4820
rect 18328 4800 18380 4820
rect 18380 4800 18382 4820
rect 19522 6432 19578 6488
rect 19916 8186 19972 8188
rect 19996 8186 20052 8188
rect 20076 8186 20132 8188
rect 20156 8186 20212 8188
rect 20236 8186 20292 8188
rect 19916 8134 19918 8186
rect 19918 8134 19970 8186
rect 19970 8134 19972 8186
rect 19996 8134 20034 8186
rect 20034 8134 20046 8186
rect 20046 8134 20052 8186
rect 20076 8134 20098 8186
rect 20098 8134 20110 8186
rect 20110 8134 20132 8186
rect 20156 8134 20162 8186
rect 20162 8134 20174 8186
rect 20174 8134 20212 8186
rect 20236 8134 20238 8186
rect 20238 8134 20290 8186
rect 20290 8134 20292 8186
rect 19916 8132 19972 8134
rect 19996 8132 20052 8134
rect 20076 8132 20132 8134
rect 20156 8132 20212 8134
rect 20236 8132 20292 8134
rect 19706 8064 19762 8120
rect 19916 7098 19972 7100
rect 19996 7098 20052 7100
rect 20076 7098 20132 7100
rect 20156 7098 20212 7100
rect 20236 7098 20292 7100
rect 19916 7046 19918 7098
rect 19918 7046 19970 7098
rect 19970 7046 19972 7098
rect 19996 7046 20034 7098
rect 20034 7046 20046 7098
rect 20046 7046 20052 7098
rect 20076 7046 20098 7098
rect 20098 7046 20110 7098
rect 20110 7046 20132 7098
rect 20156 7046 20162 7098
rect 20162 7046 20174 7098
rect 20174 7046 20212 7098
rect 20236 7046 20238 7098
rect 20238 7046 20290 7098
rect 20290 7046 20292 7098
rect 19916 7044 19972 7046
rect 19996 7044 20052 7046
rect 20076 7044 20132 7046
rect 20156 7044 20212 7046
rect 20236 7044 20292 7046
rect 21546 10240 21602 10296
rect 21546 9832 21602 9888
rect 20442 8608 20498 8664
rect 20442 8200 20498 8256
rect 20656 8730 20712 8732
rect 20736 8730 20792 8732
rect 20816 8730 20872 8732
rect 20896 8730 20952 8732
rect 20976 8730 21032 8732
rect 20656 8678 20658 8730
rect 20658 8678 20710 8730
rect 20710 8678 20712 8730
rect 20736 8678 20774 8730
rect 20774 8678 20786 8730
rect 20786 8678 20792 8730
rect 20816 8678 20838 8730
rect 20838 8678 20850 8730
rect 20850 8678 20872 8730
rect 20896 8678 20902 8730
rect 20902 8678 20914 8730
rect 20914 8678 20952 8730
rect 20976 8678 20978 8730
rect 20978 8678 21030 8730
rect 21030 8678 21032 8730
rect 20656 8676 20712 8678
rect 20736 8676 20792 8678
rect 20816 8676 20872 8678
rect 20896 8676 20952 8678
rect 20976 8676 21032 8678
rect 20718 8372 20720 8392
rect 20720 8372 20772 8392
rect 20772 8372 20774 8392
rect 20718 8336 20774 8372
rect 20656 7642 20712 7644
rect 20736 7642 20792 7644
rect 20816 7642 20872 7644
rect 20896 7642 20952 7644
rect 20976 7642 21032 7644
rect 20656 7590 20658 7642
rect 20658 7590 20710 7642
rect 20710 7590 20712 7642
rect 20736 7590 20774 7642
rect 20774 7590 20786 7642
rect 20786 7590 20792 7642
rect 20816 7590 20838 7642
rect 20838 7590 20850 7642
rect 20850 7590 20872 7642
rect 20896 7590 20902 7642
rect 20902 7590 20914 7642
rect 20914 7590 20952 7642
rect 20976 7590 20978 7642
rect 20978 7590 21030 7642
rect 21030 7590 21032 7642
rect 20656 7588 20712 7590
rect 20736 7588 20792 7590
rect 20816 7588 20872 7590
rect 20896 7588 20952 7590
rect 20976 7588 21032 7590
rect 20626 7112 20682 7168
rect 19706 6024 19762 6080
rect 20656 6554 20712 6556
rect 20736 6554 20792 6556
rect 20816 6554 20872 6556
rect 20896 6554 20952 6556
rect 20976 6554 21032 6556
rect 20656 6502 20658 6554
rect 20658 6502 20710 6554
rect 20710 6502 20712 6554
rect 20736 6502 20774 6554
rect 20774 6502 20786 6554
rect 20786 6502 20792 6554
rect 20816 6502 20838 6554
rect 20838 6502 20850 6554
rect 20850 6502 20872 6554
rect 20896 6502 20902 6554
rect 20902 6502 20914 6554
rect 20914 6502 20952 6554
rect 20976 6502 20978 6554
rect 20978 6502 21030 6554
rect 21030 6502 21032 6554
rect 20656 6500 20712 6502
rect 20736 6500 20792 6502
rect 20816 6500 20872 6502
rect 20896 6500 20952 6502
rect 20976 6500 21032 6502
rect 19614 5908 19670 5944
rect 19614 5888 19616 5908
rect 19616 5888 19668 5908
rect 19668 5888 19670 5908
rect 19916 6010 19972 6012
rect 19996 6010 20052 6012
rect 20076 6010 20132 6012
rect 20156 6010 20212 6012
rect 20236 6010 20292 6012
rect 19916 5958 19918 6010
rect 19918 5958 19970 6010
rect 19970 5958 19972 6010
rect 19996 5958 20034 6010
rect 20034 5958 20046 6010
rect 20046 5958 20052 6010
rect 20076 5958 20098 6010
rect 20098 5958 20110 6010
rect 20110 5958 20132 6010
rect 20156 5958 20162 6010
rect 20162 5958 20174 6010
rect 20174 5958 20212 6010
rect 20236 5958 20238 6010
rect 20238 5958 20290 6010
rect 20290 5958 20292 6010
rect 19916 5956 19972 5958
rect 19996 5956 20052 5958
rect 20076 5956 20132 5958
rect 20156 5956 20212 5958
rect 20236 5956 20292 5958
rect 19614 5652 19616 5672
rect 19616 5652 19668 5672
rect 19668 5652 19670 5672
rect 19614 5616 19670 5652
rect 19338 5344 19394 5400
rect 18510 4800 18566 4856
rect 17866 2760 17922 2816
rect 18234 4528 18290 4584
rect 18142 3712 18198 3768
rect 18602 4392 18658 4448
rect 19798 5344 19854 5400
rect 20902 5908 20958 5944
rect 20902 5888 20904 5908
rect 20904 5888 20956 5908
rect 20956 5888 20958 5908
rect 19430 4800 19486 4856
rect 18970 4392 19026 4448
rect 18878 4120 18934 4176
rect 19338 4256 19394 4312
rect 18418 2932 18420 2952
rect 18420 2932 18472 2952
rect 18472 2932 18474 2952
rect 18418 2896 18474 2932
rect 18786 2644 18842 2680
rect 18786 2624 18788 2644
rect 18788 2624 18840 2644
rect 18840 2624 18842 2644
rect 18234 1808 18290 1864
rect 19430 3848 19486 3904
rect 19062 3576 19118 3632
rect 19154 3168 19210 3224
rect 19706 4936 19762 4992
rect 19916 4922 19972 4924
rect 19996 4922 20052 4924
rect 20076 4922 20132 4924
rect 20156 4922 20212 4924
rect 20236 4922 20292 4924
rect 19916 4870 19918 4922
rect 19918 4870 19970 4922
rect 19970 4870 19972 4922
rect 19996 4870 20034 4922
rect 20034 4870 20046 4922
rect 20046 4870 20052 4922
rect 20076 4870 20098 4922
rect 20098 4870 20110 4922
rect 20110 4870 20132 4922
rect 20156 4870 20162 4922
rect 20162 4870 20174 4922
rect 20174 4870 20212 4922
rect 20236 4870 20238 4922
rect 20238 4870 20290 4922
rect 20290 4870 20292 4922
rect 19916 4868 19972 4870
rect 19996 4868 20052 4870
rect 20076 4868 20132 4870
rect 20156 4868 20212 4870
rect 20236 4868 20292 4870
rect 20656 5466 20712 5468
rect 20736 5466 20792 5468
rect 20816 5466 20872 5468
rect 20896 5466 20952 5468
rect 20976 5466 21032 5468
rect 20656 5414 20658 5466
rect 20658 5414 20710 5466
rect 20710 5414 20712 5466
rect 20736 5414 20774 5466
rect 20774 5414 20786 5466
rect 20786 5414 20792 5466
rect 20816 5414 20838 5466
rect 20838 5414 20850 5466
rect 20850 5414 20872 5466
rect 20896 5414 20902 5466
rect 20902 5414 20914 5466
rect 20914 5414 20952 5466
rect 20976 5414 20978 5466
rect 20978 5414 21030 5466
rect 21030 5414 21032 5466
rect 20656 5412 20712 5414
rect 20736 5412 20792 5414
rect 20816 5412 20872 5414
rect 20896 5412 20952 5414
rect 20976 5412 21032 5414
rect 20626 5072 20682 5128
rect 20626 4936 20682 4992
rect 19890 4120 19946 4176
rect 20656 4378 20712 4380
rect 20736 4378 20792 4380
rect 20816 4378 20872 4380
rect 20896 4378 20952 4380
rect 20976 4378 21032 4380
rect 20656 4326 20658 4378
rect 20658 4326 20710 4378
rect 20710 4326 20712 4378
rect 20736 4326 20774 4378
rect 20774 4326 20786 4378
rect 20786 4326 20792 4378
rect 20816 4326 20838 4378
rect 20838 4326 20850 4378
rect 20850 4326 20872 4378
rect 20896 4326 20902 4378
rect 20902 4326 20914 4378
rect 20914 4326 20952 4378
rect 20976 4326 20978 4378
rect 20978 4326 21030 4378
rect 21030 4326 21032 4378
rect 20656 4324 20712 4326
rect 20736 4324 20792 4326
rect 20816 4324 20872 4326
rect 20896 4324 20952 4326
rect 20976 4324 21032 4326
rect 21178 4256 21234 4312
rect 20534 3848 20590 3904
rect 19916 3834 19972 3836
rect 19996 3834 20052 3836
rect 20076 3834 20132 3836
rect 20156 3834 20212 3836
rect 20236 3834 20292 3836
rect 19916 3782 19918 3834
rect 19918 3782 19970 3834
rect 19970 3782 19972 3834
rect 19996 3782 20034 3834
rect 20034 3782 20046 3834
rect 20046 3782 20052 3834
rect 20076 3782 20098 3834
rect 20098 3782 20110 3834
rect 20110 3782 20132 3834
rect 20156 3782 20162 3834
rect 20162 3782 20174 3834
rect 20174 3782 20212 3834
rect 20236 3782 20238 3834
rect 20238 3782 20290 3834
rect 20290 3782 20292 3834
rect 19916 3780 19972 3782
rect 19996 3780 20052 3782
rect 20076 3780 20132 3782
rect 20156 3780 20212 3782
rect 20236 3780 20292 3782
rect 19890 3476 19892 3496
rect 19892 3476 19944 3496
rect 19944 3476 19946 3496
rect 19890 3440 19946 3476
rect 19916 2746 19972 2748
rect 19996 2746 20052 2748
rect 20076 2746 20132 2748
rect 20156 2746 20212 2748
rect 20236 2746 20292 2748
rect 19916 2694 19918 2746
rect 19918 2694 19970 2746
rect 19970 2694 19972 2746
rect 19996 2694 20034 2746
rect 20034 2694 20046 2746
rect 20046 2694 20052 2746
rect 20076 2694 20098 2746
rect 20098 2694 20110 2746
rect 20110 2694 20132 2746
rect 20156 2694 20162 2746
rect 20162 2694 20174 2746
rect 20174 2694 20212 2746
rect 20236 2694 20238 2746
rect 20238 2694 20290 2746
rect 20290 2694 20292 2746
rect 19916 2692 19972 2694
rect 19996 2692 20052 2694
rect 20076 2692 20132 2694
rect 20156 2692 20212 2694
rect 20236 2692 20292 2694
rect 20442 2760 20498 2816
rect 20656 3290 20712 3292
rect 20736 3290 20792 3292
rect 20816 3290 20872 3292
rect 20896 3290 20952 3292
rect 20976 3290 21032 3292
rect 20656 3238 20658 3290
rect 20658 3238 20710 3290
rect 20710 3238 20712 3290
rect 20736 3238 20774 3290
rect 20774 3238 20786 3290
rect 20786 3238 20792 3290
rect 20816 3238 20838 3290
rect 20838 3238 20850 3290
rect 20850 3238 20872 3290
rect 20896 3238 20902 3290
rect 20902 3238 20914 3290
rect 20914 3238 20952 3290
rect 20976 3238 20978 3290
rect 20978 3238 21030 3290
rect 21030 3238 21032 3290
rect 20656 3236 20712 3238
rect 20736 3236 20792 3238
rect 20816 3236 20872 3238
rect 20896 3236 20952 3238
rect 20976 3236 21032 3238
rect 20656 2202 20712 2204
rect 20736 2202 20792 2204
rect 20816 2202 20872 2204
rect 20896 2202 20952 2204
rect 20976 2202 21032 2204
rect 20656 2150 20658 2202
rect 20658 2150 20710 2202
rect 20710 2150 20712 2202
rect 20736 2150 20774 2202
rect 20774 2150 20786 2202
rect 20786 2150 20792 2202
rect 20816 2150 20838 2202
rect 20838 2150 20850 2202
rect 20850 2150 20872 2202
rect 20896 2150 20902 2202
rect 20902 2150 20914 2202
rect 20914 2150 20952 2202
rect 20976 2150 20978 2202
rect 20978 2150 21030 2202
rect 21030 2150 21032 2202
rect 20656 2148 20712 2150
rect 20736 2148 20792 2150
rect 20816 2148 20872 2150
rect 20896 2148 20952 2150
rect 20976 2148 21032 2150
rect 21546 6976 21602 7032
rect 21546 6568 21602 6624
rect 21454 6296 21510 6352
rect 21454 6024 21510 6080
rect 21914 8608 21970 8664
rect 22006 8236 22008 8256
rect 22008 8236 22060 8256
rect 22060 8236 22062 8256
rect 22006 8200 22062 8236
rect 21914 7928 21970 7984
rect 21914 6976 21970 7032
rect 21914 6840 21970 6896
rect 22190 8608 22246 8664
rect 22466 6860 22522 6896
rect 22466 6840 22468 6860
rect 22468 6840 22520 6860
rect 22520 6840 22522 6860
rect 22374 6432 22430 6488
rect 21822 5208 21878 5264
rect 22098 5480 22154 5536
rect 21730 4936 21786 4992
rect 22006 4936 22062 4992
rect 21454 4528 21510 4584
rect 21546 4256 21602 4312
rect 22098 3576 22154 3632
rect 21454 3440 21510 3496
rect 21270 2644 21326 2680
rect 21270 2624 21272 2644
rect 21272 2624 21324 2644
rect 21324 2624 21326 2644
rect 22190 2896 22246 2952
rect 22558 4256 22614 4312
rect 22742 7112 22798 7168
rect 22742 6976 22798 7032
rect 23294 7384 23350 7440
rect 23386 6840 23442 6896
rect 23754 8200 23810 8256
rect 23846 5480 23902 5536
rect 23846 5344 23902 5400
rect 23570 4936 23626 4992
rect 23202 3848 23258 3904
rect 23202 3576 23258 3632
rect 23754 4528 23810 4584
rect 22190 1808 22246 1864
rect 24122 5228 24178 5264
rect 24122 5208 24124 5228
rect 24124 5208 24176 5228
rect 24176 5208 24178 5228
rect 24030 4392 24086 4448
rect 24674 10124 24730 10160
rect 24674 10104 24676 10124
rect 24676 10104 24728 10124
rect 24728 10104 24730 10124
rect 24122 3052 24178 3088
rect 24122 3032 24124 3052
rect 24124 3032 24176 3052
rect 24176 3032 24178 3052
rect 24858 6568 24914 6624
rect 24950 6432 25006 6488
rect 25134 6432 25190 6488
rect 24490 5480 24546 5536
rect 24582 5208 24638 5264
rect 24582 4120 24638 4176
rect 24766 3576 24822 3632
rect 25916 8186 25972 8188
rect 25996 8186 26052 8188
rect 26076 8186 26132 8188
rect 26156 8186 26212 8188
rect 26236 8186 26292 8188
rect 25916 8134 25918 8186
rect 25918 8134 25970 8186
rect 25970 8134 25972 8186
rect 25996 8134 26034 8186
rect 26034 8134 26046 8186
rect 26046 8134 26052 8186
rect 26076 8134 26098 8186
rect 26098 8134 26110 8186
rect 26110 8134 26132 8186
rect 26156 8134 26162 8186
rect 26162 8134 26174 8186
rect 26174 8134 26212 8186
rect 26236 8134 26238 8186
rect 26238 8134 26290 8186
rect 26290 8134 26292 8186
rect 25916 8132 25972 8134
rect 25996 8132 26052 8134
rect 26076 8132 26132 8134
rect 26156 8132 26212 8134
rect 26236 8132 26292 8134
rect 25962 7656 26018 7712
rect 26656 8730 26712 8732
rect 26736 8730 26792 8732
rect 26816 8730 26872 8732
rect 26896 8730 26952 8732
rect 26976 8730 27032 8732
rect 26656 8678 26658 8730
rect 26658 8678 26710 8730
rect 26710 8678 26712 8730
rect 26736 8678 26774 8730
rect 26774 8678 26786 8730
rect 26786 8678 26792 8730
rect 26816 8678 26838 8730
rect 26838 8678 26850 8730
rect 26850 8678 26872 8730
rect 26896 8678 26902 8730
rect 26902 8678 26914 8730
rect 26914 8678 26952 8730
rect 26976 8678 26978 8730
rect 26978 8678 27030 8730
rect 27030 8678 27032 8730
rect 26656 8676 26712 8678
rect 26736 8676 26792 8678
rect 26816 8676 26872 8678
rect 26896 8676 26952 8678
rect 26976 8676 27032 8678
rect 26882 7792 26938 7848
rect 26656 7642 26712 7644
rect 26736 7642 26792 7644
rect 26816 7642 26872 7644
rect 26896 7642 26952 7644
rect 26976 7642 27032 7644
rect 26656 7590 26658 7642
rect 26658 7590 26710 7642
rect 26710 7590 26712 7642
rect 26736 7590 26774 7642
rect 26774 7590 26786 7642
rect 26786 7590 26792 7642
rect 26816 7590 26838 7642
rect 26838 7590 26850 7642
rect 26850 7590 26872 7642
rect 26896 7590 26902 7642
rect 26902 7590 26914 7642
rect 26914 7590 26952 7642
rect 26976 7590 26978 7642
rect 26978 7590 27030 7642
rect 27030 7590 27032 7642
rect 26656 7588 26712 7590
rect 26736 7588 26792 7590
rect 26816 7588 26872 7590
rect 26896 7588 26952 7590
rect 26976 7588 27032 7590
rect 25916 7098 25972 7100
rect 25996 7098 26052 7100
rect 26076 7098 26132 7100
rect 26156 7098 26212 7100
rect 26236 7098 26292 7100
rect 25916 7046 25918 7098
rect 25918 7046 25970 7098
rect 25970 7046 25972 7098
rect 25996 7046 26034 7098
rect 26034 7046 26046 7098
rect 26046 7046 26052 7098
rect 26076 7046 26098 7098
rect 26098 7046 26110 7098
rect 26110 7046 26132 7098
rect 26156 7046 26162 7098
rect 26162 7046 26174 7098
rect 26174 7046 26212 7098
rect 26236 7046 26238 7098
rect 26238 7046 26290 7098
rect 26290 7046 26292 7098
rect 25916 7044 25972 7046
rect 25996 7044 26052 7046
rect 26076 7044 26132 7046
rect 26156 7044 26212 7046
rect 26236 7044 26292 7046
rect 26146 6840 26202 6896
rect 26656 6554 26712 6556
rect 26736 6554 26792 6556
rect 26816 6554 26872 6556
rect 26896 6554 26952 6556
rect 26976 6554 27032 6556
rect 26656 6502 26658 6554
rect 26658 6502 26710 6554
rect 26710 6502 26712 6554
rect 26736 6502 26774 6554
rect 26774 6502 26786 6554
rect 26786 6502 26792 6554
rect 26816 6502 26838 6554
rect 26838 6502 26850 6554
rect 26850 6502 26872 6554
rect 26896 6502 26902 6554
rect 26902 6502 26914 6554
rect 26914 6502 26952 6554
rect 26976 6502 26978 6554
rect 26978 6502 27030 6554
rect 27030 6502 27032 6554
rect 26656 6500 26712 6502
rect 26736 6500 26792 6502
rect 26816 6500 26872 6502
rect 26896 6500 26952 6502
rect 26976 6500 27032 6502
rect 27342 9696 27398 9752
rect 27434 7792 27490 7848
rect 27250 7656 27306 7712
rect 25916 6010 25972 6012
rect 25996 6010 26052 6012
rect 26076 6010 26132 6012
rect 26156 6010 26212 6012
rect 26236 6010 26292 6012
rect 25916 5958 25918 6010
rect 25918 5958 25970 6010
rect 25970 5958 25972 6010
rect 25996 5958 26034 6010
rect 26034 5958 26046 6010
rect 26046 5958 26052 6010
rect 26076 5958 26098 6010
rect 26098 5958 26110 6010
rect 26110 5958 26132 6010
rect 26156 5958 26162 6010
rect 26162 5958 26174 6010
rect 26174 5958 26212 6010
rect 26236 5958 26238 6010
rect 26238 5958 26290 6010
rect 26290 5958 26292 6010
rect 25916 5956 25972 5958
rect 25996 5956 26052 5958
rect 26076 5956 26132 5958
rect 26156 5956 26212 5958
rect 26236 5956 26292 5958
rect 26698 5888 26754 5944
rect 25226 5344 25282 5400
rect 25134 4800 25190 4856
rect 25594 3712 25650 3768
rect 25870 5480 25926 5536
rect 26054 5480 26110 5536
rect 25962 5344 26018 5400
rect 26606 5788 26608 5808
rect 26608 5788 26660 5808
rect 26660 5788 26662 5808
rect 26606 5752 26662 5788
rect 27342 6704 27398 6760
rect 27250 6024 27306 6080
rect 26656 5466 26712 5468
rect 26736 5466 26792 5468
rect 26816 5466 26872 5468
rect 26896 5466 26952 5468
rect 26976 5466 27032 5468
rect 26656 5414 26658 5466
rect 26658 5414 26710 5466
rect 26710 5414 26712 5466
rect 26736 5414 26774 5466
rect 26774 5414 26786 5466
rect 26786 5414 26792 5466
rect 26816 5414 26838 5466
rect 26838 5414 26850 5466
rect 26850 5414 26872 5466
rect 26896 5414 26902 5466
rect 26902 5414 26914 5466
rect 26914 5414 26952 5466
rect 26976 5414 26978 5466
rect 26978 5414 27030 5466
rect 27030 5414 27032 5466
rect 26656 5412 26712 5414
rect 26736 5412 26792 5414
rect 26816 5412 26872 5414
rect 26896 5412 26952 5414
rect 26976 5412 27032 5414
rect 26514 5344 26570 5400
rect 26698 5208 26754 5264
rect 26974 5228 27030 5264
rect 26974 5208 26976 5228
rect 26976 5208 27028 5228
rect 27028 5208 27030 5228
rect 25916 4922 25972 4924
rect 25996 4922 26052 4924
rect 26076 4922 26132 4924
rect 26156 4922 26212 4924
rect 26236 4922 26292 4924
rect 25916 4870 25918 4922
rect 25918 4870 25970 4922
rect 25970 4870 25972 4922
rect 25996 4870 26034 4922
rect 26034 4870 26046 4922
rect 26046 4870 26052 4922
rect 26076 4870 26098 4922
rect 26098 4870 26110 4922
rect 26110 4870 26132 4922
rect 26156 4870 26162 4922
rect 26162 4870 26174 4922
rect 26174 4870 26212 4922
rect 26236 4870 26238 4922
rect 26238 4870 26290 4922
rect 26290 4870 26292 4922
rect 25916 4868 25972 4870
rect 25996 4868 26052 4870
rect 26076 4868 26132 4870
rect 26156 4868 26212 4870
rect 26236 4868 26292 4870
rect 25962 4664 26018 4720
rect 25870 4256 25926 4312
rect 26606 4800 26662 4856
rect 26656 4378 26712 4380
rect 26736 4378 26792 4380
rect 26816 4378 26872 4380
rect 26896 4378 26952 4380
rect 26976 4378 27032 4380
rect 26656 4326 26658 4378
rect 26658 4326 26710 4378
rect 26710 4326 26712 4378
rect 26736 4326 26774 4378
rect 26774 4326 26786 4378
rect 26786 4326 26792 4378
rect 26816 4326 26838 4378
rect 26838 4326 26850 4378
rect 26850 4326 26872 4378
rect 26896 4326 26902 4378
rect 26902 4326 26914 4378
rect 26914 4326 26952 4378
rect 26976 4326 26978 4378
rect 26978 4326 27030 4378
rect 27030 4326 27032 4378
rect 26656 4324 26712 4326
rect 26736 4324 26792 4326
rect 26816 4324 26872 4326
rect 26896 4324 26952 4326
rect 26976 4324 27032 4326
rect 26330 3984 26386 4040
rect 26514 3984 26570 4040
rect 25916 3834 25972 3836
rect 25996 3834 26052 3836
rect 26076 3834 26132 3836
rect 26156 3834 26212 3836
rect 26236 3834 26292 3836
rect 25916 3782 25918 3834
rect 25918 3782 25970 3834
rect 25970 3782 25972 3834
rect 25996 3782 26034 3834
rect 26034 3782 26046 3834
rect 26046 3782 26052 3834
rect 26076 3782 26098 3834
rect 26098 3782 26110 3834
rect 26110 3782 26132 3834
rect 26156 3782 26162 3834
rect 26162 3782 26174 3834
rect 26174 3782 26212 3834
rect 26236 3782 26238 3834
rect 26238 3782 26290 3834
rect 26290 3782 26292 3834
rect 25916 3780 25972 3782
rect 25996 3780 26052 3782
rect 26076 3780 26132 3782
rect 26156 3780 26212 3782
rect 26236 3780 26292 3782
rect 26422 3712 26478 3768
rect 25410 2760 25466 2816
rect 25916 2746 25972 2748
rect 25996 2746 26052 2748
rect 26076 2746 26132 2748
rect 26156 2746 26212 2748
rect 26236 2746 26292 2748
rect 25916 2694 25918 2746
rect 25918 2694 25970 2746
rect 25970 2694 25972 2746
rect 25996 2694 26034 2746
rect 26034 2694 26046 2746
rect 26046 2694 26052 2746
rect 26076 2694 26098 2746
rect 26098 2694 26110 2746
rect 26110 2694 26132 2746
rect 26156 2694 26162 2746
rect 26162 2694 26174 2746
rect 26174 2694 26212 2746
rect 26236 2694 26238 2746
rect 26238 2694 26290 2746
rect 26290 2694 26292 2746
rect 25916 2692 25972 2694
rect 25996 2692 26052 2694
rect 26076 2692 26132 2694
rect 26156 2692 26212 2694
rect 26236 2692 26292 2694
rect 25778 2624 25834 2680
rect 26606 3848 26662 3904
rect 27526 6860 27582 6896
rect 27526 6840 27528 6860
rect 27528 6840 27580 6860
rect 27580 6840 27582 6860
rect 27434 6432 27490 6488
rect 27434 5616 27490 5672
rect 27342 4800 27398 4856
rect 27618 4664 27674 4720
rect 27158 3848 27214 3904
rect 26882 3712 26938 3768
rect 26656 3290 26712 3292
rect 26736 3290 26792 3292
rect 26816 3290 26872 3292
rect 26896 3290 26952 3292
rect 26976 3290 27032 3292
rect 26656 3238 26658 3290
rect 26658 3238 26710 3290
rect 26710 3238 26712 3290
rect 26736 3238 26774 3290
rect 26774 3238 26786 3290
rect 26786 3238 26792 3290
rect 26816 3238 26838 3290
rect 26838 3238 26850 3290
rect 26850 3238 26872 3290
rect 26896 3238 26902 3290
rect 26902 3238 26914 3290
rect 26914 3238 26952 3290
rect 26976 3238 26978 3290
rect 26978 3238 27030 3290
rect 27030 3238 27032 3290
rect 26656 3236 26712 3238
rect 26736 3236 26792 3238
rect 26816 3236 26872 3238
rect 26896 3236 26952 3238
rect 26976 3236 27032 3238
rect 27158 2916 27214 2952
rect 27158 2896 27160 2916
rect 27160 2896 27212 2916
rect 27212 2896 27214 2916
rect 26656 2202 26712 2204
rect 26736 2202 26792 2204
rect 26816 2202 26872 2204
rect 26896 2202 26952 2204
rect 26976 2202 27032 2204
rect 26656 2150 26658 2202
rect 26658 2150 26710 2202
rect 26710 2150 26712 2202
rect 26736 2150 26774 2202
rect 26774 2150 26786 2202
rect 26786 2150 26792 2202
rect 26816 2150 26838 2202
rect 26838 2150 26850 2202
rect 26850 2150 26872 2202
rect 26896 2150 26902 2202
rect 26902 2150 26914 2202
rect 26914 2150 26952 2202
rect 26976 2150 26978 2202
rect 26978 2150 27030 2202
rect 27030 2150 27032 2202
rect 26656 2148 26712 2150
rect 26736 2148 26792 2150
rect 26816 2148 26872 2150
rect 26896 2148 26952 2150
rect 26976 2148 27032 2150
rect 26238 1808 26294 1864
rect 28170 8064 28226 8120
rect 28078 6976 28134 7032
rect 28262 6296 28318 6352
rect 28354 5752 28410 5808
rect 28170 5344 28226 5400
rect 28078 5072 28134 5128
rect 28262 4684 28318 4720
rect 28262 4664 28264 4684
rect 28264 4664 28316 4684
rect 28316 4664 28318 4684
rect 28722 9424 28778 9480
rect 28630 6568 28686 6624
rect 28906 6976 28962 7032
rect 29366 7384 29422 7440
rect 28814 6568 28870 6624
rect 28906 6160 28962 6216
rect 28722 5344 28778 5400
rect 28538 4664 28594 4720
rect 28538 4120 28594 4176
rect 28170 3576 28226 3632
rect 28446 3576 28502 3632
rect 29182 5752 29238 5808
rect 29366 5888 29422 5944
rect 29458 5208 29514 5264
rect 29366 5072 29422 5128
rect 29182 4528 29238 4584
rect 28906 3712 28962 3768
rect 29458 1400 29514 1456
rect 29642 5752 29698 5808
rect 29918 7928 29974 7984
rect 30654 10512 30710 10568
rect 30470 7928 30526 7984
rect 31298 9560 31354 9616
rect 30930 8880 30986 8936
rect 30746 7656 30802 7712
rect 30286 5908 30342 5944
rect 30286 5888 30288 5908
rect 30288 5888 30340 5908
rect 30340 5888 30342 5908
rect 30470 5888 30526 5944
rect 30286 5752 30342 5808
rect 30102 3304 30158 3360
rect 31114 7112 31170 7168
rect 30930 6296 30986 6352
rect 30930 4936 30986 4992
rect 30746 3052 30802 3088
rect 30746 3032 30748 3052
rect 30748 3032 30800 3052
rect 30800 3032 30802 3052
rect 30194 2896 30250 2952
rect 30930 4120 30986 4176
rect 31758 9152 31814 9208
rect 32310 8608 32366 8664
rect 31916 8186 31972 8188
rect 31996 8186 32052 8188
rect 32076 8186 32132 8188
rect 32156 8186 32212 8188
rect 32236 8186 32292 8188
rect 31916 8134 31918 8186
rect 31918 8134 31970 8186
rect 31970 8134 31972 8186
rect 31996 8134 32034 8186
rect 32034 8134 32046 8186
rect 32046 8134 32052 8186
rect 32076 8134 32098 8186
rect 32098 8134 32110 8186
rect 32110 8134 32132 8186
rect 32156 8134 32162 8186
rect 32162 8134 32174 8186
rect 32174 8134 32212 8186
rect 32236 8134 32238 8186
rect 32238 8134 32290 8186
rect 32290 8134 32292 8186
rect 31916 8132 31972 8134
rect 31996 8132 32052 8134
rect 32076 8132 32132 8134
rect 32156 8132 32212 8134
rect 32236 8132 32292 8134
rect 31298 6316 31354 6352
rect 31298 6296 31300 6316
rect 31300 6296 31352 6316
rect 31352 6296 31354 6316
rect 31666 6568 31722 6624
rect 31942 7384 31998 7440
rect 31916 7098 31972 7100
rect 31996 7098 32052 7100
rect 32076 7098 32132 7100
rect 32156 7098 32212 7100
rect 32236 7098 32292 7100
rect 31916 7046 31918 7098
rect 31918 7046 31970 7098
rect 31970 7046 31972 7098
rect 31996 7046 32034 7098
rect 32034 7046 32046 7098
rect 32046 7046 32052 7098
rect 32076 7046 32098 7098
rect 32098 7046 32110 7098
rect 32110 7046 32132 7098
rect 32156 7046 32162 7098
rect 32162 7046 32174 7098
rect 32174 7046 32212 7098
rect 32236 7046 32238 7098
rect 32238 7046 32290 7098
rect 32290 7046 32292 7098
rect 31916 7044 31972 7046
rect 31996 7044 32052 7046
rect 32076 7044 32132 7046
rect 32156 7044 32212 7046
rect 32236 7044 32292 7046
rect 31850 6568 31906 6624
rect 32656 8730 32712 8732
rect 32736 8730 32792 8732
rect 32816 8730 32872 8732
rect 32896 8730 32952 8732
rect 32976 8730 33032 8732
rect 32656 8678 32658 8730
rect 32658 8678 32710 8730
rect 32710 8678 32712 8730
rect 32736 8678 32774 8730
rect 32774 8678 32786 8730
rect 32786 8678 32792 8730
rect 32816 8678 32838 8730
rect 32838 8678 32850 8730
rect 32850 8678 32872 8730
rect 32896 8678 32902 8730
rect 32902 8678 32914 8730
rect 32914 8678 32952 8730
rect 32976 8678 32978 8730
rect 32978 8678 33030 8730
rect 33030 8678 33032 8730
rect 32656 8676 32712 8678
rect 32736 8676 32792 8678
rect 32816 8676 32872 8678
rect 32896 8676 32952 8678
rect 32976 8676 33032 8678
rect 32954 8064 33010 8120
rect 32656 7642 32712 7644
rect 32736 7642 32792 7644
rect 32816 7642 32872 7644
rect 32896 7642 32952 7644
rect 32976 7642 33032 7644
rect 32656 7590 32658 7642
rect 32658 7590 32710 7642
rect 32710 7590 32712 7642
rect 32736 7590 32774 7642
rect 32774 7590 32786 7642
rect 32786 7590 32792 7642
rect 32816 7590 32838 7642
rect 32838 7590 32850 7642
rect 32850 7590 32872 7642
rect 32896 7590 32902 7642
rect 32902 7590 32914 7642
rect 32914 7590 32952 7642
rect 32976 7590 32978 7642
rect 32978 7590 33030 7642
rect 33030 7590 33032 7642
rect 32656 7588 32712 7590
rect 32736 7588 32792 7590
rect 32816 7588 32872 7590
rect 32896 7588 32952 7590
rect 32976 7588 33032 7590
rect 32494 7112 32550 7168
rect 32586 6996 32642 7032
rect 32586 6976 32588 6996
rect 32588 6976 32640 6996
rect 32640 6976 32642 6996
rect 32586 6860 32642 6896
rect 32586 6840 32588 6860
rect 32588 6840 32640 6860
rect 32640 6840 32642 6860
rect 31916 6010 31972 6012
rect 31996 6010 32052 6012
rect 32076 6010 32132 6012
rect 32156 6010 32212 6012
rect 32236 6010 32292 6012
rect 31916 5958 31918 6010
rect 31918 5958 31970 6010
rect 31970 5958 31972 6010
rect 31996 5958 32034 6010
rect 32034 5958 32046 6010
rect 32046 5958 32052 6010
rect 32076 5958 32098 6010
rect 32098 5958 32110 6010
rect 32110 5958 32132 6010
rect 32156 5958 32162 6010
rect 32162 5958 32174 6010
rect 32174 5958 32212 6010
rect 32236 5958 32238 6010
rect 32238 5958 32290 6010
rect 32290 5958 32292 6010
rect 31916 5956 31972 5958
rect 31996 5956 32052 5958
rect 32076 5956 32132 5958
rect 32156 5956 32212 5958
rect 32236 5956 32292 5958
rect 31666 5888 31722 5944
rect 31482 5072 31538 5128
rect 31298 4548 31354 4584
rect 31298 4528 31300 4548
rect 31300 4528 31352 4548
rect 31352 4528 31354 4548
rect 31758 5480 31814 5536
rect 31758 5364 31814 5400
rect 31758 5344 31760 5364
rect 31760 5344 31812 5364
rect 31812 5344 31814 5364
rect 32034 5480 32090 5536
rect 31916 4922 31972 4924
rect 31996 4922 32052 4924
rect 32076 4922 32132 4924
rect 32156 4922 32212 4924
rect 32236 4922 32292 4924
rect 31916 4870 31918 4922
rect 31918 4870 31970 4922
rect 31970 4870 31972 4922
rect 31996 4870 32034 4922
rect 32034 4870 32046 4922
rect 32046 4870 32052 4922
rect 32076 4870 32098 4922
rect 32098 4870 32110 4922
rect 32110 4870 32132 4922
rect 32156 4870 32162 4922
rect 32162 4870 32174 4922
rect 32174 4870 32212 4922
rect 32236 4870 32238 4922
rect 32238 4870 32290 4922
rect 32290 4870 32292 4922
rect 31916 4868 31972 4870
rect 31996 4868 32052 4870
rect 32076 4868 32132 4870
rect 32156 4868 32212 4870
rect 32236 4868 32292 4870
rect 31916 3834 31972 3836
rect 31996 3834 32052 3836
rect 32076 3834 32132 3836
rect 32156 3834 32212 3836
rect 32236 3834 32292 3836
rect 31916 3782 31918 3834
rect 31918 3782 31970 3834
rect 31970 3782 31972 3834
rect 31996 3782 32034 3834
rect 32034 3782 32046 3834
rect 32046 3782 32052 3834
rect 32076 3782 32098 3834
rect 32098 3782 32110 3834
rect 32110 3782 32132 3834
rect 32156 3782 32162 3834
rect 32162 3782 32174 3834
rect 32174 3782 32212 3834
rect 32236 3782 32238 3834
rect 32238 3782 32290 3834
rect 32290 3782 32292 3834
rect 31916 3780 31972 3782
rect 31996 3780 32052 3782
rect 32076 3780 32132 3782
rect 32156 3780 32212 3782
rect 32236 3780 32292 3782
rect 32656 6554 32712 6556
rect 32736 6554 32792 6556
rect 32816 6554 32872 6556
rect 32896 6554 32952 6556
rect 32976 6554 33032 6556
rect 32656 6502 32658 6554
rect 32658 6502 32710 6554
rect 32710 6502 32712 6554
rect 32736 6502 32774 6554
rect 32774 6502 32786 6554
rect 32786 6502 32792 6554
rect 32816 6502 32838 6554
rect 32838 6502 32850 6554
rect 32850 6502 32872 6554
rect 32896 6502 32902 6554
rect 32902 6502 32914 6554
rect 32914 6502 32952 6554
rect 32976 6502 32978 6554
rect 32978 6502 33030 6554
rect 33030 6502 33032 6554
rect 32656 6500 32712 6502
rect 32736 6500 32792 6502
rect 32816 6500 32872 6502
rect 32896 6500 32952 6502
rect 32976 6500 33032 6502
rect 32678 6024 32734 6080
rect 32862 6316 32918 6352
rect 32862 6296 32864 6316
rect 32864 6296 32916 6316
rect 32916 6296 32918 6316
rect 32656 5466 32712 5468
rect 32736 5466 32792 5468
rect 32816 5466 32872 5468
rect 32896 5466 32952 5468
rect 32976 5466 33032 5468
rect 32656 5414 32658 5466
rect 32658 5414 32710 5466
rect 32710 5414 32712 5466
rect 32736 5414 32774 5466
rect 32774 5414 32786 5466
rect 32786 5414 32792 5466
rect 32816 5414 32838 5466
rect 32838 5414 32850 5466
rect 32850 5414 32872 5466
rect 32896 5414 32902 5466
rect 32902 5414 32914 5466
rect 32914 5414 32952 5466
rect 32976 5414 32978 5466
rect 32978 5414 33030 5466
rect 33030 5414 33032 5466
rect 32656 5412 32712 5414
rect 32736 5412 32792 5414
rect 32816 5412 32872 5414
rect 32896 5412 32952 5414
rect 32976 5412 33032 5414
rect 32494 4936 32550 4992
rect 32402 4800 32458 4856
rect 32954 4664 33010 4720
rect 32656 4378 32712 4380
rect 32736 4378 32792 4380
rect 32816 4378 32872 4380
rect 32896 4378 32952 4380
rect 32976 4378 33032 4380
rect 32656 4326 32658 4378
rect 32658 4326 32710 4378
rect 32710 4326 32712 4378
rect 32736 4326 32774 4378
rect 32774 4326 32786 4378
rect 32786 4326 32792 4378
rect 32816 4326 32838 4378
rect 32838 4326 32850 4378
rect 32850 4326 32872 4378
rect 32896 4326 32902 4378
rect 32902 4326 32914 4378
rect 32914 4326 32952 4378
rect 32976 4326 32978 4378
rect 32978 4326 33030 4378
rect 33030 4326 33032 4378
rect 32656 4324 32712 4326
rect 32736 4324 32792 4326
rect 32816 4324 32872 4326
rect 32896 4324 32952 4326
rect 32976 4324 33032 4326
rect 32402 3168 32458 3224
rect 32586 4140 32642 4176
rect 32586 4120 32588 4140
rect 32588 4120 32640 4140
rect 32640 4120 32642 4140
rect 33506 9968 33562 10024
rect 33598 7384 33654 7440
rect 33506 6840 33562 6896
rect 32770 3848 32826 3904
rect 32586 3712 32642 3768
rect 32310 3032 32366 3088
rect 32954 3576 33010 3632
rect 32656 3290 32712 3292
rect 32736 3290 32792 3292
rect 32816 3290 32872 3292
rect 32896 3290 32952 3292
rect 32976 3290 33032 3292
rect 32656 3238 32658 3290
rect 32658 3238 32710 3290
rect 32710 3238 32712 3290
rect 32736 3238 32774 3290
rect 32774 3238 32786 3290
rect 32786 3238 32792 3290
rect 32816 3238 32838 3290
rect 32838 3238 32850 3290
rect 32850 3238 32872 3290
rect 32896 3238 32902 3290
rect 32902 3238 32914 3290
rect 32914 3238 32952 3290
rect 32976 3238 32978 3290
rect 32978 3238 33030 3290
rect 33030 3238 33032 3290
rect 32656 3236 32712 3238
rect 32736 3236 32792 3238
rect 32816 3236 32872 3238
rect 32896 3236 32952 3238
rect 32976 3236 33032 3238
rect 31916 2746 31972 2748
rect 31996 2746 32052 2748
rect 32076 2746 32132 2748
rect 32156 2746 32212 2748
rect 32236 2746 32292 2748
rect 31916 2694 31918 2746
rect 31918 2694 31970 2746
rect 31970 2694 31972 2746
rect 31996 2694 32034 2746
rect 32034 2694 32046 2746
rect 32046 2694 32052 2746
rect 32076 2694 32098 2746
rect 32098 2694 32110 2746
rect 32110 2694 32132 2746
rect 32156 2694 32162 2746
rect 32162 2694 32174 2746
rect 32174 2694 32212 2746
rect 32236 2694 32238 2746
rect 32238 2694 32290 2746
rect 32290 2694 32292 2746
rect 31916 2692 31972 2694
rect 31996 2692 32052 2694
rect 32076 2692 32132 2694
rect 32156 2692 32212 2694
rect 32236 2692 32292 2694
rect 32656 2202 32712 2204
rect 32736 2202 32792 2204
rect 32816 2202 32872 2204
rect 32896 2202 32952 2204
rect 32976 2202 33032 2204
rect 32656 2150 32658 2202
rect 32658 2150 32710 2202
rect 32710 2150 32712 2202
rect 32736 2150 32774 2202
rect 32774 2150 32786 2202
rect 32786 2150 32792 2202
rect 32816 2150 32838 2202
rect 32838 2150 32850 2202
rect 32850 2150 32872 2202
rect 32896 2150 32902 2202
rect 32902 2150 32914 2202
rect 32914 2150 32952 2202
rect 32976 2150 32978 2202
rect 32978 2150 33030 2202
rect 33030 2150 33032 2202
rect 32656 2148 32712 2150
rect 32736 2148 32792 2150
rect 32816 2148 32872 2150
rect 32896 2148 32952 2150
rect 32976 2148 33032 2150
rect 29090 856 29146 912
rect 32770 1264 32826 1320
rect 33046 584 33102 640
rect 33414 4140 33470 4176
rect 33414 4120 33416 4140
rect 33416 4120 33468 4140
rect 33468 4120 33470 4140
rect 33506 3848 33562 3904
rect 33874 8200 33930 8256
rect 34426 9288 34482 9344
rect 34242 6996 34298 7032
rect 34242 6976 34244 6996
rect 34244 6976 34296 6996
rect 34296 6976 34298 6996
rect 33874 6196 33876 6216
rect 33876 6196 33928 6216
rect 33928 6196 33930 6216
rect 33874 6160 33930 6196
rect 33966 3848 34022 3904
rect 33966 1672 34022 1728
rect 35438 10376 35494 10432
rect 35714 10240 35770 10296
rect 34978 8372 34980 8392
rect 34980 8372 35032 8392
rect 35032 8372 35034 8392
rect 34978 8336 35034 8372
rect 34426 4936 34482 4992
rect 34242 4120 34298 4176
rect 34334 3712 34390 3768
rect 35070 5616 35126 5672
rect 35070 4800 35126 4856
rect 35254 6704 35310 6760
rect 35438 6704 35494 6760
rect 35622 6432 35678 6488
rect 36542 8880 36598 8936
rect 36358 8064 36414 8120
rect 35806 7384 35862 7440
rect 35346 4140 35402 4176
rect 35346 4120 35348 4140
rect 35348 4120 35400 4140
rect 35400 4120 35402 4140
rect 35254 3984 35310 4040
rect 34702 3032 34758 3088
rect 35438 3440 35494 3496
rect 34518 1944 34574 2000
rect 36082 7248 36138 7304
rect 35898 3476 35900 3496
rect 35900 3476 35952 3496
rect 35952 3476 35954 3496
rect 35898 3440 35954 3476
rect 36358 4664 36414 4720
rect 33690 720 33746 776
rect 36634 4664 36690 4720
rect 37370 8472 37426 8528
rect 38656 8730 38712 8732
rect 38736 8730 38792 8732
rect 38816 8730 38872 8732
rect 38896 8730 38952 8732
rect 38976 8730 39032 8732
rect 38656 8678 38658 8730
rect 38658 8678 38710 8730
rect 38710 8678 38712 8730
rect 38736 8678 38774 8730
rect 38774 8678 38786 8730
rect 38786 8678 38792 8730
rect 38816 8678 38838 8730
rect 38838 8678 38850 8730
rect 38850 8678 38872 8730
rect 38896 8678 38902 8730
rect 38902 8678 38914 8730
rect 38914 8678 38952 8730
rect 38976 8678 38978 8730
rect 38978 8678 39030 8730
rect 39030 8678 39032 8730
rect 38656 8676 38712 8678
rect 38736 8676 38792 8678
rect 38816 8676 38872 8678
rect 38896 8676 38952 8678
rect 38976 8676 39032 8678
rect 37916 8186 37972 8188
rect 37996 8186 38052 8188
rect 38076 8186 38132 8188
rect 38156 8186 38212 8188
rect 38236 8186 38292 8188
rect 37916 8134 37918 8186
rect 37918 8134 37970 8186
rect 37970 8134 37972 8186
rect 37996 8134 38034 8186
rect 38034 8134 38046 8186
rect 38046 8134 38052 8186
rect 38076 8134 38098 8186
rect 38098 8134 38110 8186
rect 38110 8134 38132 8186
rect 38156 8134 38162 8186
rect 38162 8134 38174 8186
rect 38174 8134 38212 8186
rect 38236 8134 38238 8186
rect 38238 8134 38290 8186
rect 38290 8134 38292 8186
rect 37916 8132 37972 8134
rect 37996 8132 38052 8134
rect 38076 8132 38132 8134
rect 38156 8132 38212 8134
rect 38236 8132 38292 8134
rect 37462 6024 37518 6080
rect 37738 6432 37794 6488
rect 36542 2896 36598 2952
rect 37002 1128 37058 1184
rect 37278 1536 37334 1592
rect 37186 992 37242 1048
rect 37916 7098 37972 7100
rect 37996 7098 38052 7100
rect 38076 7098 38132 7100
rect 38156 7098 38212 7100
rect 38236 7098 38292 7100
rect 37916 7046 37918 7098
rect 37918 7046 37970 7098
rect 37970 7046 37972 7098
rect 37996 7046 38034 7098
rect 38034 7046 38046 7098
rect 38046 7046 38052 7098
rect 38076 7046 38098 7098
rect 38098 7046 38110 7098
rect 38110 7046 38132 7098
rect 38156 7046 38162 7098
rect 38162 7046 38174 7098
rect 38174 7046 38212 7098
rect 38236 7046 38238 7098
rect 38238 7046 38290 7098
rect 38290 7046 38292 7098
rect 37916 7044 37972 7046
rect 37996 7044 38052 7046
rect 38076 7044 38132 7046
rect 38156 7044 38212 7046
rect 38236 7044 38292 7046
rect 37916 6010 37972 6012
rect 37996 6010 38052 6012
rect 38076 6010 38132 6012
rect 38156 6010 38212 6012
rect 38236 6010 38292 6012
rect 37916 5958 37918 6010
rect 37918 5958 37970 6010
rect 37970 5958 37972 6010
rect 37996 5958 38034 6010
rect 38034 5958 38046 6010
rect 38046 5958 38052 6010
rect 38076 5958 38098 6010
rect 38098 5958 38110 6010
rect 38110 5958 38132 6010
rect 38156 5958 38162 6010
rect 38162 5958 38174 6010
rect 38174 5958 38212 6010
rect 38236 5958 38238 6010
rect 38238 5958 38290 6010
rect 38290 5958 38292 6010
rect 37916 5956 37972 5958
rect 37996 5956 38052 5958
rect 38076 5956 38132 5958
rect 38156 5956 38212 5958
rect 38236 5956 38292 5958
rect 37916 4922 37972 4924
rect 37996 4922 38052 4924
rect 38076 4922 38132 4924
rect 38156 4922 38212 4924
rect 38236 4922 38292 4924
rect 37916 4870 37918 4922
rect 37918 4870 37970 4922
rect 37970 4870 37972 4922
rect 37996 4870 38034 4922
rect 38034 4870 38046 4922
rect 38046 4870 38052 4922
rect 38076 4870 38098 4922
rect 38098 4870 38110 4922
rect 38110 4870 38132 4922
rect 38156 4870 38162 4922
rect 38162 4870 38174 4922
rect 38174 4870 38212 4922
rect 38236 4870 38238 4922
rect 38238 4870 38290 4922
rect 38290 4870 38292 4922
rect 37916 4868 37972 4870
rect 37996 4868 38052 4870
rect 38076 4868 38132 4870
rect 38156 4868 38212 4870
rect 38236 4868 38292 4870
rect 38656 7642 38712 7644
rect 38736 7642 38792 7644
rect 38816 7642 38872 7644
rect 38896 7642 38952 7644
rect 38976 7642 39032 7644
rect 38656 7590 38658 7642
rect 38658 7590 38710 7642
rect 38710 7590 38712 7642
rect 38736 7590 38774 7642
rect 38774 7590 38786 7642
rect 38786 7590 38792 7642
rect 38816 7590 38838 7642
rect 38838 7590 38850 7642
rect 38850 7590 38872 7642
rect 38896 7590 38902 7642
rect 38902 7590 38914 7642
rect 38914 7590 38952 7642
rect 38976 7590 38978 7642
rect 38978 7590 39030 7642
rect 39030 7590 39032 7642
rect 38656 7588 38712 7590
rect 38736 7588 38792 7590
rect 38816 7588 38872 7590
rect 38896 7588 38952 7590
rect 38976 7588 39032 7590
rect 38750 6704 38806 6760
rect 38656 6554 38712 6556
rect 38736 6554 38792 6556
rect 38816 6554 38872 6556
rect 38896 6554 38952 6556
rect 38976 6554 39032 6556
rect 38656 6502 38658 6554
rect 38658 6502 38710 6554
rect 38710 6502 38712 6554
rect 38736 6502 38774 6554
rect 38774 6502 38786 6554
rect 38786 6502 38792 6554
rect 38816 6502 38838 6554
rect 38838 6502 38850 6554
rect 38850 6502 38872 6554
rect 38896 6502 38902 6554
rect 38902 6502 38914 6554
rect 38914 6502 38952 6554
rect 38976 6502 38978 6554
rect 38978 6502 39030 6554
rect 39030 6502 39032 6554
rect 38656 6500 38712 6502
rect 38736 6500 38792 6502
rect 38816 6500 38872 6502
rect 38896 6500 38952 6502
rect 38976 6500 39032 6502
rect 38656 5466 38712 5468
rect 38736 5466 38792 5468
rect 38816 5466 38872 5468
rect 38896 5466 38952 5468
rect 38976 5466 39032 5468
rect 38656 5414 38658 5466
rect 38658 5414 38710 5466
rect 38710 5414 38712 5466
rect 38736 5414 38774 5466
rect 38774 5414 38786 5466
rect 38786 5414 38792 5466
rect 38816 5414 38838 5466
rect 38838 5414 38850 5466
rect 38850 5414 38872 5466
rect 38896 5414 38902 5466
rect 38902 5414 38914 5466
rect 38914 5414 38952 5466
rect 38976 5414 38978 5466
rect 38978 5414 39030 5466
rect 39030 5414 39032 5466
rect 38656 5412 38712 5414
rect 38736 5412 38792 5414
rect 38816 5412 38872 5414
rect 38896 5412 38952 5414
rect 38976 5412 39032 5414
rect 38474 5092 38530 5128
rect 38474 5072 38476 5092
rect 38476 5072 38528 5092
rect 38528 5072 38530 5092
rect 38290 4664 38346 4720
rect 37916 3834 37972 3836
rect 37996 3834 38052 3836
rect 38076 3834 38132 3836
rect 38156 3834 38212 3836
rect 38236 3834 38292 3836
rect 37916 3782 37918 3834
rect 37918 3782 37970 3834
rect 37970 3782 37972 3834
rect 37996 3782 38034 3834
rect 38034 3782 38046 3834
rect 38046 3782 38052 3834
rect 38076 3782 38098 3834
rect 38098 3782 38110 3834
rect 38110 3782 38132 3834
rect 38156 3782 38162 3834
rect 38162 3782 38174 3834
rect 38174 3782 38212 3834
rect 38236 3782 38238 3834
rect 38238 3782 38290 3834
rect 38290 3782 38292 3834
rect 37916 3780 37972 3782
rect 37996 3780 38052 3782
rect 38076 3780 38132 3782
rect 38156 3780 38212 3782
rect 38236 3780 38292 3782
rect 37916 2746 37972 2748
rect 37996 2746 38052 2748
rect 38076 2746 38132 2748
rect 38156 2746 38212 2748
rect 38236 2746 38292 2748
rect 37916 2694 37918 2746
rect 37918 2694 37970 2746
rect 37970 2694 37972 2746
rect 37996 2694 38034 2746
rect 38034 2694 38046 2746
rect 38046 2694 38052 2746
rect 38076 2694 38098 2746
rect 38098 2694 38110 2746
rect 38110 2694 38132 2746
rect 38156 2694 38162 2746
rect 38162 2694 38174 2746
rect 38174 2694 38212 2746
rect 38236 2694 38238 2746
rect 38238 2694 38290 2746
rect 38290 2694 38292 2746
rect 37916 2692 37972 2694
rect 37996 2692 38052 2694
rect 38076 2692 38132 2694
rect 38156 2692 38212 2694
rect 38236 2692 38292 2694
rect 38656 4378 38712 4380
rect 38736 4378 38792 4380
rect 38816 4378 38872 4380
rect 38896 4378 38952 4380
rect 38976 4378 39032 4380
rect 38656 4326 38658 4378
rect 38658 4326 38710 4378
rect 38710 4326 38712 4378
rect 38736 4326 38774 4378
rect 38774 4326 38786 4378
rect 38786 4326 38792 4378
rect 38816 4326 38838 4378
rect 38838 4326 38850 4378
rect 38850 4326 38872 4378
rect 38896 4326 38902 4378
rect 38902 4326 38914 4378
rect 38914 4326 38952 4378
rect 38976 4326 38978 4378
rect 38978 4326 39030 4378
rect 39030 4326 39032 4378
rect 38656 4324 38712 4326
rect 38736 4324 38792 4326
rect 38816 4324 38872 4326
rect 38896 4324 38952 4326
rect 38976 4324 39032 4326
rect 38656 3290 38712 3292
rect 38736 3290 38792 3292
rect 38816 3290 38872 3292
rect 38896 3290 38952 3292
rect 38976 3290 39032 3292
rect 38656 3238 38658 3290
rect 38658 3238 38710 3290
rect 38710 3238 38712 3290
rect 38736 3238 38774 3290
rect 38774 3238 38786 3290
rect 38786 3238 38792 3290
rect 38816 3238 38838 3290
rect 38838 3238 38850 3290
rect 38850 3238 38872 3290
rect 38896 3238 38902 3290
rect 38902 3238 38914 3290
rect 38914 3238 38952 3290
rect 38976 3238 38978 3290
rect 38978 3238 39030 3290
rect 39030 3238 39032 3290
rect 38656 3236 38712 3238
rect 38736 3236 38792 3238
rect 38816 3236 38872 3238
rect 38896 3236 38952 3238
rect 38976 3236 39032 3238
rect 39578 6704 39634 6760
rect 38656 2202 38712 2204
rect 38736 2202 38792 2204
rect 38816 2202 38872 2204
rect 38896 2202 38952 2204
rect 38976 2202 39032 2204
rect 38656 2150 38658 2202
rect 38658 2150 38710 2202
rect 38710 2150 38712 2202
rect 38736 2150 38774 2202
rect 38774 2150 38786 2202
rect 38786 2150 38792 2202
rect 38816 2150 38838 2202
rect 38838 2150 38850 2202
rect 38850 2150 38872 2202
rect 38896 2150 38902 2202
rect 38902 2150 38914 2202
rect 38914 2150 38952 2202
rect 38976 2150 38978 2202
rect 38978 2150 39030 2202
rect 39030 2150 39032 2202
rect 38656 2148 38712 2150
rect 38736 2148 38792 2150
rect 38816 2148 38872 2150
rect 38896 2148 38952 2150
rect 38976 2148 39032 2150
rect 39394 2488 39450 2544
rect 40682 7792 40738 7848
rect 40958 3440 41014 3496
rect 39946 2352 40002 2408
rect 39486 448 39542 504
rect 42154 7928 42210 7984
rect 43534 9832 43590 9888
rect 43350 9560 43406 9616
rect 43258 9288 43314 9344
rect 43166 9016 43222 9072
rect 42798 8744 42854 8800
rect 43074 8200 43130 8256
rect 42890 7928 42946 7984
rect 42890 7404 42946 7440
rect 42890 7384 42892 7404
rect 42892 7384 42944 7404
rect 42944 7384 42946 7404
rect 43442 8472 43498 8528
rect 43442 7692 43444 7712
rect 43444 7692 43496 7712
rect 43496 7692 43498 7712
rect 43442 7656 43498 7692
rect 43074 7384 43130 7440
rect 43442 7148 43444 7168
rect 43444 7148 43496 7168
rect 43496 7148 43498 7168
rect 43442 7112 43498 7148
rect 43442 6840 43498 6896
rect 43074 6724 43130 6760
rect 43074 6704 43076 6724
rect 43076 6704 43128 6724
rect 43128 6704 43130 6724
rect 42890 6604 42892 6624
rect 42892 6604 42944 6624
rect 42944 6604 42946 6624
rect 42890 6568 42946 6604
rect 43442 6296 43498 6352
rect 42706 5752 42762 5808
rect 43074 6060 43076 6080
rect 43076 6060 43128 6080
rect 43128 6060 43130 6080
rect 43074 6024 43130 6060
rect 43074 5516 43076 5536
rect 43076 5516 43128 5536
rect 43128 5516 43130 5536
rect 43074 5480 43130 5516
rect 43074 4972 43076 4992
rect 43076 4972 43128 4992
rect 43128 4972 43130 4992
rect 43074 4936 43130 4972
rect 43258 5228 43314 5264
rect 43258 5208 43260 5228
rect 43260 5208 43312 5228
rect 43312 5208 43314 5228
rect 43258 4664 43314 4720
rect 43442 5788 43444 5808
rect 43444 5788 43496 5808
rect 43496 5788 43498 5808
rect 43442 5752 43498 5788
rect 43442 5208 43498 5264
rect 43442 4700 43444 4720
rect 43444 4700 43496 4720
rect 43496 4700 43498 4720
rect 43442 4664 43498 4700
rect 43074 4428 43076 4448
rect 43076 4428 43128 4448
rect 43128 4428 43130 4448
rect 43074 4392 43130 4428
rect 43442 4120 43498 4176
rect 43074 3884 43076 3904
rect 43076 3884 43128 3904
rect 43128 3884 43130 3904
rect 43074 3848 43130 3884
rect 43442 3612 43444 3632
rect 43444 3612 43496 3632
rect 43496 3612 43498 3632
rect 43442 3576 43498 3612
rect 43258 3476 43260 3496
rect 43260 3476 43312 3496
rect 43312 3476 43314 3496
rect 43258 3440 43314 3476
rect 42890 2352 42946 2408
rect 42798 1672 42854 1728
rect 42890 1400 42946 1456
rect 43074 3340 43076 3360
rect 43076 3340 43128 3360
rect 43128 3340 43130 3360
rect 43074 3304 43130 3340
rect 43074 2796 43076 2816
rect 43076 2796 43128 2816
rect 43128 2796 43130 2816
rect 43074 2760 43130 2796
rect 43074 2252 43076 2272
rect 43076 2252 43128 2272
rect 43128 2252 43130 2272
rect 43074 2216 43130 2252
rect 43442 3032 43498 3088
rect 43442 2524 43444 2544
rect 43444 2524 43496 2544
rect 43496 2524 43498 2544
rect 43442 2488 43498 2524
<< metal3 >>
rect 6310 10508 6316 10572
rect 6380 10570 6386 10572
rect 30649 10570 30715 10573
rect 6380 10568 30715 10570
rect 6380 10512 30654 10568
rect 30710 10512 30715 10568
rect 6380 10510 30715 10512
rect 6380 10508 6386 10510
rect 30649 10507 30715 10510
rect 10358 10372 10364 10436
rect 10428 10434 10434 10436
rect 35433 10434 35499 10437
rect 10428 10432 35499 10434
rect 10428 10376 35438 10432
rect 35494 10376 35499 10432
rect 10428 10374 35499 10376
rect 10428 10372 10434 10374
rect 35433 10371 35499 10374
rect 19149 10298 19215 10301
rect 21214 10298 21220 10300
rect 19149 10296 21220 10298
rect 19149 10240 19154 10296
rect 19210 10240 21220 10296
rect 19149 10238 21220 10240
rect 19149 10235 19215 10238
rect 21214 10236 21220 10238
rect 21284 10236 21290 10300
rect 21541 10298 21607 10301
rect 35709 10298 35775 10301
rect 21541 10296 35775 10298
rect 21541 10240 21546 10296
rect 21602 10240 35714 10296
rect 35770 10240 35775 10296
rect 21541 10238 35775 10240
rect 21541 10235 21607 10238
rect 35709 10235 35775 10238
rect 5942 10100 5948 10164
rect 6012 10162 6018 10164
rect 24669 10162 24735 10165
rect 6012 10160 24735 10162
rect 6012 10104 24674 10160
rect 24730 10104 24735 10160
rect 6012 10102 24735 10104
rect 6012 10100 6018 10102
rect 24669 10099 24735 10102
rect 11697 10026 11763 10029
rect 33501 10026 33567 10029
rect 11697 10024 33567 10026
rect 11697 9968 11702 10024
rect 11758 9968 33506 10024
rect 33562 9968 33567 10024
rect 11697 9966 33567 9968
rect 11697 9963 11763 9966
rect 33501 9963 33567 9966
rect 0 9890 800 9920
rect 3417 9890 3483 9893
rect 0 9888 3483 9890
rect 0 9832 3422 9888
rect 3478 9832 3483 9888
rect 0 9830 3483 9832
rect 0 9800 800 9830
rect 3417 9827 3483 9830
rect 10041 9890 10107 9893
rect 17125 9890 17191 9893
rect 10041 9888 17191 9890
rect 10041 9832 10046 9888
rect 10102 9832 17130 9888
rect 17186 9832 17191 9888
rect 10041 9830 17191 9832
rect 10041 9827 10107 9830
rect 17125 9827 17191 9830
rect 17350 9828 17356 9892
rect 17420 9890 17426 9892
rect 21541 9890 21607 9893
rect 17420 9888 21607 9890
rect 17420 9832 21546 9888
rect 21602 9832 21607 9888
rect 17420 9830 21607 9832
rect 17420 9828 17426 9830
rect 21541 9827 21607 9830
rect 43529 9890 43595 9893
rect 44200 9890 45000 9920
rect 43529 9888 45000 9890
rect 43529 9832 43534 9888
rect 43590 9832 45000 9888
rect 43529 9830 45000 9832
rect 43529 9827 43595 9830
rect 44200 9800 45000 9830
rect 16982 9692 16988 9756
rect 17052 9754 17058 9756
rect 27337 9754 27403 9757
rect 17052 9752 27403 9754
rect 17052 9696 27342 9752
rect 27398 9696 27403 9752
rect 17052 9694 27403 9696
rect 17052 9692 17058 9694
rect 27337 9691 27403 9694
rect 0 9618 800 9648
rect 3049 9618 3115 9621
rect 0 9616 3115 9618
rect 0 9560 3054 9616
rect 3110 9560 3115 9616
rect 0 9558 3115 9560
rect 0 9528 800 9558
rect 3049 9555 3115 9558
rect 9305 9618 9371 9621
rect 31293 9618 31359 9621
rect 9305 9616 31359 9618
rect 9305 9560 9310 9616
rect 9366 9560 31298 9616
rect 31354 9560 31359 9616
rect 9305 9558 31359 9560
rect 9305 9555 9371 9558
rect 31293 9555 31359 9558
rect 43345 9618 43411 9621
rect 44200 9618 45000 9648
rect 43345 9616 45000 9618
rect 43345 9560 43350 9616
rect 43406 9560 45000 9616
rect 43345 9558 45000 9560
rect 43345 9555 43411 9558
rect 44200 9528 45000 9558
rect 3325 9482 3391 9485
rect 15142 9482 15148 9484
rect 3325 9480 15148 9482
rect 3325 9424 3330 9480
rect 3386 9424 15148 9480
rect 3325 9422 15148 9424
rect 3325 9419 3391 9422
rect 15142 9420 15148 9422
rect 15212 9420 15218 9484
rect 21214 9420 21220 9484
rect 21284 9482 21290 9484
rect 28717 9482 28783 9485
rect 21284 9480 28783 9482
rect 21284 9424 28722 9480
rect 28778 9424 28783 9480
rect 21284 9422 28783 9424
rect 21284 9420 21290 9422
rect 28717 9419 28783 9422
rect 0 9346 800 9376
rect 1393 9346 1459 9349
rect 0 9344 1459 9346
rect 0 9288 1398 9344
rect 1454 9288 1459 9344
rect 0 9286 1459 9288
rect 0 9256 800 9286
rect 1393 9283 1459 9286
rect 10317 9346 10383 9349
rect 34421 9346 34487 9349
rect 10317 9344 34487 9346
rect 10317 9288 10322 9344
rect 10378 9288 34426 9344
rect 34482 9288 34487 9344
rect 10317 9286 34487 9288
rect 10317 9283 10383 9286
rect 34421 9283 34487 9286
rect 43253 9346 43319 9349
rect 44200 9346 45000 9376
rect 43253 9344 45000 9346
rect 43253 9288 43258 9344
rect 43314 9288 45000 9344
rect 43253 9286 45000 9288
rect 43253 9283 43319 9286
rect 44200 9256 45000 9286
rect 9397 9210 9463 9213
rect 31753 9210 31819 9213
rect 9397 9208 31819 9210
rect 9397 9152 9402 9208
rect 9458 9152 31758 9208
rect 31814 9152 31819 9208
rect 9397 9150 31819 9152
rect 9397 9147 9463 9150
rect 31753 9147 31819 9150
rect 0 9074 800 9104
rect 3141 9074 3207 9077
rect 0 9072 3207 9074
rect 0 9016 3146 9072
rect 3202 9016 3207 9072
rect 0 9014 3207 9016
rect 0 8984 800 9014
rect 3141 9011 3207 9014
rect 8017 9074 8083 9077
rect 17718 9074 17724 9076
rect 8017 9072 17724 9074
rect 8017 9016 8022 9072
rect 8078 9016 17724 9072
rect 8017 9014 17724 9016
rect 8017 9011 8083 9014
rect 17718 9012 17724 9014
rect 17788 9012 17794 9076
rect 17953 9074 18019 9077
rect 35014 9074 35020 9076
rect 17953 9072 35020 9074
rect 17953 9016 17958 9072
rect 18014 9016 35020 9072
rect 17953 9014 35020 9016
rect 17953 9011 18019 9014
rect 35014 9012 35020 9014
rect 35084 9012 35090 9076
rect 43161 9074 43227 9077
rect 44200 9074 45000 9104
rect 43161 9072 45000 9074
rect 43161 9016 43166 9072
rect 43222 9016 45000 9072
rect 43161 9014 45000 9016
rect 43161 9011 43227 9014
rect 44200 8984 45000 9014
rect 8385 8938 8451 8941
rect 27654 8938 27660 8940
rect 8385 8936 27660 8938
rect 8385 8880 8390 8936
rect 8446 8880 27660 8936
rect 8385 8878 27660 8880
rect 8385 8875 8451 8878
rect 27654 8876 27660 8878
rect 27724 8876 27730 8940
rect 30925 8938 30991 8941
rect 36537 8938 36603 8941
rect 30925 8936 36603 8938
rect 30925 8880 30930 8936
rect 30986 8880 36542 8936
rect 36598 8880 36603 8936
rect 30925 8878 36603 8880
rect 30925 8875 30991 8878
rect 36537 8875 36603 8878
rect 0 8802 800 8832
rect 2313 8802 2379 8805
rect 0 8800 2379 8802
rect 0 8744 2318 8800
rect 2374 8744 2379 8800
rect 0 8742 2379 8744
rect 0 8712 800 8742
rect 2313 8739 2379 8742
rect 19558 8740 19564 8804
rect 19628 8802 19634 8804
rect 19793 8802 19859 8805
rect 19628 8800 19859 8802
rect 19628 8744 19798 8800
rect 19854 8744 19859 8800
rect 19628 8742 19859 8744
rect 19628 8740 19634 8742
rect 19793 8739 19859 8742
rect 42793 8802 42859 8805
rect 44200 8802 45000 8832
rect 42793 8800 45000 8802
rect 42793 8744 42798 8800
rect 42854 8744 45000 8800
rect 42793 8742 45000 8744
rect 42793 8739 42859 8742
rect 2646 8736 3042 8737
rect 2646 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3042 8736
rect 2646 8671 3042 8672
rect 8646 8736 9042 8737
rect 8646 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9042 8736
rect 8646 8671 9042 8672
rect 14646 8736 15042 8737
rect 14646 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15042 8736
rect 14646 8671 15042 8672
rect 20646 8736 21042 8737
rect 20646 8672 20652 8736
rect 20716 8672 20732 8736
rect 20796 8672 20812 8736
rect 20876 8672 20892 8736
rect 20956 8672 20972 8736
rect 21036 8672 21042 8736
rect 20646 8671 21042 8672
rect 26646 8736 27042 8737
rect 26646 8672 26652 8736
rect 26716 8672 26732 8736
rect 26796 8672 26812 8736
rect 26876 8672 26892 8736
rect 26956 8672 26972 8736
rect 27036 8672 27042 8736
rect 26646 8671 27042 8672
rect 32646 8736 33042 8737
rect 32646 8672 32652 8736
rect 32716 8672 32732 8736
rect 32796 8672 32812 8736
rect 32876 8672 32892 8736
rect 32956 8672 32972 8736
rect 33036 8672 33042 8736
rect 32646 8671 33042 8672
rect 38646 8736 39042 8737
rect 38646 8672 38652 8736
rect 38716 8672 38732 8736
rect 38796 8672 38812 8736
rect 38876 8672 38892 8736
rect 38956 8672 38972 8736
rect 39036 8672 39042 8736
rect 44200 8712 45000 8742
rect 38646 8671 39042 8672
rect 7097 8666 7163 8669
rect 5030 8664 7163 8666
rect 5030 8608 7102 8664
rect 7158 8608 7163 8664
rect 5030 8606 7163 8608
rect 0 8530 800 8560
rect 1669 8530 1735 8533
rect 0 8528 1735 8530
rect 0 8472 1674 8528
rect 1730 8472 1735 8528
rect 0 8470 1735 8472
rect 0 8440 800 8470
rect 1669 8467 1735 8470
rect 5030 8397 5090 8606
rect 7097 8603 7163 8606
rect 15326 8604 15332 8668
rect 15396 8666 15402 8668
rect 20437 8666 20503 8669
rect 15396 8664 20503 8666
rect 15396 8608 20442 8664
rect 20498 8608 20503 8664
rect 15396 8606 20503 8608
rect 15396 8604 15402 8606
rect 20437 8603 20503 8606
rect 21909 8666 21975 8669
rect 22185 8666 22251 8669
rect 21909 8664 22251 8666
rect 21909 8608 21914 8664
rect 21970 8608 22190 8664
rect 22246 8608 22251 8664
rect 21909 8606 22251 8608
rect 21909 8603 21975 8606
rect 22185 8603 22251 8606
rect 32305 8666 32371 8669
rect 32438 8666 32444 8668
rect 32305 8664 32444 8666
rect 32305 8608 32310 8664
rect 32366 8608 32444 8664
rect 32305 8606 32444 8608
rect 32305 8603 32371 8606
rect 32438 8604 32444 8606
rect 32508 8604 32514 8668
rect 10409 8530 10475 8533
rect 37365 8530 37431 8533
rect 10409 8528 37431 8530
rect 10409 8472 10414 8528
rect 10470 8472 37370 8528
rect 37426 8472 37431 8528
rect 10409 8470 37431 8472
rect 10409 8467 10475 8470
rect 37365 8467 37431 8470
rect 43437 8530 43503 8533
rect 44200 8530 45000 8560
rect 43437 8528 45000 8530
rect 43437 8472 43442 8528
rect 43498 8472 45000 8528
rect 43437 8470 45000 8472
rect 43437 8467 43503 8470
rect 44200 8440 45000 8470
rect 4981 8392 5090 8397
rect 4981 8336 4986 8392
rect 5042 8336 5090 8392
rect 4981 8334 5090 8336
rect 5349 8394 5415 8397
rect 10501 8394 10567 8397
rect 5349 8392 10567 8394
rect 5349 8336 5354 8392
rect 5410 8336 10506 8392
rect 10562 8336 10567 8392
rect 5349 8334 10567 8336
rect 4981 8331 5047 8334
rect 5349 8331 5415 8334
rect 10501 8331 10567 8334
rect 10726 8332 10732 8396
rect 10796 8394 10802 8396
rect 10869 8394 10935 8397
rect 12249 8394 12315 8397
rect 15510 8394 15516 8396
rect 10796 8392 12315 8394
rect 10796 8336 10874 8392
rect 10930 8336 12254 8392
rect 12310 8336 12315 8392
rect 10796 8334 12315 8336
rect 10796 8332 10802 8334
rect 10869 8331 10935 8334
rect 12249 8331 12315 8334
rect 13678 8334 15516 8394
rect 0 8258 800 8288
rect 3049 8258 3115 8261
rect 7649 8258 7715 8261
rect 0 8198 1778 8258
rect 0 8168 800 8198
rect 0 7986 800 8016
rect 1485 7986 1551 7989
rect 0 7984 1551 7986
rect 0 7928 1490 7984
rect 1546 7928 1551 7984
rect 0 7926 1551 7928
rect 1718 7986 1778 8198
rect 3049 8256 7715 8258
rect 3049 8200 3054 8256
rect 3110 8200 7654 8256
rect 7710 8200 7715 8256
rect 3049 8198 7715 8200
rect 3049 8195 3115 8198
rect 7649 8195 7715 8198
rect 12801 8258 12867 8261
rect 13486 8258 13492 8260
rect 12801 8256 13492 8258
rect 12801 8200 12806 8256
rect 12862 8200 13492 8256
rect 12801 8198 13492 8200
rect 12801 8195 12867 8198
rect 13486 8196 13492 8198
rect 13556 8196 13562 8260
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 5073 8122 5139 8125
rect 7005 8122 7071 8125
rect 5073 8120 7071 8122
rect 5073 8064 5078 8120
rect 5134 8064 7010 8120
rect 7066 8064 7071 8120
rect 5073 8062 7071 8064
rect 5073 8059 5139 8062
rect 7005 8059 7071 8062
rect 8661 8122 8727 8125
rect 13678 8122 13738 8334
rect 15510 8332 15516 8334
rect 15580 8332 15586 8396
rect 16113 8394 16179 8397
rect 20713 8394 20779 8397
rect 34973 8394 35039 8397
rect 16113 8392 20779 8394
rect 16113 8336 16118 8392
rect 16174 8336 20718 8392
rect 20774 8336 20779 8392
rect 16113 8334 20779 8336
rect 16113 8331 16179 8334
rect 20713 8331 20779 8334
rect 20854 8392 35039 8394
rect 20854 8336 34978 8392
rect 35034 8336 35039 8392
rect 20854 8334 35039 8336
rect 20437 8258 20503 8261
rect 20854 8258 20914 8334
rect 34973 8331 35039 8334
rect 20437 8256 20914 8258
rect 20437 8200 20442 8256
rect 20498 8200 20914 8256
rect 20437 8198 20914 8200
rect 22001 8258 22067 8261
rect 23749 8258 23815 8261
rect 33869 8260 33935 8261
rect 33869 8258 33916 8260
rect 22001 8256 23815 8258
rect 22001 8200 22006 8256
rect 22062 8200 23754 8256
rect 23810 8200 23815 8256
rect 22001 8198 23815 8200
rect 33824 8256 33916 8258
rect 33824 8200 33874 8256
rect 33824 8198 33916 8200
rect 20437 8195 20503 8198
rect 22001 8195 22067 8198
rect 23749 8195 23815 8198
rect 33869 8196 33916 8198
rect 33980 8196 33986 8260
rect 43069 8258 43135 8261
rect 44200 8258 45000 8288
rect 43069 8256 45000 8258
rect 43069 8200 43074 8256
rect 43130 8200 45000 8256
rect 43069 8198 45000 8200
rect 33869 8195 33935 8196
rect 43069 8195 43135 8198
rect 13906 8192 14302 8193
rect 13906 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14302 8192
rect 13906 8127 14302 8128
rect 19906 8192 20302 8193
rect 19906 8128 19912 8192
rect 19976 8128 19992 8192
rect 20056 8128 20072 8192
rect 20136 8128 20152 8192
rect 20216 8128 20232 8192
rect 20296 8128 20302 8192
rect 19906 8127 20302 8128
rect 25906 8192 26302 8193
rect 25906 8128 25912 8192
rect 25976 8128 25992 8192
rect 26056 8128 26072 8192
rect 26136 8128 26152 8192
rect 26216 8128 26232 8192
rect 26296 8128 26302 8192
rect 25906 8127 26302 8128
rect 31906 8192 32302 8193
rect 31906 8128 31912 8192
rect 31976 8128 31992 8192
rect 32056 8128 32072 8192
rect 32136 8128 32152 8192
rect 32216 8128 32232 8192
rect 32296 8128 32302 8192
rect 31906 8127 32302 8128
rect 37906 8192 38302 8193
rect 37906 8128 37912 8192
rect 37976 8128 37992 8192
rect 38056 8128 38072 8192
rect 38136 8128 38152 8192
rect 38216 8128 38232 8192
rect 38296 8128 38302 8192
rect 44200 8168 45000 8198
rect 37906 8127 38302 8128
rect 8661 8120 13738 8122
rect 8661 8064 8666 8120
rect 8722 8064 13738 8120
rect 8661 8062 13738 8064
rect 18045 8122 18111 8125
rect 19701 8122 19767 8125
rect 18045 8120 19767 8122
rect 18045 8064 18050 8120
rect 18106 8064 19706 8120
rect 19762 8064 19767 8120
rect 18045 8062 19767 8064
rect 8661 8059 8727 8062
rect 18045 8059 18111 8062
rect 19701 8059 19767 8062
rect 20478 8060 20484 8124
rect 20548 8122 20554 8124
rect 20548 8062 22110 8122
rect 20548 8060 20554 8062
rect 3049 7986 3115 7989
rect 1718 7984 3115 7986
rect 1718 7928 3054 7984
rect 3110 7928 3115 7984
rect 1718 7926 3115 7928
rect 0 7896 800 7926
rect 1485 7923 1551 7926
rect 3049 7923 3115 7926
rect 5441 7986 5507 7989
rect 13445 7986 13511 7989
rect 21909 7986 21975 7989
rect 5441 7984 9184 7986
rect 5441 7928 5446 7984
rect 5502 7928 9184 7984
rect 5441 7926 9184 7928
rect 5441 7923 5507 7926
rect 2405 7850 2471 7853
rect 8385 7850 8451 7853
rect 8661 7850 8727 7853
rect 2405 7848 8451 7850
rect 2405 7792 2410 7848
rect 2466 7792 8390 7848
rect 8446 7792 8451 7848
rect 2405 7790 8451 7792
rect 2405 7787 2471 7790
rect 8385 7787 8451 7790
rect 8526 7848 8727 7850
rect 8526 7792 8666 7848
rect 8722 7792 8727 7848
rect 8526 7790 8727 7792
rect 0 7714 800 7744
rect 4337 7716 4403 7717
rect 0 7654 2514 7714
rect 0 7624 800 7654
rect 0 7442 800 7472
rect 2313 7442 2379 7445
rect 0 7440 2379 7442
rect 0 7384 2318 7440
rect 2374 7384 2379 7440
rect 0 7382 2379 7384
rect 2454 7442 2514 7654
rect 4286 7652 4292 7716
rect 4356 7714 4403 7716
rect 5257 7714 5323 7717
rect 4356 7712 5323 7714
rect 4398 7656 5262 7712
rect 5318 7656 5323 7712
rect 4356 7654 5323 7656
rect 4356 7652 4403 7654
rect 4337 7651 4403 7652
rect 5257 7651 5323 7654
rect 5809 7714 5875 7717
rect 5942 7714 5948 7716
rect 5809 7712 5948 7714
rect 5809 7656 5814 7712
rect 5870 7656 5948 7712
rect 5809 7654 5948 7656
rect 5809 7651 5875 7654
rect 5942 7652 5948 7654
rect 6012 7652 6018 7716
rect 6177 7714 6243 7717
rect 6310 7714 6316 7716
rect 6177 7712 6316 7714
rect 6177 7656 6182 7712
rect 6238 7656 6316 7712
rect 6177 7654 6316 7656
rect 6177 7651 6243 7654
rect 6310 7652 6316 7654
rect 6380 7652 6386 7716
rect 7373 7714 7439 7717
rect 7741 7714 7807 7717
rect 7373 7712 7807 7714
rect 7373 7656 7378 7712
rect 7434 7656 7746 7712
rect 7802 7656 7807 7712
rect 7373 7654 7807 7656
rect 7373 7651 7439 7654
rect 7741 7651 7807 7654
rect 2646 7648 3042 7649
rect 2646 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3042 7648
rect 2646 7583 3042 7584
rect 3233 7578 3299 7581
rect 8526 7578 8586 7790
rect 8661 7787 8727 7790
rect 9124 7714 9184 7926
rect 13310 7984 21975 7986
rect 13310 7928 13450 7984
rect 13506 7928 21914 7984
rect 21970 7928 21975 7984
rect 13310 7926 21975 7928
rect 22050 7986 22110 8062
rect 26366 8060 26372 8124
rect 26436 8122 26442 8124
rect 28165 8122 28231 8125
rect 26436 8120 28231 8122
rect 26436 8064 28170 8120
rect 28226 8064 28231 8120
rect 26436 8062 28231 8064
rect 26436 8060 26442 8062
rect 28165 8059 28231 8062
rect 32949 8122 33015 8125
rect 36353 8122 36419 8125
rect 32949 8120 36419 8122
rect 32949 8064 32954 8120
rect 33010 8064 36358 8120
rect 36414 8064 36419 8120
rect 32949 8062 36419 8064
rect 32949 8059 33015 8062
rect 36353 8059 36419 8062
rect 29913 7986 29979 7989
rect 22050 7984 29979 7986
rect 22050 7928 29918 7984
rect 29974 7928 29979 7984
rect 22050 7926 29979 7928
rect 12065 7850 12131 7853
rect 13310 7850 13370 7926
rect 13445 7923 13511 7926
rect 21909 7923 21975 7926
rect 29913 7923 29979 7926
rect 30465 7986 30531 7989
rect 42149 7986 42215 7989
rect 30465 7984 42215 7986
rect 30465 7928 30470 7984
rect 30526 7928 42154 7984
rect 42210 7928 42215 7984
rect 30465 7926 42215 7928
rect 30465 7923 30531 7926
rect 42149 7923 42215 7926
rect 42885 7986 42951 7989
rect 44200 7986 45000 8016
rect 42885 7984 45000 7986
rect 42885 7928 42890 7984
rect 42946 7928 45000 7984
rect 42885 7926 45000 7928
rect 42885 7923 42951 7926
rect 44200 7896 45000 7926
rect 12065 7848 13370 7850
rect 12065 7792 12070 7848
rect 12126 7792 13370 7848
rect 12065 7790 13370 7792
rect 12065 7787 12131 7790
rect 13670 7788 13676 7852
rect 13740 7850 13746 7852
rect 14825 7850 14891 7853
rect 16573 7850 16639 7853
rect 17861 7850 17927 7853
rect 26366 7850 26372 7852
rect 13740 7848 15210 7850
rect 13740 7792 14830 7848
rect 14886 7792 15210 7848
rect 13740 7790 15210 7792
rect 13740 7788 13746 7790
rect 14825 7787 14891 7790
rect 9124 7654 12450 7714
rect 8646 7648 9042 7649
rect 8646 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9042 7648
rect 8646 7583 9042 7584
rect 3233 7576 8586 7578
rect 3233 7520 3238 7576
rect 3294 7520 8586 7576
rect 3233 7518 8586 7520
rect 10225 7578 10291 7581
rect 11421 7578 11487 7581
rect 10225 7576 11487 7578
rect 10225 7520 10230 7576
rect 10286 7520 11426 7576
rect 11482 7520 11487 7576
rect 10225 7518 11487 7520
rect 3233 7515 3299 7518
rect 10225 7515 10291 7518
rect 11421 7515 11487 7518
rect 2957 7442 3023 7445
rect 2454 7440 3023 7442
rect 2454 7384 2962 7440
rect 3018 7384 3023 7440
rect 2454 7382 3023 7384
rect 0 7352 800 7382
rect 2313 7379 2379 7382
rect 2957 7379 3023 7382
rect 4061 7442 4127 7445
rect 11789 7442 11855 7445
rect 4061 7440 11855 7442
rect 4061 7384 4066 7440
rect 4122 7384 11794 7440
rect 11850 7384 11855 7440
rect 4061 7382 11855 7384
rect 12390 7442 12450 7654
rect 14646 7648 15042 7649
rect 14646 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15042 7648
rect 14646 7583 15042 7584
rect 12566 7516 12572 7580
rect 12636 7578 12642 7580
rect 13905 7578 13971 7581
rect 12636 7576 13971 7578
rect 12636 7520 13910 7576
rect 13966 7520 13971 7576
rect 12636 7518 13971 7520
rect 15150 7578 15210 7790
rect 16573 7848 26372 7850
rect 16573 7792 16578 7848
rect 16634 7792 17866 7848
rect 17922 7792 26372 7848
rect 16573 7790 26372 7792
rect 16573 7787 16639 7790
rect 17861 7787 17927 7790
rect 26366 7788 26372 7790
rect 26436 7788 26442 7852
rect 26877 7850 26943 7853
rect 26512 7848 26943 7850
rect 26512 7792 26882 7848
rect 26938 7792 26943 7848
rect 26512 7790 26943 7792
rect 17033 7714 17099 7717
rect 18321 7714 18387 7717
rect 17033 7712 18387 7714
rect 17033 7656 17038 7712
rect 17094 7656 18326 7712
rect 18382 7656 18387 7712
rect 17033 7654 18387 7656
rect 17033 7651 17099 7654
rect 18321 7651 18387 7654
rect 21398 7652 21404 7716
rect 21468 7714 21474 7716
rect 25957 7714 26023 7717
rect 26512 7714 26572 7790
rect 26877 7787 26943 7790
rect 27429 7850 27495 7853
rect 40677 7850 40743 7853
rect 27429 7848 40743 7850
rect 27429 7792 27434 7848
rect 27490 7792 40682 7848
rect 40738 7792 40743 7848
rect 27429 7790 40743 7792
rect 27429 7787 27495 7790
rect 40677 7787 40743 7790
rect 21468 7712 26572 7714
rect 21468 7656 25962 7712
rect 26018 7656 26572 7712
rect 21468 7654 26572 7656
rect 27245 7714 27311 7717
rect 30741 7714 30807 7717
rect 27245 7712 30807 7714
rect 27245 7656 27250 7712
rect 27306 7656 30746 7712
rect 30802 7656 30807 7712
rect 27245 7654 30807 7656
rect 21468 7652 21474 7654
rect 25957 7651 26023 7654
rect 27245 7651 27311 7654
rect 30741 7651 30807 7654
rect 43437 7714 43503 7717
rect 44200 7714 45000 7744
rect 43437 7712 45000 7714
rect 43437 7656 43442 7712
rect 43498 7656 45000 7712
rect 43437 7654 45000 7656
rect 43437 7651 43503 7654
rect 20646 7648 21042 7649
rect 20646 7584 20652 7648
rect 20716 7584 20732 7648
rect 20796 7584 20812 7648
rect 20876 7584 20892 7648
rect 20956 7584 20972 7648
rect 21036 7584 21042 7648
rect 20646 7583 21042 7584
rect 26646 7648 27042 7649
rect 26646 7584 26652 7648
rect 26716 7584 26732 7648
rect 26796 7584 26812 7648
rect 26876 7584 26892 7648
rect 26956 7584 26972 7648
rect 27036 7584 27042 7648
rect 26646 7583 27042 7584
rect 32646 7648 33042 7649
rect 32646 7584 32652 7648
rect 32716 7584 32732 7648
rect 32796 7584 32812 7648
rect 32876 7584 32892 7648
rect 32956 7584 32972 7648
rect 33036 7584 33042 7648
rect 32646 7583 33042 7584
rect 38646 7648 39042 7649
rect 38646 7584 38652 7648
rect 38716 7584 38732 7648
rect 38796 7584 38812 7648
rect 38876 7584 38892 7648
rect 38956 7584 38972 7648
rect 39036 7584 39042 7648
rect 44200 7624 45000 7654
rect 38646 7583 39042 7584
rect 20478 7578 20484 7580
rect 15150 7518 20484 7578
rect 12636 7516 12642 7518
rect 13905 7515 13971 7518
rect 20478 7516 20484 7518
rect 20548 7516 20554 7580
rect 26366 7578 26372 7580
rect 22188 7518 26372 7578
rect 16941 7442 17007 7445
rect 22188 7442 22248 7518
rect 26366 7516 26372 7518
rect 26436 7516 26442 7580
rect 12390 7440 17007 7442
rect 12390 7384 16946 7440
rect 17002 7384 17007 7440
rect 12390 7382 17007 7384
rect 4061 7379 4127 7382
rect 11789 7379 11855 7382
rect 16941 7379 17007 7382
rect 17128 7382 22248 7442
rect 23289 7442 23355 7445
rect 29361 7442 29427 7445
rect 23289 7440 29427 7442
rect 23289 7384 23294 7440
rect 23350 7384 29366 7440
rect 29422 7384 29427 7440
rect 23289 7382 29427 7384
rect 3325 7306 3391 7309
rect 12249 7306 12315 7309
rect 3325 7304 12315 7306
rect 3325 7248 3330 7304
rect 3386 7248 12254 7304
rect 12310 7248 12315 7304
rect 3325 7246 12315 7248
rect 3325 7243 3391 7246
rect 12249 7243 12315 7246
rect 13261 7306 13327 7309
rect 15377 7306 15443 7309
rect 16757 7306 16823 7309
rect 17128 7306 17188 7382
rect 23289 7379 23355 7382
rect 29361 7379 29427 7382
rect 31937 7442 32003 7445
rect 33593 7442 33659 7445
rect 31937 7440 33659 7442
rect 31937 7384 31942 7440
rect 31998 7384 33598 7440
rect 33654 7384 33659 7440
rect 31937 7382 33659 7384
rect 31937 7379 32003 7382
rect 33593 7379 33659 7382
rect 35801 7442 35867 7445
rect 42885 7442 42951 7445
rect 35801 7440 42951 7442
rect 35801 7384 35806 7440
rect 35862 7384 42890 7440
rect 42946 7384 42951 7440
rect 35801 7382 42951 7384
rect 35801 7379 35867 7382
rect 42885 7379 42951 7382
rect 43069 7442 43135 7445
rect 44200 7442 45000 7472
rect 43069 7440 45000 7442
rect 43069 7384 43074 7440
rect 43130 7384 45000 7440
rect 43069 7382 45000 7384
rect 43069 7379 43135 7382
rect 44200 7352 45000 7382
rect 13261 7304 17188 7306
rect 13261 7248 13266 7304
rect 13322 7248 15382 7304
rect 15438 7248 16762 7304
rect 16818 7248 17188 7304
rect 13261 7246 17188 7248
rect 18873 7306 18939 7309
rect 36077 7306 36143 7309
rect 18873 7304 36143 7306
rect 18873 7248 18878 7304
rect 18934 7248 36082 7304
rect 36138 7248 36143 7304
rect 18873 7246 36143 7248
rect 13261 7243 13327 7246
rect 15377 7243 15443 7246
rect 16757 7243 16823 7246
rect 18873 7243 18939 7246
rect 36077 7243 36143 7246
rect 0 7170 800 7200
rect 1393 7170 1459 7173
rect 0 7168 1459 7170
rect 0 7112 1398 7168
rect 1454 7112 1459 7168
rect 0 7110 1459 7112
rect 0 7080 800 7110
rect 1393 7107 1459 7110
rect 20621 7170 20687 7173
rect 21582 7170 21588 7172
rect 20621 7168 21588 7170
rect 20621 7112 20626 7168
rect 20682 7112 21588 7168
rect 20621 7110 21588 7112
rect 20621 7107 20687 7110
rect 21582 7108 21588 7110
rect 21652 7108 21658 7172
rect 21766 7108 21772 7172
rect 21836 7170 21842 7172
rect 22737 7170 22803 7173
rect 21836 7168 22803 7170
rect 21836 7112 22742 7168
rect 22798 7112 22803 7168
rect 21836 7110 22803 7112
rect 21836 7108 21842 7110
rect 22737 7107 22803 7110
rect 26366 7108 26372 7172
rect 26436 7170 26442 7172
rect 31109 7170 31175 7173
rect 32489 7172 32555 7173
rect 26436 7168 31175 7170
rect 26436 7112 31114 7168
rect 31170 7112 31175 7168
rect 26436 7110 31175 7112
rect 26436 7108 26442 7110
rect 31109 7107 31175 7110
rect 32438 7108 32444 7172
rect 32508 7170 32555 7172
rect 43437 7170 43503 7173
rect 44200 7170 45000 7200
rect 32508 7168 32600 7170
rect 32550 7112 32600 7168
rect 32508 7110 32600 7112
rect 43437 7168 45000 7170
rect 43437 7112 43442 7168
rect 43498 7112 45000 7168
rect 43437 7110 45000 7112
rect 32508 7108 32555 7110
rect 32489 7107 32555 7108
rect 43437 7107 43503 7110
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 13906 7104 14302 7105
rect 13906 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14302 7104
rect 13906 7039 14302 7040
rect 19906 7104 20302 7105
rect 19906 7040 19912 7104
rect 19976 7040 19992 7104
rect 20056 7040 20072 7104
rect 20136 7040 20152 7104
rect 20216 7040 20232 7104
rect 20296 7040 20302 7104
rect 19906 7039 20302 7040
rect 25906 7104 26302 7105
rect 25906 7040 25912 7104
rect 25976 7040 25992 7104
rect 26056 7040 26072 7104
rect 26136 7040 26152 7104
rect 26216 7040 26232 7104
rect 26296 7040 26302 7104
rect 25906 7039 26302 7040
rect 31906 7104 32302 7105
rect 31906 7040 31912 7104
rect 31976 7040 31992 7104
rect 32056 7040 32072 7104
rect 32136 7040 32152 7104
rect 32216 7040 32232 7104
rect 32296 7040 32302 7104
rect 31906 7039 32302 7040
rect 37906 7104 38302 7105
rect 37906 7040 37912 7104
rect 37976 7040 37992 7104
rect 38056 7040 38072 7104
rect 38136 7040 38152 7104
rect 38216 7040 38232 7104
rect 38296 7040 38302 7104
rect 44200 7080 45000 7110
rect 37906 7039 38302 7040
rect 8385 7034 8451 7037
rect 13077 7034 13143 7037
rect 8385 7032 13143 7034
rect 8385 6976 8390 7032
rect 8446 6976 13082 7032
rect 13138 6976 13143 7032
rect 8385 6974 13143 6976
rect 8385 6971 8451 6974
rect 13077 6971 13143 6974
rect 19057 7034 19123 7037
rect 19190 7034 19196 7036
rect 19057 7032 19196 7034
rect 19057 6976 19062 7032
rect 19118 6976 19196 7032
rect 19057 6974 19196 6976
rect 19057 6971 19123 6974
rect 19190 6972 19196 6974
rect 19260 6972 19266 7036
rect 21214 6972 21220 7036
rect 21284 7034 21290 7036
rect 21541 7034 21607 7037
rect 21284 7032 21607 7034
rect 21284 6976 21546 7032
rect 21602 6976 21607 7032
rect 21284 6974 21607 6976
rect 21284 6972 21290 6974
rect 21541 6971 21607 6974
rect 21909 7034 21975 7037
rect 22737 7034 22803 7037
rect 21909 7032 22803 7034
rect 21909 6976 21914 7032
rect 21970 6976 22742 7032
rect 22798 6976 22803 7032
rect 21909 6974 22803 6976
rect 21909 6971 21975 6974
rect 22737 6971 22803 6974
rect 26366 6972 26372 7036
rect 26436 7034 26442 7036
rect 28073 7034 28139 7037
rect 28901 7034 28967 7037
rect 26436 7032 28967 7034
rect 26436 6976 28078 7032
rect 28134 6976 28906 7032
rect 28962 6976 28967 7032
rect 26436 6974 28967 6976
rect 26436 6972 26442 6974
rect 28073 6971 28139 6974
rect 28901 6971 28967 6974
rect 32581 7034 32647 7037
rect 34237 7034 34303 7037
rect 32581 7032 34303 7034
rect 32581 6976 32586 7032
rect 32642 6976 34242 7032
rect 34298 6976 34303 7032
rect 32581 6974 34303 6976
rect 32581 6971 32647 6974
rect 34237 6971 34303 6974
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 3417 6898 3483 6901
rect 5533 6898 5599 6901
rect 10409 6898 10475 6901
rect 3417 6896 10475 6898
rect 3417 6840 3422 6896
rect 3478 6840 5538 6896
rect 5594 6840 10414 6896
rect 10470 6840 10475 6896
rect 3417 6838 10475 6840
rect 3417 6835 3483 6838
rect 5533 6835 5599 6838
rect 10409 6835 10475 6838
rect 10869 6898 10935 6901
rect 14181 6898 14247 6901
rect 10869 6896 14247 6898
rect 10869 6840 10874 6896
rect 10930 6840 14186 6896
rect 14242 6840 14247 6896
rect 10869 6838 14247 6840
rect 10869 6835 10935 6838
rect 14181 6835 14247 6838
rect 14457 6898 14523 6901
rect 16205 6898 16271 6901
rect 14457 6896 16271 6898
rect 14457 6840 14462 6896
rect 14518 6840 16210 6896
rect 16266 6840 16271 6896
rect 14457 6838 16271 6840
rect 14457 6835 14523 6838
rect 16205 6835 16271 6838
rect 19006 6836 19012 6900
rect 19076 6898 19082 6900
rect 19241 6898 19307 6901
rect 19076 6896 19307 6898
rect 19076 6840 19246 6896
rect 19302 6840 19307 6896
rect 19076 6838 19307 6840
rect 19076 6836 19082 6838
rect 19241 6835 19307 6838
rect 19517 6898 19583 6901
rect 21909 6898 21975 6901
rect 19517 6896 21975 6898
rect 19517 6840 19522 6896
rect 19578 6840 21914 6896
rect 21970 6840 21975 6896
rect 19517 6838 21975 6840
rect 19517 6835 19583 6838
rect 21909 6835 21975 6838
rect 22461 6898 22527 6901
rect 23381 6898 23447 6901
rect 26141 6898 26207 6901
rect 22461 6896 26207 6898
rect 22461 6840 22466 6896
rect 22522 6840 23386 6896
rect 23442 6840 26146 6896
rect 26202 6840 26207 6896
rect 22461 6838 26207 6840
rect 22461 6835 22527 6838
rect 23381 6835 23447 6838
rect 26141 6835 26207 6838
rect 27521 6898 27587 6901
rect 32581 6898 32647 6901
rect 27521 6896 32647 6898
rect 27521 6840 27526 6896
rect 27582 6840 32586 6896
rect 32642 6840 32647 6896
rect 27521 6838 32647 6840
rect 27521 6835 27587 6838
rect 32581 6835 32647 6838
rect 33501 6898 33567 6901
rect 43437 6898 43503 6901
rect 44200 6898 45000 6928
rect 33501 6896 41430 6898
rect 33501 6840 33506 6896
rect 33562 6840 41430 6896
rect 33501 6838 41430 6840
rect 33501 6835 33567 6838
rect 3969 6762 4035 6765
rect 27337 6762 27403 6765
rect 35249 6762 35315 6765
rect 35433 6762 35499 6765
rect 3969 6760 35499 6762
rect 3969 6704 3974 6760
rect 4030 6704 27342 6760
rect 27398 6704 35254 6760
rect 35310 6704 35438 6760
rect 35494 6704 35499 6760
rect 3969 6702 35499 6704
rect 3969 6699 4035 6702
rect 27337 6699 27403 6702
rect 35249 6699 35315 6702
rect 35433 6699 35499 6702
rect 38745 6762 38811 6765
rect 39573 6762 39639 6765
rect 38745 6760 39639 6762
rect 38745 6704 38750 6760
rect 38806 6704 39578 6760
rect 39634 6704 39639 6760
rect 38745 6702 39639 6704
rect 41370 6762 41430 6838
rect 43437 6896 45000 6898
rect 43437 6840 43442 6896
rect 43498 6840 45000 6896
rect 43437 6838 45000 6840
rect 43437 6835 43503 6838
rect 44200 6808 45000 6838
rect 43069 6762 43135 6765
rect 41370 6760 43135 6762
rect 41370 6704 43074 6760
rect 43130 6704 43135 6760
rect 41370 6702 43135 6704
rect 38745 6699 38811 6702
rect 39573 6699 39639 6702
rect 43069 6699 43135 6702
rect 0 6626 800 6656
rect 1485 6626 1551 6629
rect 0 6624 1551 6626
rect 0 6568 1490 6624
rect 1546 6568 1551 6624
rect 0 6566 1551 6568
rect 0 6536 800 6566
rect 1485 6563 1551 6566
rect 10041 6624 10107 6629
rect 10041 6568 10046 6624
rect 10102 6568 10107 6624
rect 10041 6563 10107 6568
rect 11329 6626 11395 6629
rect 12525 6626 12591 6629
rect 11329 6624 12591 6626
rect 11329 6568 11334 6624
rect 11390 6568 12530 6624
rect 12586 6568 12591 6624
rect 11329 6566 12591 6568
rect 11329 6563 11395 6566
rect 12525 6563 12591 6566
rect 17677 6626 17743 6629
rect 20478 6626 20484 6628
rect 17677 6624 20484 6626
rect 17677 6568 17682 6624
rect 17738 6568 20484 6624
rect 17677 6566 20484 6568
rect 17677 6563 17743 6566
rect 20478 6564 20484 6566
rect 20548 6564 20554 6628
rect 21541 6626 21607 6629
rect 24853 6626 24919 6629
rect 21541 6624 24919 6626
rect 21541 6568 21546 6624
rect 21602 6568 24858 6624
rect 24914 6568 24919 6624
rect 21541 6566 24919 6568
rect 21541 6563 21607 6566
rect 24853 6563 24919 6566
rect 28625 6626 28691 6629
rect 28809 6626 28875 6629
rect 28625 6624 28875 6626
rect 28625 6568 28630 6624
rect 28686 6568 28814 6624
rect 28870 6568 28875 6624
rect 28625 6566 28875 6568
rect 28625 6563 28691 6566
rect 28809 6563 28875 6566
rect 31661 6626 31727 6629
rect 31845 6626 31911 6629
rect 31661 6624 31911 6626
rect 31661 6568 31666 6624
rect 31722 6568 31850 6624
rect 31906 6568 31911 6624
rect 31661 6566 31911 6568
rect 31661 6563 31727 6566
rect 31845 6563 31911 6566
rect 42885 6626 42951 6629
rect 44200 6626 45000 6656
rect 42885 6624 45000 6626
rect 42885 6568 42890 6624
rect 42946 6568 45000 6624
rect 42885 6566 45000 6568
rect 42885 6563 42951 6566
rect 2646 6560 3042 6561
rect 2646 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3042 6560
rect 2646 6495 3042 6496
rect 8646 6560 9042 6561
rect 8646 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9042 6560
rect 8646 6495 9042 6496
rect 3325 6490 3391 6493
rect 3785 6490 3851 6493
rect 3325 6488 3851 6490
rect 3325 6432 3330 6488
rect 3386 6432 3790 6488
rect 3846 6432 3851 6488
rect 3325 6430 3851 6432
rect 3325 6427 3391 6430
rect 3785 6427 3851 6430
rect 6729 6490 6795 6493
rect 7925 6490 7991 6493
rect 6729 6488 7991 6490
rect 6729 6432 6734 6488
rect 6790 6432 7930 6488
rect 7986 6432 7991 6488
rect 6729 6430 7991 6432
rect 6729 6427 6795 6430
rect 7925 6427 7991 6430
rect 9305 6490 9371 6493
rect 10044 6490 10104 6563
rect 14646 6560 15042 6561
rect 14646 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15042 6560
rect 14646 6495 15042 6496
rect 20646 6560 21042 6561
rect 20646 6496 20652 6560
rect 20716 6496 20732 6560
rect 20796 6496 20812 6560
rect 20876 6496 20892 6560
rect 20956 6496 20972 6560
rect 21036 6496 21042 6560
rect 20646 6495 21042 6496
rect 26646 6560 27042 6561
rect 26646 6496 26652 6560
rect 26716 6496 26732 6560
rect 26796 6496 26812 6560
rect 26876 6496 26892 6560
rect 26956 6496 26972 6560
rect 27036 6496 27042 6560
rect 26646 6495 27042 6496
rect 32646 6560 33042 6561
rect 32646 6496 32652 6560
rect 32716 6496 32732 6560
rect 32796 6496 32812 6560
rect 32876 6496 32892 6560
rect 32956 6496 32972 6560
rect 33036 6496 33042 6560
rect 32646 6495 33042 6496
rect 38646 6560 39042 6561
rect 38646 6496 38652 6560
rect 38716 6496 38732 6560
rect 38796 6496 38812 6560
rect 38876 6496 38892 6560
rect 38956 6496 38972 6560
rect 39036 6496 39042 6560
rect 44200 6536 45000 6566
rect 38646 6495 39042 6496
rect 11237 6490 11303 6493
rect 19517 6490 19583 6493
rect 22369 6490 22435 6493
rect 24945 6490 25011 6493
rect 9305 6488 11303 6490
rect 9305 6432 9310 6488
rect 9366 6432 11242 6488
rect 11298 6432 11303 6488
rect 9305 6430 11303 6432
rect 9305 6427 9371 6430
rect 11237 6427 11303 6430
rect 17358 6488 19583 6490
rect 17358 6432 19522 6488
rect 19578 6432 19583 6488
rect 17358 6430 19583 6432
rect 0 6354 800 6384
rect 2313 6354 2379 6357
rect 0 6352 2379 6354
rect 0 6296 2318 6352
rect 2374 6296 2379 6352
rect 0 6294 2379 6296
rect 0 6264 800 6294
rect 2313 6291 2379 6294
rect 2497 6354 2563 6357
rect 17125 6354 17191 6357
rect 2497 6352 17191 6354
rect 2497 6296 2502 6352
rect 2558 6296 17130 6352
rect 17186 6296 17191 6352
rect 2497 6294 17191 6296
rect 2497 6291 2563 6294
rect 17125 6291 17191 6294
rect 3417 6218 3483 6221
rect 17358 6218 17418 6430
rect 19517 6427 19583 6430
rect 21268 6488 25011 6490
rect 21268 6432 22374 6488
rect 22430 6432 24950 6488
rect 25006 6432 25011 6488
rect 21268 6430 25011 6432
rect 17585 6354 17651 6357
rect 21268 6354 21328 6430
rect 22369 6427 22435 6430
rect 24945 6427 25011 6430
rect 25129 6490 25195 6493
rect 26366 6490 26372 6492
rect 25129 6488 26372 6490
rect 25129 6432 25134 6488
rect 25190 6432 26372 6488
rect 25129 6430 26372 6432
rect 25129 6427 25195 6430
rect 26366 6428 26372 6430
rect 26436 6428 26442 6492
rect 27102 6428 27108 6492
rect 27172 6490 27178 6492
rect 27429 6490 27495 6493
rect 35617 6490 35683 6493
rect 37733 6490 37799 6493
rect 27172 6488 32506 6490
rect 27172 6432 27434 6488
rect 27490 6432 32506 6488
rect 27172 6430 32506 6432
rect 27172 6428 27178 6430
rect 27429 6427 27495 6430
rect 17585 6352 21328 6354
rect 17585 6296 17590 6352
rect 17646 6296 21328 6352
rect 17585 6294 21328 6296
rect 21449 6354 21515 6357
rect 28257 6354 28323 6357
rect 30925 6354 30991 6357
rect 31293 6354 31359 6357
rect 32446 6356 32506 6430
rect 35617 6488 37799 6490
rect 35617 6432 35622 6488
rect 35678 6432 37738 6488
rect 37794 6432 37799 6488
rect 35617 6430 37799 6432
rect 35617 6427 35683 6430
rect 37733 6427 37799 6430
rect 32438 6354 32444 6356
rect 21449 6352 31359 6354
rect 21449 6296 21454 6352
rect 21510 6296 28262 6352
rect 28318 6296 30930 6352
rect 30986 6296 31298 6352
rect 31354 6296 31359 6352
rect 21449 6294 31359 6296
rect 32356 6294 32444 6354
rect 17585 6291 17651 6294
rect 21449 6291 21515 6294
rect 28257 6291 28323 6294
rect 30925 6291 30991 6294
rect 31293 6291 31359 6294
rect 32438 6292 32444 6294
rect 32508 6354 32514 6356
rect 32857 6354 32923 6357
rect 32508 6352 32923 6354
rect 32508 6296 32862 6352
rect 32918 6296 32923 6352
rect 32508 6294 32923 6296
rect 32508 6292 32514 6294
rect 32857 6291 32923 6294
rect 43437 6354 43503 6357
rect 44200 6354 45000 6384
rect 43437 6352 45000 6354
rect 43437 6296 43442 6352
rect 43498 6296 45000 6352
rect 43437 6294 45000 6296
rect 43437 6291 43503 6294
rect 44200 6264 45000 6294
rect 3417 6216 17418 6218
rect 3417 6160 3422 6216
rect 3478 6160 17418 6216
rect 3417 6158 17418 6160
rect 17493 6218 17559 6221
rect 18689 6218 18755 6221
rect 17493 6216 18755 6218
rect 17493 6160 17498 6216
rect 17554 6160 18694 6216
rect 18750 6160 18755 6216
rect 17493 6158 18755 6160
rect 3417 6155 3483 6158
rect 17493 6155 17559 6158
rect 18689 6155 18755 6158
rect 18873 6218 18939 6221
rect 28901 6218 28967 6221
rect 33869 6218 33935 6221
rect 18873 6216 28967 6218
rect 18873 6160 18878 6216
rect 18934 6160 28906 6216
rect 28962 6160 28967 6216
rect 18873 6158 28967 6160
rect 18873 6155 18939 6158
rect 28901 6155 28967 6158
rect 31756 6216 33935 6218
rect 31756 6160 33874 6216
rect 33930 6160 33935 6216
rect 31756 6158 33935 6160
rect 0 6082 800 6112
rect 1393 6082 1459 6085
rect 0 6080 1459 6082
rect 0 6024 1398 6080
rect 1454 6024 1459 6080
rect 0 6022 1459 6024
rect 0 5992 800 6022
rect 1393 6019 1459 6022
rect 3601 6082 3667 6085
rect 3969 6082 4035 6085
rect 5349 6082 5415 6085
rect 3601 6080 5415 6082
rect 3601 6024 3606 6080
rect 3662 6024 3974 6080
rect 4030 6024 5354 6080
rect 5410 6024 5415 6080
rect 3601 6022 5415 6024
rect 3601 6019 3667 6022
rect 3969 6019 4035 6022
rect 5349 6019 5415 6022
rect 8661 6082 8727 6085
rect 10869 6082 10935 6085
rect 8661 6080 10935 6082
rect 8661 6024 8666 6080
rect 8722 6024 10874 6080
rect 10930 6024 10935 6080
rect 8661 6022 10935 6024
rect 8661 6019 8727 6022
rect 10869 6019 10935 6022
rect 11237 6082 11303 6085
rect 13445 6082 13511 6085
rect 11237 6080 13511 6082
rect 11237 6024 11242 6080
rect 11298 6024 13450 6080
rect 13506 6024 13511 6080
rect 11237 6022 13511 6024
rect 11237 6019 11303 6022
rect 13445 6019 13511 6022
rect 14641 6082 14707 6085
rect 15193 6082 15259 6085
rect 18781 6082 18847 6085
rect 14641 6080 15259 6082
rect 14641 6024 14646 6080
rect 14702 6024 15198 6080
rect 15254 6024 15259 6080
rect 14641 6022 15259 6024
rect 14641 6019 14707 6022
rect 15193 6019 15259 6022
rect 17312 6080 18847 6082
rect 17312 6024 18786 6080
rect 18842 6024 18847 6080
rect 17312 6022 18847 6024
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 13906 6016 14302 6017
rect 13906 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14302 6016
rect 13906 5951 14302 5952
rect 17312 5949 17372 6022
rect 18781 6019 18847 6022
rect 18965 6082 19031 6085
rect 19701 6082 19767 6085
rect 18965 6080 19767 6082
rect 18965 6024 18970 6080
rect 19026 6024 19706 6080
rect 19762 6024 19767 6080
rect 18965 6022 19767 6024
rect 18965 6019 19031 6022
rect 19701 6019 19767 6022
rect 20478 6020 20484 6084
rect 20548 6082 20554 6084
rect 21449 6082 21515 6085
rect 27102 6082 27108 6084
rect 20548 6080 21515 6082
rect 20548 6024 21454 6080
rect 21510 6024 21515 6080
rect 20548 6022 21515 6024
rect 20548 6020 20554 6022
rect 21449 6019 21515 6022
rect 26420 6022 27108 6082
rect 19906 6016 20302 6017
rect 19906 5952 19912 6016
rect 19976 5952 19992 6016
rect 20056 5952 20072 6016
rect 20136 5952 20152 6016
rect 20216 5952 20232 6016
rect 20296 5952 20302 6016
rect 19906 5951 20302 5952
rect 25906 6016 26302 6017
rect 25906 5952 25912 6016
rect 25976 5952 25992 6016
rect 26056 5952 26072 6016
rect 26136 5952 26152 6016
rect 26216 5952 26232 6016
rect 26296 5952 26302 6016
rect 25906 5951 26302 5952
rect 9765 5946 9831 5949
rect 10041 5946 10107 5949
rect 8388 5944 10107 5946
rect 8388 5888 9770 5944
rect 9826 5888 10046 5944
rect 10102 5888 10107 5944
rect 8388 5886 10107 5888
rect 0 5810 800 5840
rect 1669 5810 1735 5813
rect 0 5808 1735 5810
rect 0 5752 1674 5808
rect 1730 5752 1735 5808
rect 0 5750 1735 5752
rect 0 5720 800 5750
rect 1669 5747 1735 5750
rect 4613 5810 4679 5813
rect 5165 5810 5231 5813
rect 4613 5808 5231 5810
rect 4613 5752 4618 5808
rect 4674 5752 5170 5808
rect 5226 5752 5231 5808
rect 4613 5750 5231 5752
rect 4613 5747 4679 5750
rect 5165 5747 5231 5750
rect 6729 5810 6795 5813
rect 8388 5810 8448 5886
rect 9765 5883 9831 5886
rect 10041 5883 10107 5886
rect 14549 5946 14615 5949
rect 17033 5946 17099 5949
rect 14549 5944 17099 5946
rect 14549 5888 14554 5944
rect 14610 5888 17038 5944
rect 17094 5888 17099 5944
rect 14549 5886 17099 5888
rect 14549 5883 14615 5886
rect 17033 5883 17099 5886
rect 17309 5944 17375 5949
rect 17309 5888 17314 5944
rect 17370 5888 17375 5944
rect 17309 5883 17375 5888
rect 17677 5946 17743 5949
rect 19609 5946 19675 5949
rect 17677 5944 19675 5946
rect 17677 5888 17682 5944
rect 17738 5888 19614 5944
rect 19670 5888 19675 5944
rect 17677 5886 19675 5888
rect 17677 5883 17743 5886
rect 19609 5883 19675 5886
rect 20478 5884 20484 5948
rect 20548 5946 20554 5948
rect 20897 5946 20963 5949
rect 20548 5944 20963 5946
rect 20548 5888 20902 5944
rect 20958 5888 20963 5944
rect 20548 5886 20963 5888
rect 20548 5884 20554 5886
rect 20897 5883 20963 5886
rect 6729 5808 8448 5810
rect 6729 5752 6734 5808
rect 6790 5752 8448 5808
rect 6729 5750 8448 5752
rect 6729 5747 6795 5750
rect 9438 5748 9444 5812
rect 9508 5810 9514 5812
rect 9857 5810 9923 5813
rect 9508 5808 9923 5810
rect 9508 5752 9862 5808
rect 9918 5752 9923 5808
rect 9508 5750 9923 5752
rect 9508 5748 9514 5750
rect 9857 5747 9923 5750
rect 10777 5810 10843 5813
rect 26420 5810 26480 6022
rect 27102 6020 27108 6022
rect 27172 6020 27178 6084
rect 27245 6082 27311 6085
rect 31756 6082 31816 6158
rect 33869 6155 33935 6158
rect 27245 6080 31816 6082
rect 27245 6024 27250 6080
rect 27306 6024 31816 6080
rect 27245 6022 31816 6024
rect 32673 6082 32739 6085
rect 37457 6082 37523 6085
rect 32673 6080 37523 6082
rect 32673 6024 32678 6080
rect 32734 6024 37462 6080
rect 37518 6024 37523 6080
rect 32673 6022 37523 6024
rect 27245 6019 27311 6022
rect 32673 6019 32739 6022
rect 37457 6019 37523 6022
rect 43069 6082 43135 6085
rect 44200 6082 45000 6112
rect 43069 6080 45000 6082
rect 43069 6024 43074 6080
rect 43130 6024 45000 6080
rect 43069 6022 45000 6024
rect 43069 6019 43135 6022
rect 31906 6016 32302 6017
rect 31906 5952 31912 6016
rect 31976 5952 31992 6016
rect 32056 5952 32072 6016
rect 32136 5952 32152 6016
rect 32216 5952 32232 6016
rect 32296 5952 32302 6016
rect 31906 5951 32302 5952
rect 37906 6016 38302 6017
rect 37906 5952 37912 6016
rect 37976 5952 37992 6016
rect 38056 5952 38072 6016
rect 38136 5952 38152 6016
rect 38216 5952 38232 6016
rect 38296 5952 38302 6016
rect 44200 5992 45000 6022
rect 37906 5951 38302 5952
rect 26693 5946 26759 5949
rect 28022 5946 28028 5948
rect 26693 5944 28028 5946
rect 26693 5888 26698 5944
rect 26754 5888 28028 5944
rect 26693 5886 28028 5888
rect 26693 5883 26759 5886
rect 28022 5884 28028 5886
rect 28092 5884 28098 5948
rect 29361 5946 29427 5949
rect 30281 5946 30347 5949
rect 29361 5944 30347 5946
rect 29361 5888 29366 5944
rect 29422 5888 30286 5944
rect 30342 5888 30347 5944
rect 29361 5886 30347 5888
rect 29361 5883 29427 5886
rect 30281 5883 30347 5886
rect 30465 5946 30531 5949
rect 31661 5946 31727 5949
rect 30465 5944 31727 5946
rect 30465 5888 30470 5944
rect 30526 5888 31666 5944
rect 31722 5888 31727 5944
rect 30465 5886 31727 5888
rect 30465 5883 30531 5886
rect 31661 5883 31727 5886
rect 10777 5808 26480 5810
rect 10777 5752 10782 5808
rect 10838 5752 26480 5808
rect 10777 5750 26480 5752
rect 26601 5810 26667 5813
rect 28349 5810 28415 5813
rect 26601 5808 28415 5810
rect 26601 5752 26606 5808
rect 26662 5752 28354 5808
rect 28410 5752 28415 5808
rect 26601 5750 28415 5752
rect 10777 5747 10843 5750
rect 26601 5747 26667 5750
rect 28349 5747 28415 5750
rect 29177 5810 29243 5813
rect 29637 5810 29703 5813
rect 29177 5808 29703 5810
rect 29177 5752 29182 5808
rect 29238 5752 29642 5808
rect 29698 5752 29703 5808
rect 29177 5750 29703 5752
rect 29177 5747 29243 5750
rect 29637 5747 29703 5750
rect 30281 5810 30347 5813
rect 42701 5810 42767 5813
rect 30281 5808 42767 5810
rect 30281 5752 30286 5808
rect 30342 5752 42706 5808
rect 42762 5752 42767 5808
rect 30281 5750 42767 5752
rect 30281 5747 30347 5750
rect 42701 5747 42767 5750
rect 43437 5810 43503 5813
rect 44200 5810 45000 5840
rect 43437 5808 45000 5810
rect 43437 5752 43442 5808
rect 43498 5752 45000 5808
rect 43437 5750 45000 5752
rect 43437 5747 43503 5750
rect 44200 5720 45000 5750
rect 3233 5674 3299 5677
rect 4286 5674 4292 5676
rect 3233 5672 4292 5674
rect 3233 5616 3238 5672
rect 3294 5616 4292 5672
rect 3233 5614 4292 5616
rect 3233 5611 3299 5614
rect 4286 5612 4292 5614
rect 4356 5612 4362 5676
rect 4797 5674 4863 5677
rect 5257 5674 5323 5677
rect 4797 5672 5323 5674
rect 4797 5616 4802 5672
rect 4858 5616 5262 5672
rect 5318 5616 5323 5672
rect 4797 5614 5323 5616
rect 4797 5611 4863 5614
rect 5257 5611 5323 5614
rect 5533 5674 5599 5677
rect 10501 5674 10567 5677
rect 12566 5674 12572 5676
rect 5533 5672 9322 5674
rect 5533 5616 5538 5672
rect 5594 5616 9322 5672
rect 5533 5614 9322 5616
rect 5533 5611 5599 5614
rect 0 5538 800 5568
rect 2497 5538 2563 5541
rect 0 5536 2563 5538
rect 0 5480 2502 5536
rect 2558 5480 2563 5536
rect 0 5478 2563 5480
rect 0 5448 800 5478
rect 2497 5475 2563 5478
rect 3141 5538 3207 5541
rect 4153 5538 4219 5541
rect 8017 5538 8083 5541
rect 3141 5536 8083 5538
rect 3141 5480 3146 5536
rect 3202 5480 4158 5536
rect 4214 5480 8022 5536
rect 8078 5480 8083 5536
rect 3141 5478 8083 5480
rect 9262 5538 9322 5614
rect 10501 5672 12572 5674
rect 10501 5616 10506 5672
rect 10562 5616 12572 5672
rect 10501 5614 12572 5616
rect 10501 5611 10567 5614
rect 12566 5612 12572 5614
rect 12636 5612 12642 5676
rect 12985 5674 13051 5677
rect 19609 5676 19675 5677
rect 12985 5672 15762 5674
rect 12985 5616 12990 5672
rect 13046 5616 15762 5672
rect 12985 5614 15762 5616
rect 12985 5611 13051 5614
rect 15702 5541 15762 5614
rect 19558 5612 19564 5676
rect 19628 5674 19675 5676
rect 21398 5674 21404 5676
rect 19628 5672 19720 5674
rect 19670 5616 19720 5672
rect 19628 5614 19720 5616
rect 20486 5614 21404 5674
rect 19628 5612 19675 5614
rect 19609 5611 19675 5612
rect 12065 5538 12131 5541
rect 15561 5538 15627 5541
rect 9262 5536 12131 5538
rect 9262 5480 12070 5536
rect 12126 5480 12131 5536
rect 9262 5478 12131 5480
rect 3141 5475 3207 5478
rect 4153 5475 4219 5478
rect 8017 5475 8083 5478
rect 12065 5475 12131 5478
rect 15518 5536 15627 5538
rect 15518 5480 15566 5536
rect 15622 5480 15627 5536
rect 15518 5475 15627 5480
rect 15702 5536 15811 5541
rect 15702 5480 15750 5536
rect 15806 5480 15811 5536
rect 15702 5478 15811 5480
rect 15745 5475 15811 5478
rect 18137 5538 18203 5541
rect 18505 5538 18571 5541
rect 18137 5536 18571 5538
rect 18137 5480 18142 5536
rect 18198 5480 18510 5536
rect 18566 5480 18571 5536
rect 18137 5478 18571 5480
rect 18137 5475 18203 5478
rect 18505 5475 18571 5478
rect 18689 5538 18755 5541
rect 20486 5538 20546 5614
rect 21398 5612 21404 5614
rect 21468 5612 21474 5676
rect 27429 5674 27495 5677
rect 35065 5674 35131 5677
rect 21774 5672 35131 5674
rect 21774 5616 27434 5672
rect 27490 5616 35070 5672
rect 35126 5616 35131 5672
rect 21774 5614 35131 5616
rect 21774 5538 21834 5614
rect 27429 5611 27495 5614
rect 35065 5611 35131 5614
rect 18689 5536 20546 5538
rect 18689 5480 18694 5536
rect 18750 5480 20546 5536
rect 18689 5478 20546 5480
rect 21222 5478 21834 5538
rect 22093 5538 22159 5541
rect 23841 5538 23907 5541
rect 22093 5536 23907 5538
rect 22093 5480 22098 5536
rect 22154 5480 23846 5536
rect 23902 5480 23907 5536
rect 22093 5478 23907 5480
rect 18689 5475 18755 5478
rect 2646 5472 3042 5473
rect 2646 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3042 5472
rect 2646 5407 3042 5408
rect 8646 5472 9042 5473
rect 8646 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9042 5472
rect 8646 5407 9042 5408
rect 14646 5472 15042 5473
rect 14646 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15042 5472
rect 14646 5407 15042 5408
rect 3693 5402 3759 5405
rect 6637 5402 6703 5405
rect 8293 5402 8359 5405
rect 3693 5400 8359 5402
rect 3693 5344 3698 5400
rect 3754 5344 6642 5400
rect 6698 5344 8298 5400
rect 8354 5344 8359 5400
rect 3693 5342 8359 5344
rect 3693 5339 3759 5342
rect 6637 5339 6703 5342
rect 8293 5339 8359 5342
rect 9765 5402 9831 5405
rect 11605 5402 11671 5405
rect 9765 5400 11671 5402
rect 9765 5344 9770 5400
rect 9826 5344 11610 5400
rect 11666 5344 11671 5400
rect 9765 5342 11671 5344
rect 9765 5339 9831 5342
rect 11605 5339 11671 5342
rect 13353 5402 13419 5405
rect 14457 5402 14523 5405
rect 13353 5400 14523 5402
rect 13353 5344 13358 5400
rect 13414 5344 14462 5400
rect 14518 5344 14523 5400
rect 13353 5342 14523 5344
rect 13353 5339 13419 5342
rect 14457 5339 14523 5342
rect 0 5266 800 5296
rect 3417 5266 3483 5269
rect 0 5264 3483 5266
rect 0 5208 3422 5264
rect 3478 5208 3483 5264
rect 0 5206 3483 5208
rect 0 5176 800 5206
rect 3417 5203 3483 5206
rect 6269 5266 6335 5269
rect 7649 5266 7715 5269
rect 6269 5264 7715 5266
rect 6269 5208 6274 5264
rect 6330 5208 7654 5264
rect 7710 5208 7715 5264
rect 6269 5206 7715 5208
rect 6269 5203 6335 5206
rect 7649 5203 7715 5206
rect 7925 5266 7991 5269
rect 9768 5266 9828 5339
rect 15518 5269 15578 5475
rect 20646 5472 21042 5473
rect 20646 5408 20652 5472
rect 20716 5408 20732 5472
rect 20796 5408 20812 5472
rect 20876 5408 20892 5472
rect 20956 5408 20972 5472
rect 21036 5408 21042 5472
rect 20646 5407 21042 5408
rect 15929 5402 15995 5405
rect 19333 5402 19399 5405
rect 15929 5400 19399 5402
rect 15929 5344 15934 5400
rect 15990 5344 19338 5400
rect 19394 5344 19399 5400
rect 15929 5342 19399 5344
rect 15929 5339 15995 5342
rect 19333 5339 19399 5342
rect 19793 5402 19859 5405
rect 20478 5402 20484 5404
rect 19793 5400 20484 5402
rect 19793 5344 19798 5400
rect 19854 5344 20484 5400
rect 19793 5342 20484 5344
rect 19793 5339 19859 5342
rect 20478 5340 20484 5342
rect 20548 5340 20554 5404
rect 7925 5264 9828 5266
rect 7925 5208 7930 5264
rect 7986 5208 9828 5264
rect 7925 5206 9828 5208
rect 10685 5266 10751 5269
rect 12525 5266 12591 5269
rect 14825 5266 14891 5269
rect 10685 5264 14891 5266
rect 10685 5208 10690 5264
rect 10746 5208 12530 5264
rect 12586 5208 14830 5264
rect 14886 5208 14891 5264
rect 10685 5206 14891 5208
rect 15518 5264 15627 5269
rect 15518 5208 15566 5264
rect 15622 5208 15627 5264
rect 15518 5206 15627 5208
rect 7925 5203 7991 5206
rect 10685 5203 10751 5206
rect 12525 5203 12591 5206
rect 14825 5203 14891 5206
rect 15561 5203 15627 5206
rect 17125 5266 17191 5269
rect 21222 5266 21282 5478
rect 22093 5475 22159 5478
rect 23841 5475 23907 5478
rect 24485 5538 24551 5541
rect 25865 5538 25931 5541
rect 24485 5536 25931 5538
rect 24485 5480 24490 5536
rect 24546 5480 25870 5536
rect 25926 5480 25931 5536
rect 24485 5478 25931 5480
rect 24485 5475 24551 5478
rect 25865 5475 25931 5478
rect 26049 5538 26115 5541
rect 26049 5536 26572 5538
rect 26049 5480 26054 5536
rect 26110 5480 26572 5536
rect 26049 5478 26572 5480
rect 26049 5475 26115 5478
rect 26512 5405 26572 5478
rect 27654 5476 27660 5540
rect 27724 5538 27730 5540
rect 31753 5538 31819 5541
rect 32029 5538 32095 5541
rect 27724 5478 29930 5538
rect 27724 5476 27730 5478
rect 26646 5472 27042 5473
rect 26646 5408 26652 5472
rect 26716 5408 26732 5472
rect 26796 5408 26812 5472
rect 26876 5408 26892 5472
rect 26956 5408 26972 5472
rect 27036 5408 27042 5472
rect 26646 5407 27042 5408
rect 23841 5402 23907 5405
rect 25221 5402 25287 5405
rect 25957 5402 26023 5405
rect 23841 5400 26023 5402
rect 23841 5344 23846 5400
rect 23902 5344 25226 5400
rect 25282 5344 25962 5400
rect 26018 5344 26023 5400
rect 23841 5342 26023 5344
rect 23841 5339 23907 5342
rect 25221 5339 25287 5342
rect 25957 5339 26023 5342
rect 26509 5400 26575 5405
rect 28165 5402 28231 5405
rect 26509 5344 26514 5400
rect 26570 5344 26575 5400
rect 26509 5339 26575 5344
rect 27662 5400 28231 5402
rect 27662 5344 28170 5400
rect 28226 5344 28231 5400
rect 27662 5342 28231 5344
rect 17125 5264 21282 5266
rect 17125 5208 17130 5264
rect 17186 5208 21282 5264
rect 17125 5206 21282 5208
rect 21817 5266 21883 5269
rect 24117 5266 24183 5269
rect 21817 5264 24183 5266
rect 21817 5208 21822 5264
rect 21878 5208 24122 5264
rect 24178 5208 24183 5264
rect 21817 5206 24183 5208
rect 17125 5203 17191 5206
rect 21817 5203 21883 5206
rect 24117 5203 24183 5206
rect 24577 5266 24643 5269
rect 26693 5266 26759 5269
rect 24577 5264 26759 5266
rect 24577 5208 24582 5264
rect 24638 5208 26698 5264
rect 26754 5208 26759 5264
rect 24577 5206 26759 5208
rect 24577 5203 24643 5206
rect 26693 5203 26759 5206
rect 26969 5266 27035 5269
rect 27662 5266 27722 5342
rect 28165 5339 28231 5342
rect 28717 5402 28783 5405
rect 29870 5402 29930 5478
rect 31753 5536 32095 5538
rect 31753 5480 31758 5536
rect 31814 5480 32034 5536
rect 32090 5480 32095 5536
rect 31753 5478 32095 5480
rect 31753 5475 31819 5478
rect 32029 5475 32095 5478
rect 43069 5538 43135 5541
rect 44200 5538 45000 5568
rect 43069 5536 45000 5538
rect 43069 5480 43074 5536
rect 43130 5480 45000 5536
rect 43069 5478 45000 5480
rect 43069 5475 43135 5478
rect 32646 5472 33042 5473
rect 32646 5408 32652 5472
rect 32716 5408 32732 5472
rect 32796 5408 32812 5472
rect 32876 5408 32892 5472
rect 32956 5408 32972 5472
rect 33036 5408 33042 5472
rect 32646 5407 33042 5408
rect 38646 5472 39042 5473
rect 38646 5408 38652 5472
rect 38716 5408 38732 5472
rect 38796 5408 38812 5472
rect 38876 5408 38892 5472
rect 38956 5408 38972 5472
rect 39036 5408 39042 5472
rect 44200 5448 45000 5478
rect 38646 5407 39042 5408
rect 31753 5402 31819 5405
rect 28717 5400 29746 5402
rect 28717 5344 28722 5400
rect 28778 5344 29746 5400
rect 28717 5342 29746 5344
rect 29870 5400 31819 5402
rect 29870 5344 31758 5400
rect 31814 5344 31819 5400
rect 29870 5342 31819 5344
rect 28717 5339 28783 5342
rect 26969 5264 27722 5266
rect 26969 5208 26974 5264
rect 27030 5208 27722 5264
rect 26969 5206 27722 5208
rect 26969 5203 27035 5206
rect 27838 5204 27844 5268
rect 27908 5266 27914 5268
rect 29453 5266 29519 5269
rect 27908 5264 29519 5266
rect 27908 5208 29458 5264
rect 29514 5208 29519 5264
rect 27908 5206 29519 5208
rect 29686 5266 29746 5342
rect 31753 5339 31819 5342
rect 43253 5266 43319 5269
rect 29686 5264 43319 5266
rect 29686 5208 43258 5264
rect 43314 5208 43319 5264
rect 29686 5206 43319 5208
rect 27908 5204 27914 5206
rect 29453 5203 29519 5206
rect 43253 5203 43319 5206
rect 43437 5266 43503 5269
rect 44200 5266 45000 5296
rect 43437 5264 45000 5266
rect 43437 5208 43442 5264
rect 43498 5208 45000 5264
rect 43437 5206 45000 5208
rect 43437 5203 43503 5206
rect 44200 5176 45000 5206
rect 1761 5130 1827 5133
rect 5717 5130 5783 5133
rect 7557 5130 7623 5133
rect 1761 5128 7623 5130
rect 1761 5072 1766 5128
rect 1822 5072 5722 5128
rect 5778 5072 7562 5128
rect 7618 5072 7623 5128
rect 1761 5070 7623 5072
rect 1761 5067 1827 5070
rect 5717 5067 5783 5070
rect 7557 5067 7623 5070
rect 7741 5130 7807 5133
rect 9673 5130 9739 5133
rect 7741 5128 9739 5130
rect 7741 5072 7746 5128
rect 7802 5072 9678 5128
rect 9734 5072 9739 5128
rect 7741 5070 9739 5072
rect 7741 5067 7807 5070
rect 9673 5067 9739 5070
rect 10317 5130 10383 5133
rect 11053 5130 11119 5133
rect 10317 5128 11119 5130
rect 10317 5072 10322 5128
rect 10378 5072 11058 5128
rect 11114 5072 11119 5128
rect 10317 5070 11119 5072
rect 10317 5067 10383 5070
rect 11053 5067 11119 5070
rect 13077 5130 13143 5133
rect 20621 5130 20687 5133
rect 28073 5130 28139 5133
rect 13077 5128 20546 5130
rect 13077 5072 13082 5128
rect 13138 5072 20546 5128
rect 13077 5070 20546 5072
rect 13077 5067 13143 5070
rect 0 4994 800 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 800 4934
rect 1485 4931 1551 4934
rect 12341 4994 12407 4997
rect 13670 4994 13676 4996
rect 12341 4992 13676 4994
rect 12341 4936 12346 4992
rect 12402 4936 13676 4992
rect 12341 4934 13676 4936
rect 12341 4931 12407 4934
rect 13670 4932 13676 4934
rect 13740 4932 13746 4996
rect 14825 4994 14891 4997
rect 19701 4994 19767 4997
rect 14825 4992 19767 4994
rect 14825 4936 14830 4992
rect 14886 4936 19706 4992
rect 19762 4936 19767 4992
rect 14825 4934 19767 4936
rect 14825 4931 14891 4934
rect 19701 4931 19767 4934
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 13906 4928 14302 4929
rect 13906 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14302 4928
rect 13906 4863 14302 4864
rect 19906 4928 20302 4929
rect 19906 4864 19912 4928
rect 19976 4864 19992 4928
rect 20056 4864 20072 4928
rect 20136 4864 20152 4928
rect 20216 4864 20232 4928
rect 20296 4864 20302 4928
rect 19906 4863 20302 4864
rect 9029 4858 9095 4861
rect 9949 4858 10015 4861
rect 13629 4858 13695 4861
rect 9029 4856 13695 4858
rect 9029 4800 9034 4856
rect 9090 4800 9954 4856
rect 10010 4800 13634 4856
rect 13690 4800 13695 4856
rect 9029 4798 13695 4800
rect 9029 4795 9095 4798
rect 9949 4795 10015 4798
rect 13629 4795 13695 4798
rect 15142 4796 15148 4860
rect 15212 4858 15218 4860
rect 15377 4858 15443 4861
rect 15212 4856 15443 4858
rect 15212 4800 15382 4856
rect 15438 4800 15443 4856
rect 15212 4798 15443 4800
rect 15212 4796 15218 4798
rect 15377 4795 15443 4798
rect 17493 4858 17559 4861
rect 18321 4858 18387 4861
rect 17493 4856 18387 4858
rect 17493 4800 17498 4856
rect 17554 4800 18326 4856
rect 18382 4800 18387 4856
rect 17493 4798 18387 4800
rect 17493 4795 17559 4798
rect 18321 4795 18387 4798
rect 18505 4858 18571 4861
rect 19425 4858 19491 4861
rect 18505 4856 19491 4858
rect 18505 4800 18510 4856
rect 18566 4800 19430 4856
rect 19486 4800 19491 4856
rect 18505 4798 19491 4800
rect 20486 4858 20546 5070
rect 20621 5128 28139 5130
rect 20621 5072 20626 5128
rect 20682 5072 28078 5128
rect 28134 5072 28139 5128
rect 20621 5070 28139 5072
rect 20621 5067 20687 5070
rect 28073 5067 28139 5070
rect 29361 5130 29427 5133
rect 31477 5130 31543 5133
rect 38469 5130 38535 5133
rect 29361 5128 31543 5130
rect 29361 5072 29366 5128
rect 29422 5072 31482 5128
rect 31538 5072 31543 5128
rect 29361 5070 31543 5072
rect 29361 5067 29427 5070
rect 31477 5067 31543 5070
rect 31710 5128 38535 5130
rect 31710 5072 38474 5128
rect 38530 5072 38535 5128
rect 31710 5070 38535 5072
rect 20621 4994 20687 4997
rect 21725 4994 21791 4997
rect 20621 4992 21791 4994
rect 20621 4936 20626 4992
rect 20682 4936 21730 4992
rect 21786 4936 21791 4992
rect 20621 4934 21791 4936
rect 20621 4931 20687 4934
rect 21725 4931 21791 4934
rect 22001 4994 22067 4997
rect 23565 4994 23631 4997
rect 22001 4992 23631 4994
rect 22001 4936 22006 4992
rect 22062 4936 23570 4992
rect 23626 4936 23631 4992
rect 22001 4934 23631 4936
rect 22001 4931 22067 4934
rect 23565 4931 23631 4934
rect 26366 4932 26372 4996
rect 26436 4994 26442 4996
rect 30925 4994 30991 4997
rect 26436 4992 30991 4994
rect 26436 4936 30930 4992
rect 30986 4936 30991 4992
rect 26436 4934 30991 4936
rect 26436 4932 26442 4934
rect 30925 4931 30991 4934
rect 25906 4928 26302 4929
rect 25906 4864 25912 4928
rect 25976 4864 25992 4928
rect 26056 4864 26072 4928
rect 26136 4864 26152 4928
rect 26216 4864 26232 4928
rect 26296 4864 26302 4928
rect 25906 4863 26302 4864
rect 25129 4858 25195 4861
rect 20486 4856 25195 4858
rect 20486 4800 25134 4856
rect 25190 4800 25195 4856
rect 20486 4798 25195 4800
rect 18505 4795 18571 4798
rect 19425 4795 19491 4798
rect 25129 4795 25195 4798
rect 26601 4858 26667 4861
rect 27337 4858 27403 4861
rect 31710 4858 31770 5070
rect 38469 5067 38535 5070
rect 32489 4994 32555 4997
rect 34421 4994 34487 4997
rect 32489 4992 34487 4994
rect 32489 4936 32494 4992
rect 32550 4936 34426 4992
rect 34482 4936 34487 4992
rect 32489 4934 34487 4936
rect 32489 4931 32555 4934
rect 34421 4931 34487 4934
rect 43069 4994 43135 4997
rect 44200 4994 45000 5024
rect 43069 4992 45000 4994
rect 43069 4936 43074 4992
rect 43130 4936 45000 4992
rect 43069 4934 45000 4936
rect 43069 4931 43135 4934
rect 31906 4928 32302 4929
rect 31906 4864 31912 4928
rect 31976 4864 31992 4928
rect 32056 4864 32072 4928
rect 32136 4864 32152 4928
rect 32216 4864 32232 4928
rect 32296 4864 32302 4928
rect 31906 4863 32302 4864
rect 37906 4928 38302 4929
rect 37906 4864 37912 4928
rect 37976 4864 37992 4928
rect 38056 4864 38072 4928
rect 38136 4864 38152 4928
rect 38216 4864 38232 4928
rect 38296 4864 38302 4928
rect 44200 4904 45000 4934
rect 37906 4863 38302 4864
rect 26601 4856 27403 4858
rect 26601 4800 26606 4856
rect 26662 4800 27342 4856
rect 27398 4800 27403 4856
rect 26601 4798 27403 4800
rect 26601 4795 26667 4798
rect 27337 4795 27403 4798
rect 27846 4798 31770 4858
rect 32397 4856 32463 4861
rect 35065 4860 35131 4861
rect 32397 4800 32402 4856
rect 32458 4800 32463 4856
rect 0 4722 800 4752
rect 1853 4722 1919 4725
rect 0 4720 1919 4722
rect 0 4664 1858 4720
rect 1914 4664 1919 4720
rect 0 4662 1919 4664
rect 0 4632 800 4662
rect 1853 4659 1919 4662
rect 6177 4722 6243 4725
rect 10685 4722 10751 4725
rect 6177 4720 10751 4722
rect 6177 4664 6182 4720
rect 6238 4664 10690 4720
rect 10746 4664 10751 4720
rect 6177 4662 10751 4664
rect 6177 4659 6243 4662
rect 10685 4659 10751 4662
rect 12065 4722 12131 4725
rect 25957 4722 26023 4725
rect 27613 4722 27679 4725
rect 12065 4720 27679 4722
rect 12065 4664 12070 4720
rect 12126 4664 25962 4720
rect 26018 4664 27618 4720
rect 27674 4664 27679 4720
rect 12065 4662 27679 4664
rect 12065 4659 12131 4662
rect 25957 4659 26023 4662
rect 27613 4659 27679 4662
rect 2037 4586 2103 4589
rect 14089 4586 14155 4589
rect 2037 4584 14155 4586
rect 2037 4528 2042 4584
rect 2098 4528 14094 4584
rect 14150 4528 14155 4584
rect 2037 4526 14155 4528
rect 2037 4523 2103 4526
rect 14089 4523 14155 4526
rect 14273 4586 14339 4589
rect 17769 4586 17835 4589
rect 14273 4584 17835 4586
rect 14273 4528 14278 4584
rect 14334 4528 17774 4584
rect 17830 4528 17835 4584
rect 14273 4526 17835 4528
rect 14273 4523 14339 4526
rect 17769 4523 17835 4526
rect 18229 4586 18295 4589
rect 21449 4586 21515 4589
rect 18229 4584 21515 4586
rect 18229 4528 18234 4584
rect 18290 4528 21454 4584
rect 21510 4528 21515 4584
rect 18229 4526 21515 4528
rect 18229 4523 18295 4526
rect 21449 4523 21515 4526
rect 23749 4586 23815 4589
rect 27846 4586 27906 4798
rect 32397 4795 32463 4800
rect 35014 4796 35020 4860
rect 35084 4858 35131 4860
rect 35084 4856 35176 4858
rect 35126 4800 35176 4856
rect 35084 4798 35176 4800
rect 35084 4796 35131 4798
rect 35065 4795 35131 4796
rect 28022 4660 28028 4724
rect 28092 4722 28098 4724
rect 28257 4722 28323 4725
rect 28092 4720 28323 4722
rect 28092 4664 28262 4720
rect 28318 4664 28323 4720
rect 28092 4662 28323 4664
rect 28092 4660 28098 4662
rect 28257 4659 28323 4662
rect 28533 4722 28599 4725
rect 32400 4722 32460 4795
rect 28533 4720 32460 4722
rect 28533 4664 28538 4720
rect 28594 4664 32460 4720
rect 28533 4662 32460 4664
rect 32949 4722 33015 4725
rect 36353 4722 36419 4725
rect 32949 4720 36419 4722
rect 32949 4664 32954 4720
rect 33010 4664 36358 4720
rect 36414 4664 36419 4720
rect 32949 4662 36419 4664
rect 28533 4659 28599 4662
rect 32949 4659 33015 4662
rect 36353 4659 36419 4662
rect 36629 4722 36695 4725
rect 38285 4722 38351 4725
rect 43253 4722 43319 4725
rect 36629 4720 38351 4722
rect 36629 4664 36634 4720
rect 36690 4664 38290 4720
rect 38346 4664 38351 4720
rect 36629 4662 38351 4664
rect 36629 4659 36695 4662
rect 38285 4659 38351 4662
rect 41370 4720 43319 4722
rect 41370 4664 43258 4720
rect 43314 4664 43319 4720
rect 41370 4662 43319 4664
rect 23749 4584 27906 4586
rect 23749 4528 23754 4584
rect 23810 4528 27906 4584
rect 23749 4526 27906 4528
rect 29177 4586 29243 4589
rect 31293 4586 31359 4589
rect 41370 4586 41430 4662
rect 43253 4659 43319 4662
rect 43437 4722 43503 4725
rect 44200 4722 45000 4752
rect 43437 4720 45000 4722
rect 43437 4664 43442 4720
rect 43498 4664 45000 4720
rect 43437 4662 45000 4664
rect 43437 4659 43503 4662
rect 44200 4632 45000 4662
rect 29177 4584 31359 4586
rect 29177 4528 29182 4584
rect 29238 4528 31298 4584
rect 31354 4528 31359 4584
rect 29177 4526 31359 4528
rect 23749 4523 23815 4526
rect 29177 4523 29243 4526
rect 31293 4523 31359 4526
rect 31710 4526 41430 4586
rect 0 4450 800 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 800 4390
rect 1393 4387 1459 4390
rect 5073 4450 5139 4453
rect 6269 4450 6335 4453
rect 5073 4448 6335 4450
rect 5073 4392 5078 4448
rect 5134 4392 6274 4448
rect 6330 4392 6335 4448
rect 5073 4390 6335 4392
rect 5073 4387 5139 4390
rect 6269 4387 6335 4390
rect 9949 4450 10015 4453
rect 13077 4450 13143 4453
rect 9949 4448 13143 4450
rect 9949 4392 9954 4448
rect 10010 4392 13082 4448
rect 13138 4392 13143 4448
rect 9949 4390 13143 4392
rect 9949 4387 10015 4390
rect 13077 4387 13143 4390
rect 13486 4388 13492 4452
rect 13556 4450 13562 4452
rect 13997 4450 14063 4453
rect 13556 4448 14063 4450
rect 13556 4392 14002 4448
rect 14058 4392 14063 4448
rect 13556 4390 14063 4392
rect 13556 4388 13562 4390
rect 13997 4387 14063 4390
rect 16849 4450 16915 4453
rect 18597 4450 18663 4453
rect 18965 4450 19031 4453
rect 16849 4448 19031 4450
rect 16849 4392 16854 4448
rect 16910 4392 18602 4448
rect 18658 4392 18970 4448
rect 19026 4392 19031 4448
rect 16849 4390 19031 4392
rect 16849 4387 16915 4390
rect 18597 4387 18663 4390
rect 18965 4387 19031 4390
rect 24025 4450 24091 4453
rect 26366 4450 26372 4452
rect 24025 4448 26372 4450
rect 24025 4392 24030 4448
rect 24086 4392 26372 4448
rect 24025 4390 26372 4392
rect 24025 4387 24091 4390
rect 26366 4388 26372 4390
rect 26436 4388 26442 4452
rect 2646 4384 3042 4385
rect 2646 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3042 4384
rect 2646 4319 3042 4320
rect 8646 4384 9042 4385
rect 8646 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9042 4384
rect 8646 4319 9042 4320
rect 14646 4384 15042 4385
rect 14646 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15042 4384
rect 14646 4319 15042 4320
rect 20646 4384 21042 4385
rect 20646 4320 20652 4384
rect 20716 4320 20732 4384
rect 20796 4320 20812 4384
rect 20876 4320 20892 4384
rect 20956 4320 20972 4384
rect 21036 4320 21042 4384
rect 20646 4319 21042 4320
rect 26646 4384 27042 4385
rect 26646 4320 26652 4384
rect 26716 4320 26732 4384
rect 26796 4320 26812 4384
rect 26876 4320 26892 4384
rect 26956 4320 26972 4384
rect 27036 4320 27042 4384
rect 26646 4319 27042 4320
rect 9397 4314 9463 4317
rect 12433 4314 12499 4317
rect 14273 4314 14339 4317
rect 9397 4312 12499 4314
rect 9397 4256 9402 4312
rect 9458 4256 12438 4312
rect 12494 4256 12499 4312
rect 9397 4254 12499 4256
rect 9397 4251 9463 4254
rect 12433 4251 12499 4254
rect 13494 4312 14339 4314
rect 13494 4256 14278 4312
rect 14334 4256 14339 4312
rect 13494 4254 14339 4256
rect 0 4178 800 4208
rect 2221 4178 2287 4181
rect 0 4176 2287 4178
rect 0 4120 2226 4176
rect 2282 4120 2287 4176
rect 0 4118 2287 4120
rect 0 4088 800 4118
rect 2221 4115 2287 4118
rect 8385 4178 8451 4181
rect 13494 4178 13554 4254
rect 14273 4251 14339 4254
rect 16297 4314 16363 4317
rect 17769 4314 17835 4317
rect 16297 4312 17835 4314
rect 16297 4256 16302 4312
rect 16358 4256 17774 4312
rect 17830 4256 17835 4312
rect 16297 4254 17835 4256
rect 16297 4251 16363 4254
rect 17769 4251 17835 4254
rect 17902 4252 17908 4316
rect 17972 4314 17978 4316
rect 19333 4314 19399 4317
rect 17972 4312 19399 4314
rect 17972 4256 19338 4312
rect 19394 4256 19399 4312
rect 17972 4254 19399 4256
rect 17972 4252 17978 4254
rect 19333 4251 19399 4254
rect 21173 4316 21239 4317
rect 21173 4312 21220 4316
rect 21284 4314 21290 4316
rect 21541 4314 21607 4317
rect 22553 4314 22619 4317
rect 25865 4314 25931 4317
rect 31710 4314 31770 4526
rect 43069 4450 43135 4453
rect 44200 4450 45000 4480
rect 43069 4448 45000 4450
rect 43069 4392 43074 4448
rect 43130 4392 45000 4448
rect 43069 4390 45000 4392
rect 43069 4387 43135 4390
rect 32646 4384 33042 4385
rect 32646 4320 32652 4384
rect 32716 4320 32732 4384
rect 32796 4320 32812 4384
rect 32876 4320 32892 4384
rect 32956 4320 32972 4384
rect 33036 4320 33042 4384
rect 32646 4319 33042 4320
rect 38646 4384 39042 4385
rect 38646 4320 38652 4384
rect 38716 4320 38732 4384
rect 38796 4320 38812 4384
rect 38876 4320 38892 4384
rect 38956 4320 38972 4384
rect 39036 4320 39042 4384
rect 44200 4360 45000 4390
rect 38646 4319 39042 4320
rect 21173 4256 21178 4312
rect 21173 4252 21220 4256
rect 21284 4254 21330 4314
rect 21541 4312 25931 4314
rect 21541 4256 21546 4312
rect 21602 4256 22558 4312
rect 22614 4256 25870 4312
rect 25926 4256 25931 4312
rect 21541 4254 25931 4256
rect 21284 4252 21290 4254
rect 21173 4251 21239 4252
rect 21541 4251 21607 4254
rect 22553 4251 22619 4254
rect 25865 4251 25931 4254
rect 30422 4254 31770 4314
rect 8385 4176 13554 4178
rect 8385 4120 8390 4176
rect 8446 4120 13554 4176
rect 8385 4118 13554 4120
rect 13905 4178 13971 4181
rect 18873 4178 18939 4181
rect 13905 4176 18939 4178
rect 13905 4120 13910 4176
rect 13966 4120 18878 4176
rect 18934 4120 18939 4176
rect 13905 4118 18939 4120
rect 8385 4115 8451 4118
rect 13905 4115 13971 4118
rect 18873 4115 18939 4118
rect 19885 4178 19951 4181
rect 21766 4178 21772 4180
rect 19885 4176 21772 4178
rect 19885 4120 19890 4176
rect 19946 4120 21772 4176
rect 19885 4118 21772 4120
rect 19885 4115 19951 4118
rect 21766 4116 21772 4118
rect 21836 4116 21842 4180
rect 24577 4178 24643 4181
rect 28533 4178 28599 4181
rect 24577 4176 28599 4178
rect 24577 4120 24582 4176
rect 24638 4120 28538 4176
rect 28594 4120 28599 4176
rect 24577 4118 28599 4120
rect 24577 4115 24643 4118
rect 28533 4115 28599 4118
rect 7833 4042 7899 4045
rect 13261 4042 13327 4045
rect 14641 4042 14707 4045
rect 26325 4042 26391 4045
rect 7833 4040 14428 4042
rect 7833 3984 7838 4040
rect 7894 3984 13266 4040
rect 13322 3984 14428 4040
rect 7833 3982 14428 3984
rect 7833 3979 7899 3982
rect 13261 3979 13327 3982
rect 0 3906 800 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 800 3846
rect 1485 3843 1551 3846
rect 9765 3906 9831 3909
rect 10869 3906 10935 3909
rect 9765 3904 10935 3906
rect 9765 3848 9770 3904
rect 9826 3848 10874 3904
rect 10930 3848 10935 3904
rect 9765 3846 10935 3848
rect 9765 3843 9831 3846
rect 10869 3843 10935 3846
rect 13353 3906 13419 3909
rect 13629 3906 13695 3909
rect 13353 3904 13695 3906
rect 13353 3848 13358 3904
rect 13414 3848 13634 3904
rect 13690 3848 13695 3904
rect 13353 3846 13695 3848
rect 13353 3843 13419 3846
rect 13629 3843 13695 3846
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 13906 3840 14302 3841
rect 13906 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14302 3840
rect 13906 3775 14302 3776
rect 8937 3770 9003 3773
rect 10409 3770 10475 3773
rect 8937 3768 10475 3770
rect 8937 3712 8942 3768
rect 8998 3712 10414 3768
rect 10470 3712 10475 3768
rect 8937 3710 10475 3712
rect 8937 3707 9003 3710
rect 10409 3707 10475 3710
rect 11605 3770 11671 3773
rect 13261 3770 13327 3773
rect 11605 3768 13327 3770
rect 11605 3712 11610 3768
rect 11666 3712 13266 3768
rect 13322 3712 13327 3768
rect 11605 3710 13327 3712
rect 14368 3770 14428 3982
rect 14641 4040 26391 4042
rect 14641 3984 14646 4040
rect 14702 3984 26330 4040
rect 26386 3984 26391 4040
rect 14641 3982 26391 3984
rect 14641 3979 14707 3982
rect 26325 3979 26391 3982
rect 26509 4042 26575 4045
rect 30422 4042 30482 4254
rect 30925 4178 30991 4181
rect 32581 4178 32647 4181
rect 30925 4176 32647 4178
rect 30925 4120 30930 4176
rect 30986 4120 32586 4176
rect 32642 4120 32647 4176
rect 30925 4118 32647 4120
rect 30925 4115 30991 4118
rect 32581 4115 32647 4118
rect 33409 4178 33475 4181
rect 34237 4178 34303 4181
rect 35341 4178 35407 4181
rect 33409 4176 35407 4178
rect 33409 4120 33414 4176
rect 33470 4120 34242 4176
rect 34298 4120 35346 4176
rect 35402 4120 35407 4176
rect 33409 4118 35407 4120
rect 33409 4115 33475 4118
rect 34237 4115 34303 4118
rect 35341 4115 35407 4118
rect 43437 4178 43503 4181
rect 44200 4178 45000 4208
rect 43437 4176 45000 4178
rect 43437 4120 43442 4176
rect 43498 4120 45000 4176
rect 43437 4118 45000 4120
rect 43437 4115 43503 4118
rect 44200 4088 45000 4118
rect 35249 4042 35315 4045
rect 26509 4040 30482 4042
rect 26509 3984 26514 4040
rect 26570 3984 30482 4040
rect 26509 3982 30482 3984
rect 31756 4040 35315 4042
rect 31756 3984 35254 4040
rect 35310 3984 35315 4040
rect 31756 3982 35315 3984
rect 26509 3979 26575 3982
rect 17309 3906 17375 3909
rect 19425 3906 19491 3909
rect 17309 3904 19491 3906
rect 17309 3848 17314 3904
rect 17370 3848 19430 3904
rect 19486 3848 19491 3904
rect 17309 3846 19491 3848
rect 17309 3843 17375 3846
rect 19425 3843 19491 3846
rect 20529 3906 20595 3909
rect 23197 3906 23263 3909
rect 20529 3904 23263 3906
rect 20529 3848 20534 3904
rect 20590 3848 23202 3904
rect 23258 3848 23263 3904
rect 20529 3846 23263 3848
rect 20529 3843 20595 3846
rect 23197 3843 23263 3846
rect 26601 3906 26667 3909
rect 27153 3906 27219 3909
rect 31756 3906 31816 3982
rect 35249 3979 35315 3982
rect 26601 3904 31816 3906
rect 26601 3848 26606 3904
rect 26662 3848 27158 3904
rect 27214 3848 31816 3904
rect 26601 3846 31816 3848
rect 32765 3906 32831 3909
rect 33501 3906 33567 3909
rect 33961 3908 34027 3909
rect 33910 3906 33916 3908
rect 32765 3904 33567 3906
rect 32765 3848 32770 3904
rect 32826 3848 33506 3904
rect 33562 3848 33567 3904
rect 32765 3846 33567 3848
rect 33870 3846 33916 3906
rect 33980 3904 34027 3908
rect 34022 3848 34027 3904
rect 26601 3843 26667 3846
rect 27153 3843 27219 3846
rect 32765 3843 32831 3846
rect 33501 3843 33567 3846
rect 33910 3844 33916 3846
rect 33980 3844 34027 3848
rect 33961 3843 34027 3844
rect 43069 3906 43135 3909
rect 44200 3906 45000 3936
rect 43069 3904 45000 3906
rect 43069 3848 43074 3904
rect 43130 3848 45000 3904
rect 43069 3846 45000 3848
rect 43069 3843 43135 3846
rect 19906 3840 20302 3841
rect 19906 3776 19912 3840
rect 19976 3776 19992 3840
rect 20056 3776 20072 3840
rect 20136 3776 20152 3840
rect 20216 3776 20232 3840
rect 20296 3776 20302 3840
rect 19906 3775 20302 3776
rect 25906 3840 26302 3841
rect 25906 3776 25912 3840
rect 25976 3776 25992 3840
rect 26056 3776 26072 3840
rect 26136 3776 26152 3840
rect 26216 3776 26232 3840
rect 26296 3776 26302 3840
rect 25906 3775 26302 3776
rect 31906 3840 32302 3841
rect 31906 3776 31912 3840
rect 31976 3776 31992 3840
rect 32056 3776 32072 3840
rect 32136 3776 32152 3840
rect 32216 3776 32232 3840
rect 32296 3776 32302 3840
rect 31906 3775 32302 3776
rect 37906 3840 38302 3841
rect 37906 3776 37912 3840
rect 37976 3776 37992 3840
rect 38056 3776 38072 3840
rect 38136 3776 38152 3840
rect 38216 3776 38232 3840
rect 38296 3776 38302 3840
rect 44200 3816 45000 3846
rect 37906 3775 38302 3776
rect 15326 3770 15332 3772
rect 14368 3710 15332 3770
rect 11605 3707 11671 3710
rect 13261 3707 13327 3710
rect 15326 3708 15332 3710
rect 15396 3708 15402 3772
rect 15510 3708 15516 3772
rect 15580 3770 15586 3772
rect 18137 3770 18203 3773
rect 25589 3770 25655 3773
rect 15580 3768 18203 3770
rect 15580 3712 18142 3768
rect 18198 3712 18203 3768
rect 15580 3710 18203 3712
rect 15580 3708 15586 3710
rect 18137 3707 18203 3710
rect 20532 3768 25655 3770
rect 20532 3712 25594 3768
rect 25650 3712 25655 3768
rect 20532 3710 25655 3712
rect 0 3634 800 3664
rect 1577 3634 1643 3637
rect 0 3632 1643 3634
rect 0 3576 1582 3632
rect 1638 3576 1643 3632
rect 0 3574 1643 3576
rect 0 3544 800 3574
rect 1577 3571 1643 3574
rect 2497 3634 2563 3637
rect 9121 3634 9187 3637
rect 2497 3632 9187 3634
rect 2497 3576 2502 3632
rect 2558 3576 9126 3632
rect 9182 3576 9187 3632
rect 2497 3574 9187 3576
rect 2497 3571 2563 3574
rect 9121 3571 9187 3574
rect 9857 3634 9923 3637
rect 19057 3634 19123 3637
rect 20532 3634 20592 3710
rect 25589 3707 25655 3710
rect 26417 3770 26483 3773
rect 26877 3770 26943 3773
rect 26417 3768 26943 3770
rect 26417 3712 26422 3768
rect 26478 3712 26882 3768
rect 26938 3712 26943 3768
rect 26417 3710 26943 3712
rect 26417 3707 26483 3710
rect 26877 3707 26943 3710
rect 28901 3770 28967 3773
rect 32581 3770 32647 3773
rect 34329 3770 34395 3773
rect 28901 3768 31770 3770
rect 28901 3712 28906 3768
rect 28962 3712 31770 3768
rect 28901 3710 31770 3712
rect 28901 3707 28967 3710
rect 22093 3634 22159 3637
rect 9857 3632 18890 3634
rect 9857 3576 9862 3632
rect 9918 3576 18890 3632
rect 9857 3574 18890 3576
rect 9857 3571 9923 3574
rect 6821 3498 6887 3501
rect 12617 3498 12683 3501
rect 13353 3498 13419 3501
rect 18830 3498 18890 3574
rect 19057 3632 20592 3634
rect 19057 3576 19062 3632
rect 19118 3576 20592 3632
rect 19057 3574 20592 3576
rect 20670 3632 22159 3634
rect 20670 3576 22098 3632
rect 22154 3576 22159 3632
rect 20670 3574 22159 3576
rect 19057 3571 19123 3574
rect 19885 3498 19951 3501
rect 20670 3498 20730 3574
rect 22093 3571 22159 3574
rect 23197 3634 23263 3637
rect 24761 3634 24827 3637
rect 28165 3634 28231 3637
rect 23197 3632 28231 3634
rect 23197 3576 23202 3632
rect 23258 3576 24766 3632
rect 24822 3576 28170 3632
rect 28226 3576 28231 3632
rect 23197 3574 28231 3576
rect 23197 3571 23263 3574
rect 24761 3571 24827 3574
rect 28165 3571 28231 3574
rect 28441 3634 28507 3637
rect 31710 3634 31770 3710
rect 32581 3768 34395 3770
rect 32581 3712 32586 3768
rect 32642 3712 34334 3768
rect 34390 3712 34395 3768
rect 32581 3710 34395 3712
rect 32581 3707 32647 3710
rect 34329 3707 34395 3710
rect 32949 3634 33015 3637
rect 28441 3632 30114 3634
rect 28441 3576 28446 3632
rect 28502 3576 30114 3632
rect 28441 3574 30114 3576
rect 31710 3632 33015 3634
rect 31710 3576 32954 3632
rect 33010 3576 33015 3632
rect 31710 3574 33015 3576
rect 28441 3571 28507 3574
rect 6821 3496 15210 3498
rect 6821 3440 6826 3496
rect 6882 3440 12622 3496
rect 12678 3440 13358 3496
rect 13414 3440 15210 3496
rect 6821 3438 15210 3440
rect 18830 3496 19951 3498
rect 18830 3440 19890 3496
rect 19946 3440 19951 3496
rect 18830 3438 19951 3440
rect 6821 3435 6887 3438
rect 12617 3435 12683 3438
rect 13353 3435 13419 3438
rect 0 3362 800 3392
rect 1853 3362 1919 3365
rect 0 3360 1919 3362
rect 0 3304 1858 3360
rect 1914 3304 1919 3360
rect 0 3302 1919 3304
rect 0 3272 800 3302
rect 1853 3299 1919 3302
rect 5809 3362 5875 3365
rect 8293 3362 8359 3365
rect 5809 3360 8359 3362
rect 5809 3304 5814 3360
rect 5870 3304 8298 3360
rect 8354 3304 8359 3360
rect 5809 3302 8359 3304
rect 5809 3299 5875 3302
rect 8293 3299 8359 3302
rect 9121 3362 9187 3365
rect 13813 3362 13879 3365
rect 9121 3360 13879 3362
rect 9121 3304 9126 3360
rect 9182 3304 13818 3360
rect 13874 3304 13879 3360
rect 9121 3302 13879 3304
rect 15150 3362 15210 3438
rect 19885 3435 19951 3438
rect 20118 3438 20730 3498
rect 21449 3498 21515 3501
rect 21582 3498 21588 3500
rect 21449 3496 21588 3498
rect 21449 3440 21454 3496
rect 21510 3440 21588 3496
rect 21449 3438 21588 3440
rect 20118 3362 20178 3438
rect 21449 3435 21515 3438
rect 21582 3436 21588 3438
rect 21652 3436 21658 3500
rect 30054 3498 30114 3574
rect 32949 3571 33015 3574
rect 43437 3634 43503 3637
rect 44200 3634 45000 3664
rect 43437 3632 45000 3634
rect 43437 3576 43442 3632
rect 43498 3576 45000 3632
rect 43437 3574 45000 3576
rect 43437 3571 43503 3574
rect 44200 3544 45000 3574
rect 35433 3498 35499 3501
rect 35893 3498 35959 3501
rect 22050 3438 29010 3498
rect 30054 3496 35959 3498
rect 30054 3440 35438 3496
rect 35494 3440 35898 3496
rect 35954 3440 35959 3496
rect 30054 3438 35959 3440
rect 15150 3302 20178 3362
rect 9121 3299 9187 3302
rect 13813 3299 13879 3302
rect 2646 3296 3042 3297
rect 2646 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3042 3296
rect 2646 3231 3042 3232
rect 8646 3296 9042 3297
rect 8646 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9042 3296
rect 8646 3231 9042 3232
rect 14646 3296 15042 3297
rect 14646 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15042 3296
rect 14646 3231 15042 3232
rect 20646 3296 21042 3297
rect 20646 3232 20652 3296
rect 20716 3232 20732 3296
rect 20796 3232 20812 3296
rect 20876 3232 20892 3296
rect 20956 3232 20972 3296
rect 21036 3232 21042 3296
rect 20646 3231 21042 3232
rect 2221 3226 2287 3229
rect 1166 3224 2287 3226
rect 1166 3168 2226 3224
rect 2282 3168 2287 3224
rect 1166 3166 2287 3168
rect 0 3090 800 3120
rect 1166 3090 1226 3166
rect 2221 3163 2287 3166
rect 9121 3226 9187 3229
rect 12249 3226 12315 3229
rect 14181 3226 14247 3229
rect 9121 3224 10794 3226
rect 9121 3168 9126 3224
rect 9182 3168 10794 3224
rect 9121 3166 10794 3168
rect 9121 3163 9187 3166
rect 2773 3090 2839 3093
rect 0 3030 1226 3090
rect 1396 3088 2839 3090
rect 1396 3032 2778 3088
rect 2834 3032 2839 3088
rect 1396 3030 2839 3032
rect 0 3000 800 3030
rect 0 2818 800 2848
rect 1396 2818 1456 3030
rect 2773 3027 2839 3030
rect 3509 3090 3575 3093
rect 9857 3090 9923 3093
rect 3509 3088 9923 3090
rect 3509 3032 3514 3088
rect 3570 3032 9862 3088
rect 9918 3032 9923 3088
rect 3509 3030 9923 3032
rect 10734 3090 10794 3166
rect 12249 3224 14247 3226
rect 12249 3168 12254 3224
rect 12310 3168 14186 3224
rect 14242 3168 14247 3224
rect 12249 3166 14247 3168
rect 12249 3163 12315 3166
rect 14181 3163 14247 3166
rect 16849 3226 16915 3229
rect 16982 3226 16988 3228
rect 16849 3224 16988 3226
rect 16849 3168 16854 3224
rect 16910 3168 16988 3224
rect 16849 3166 16988 3168
rect 16849 3163 16915 3166
rect 16982 3164 16988 3166
rect 17052 3164 17058 3228
rect 17217 3226 17283 3229
rect 17350 3226 17356 3228
rect 17217 3224 17356 3226
rect 17217 3168 17222 3224
rect 17278 3168 17356 3224
rect 17217 3166 17356 3168
rect 17217 3163 17283 3166
rect 17350 3164 17356 3166
rect 17420 3164 17426 3228
rect 19006 3164 19012 3228
rect 19076 3226 19082 3228
rect 19149 3226 19215 3229
rect 22050 3226 22110 3438
rect 28950 3362 29010 3438
rect 35433 3435 35499 3438
rect 35893 3435 35959 3438
rect 40953 3498 41019 3501
rect 43253 3498 43319 3501
rect 40953 3496 43319 3498
rect 40953 3440 40958 3496
rect 41014 3440 43258 3496
rect 43314 3440 43319 3496
rect 40953 3438 43319 3440
rect 40953 3435 41019 3438
rect 43253 3435 43319 3438
rect 30097 3362 30163 3365
rect 28950 3360 30163 3362
rect 28950 3304 30102 3360
rect 30158 3304 30163 3360
rect 28950 3302 30163 3304
rect 30097 3299 30163 3302
rect 43069 3362 43135 3365
rect 44200 3362 45000 3392
rect 43069 3360 45000 3362
rect 43069 3304 43074 3360
rect 43130 3304 45000 3360
rect 43069 3302 45000 3304
rect 43069 3299 43135 3302
rect 26646 3296 27042 3297
rect 26646 3232 26652 3296
rect 26716 3232 26732 3296
rect 26796 3232 26812 3296
rect 26876 3232 26892 3296
rect 26956 3232 26972 3296
rect 27036 3232 27042 3296
rect 26646 3231 27042 3232
rect 32646 3296 33042 3297
rect 32646 3232 32652 3296
rect 32716 3232 32732 3296
rect 32796 3232 32812 3296
rect 32876 3232 32892 3296
rect 32956 3232 32972 3296
rect 33036 3232 33042 3296
rect 32646 3231 33042 3232
rect 38646 3296 39042 3297
rect 38646 3232 38652 3296
rect 38716 3232 38732 3296
rect 38796 3232 38812 3296
rect 38876 3232 38892 3296
rect 38956 3232 38972 3296
rect 39036 3232 39042 3296
rect 44200 3272 45000 3302
rect 38646 3231 39042 3232
rect 32397 3228 32463 3229
rect 32397 3226 32444 3228
rect 19076 3224 19215 3226
rect 19076 3168 19154 3224
rect 19210 3168 19215 3224
rect 19076 3166 19215 3168
rect 19076 3164 19082 3166
rect 19149 3163 19215 3166
rect 21222 3166 22110 3226
rect 32352 3224 32444 3226
rect 32352 3168 32402 3224
rect 32352 3166 32444 3168
rect 13077 3090 13143 3093
rect 10734 3088 13143 3090
rect 10734 3032 13082 3088
rect 13138 3032 13143 3088
rect 10734 3030 13143 3032
rect 3509 3027 3575 3030
rect 9857 3027 9923 3030
rect 13077 3027 13143 3030
rect 13261 3090 13327 3093
rect 14273 3090 14339 3093
rect 13261 3088 14339 3090
rect 13261 3032 13266 3088
rect 13322 3032 14278 3088
rect 14334 3032 14339 3088
rect 13261 3030 14339 3032
rect 13261 3027 13327 3030
rect 14273 3027 14339 3030
rect 14457 3090 14523 3093
rect 21222 3090 21282 3166
rect 32397 3164 32444 3166
rect 32508 3164 32514 3228
rect 32397 3163 32463 3164
rect 24117 3090 24183 3093
rect 30741 3090 30807 3093
rect 14457 3088 21282 3090
rect 14457 3032 14462 3088
rect 14518 3032 21282 3088
rect 14457 3030 21282 3032
rect 22050 3088 30807 3090
rect 22050 3032 24122 3088
rect 24178 3032 30746 3088
rect 30802 3032 30807 3088
rect 22050 3030 30807 3032
rect 14457 3027 14523 3030
rect 2497 2954 2563 2957
rect 7925 2954 7991 2957
rect 8661 2954 8727 2957
rect 9438 2954 9444 2956
rect 2497 2952 7666 2954
rect 2497 2896 2502 2952
rect 2558 2896 7666 2952
rect 2497 2894 7666 2896
rect 2497 2891 2563 2894
rect 0 2758 1456 2818
rect 0 2728 800 2758
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 7606 2546 7666 2894
rect 7925 2952 8586 2954
rect 7925 2896 7930 2952
rect 7986 2896 8586 2952
rect 7925 2894 8586 2896
rect 7925 2891 7991 2894
rect 8526 2818 8586 2894
rect 8661 2952 9444 2954
rect 8661 2896 8666 2952
rect 8722 2896 9444 2952
rect 8661 2894 9444 2896
rect 8661 2891 8727 2894
rect 9438 2892 9444 2894
rect 9508 2954 9514 2956
rect 10685 2954 10751 2957
rect 9508 2952 10751 2954
rect 9508 2896 10690 2952
rect 10746 2896 10751 2952
rect 9508 2894 10751 2896
rect 9508 2892 9514 2894
rect 10685 2891 10751 2894
rect 10910 2892 10916 2956
rect 10980 2954 10986 2956
rect 18413 2954 18479 2957
rect 22050 2954 22110 3030
rect 24117 3027 24183 3030
rect 30741 3027 30807 3030
rect 32305 3090 32371 3093
rect 34697 3090 34763 3093
rect 32305 3088 34763 3090
rect 32305 3032 32310 3088
rect 32366 3032 34702 3088
rect 34758 3032 34763 3088
rect 32305 3030 34763 3032
rect 32305 3027 32371 3030
rect 34697 3027 34763 3030
rect 43437 3090 43503 3093
rect 44200 3090 45000 3120
rect 43437 3088 45000 3090
rect 43437 3032 43442 3088
rect 43498 3032 45000 3088
rect 43437 3030 45000 3032
rect 43437 3027 43503 3030
rect 44200 3000 45000 3030
rect 10980 2952 18479 2954
rect 10980 2896 18418 2952
rect 18474 2896 18479 2952
rect 10980 2894 18479 2896
rect 10980 2892 10986 2894
rect 18413 2891 18479 2894
rect 19750 2894 22110 2954
rect 22185 2954 22251 2957
rect 27153 2954 27219 2957
rect 22185 2952 27219 2954
rect 22185 2896 22190 2952
rect 22246 2896 27158 2952
rect 27214 2896 27219 2952
rect 22185 2894 27219 2896
rect 8937 2818 9003 2821
rect 8526 2816 9003 2818
rect 8526 2760 8942 2816
rect 8998 2760 9003 2816
rect 8526 2758 9003 2760
rect 8937 2755 9003 2758
rect 14365 2818 14431 2821
rect 17861 2818 17927 2821
rect 19750 2818 19810 2894
rect 22185 2891 22251 2894
rect 27153 2891 27219 2894
rect 30189 2954 30255 2957
rect 36537 2954 36603 2957
rect 30189 2952 36603 2954
rect 30189 2896 30194 2952
rect 30250 2896 36542 2952
rect 36598 2896 36603 2952
rect 30189 2894 36603 2896
rect 30189 2891 30255 2894
rect 36537 2891 36603 2894
rect 14365 2816 16498 2818
rect 14365 2760 14370 2816
rect 14426 2760 16498 2816
rect 14365 2758 16498 2760
rect 14365 2755 14431 2758
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 13906 2752 14302 2753
rect 13906 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14302 2752
rect 13906 2687 14302 2688
rect 14365 2682 14431 2685
rect 16297 2682 16363 2685
rect 14365 2680 16363 2682
rect 14365 2624 14370 2680
rect 14426 2624 16302 2680
rect 16358 2624 16363 2680
rect 14365 2622 16363 2624
rect 16438 2682 16498 2758
rect 17861 2816 19810 2818
rect 17861 2760 17866 2816
rect 17922 2760 19810 2816
rect 17861 2758 19810 2760
rect 20437 2818 20503 2821
rect 25405 2818 25471 2821
rect 20437 2816 25471 2818
rect 20437 2760 20442 2816
rect 20498 2760 25410 2816
rect 25466 2760 25471 2816
rect 20437 2758 25471 2760
rect 17861 2755 17927 2758
rect 20437 2755 20503 2758
rect 25405 2755 25471 2758
rect 43069 2818 43135 2821
rect 44200 2818 45000 2848
rect 43069 2816 45000 2818
rect 43069 2760 43074 2816
rect 43130 2760 45000 2816
rect 43069 2758 45000 2760
rect 43069 2755 43135 2758
rect 19906 2752 20302 2753
rect 19906 2688 19912 2752
rect 19976 2688 19992 2752
rect 20056 2688 20072 2752
rect 20136 2688 20152 2752
rect 20216 2688 20232 2752
rect 20296 2688 20302 2752
rect 19906 2687 20302 2688
rect 25906 2752 26302 2753
rect 25906 2688 25912 2752
rect 25976 2688 25992 2752
rect 26056 2688 26072 2752
rect 26136 2688 26152 2752
rect 26216 2688 26232 2752
rect 26296 2688 26302 2752
rect 25906 2687 26302 2688
rect 31906 2752 32302 2753
rect 31906 2688 31912 2752
rect 31976 2688 31992 2752
rect 32056 2688 32072 2752
rect 32136 2688 32152 2752
rect 32216 2688 32232 2752
rect 32296 2688 32302 2752
rect 31906 2687 32302 2688
rect 37906 2752 38302 2753
rect 37906 2688 37912 2752
rect 37976 2688 37992 2752
rect 38056 2688 38072 2752
rect 38136 2688 38152 2752
rect 38216 2688 38232 2752
rect 38296 2688 38302 2752
rect 44200 2728 45000 2758
rect 37906 2687 38302 2688
rect 18781 2682 18847 2685
rect 16438 2680 18847 2682
rect 16438 2624 18786 2680
rect 18842 2624 18847 2680
rect 16438 2622 18847 2624
rect 14365 2619 14431 2622
rect 16297 2619 16363 2622
rect 18781 2619 18847 2622
rect 21265 2682 21331 2685
rect 25773 2682 25839 2685
rect 21265 2680 25839 2682
rect 21265 2624 21270 2680
rect 21326 2624 25778 2680
rect 25834 2624 25839 2680
rect 21265 2622 25839 2624
rect 21265 2619 21331 2622
rect 25773 2619 25839 2622
rect 10726 2546 10732 2548
rect 7606 2486 10732 2546
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 10726 2484 10732 2486
rect 10796 2484 10802 2548
rect 12985 2546 13051 2549
rect 39389 2546 39455 2549
rect 12985 2544 39455 2546
rect 12985 2488 12990 2544
rect 13046 2488 39394 2544
rect 39450 2488 39455 2544
rect 12985 2486 39455 2488
rect 12985 2483 13051 2486
rect 39389 2483 39455 2486
rect 43437 2546 43503 2549
rect 44200 2546 45000 2576
rect 43437 2544 45000 2546
rect 43437 2488 43442 2544
rect 43498 2488 45000 2544
rect 43437 2486 45000 2488
rect 43437 2483 43503 2486
rect 44200 2456 45000 2486
rect 6177 2410 6243 2413
rect 14181 2410 14247 2413
rect 6177 2408 14247 2410
rect 6177 2352 6182 2408
rect 6238 2352 14186 2408
rect 14242 2352 14247 2408
rect 6177 2350 14247 2352
rect 6177 2347 6243 2350
rect 14181 2347 14247 2350
rect 14365 2410 14431 2413
rect 39941 2410 40007 2413
rect 14365 2408 40007 2410
rect 14365 2352 14370 2408
rect 14426 2352 39946 2408
rect 40002 2352 40007 2408
rect 14365 2350 40007 2352
rect 14365 2347 14431 2350
rect 39941 2347 40007 2350
rect 42885 2410 42951 2413
rect 42885 2408 42994 2410
rect 42885 2352 42890 2408
rect 42946 2352 42994 2408
rect 42885 2347 42994 2352
rect 0 2274 800 2304
rect 1393 2274 1459 2277
rect 0 2272 1459 2274
rect 0 2216 1398 2272
rect 1454 2216 1459 2272
rect 0 2214 1459 2216
rect 0 2184 800 2214
rect 1393 2211 1459 2214
rect 9581 2274 9647 2277
rect 14365 2274 14431 2277
rect 9581 2272 14431 2274
rect 9581 2216 9586 2272
rect 9642 2216 14370 2272
rect 14426 2216 14431 2272
rect 9581 2214 14431 2216
rect 9581 2211 9647 2214
rect 14365 2211 14431 2214
rect 2646 2208 3042 2209
rect 2646 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3042 2208
rect 2646 2143 3042 2144
rect 8646 2208 9042 2209
rect 8646 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9042 2208
rect 8646 2143 9042 2144
rect 14646 2208 15042 2209
rect 14646 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15042 2208
rect 14646 2143 15042 2144
rect 20646 2208 21042 2209
rect 20646 2144 20652 2208
rect 20716 2144 20732 2208
rect 20796 2144 20812 2208
rect 20876 2144 20892 2208
rect 20956 2144 20972 2208
rect 21036 2144 21042 2208
rect 20646 2143 21042 2144
rect 26646 2208 27042 2209
rect 26646 2144 26652 2208
rect 26716 2144 26732 2208
rect 26796 2144 26812 2208
rect 26876 2144 26892 2208
rect 26956 2144 26972 2208
rect 27036 2144 27042 2208
rect 26646 2143 27042 2144
rect 32646 2208 33042 2209
rect 32646 2144 32652 2208
rect 32716 2144 32732 2208
rect 32796 2144 32812 2208
rect 32876 2144 32892 2208
rect 32956 2144 32972 2208
rect 33036 2144 33042 2208
rect 32646 2143 33042 2144
rect 38646 2208 39042 2209
rect 38646 2144 38652 2208
rect 38716 2144 38732 2208
rect 38796 2144 38812 2208
rect 38876 2144 38892 2208
rect 38956 2144 38972 2208
rect 39036 2144 39042 2208
rect 38646 2143 39042 2144
rect 11329 2138 11395 2141
rect 12709 2138 12775 2141
rect 11329 2136 12775 2138
rect 11329 2080 11334 2136
rect 11390 2080 12714 2136
rect 12770 2080 12775 2136
rect 11329 2078 12775 2080
rect 11329 2075 11395 2078
rect 12709 2075 12775 2078
rect 0 2002 800 2032
rect 1761 2002 1827 2005
rect 0 2000 1827 2002
rect 0 1944 1766 2000
rect 1822 1944 1827 2000
rect 0 1942 1827 1944
rect 0 1912 800 1942
rect 1761 1939 1827 1942
rect 9489 2002 9555 2005
rect 34513 2002 34579 2005
rect 9489 2000 34579 2002
rect 9489 1944 9494 2000
rect 9550 1944 34518 2000
rect 34574 1944 34579 2000
rect 9489 1942 34579 1944
rect 42934 2002 42994 2347
rect 43069 2274 43135 2277
rect 44200 2274 45000 2304
rect 43069 2272 45000 2274
rect 43069 2216 43074 2272
rect 43130 2216 45000 2272
rect 43069 2214 45000 2216
rect 43069 2211 43135 2214
rect 44200 2184 45000 2214
rect 44200 2002 45000 2032
rect 42934 1942 45000 2002
rect 9489 1939 9555 1942
rect 34513 1939 34579 1942
rect 44200 1912 45000 1942
rect 11145 1866 11211 1869
rect 18229 1866 18295 1869
rect 11145 1864 18295 1866
rect 11145 1808 11150 1864
rect 11206 1808 18234 1864
rect 18290 1808 18295 1864
rect 11145 1806 18295 1808
rect 11145 1803 11211 1806
rect 18229 1803 18295 1806
rect 19190 1804 19196 1868
rect 19260 1866 19266 1868
rect 22185 1866 22251 1869
rect 19260 1864 22251 1866
rect 19260 1808 22190 1864
rect 22246 1808 22251 1864
rect 19260 1806 22251 1808
rect 19260 1804 19266 1806
rect 22185 1803 22251 1806
rect 26233 1866 26299 1869
rect 27838 1866 27844 1868
rect 26233 1864 27844 1866
rect 26233 1808 26238 1864
rect 26294 1808 27844 1864
rect 26233 1806 27844 1808
rect 26233 1803 26299 1806
rect 27838 1804 27844 1806
rect 27908 1804 27914 1868
rect 0 1730 800 1760
rect 3325 1730 3391 1733
rect 0 1728 3391 1730
rect 0 1672 3330 1728
rect 3386 1672 3391 1728
rect 0 1670 3391 1672
rect 0 1640 800 1670
rect 3325 1667 3391 1670
rect 12985 1730 13051 1733
rect 33961 1730 34027 1733
rect 12985 1728 34027 1730
rect 12985 1672 12990 1728
rect 13046 1672 33966 1728
rect 34022 1672 34027 1728
rect 12985 1670 34027 1672
rect 12985 1667 13051 1670
rect 33961 1667 34027 1670
rect 42793 1730 42859 1733
rect 44200 1730 45000 1760
rect 42793 1728 45000 1730
rect 42793 1672 42798 1728
rect 42854 1672 45000 1728
rect 42793 1670 45000 1672
rect 42793 1667 42859 1670
rect 44200 1640 45000 1670
rect 9213 1594 9279 1597
rect 37273 1594 37339 1597
rect 9213 1592 37339 1594
rect 9213 1536 9218 1592
rect 9274 1536 37278 1592
rect 37334 1536 37339 1592
rect 9213 1534 37339 1536
rect 9213 1531 9279 1534
rect 37273 1531 37339 1534
rect 0 1458 800 1488
rect 2405 1458 2471 1461
rect 0 1456 2471 1458
rect 0 1400 2410 1456
rect 2466 1400 2471 1456
rect 0 1398 2471 1400
rect 0 1368 800 1398
rect 2405 1395 2471 1398
rect 5993 1458 6059 1461
rect 29453 1458 29519 1461
rect 5993 1456 29519 1458
rect 5993 1400 5998 1456
rect 6054 1400 29458 1456
rect 29514 1400 29519 1456
rect 5993 1398 29519 1400
rect 5993 1395 6059 1398
rect 29453 1395 29519 1398
rect 42885 1458 42951 1461
rect 44200 1458 45000 1488
rect 42885 1456 45000 1458
rect 42885 1400 42890 1456
rect 42946 1400 45000 1456
rect 42885 1398 45000 1400
rect 42885 1395 42951 1398
rect 44200 1368 45000 1398
rect 4337 1322 4403 1325
rect 10358 1322 10364 1324
rect 4337 1320 10364 1322
rect 4337 1264 4342 1320
rect 4398 1264 10364 1320
rect 4337 1262 10364 1264
rect 4337 1259 4403 1262
rect 10358 1260 10364 1262
rect 10428 1260 10434 1324
rect 14365 1322 14431 1325
rect 32765 1322 32831 1325
rect 14365 1320 32831 1322
rect 14365 1264 14370 1320
rect 14426 1264 32770 1320
rect 32826 1264 32831 1320
rect 14365 1262 32831 1264
rect 14365 1259 14431 1262
rect 32765 1259 32831 1262
rect 3877 1186 3943 1189
rect 36997 1186 37063 1189
rect 3877 1184 37063 1186
rect 3877 1128 3882 1184
rect 3938 1128 37002 1184
rect 37058 1128 37063 1184
rect 3877 1126 37063 1128
rect 3877 1123 3943 1126
rect 36997 1123 37063 1126
rect 7649 1050 7715 1053
rect 37181 1050 37247 1053
rect 7649 1048 37247 1050
rect 7649 992 7654 1048
rect 7710 992 37186 1048
rect 37242 992 37247 1048
rect 7649 990 37247 992
rect 7649 987 7715 990
rect 37181 987 37247 990
rect 3969 914 4035 917
rect 29085 914 29151 917
rect 3969 912 29151 914
rect 3969 856 3974 912
rect 4030 856 29090 912
rect 29146 856 29151 912
rect 3969 854 29151 856
rect 3969 851 4035 854
rect 29085 851 29151 854
rect 7005 778 7071 781
rect 33685 778 33751 781
rect 7005 776 33751 778
rect 7005 720 7010 776
rect 7066 720 33690 776
rect 33746 720 33751 776
rect 7005 718 33751 720
rect 7005 715 7071 718
rect 33685 715 33751 718
rect 7465 642 7531 645
rect 33041 642 33107 645
rect 7465 640 33107 642
rect 7465 584 7470 640
rect 7526 584 33046 640
rect 33102 584 33107 640
rect 7465 582 33107 584
rect 7465 579 7531 582
rect 33041 579 33107 582
rect 10777 506 10843 509
rect 39481 506 39547 509
rect 10777 504 39547 506
rect 10777 448 10782 504
rect 10838 448 39486 504
rect 39542 448 39547 504
rect 10777 446 39547 448
rect 10777 443 10843 446
rect 39481 443 39547 446
<< via3 >>
rect 6316 10508 6380 10572
rect 10364 10372 10428 10436
rect 21220 10236 21284 10300
rect 5948 10100 6012 10164
rect 17356 9828 17420 9892
rect 16988 9692 17052 9756
rect 15148 9420 15212 9484
rect 21220 9420 21284 9484
rect 17724 9012 17788 9076
rect 35020 9012 35084 9076
rect 27660 8876 27724 8940
rect 19564 8740 19628 8804
rect 2652 8732 2716 8736
rect 2652 8676 2656 8732
rect 2656 8676 2712 8732
rect 2712 8676 2716 8732
rect 2652 8672 2716 8676
rect 2732 8732 2796 8736
rect 2732 8676 2736 8732
rect 2736 8676 2792 8732
rect 2792 8676 2796 8732
rect 2732 8672 2796 8676
rect 2812 8732 2876 8736
rect 2812 8676 2816 8732
rect 2816 8676 2872 8732
rect 2872 8676 2876 8732
rect 2812 8672 2876 8676
rect 2892 8732 2956 8736
rect 2892 8676 2896 8732
rect 2896 8676 2952 8732
rect 2952 8676 2956 8732
rect 2892 8672 2956 8676
rect 2972 8732 3036 8736
rect 2972 8676 2976 8732
rect 2976 8676 3032 8732
rect 3032 8676 3036 8732
rect 2972 8672 3036 8676
rect 8652 8732 8716 8736
rect 8652 8676 8656 8732
rect 8656 8676 8712 8732
rect 8712 8676 8716 8732
rect 8652 8672 8716 8676
rect 8732 8732 8796 8736
rect 8732 8676 8736 8732
rect 8736 8676 8792 8732
rect 8792 8676 8796 8732
rect 8732 8672 8796 8676
rect 8812 8732 8876 8736
rect 8812 8676 8816 8732
rect 8816 8676 8872 8732
rect 8872 8676 8876 8732
rect 8812 8672 8876 8676
rect 8892 8732 8956 8736
rect 8892 8676 8896 8732
rect 8896 8676 8952 8732
rect 8952 8676 8956 8732
rect 8892 8672 8956 8676
rect 8972 8732 9036 8736
rect 8972 8676 8976 8732
rect 8976 8676 9032 8732
rect 9032 8676 9036 8732
rect 8972 8672 9036 8676
rect 14652 8732 14716 8736
rect 14652 8676 14656 8732
rect 14656 8676 14712 8732
rect 14712 8676 14716 8732
rect 14652 8672 14716 8676
rect 14732 8732 14796 8736
rect 14732 8676 14736 8732
rect 14736 8676 14792 8732
rect 14792 8676 14796 8732
rect 14732 8672 14796 8676
rect 14812 8732 14876 8736
rect 14812 8676 14816 8732
rect 14816 8676 14872 8732
rect 14872 8676 14876 8732
rect 14812 8672 14876 8676
rect 14892 8732 14956 8736
rect 14892 8676 14896 8732
rect 14896 8676 14952 8732
rect 14952 8676 14956 8732
rect 14892 8672 14956 8676
rect 14972 8732 15036 8736
rect 14972 8676 14976 8732
rect 14976 8676 15032 8732
rect 15032 8676 15036 8732
rect 14972 8672 15036 8676
rect 20652 8732 20716 8736
rect 20652 8676 20656 8732
rect 20656 8676 20712 8732
rect 20712 8676 20716 8732
rect 20652 8672 20716 8676
rect 20732 8732 20796 8736
rect 20732 8676 20736 8732
rect 20736 8676 20792 8732
rect 20792 8676 20796 8732
rect 20732 8672 20796 8676
rect 20812 8732 20876 8736
rect 20812 8676 20816 8732
rect 20816 8676 20872 8732
rect 20872 8676 20876 8732
rect 20812 8672 20876 8676
rect 20892 8732 20956 8736
rect 20892 8676 20896 8732
rect 20896 8676 20952 8732
rect 20952 8676 20956 8732
rect 20892 8672 20956 8676
rect 20972 8732 21036 8736
rect 20972 8676 20976 8732
rect 20976 8676 21032 8732
rect 21032 8676 21036 8732
rect 20972 8672 21036 8676
rect 26652 8732 26716 8736
rect 26652 8676 26656 8732
rect 26656 8676 26712 8732
rect 26712 8676 26716 8732
rect 26652 8672 26716 8676
rect 26732 8732 26796 8736
rect 26732 8676 26736 8732
rect 26736 8676 26792 8732
rect 26792 8676 26796 8732
rect 26732 8672 26796 8676
rect 26812 8732 26876 8736
rect 26812 8676 26816 8732
rect 26816 8676 26872 8732
rect 26872 8676 26876 8732
rect 26812 8672 26876 8676
rect 26892 8732 26956 8736
rect 26892 8676 26896 8732
rect 26896 8676 26952 8732
rect 26952 8676 26956 8732
rect 26892 8672 26956 8676
rect 26972 8732 27036 8736
rect 26972 8676 26976 8732
rect 26976 8676 27032 8732
rect 27032 8676 27036 8732
rect 26972 8672 27036 8676
rect 32652 8732 32716 8736
rect 32652 8676 32656 8732
rect 32656 8676 32712 8732
rect 32712 8676 32716 8732
rect 32652 8672 32716 8676
rect 32732 8732 32796 8736
rect 32732 8676 32736 8732
rect 32736 8676 32792 8732
rect 32792 8676 32796 8732
rect 32732 8672 32796 8676
rect 32812 8732 32876 8736
rect 32812 8676 32816 8732
rect 32816 8676 32872 8732
rect 32872 8676 32876 8732
rect 32812 8672 32876 8676
rect 32892 8732 32956 8736
rect 32892 8676 32896 8732
rect 32896 8676 32952 8732
rect 32952 8676 32956 8732
rect 32892 8672 32956 8676
rect 32972 8732 33036 8736
rect 32972 8676 32976 8732
rect 32976 8676 33032 8732
rect 33032 8676 33036 8732
rect 32972 8672 33036 8676
rect 38652 8732 38716 8736
rect 38652 8676 38656 8732
rect 38656 8676 38712 8732
rect 38712 8676 38716 8732
rect 38652 8672 38716 8676
rect 38732 8732 38796 8736
rect 38732 8676 38736 8732
rect 38736 8676 38792 8732
rect 38792 8676 38796 8732
rect 38732 8672 38796 8676
rect 38812 8732 38876 8736
rect 38812 8676 38816 8732
rect 38816 8676 38872 8732
rect 38872 8676 38876 8732
rect 38812 8672 38876 8676
rect 38892 8732 38956 8736
rect 38892 8676 38896 8732
rect 38896 8676 38952 8732
rect 38952 8676 38956 8732
rect 38892 8672 38956 8676
rect 38972 8732 39036 8736
rect 38972 8676 38976 8732
rect 38976 8676 39032 8732
rect 39032 8676 39036 8732
rect 38972 8672 39036 8676
rect 15332 8604 15396 8668
rect 32444 8604 32508 8668
rect 10732 8332 10796 8396
rect 13492 8196 13556 8260
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 15516 8332 15580 8396
rect 33916 8256 33980 8260
rect 33916 8200 33930 8256
rect 33930 8200 33980 8256
rect 33916 8196 33980 8200
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 14152 8188 14216 8192
rect 14152 8132 14156 8188
rect 14156 8132 14212 8188
rect 14212 8132 14216 8188
rect 14152 8128 14216 8132
rect 14232 8188 14296 8192
rect 14232 8132 14236 8188
rect 14236 8132 14292 8188
rect 14292 8132 14296 8188
rect 14232 8128 14296 8132
rect 19912 8188 19976 8192
rect 19912 8132 19916 8188
rect 19916 8132 19972 8188
rect 19972 8132 19976 8188
rect 19912 8128 19976 8132
rect 19992 8188 20056 8192
rect 19992 8132 19996 8188
rect 19996 8132 20052 8188
rect 20052 8132 20056 8188
rect 19992 8128 20056 8132
rect 20072 8188 20136 8192
rect 20072 8132 20076 8188
rect 20076 8132 20132 8188
rect 20132 8132 20136 8188
rect 20072 8128 20136 8132
rect 20152 8188 20216 8192
rect 20152 8132 20156 8188
rect 20156 8132 20212 8188
rect 20212 8132 20216 8188
rect 20152 8128 20216 8132
rect 20232 8188 20296 8192
rect 20232 8132 20236 8188
rect 20236 8132 20292 8188
rect 20292 8132 20296 8188
rect 20232 8128 20296 8132
rect 25912 8188 25976 8192
rect 25912 8132 25916 8188
rect 25916 8132 25972 8188
rect 25972 8132 25976 8188
rect 25912 8128 25976 8132
rect 25992 8188 26056 8192
rect 25992 8132 25996 8188
rect 25996 8132 26052 8188
rect 26052 8132 26056 8188
rect 25992 8128 26056 8132
rect 26072 8188 26136 8192
rect 26072 8132 26076 8188
rect 26076 8132 26132 8188
rect 26132 8132 26136 8188
rect 26072 8128 26136 8132
rect 26152 8188 26216 8192
rect 26152 8132 26156 8188
rect 26156 8132 26212 8188
rect 26212 8132 26216 8188
rect 26152 8128 26216 8132
rect 26232 8188 26296 8192
rect 26232 8132 26236 8188
rect 26236 8132 26292 8188
rect 26292 8132 26296 8188
rect 26232 8128 26296 8132
rect 31912 8188 31976 8192
rect 31912 8132 31916 8188
rect 31916 8132 31972 8188
rect 31972 8132 31976 8188
rect 31912 8128 31976 8132
rect 31992 8188 32056 8192
rect 31992 8132 31996 8188
rect 31996 8132 32052 8188
rect 32052 8132 32056 8188
rect 31992 8128 32056 8132
rect 32072 8188 32136 8192
rect 32072 8132 32076 8188
rect 32076 8132 32132 8188
rect 32132 8132 32136 8188
rect 32072 8128 32136 8132
rect 32152 8188 32216 8192
rect 32152 8132 32156 8188
rect 32156 8132 32212 8188
rect 32212 8132 32216 8188
rect 32152 8128 32216 8132
rect 32232 8188 32296 8192
rect 32232 8132 32236 8188
rect 32236 8132 32292 8188
rect 32292 8132 32296 8188
rect 32232 8128 32296 8132
rect 37912 8188 37976 8192
rect 37912 8132 37916 8188
rect 37916 8132 37972 8188
rect 37972 8132 37976 8188
rect 37912 8128 37976 8132
rect 37992 8188 38056 8192
rect 37992 8132 37996 8188
rect 37996 8132 38052 8188
rect 38052 8132 38056 8188
rect 37992 8128 38056 8132
rect 38072 8188 38136 8192
rect 38072 8132 38076 8188
rect 38076 8132 38132 8188
rect 38132 8132 38136 8188
rect 38072 8128 38136 8132
rect 38152 8188 38216 8192
rect 38152 8132 38156 8188
rect 38156 8132 38212 8188
rect 38212 8132 38216 8188
rect 38152 8128 38216 8132
rect 38232 8188 38296 8192
rect 38232 8132 38236 8188
rect 38236 8132 38292 8188
rect 38292 8132 38296 8188
rect 38232 8128 38296 8132
rect 20484 8060 20548 8124
rect 4292 7712 4356 7716
rect 4292 7656 4342 7712
rect 4342 7656 4356 7712
rect 4292 7652 4356 7656
rect 5948 7652 6012 7716
rect 6316 7652 6380 7716
rect 2652 7644 2716 7648
rect 2652 7588 2656 7644
rect 2656 7588 2712 7644
rect 2712 7588 2716 7644
rect 2652 7584 2716 7588
rect 2732 7644 2796 7648
rect 2732 7588 2736 7644
rect 2736 7588 2792 7644
rect 2792 7588 2796 7644
rect 2732 7584 2796 7588
rect 2812 7644 2876 7648
rect 2812 7588 2816 7644
rect 2816 7588 2872 7644
rect 2872 7588 2876 7644
rect 2812 7584 2876 7588
rect 2892 7644 2956 7648
rect 2892 7588 2896 7644
rect 2896 7588 2952 7644
rect 2952 7588 2956 7644
rect 2892 7584 2956 7588
rect 2972 7644 3036 7648
rect 2972 7588 2976 7644
rect 2976 7588 3032 7644
rect 3032 7588 3036 7644
rect 2972 7584 3036 7588
rect 26372 8060 26436 8124
rect 13676 7788 13740 7852
rect 8652 7644 8716 7648
rect 8652 7588 8656 7644
rect 8656 7588 8712 7644
rect 8712 7588 8716 7644
rect 8652 7584 8716 7588
rect 8732 7644 8796 7648
rect 8732 7588 8736 7644
rect 8736 7588 8792 7644
rect 8792 7588 8796 7644
rect 8732 7584 8796 7588
rect 8812 7644 8876 7648
rect 8812 7588 8816 7644
rect 8816 7588 8872 7644
rect 8872 7588 8876 7644
rect 8812 7584 8876 7588
rect 8892 7644 8956 7648
rect 8892 7588 8896 7644
rect 8896 7588 8952 7644
rect 8952 7588 8956 7644
rect 8892 7584 8956 7588
rect 8972 7644 9036 7648
rect 8972 7588 8976 7644
rect 8976 7588 9032 7644
rect 9032 7588 9036 7644
rect 8972 7584 9036 7588
rect 14652 7644 14716 7648
rect 14652 7588 14656 7644
rect 14656 7588 14712 7644
rect 14712 7588 14716 7644
rect 14652 7584 14716 7588
rect 14732 7644 14796 7648
rect 14732 7588 14736 7644
rect 14736 7588 14792 7644
rect 14792 7588 14796 7644
rect 14732 7584 14796 7588
rect 14812 7644 14876 7648
rect 14812 7588 14816 7644
rect 14816 7588 14872 7644
rect 14872 7588 14876 7644
rect 14812 7584 14876 7588
rect 14892 7644 14956 7648
rect 14892 7588 14896 7644
rect 14896 7588 14952 7644
rect 14952 7588 14956 7644
rect 14892 7584 14956 7588
rect 14972 7644 15036 7648
rect 14972 7588 14976 7644
rect 14976 7588 15032 7644
rect 15032 7588 15036 7644
rect 14972 7584 15036 7588
rect 12572 7516 12636 7580
rect 26372 7788 26436 7852
rect 21404 7652 21468 7716
rect 20652 7644 20716 7648
rect 20652 7588 20656 7644
rect 20656 7588 20712 7644
rect 20712 7588 20716 7644
rect 20652 7584 20716 7588
rect 20732 7644 20796 7648
rect 20732 7588 20736 7644
rect 20736 7588 20792 7644
rect 20792 7588 20796 7644
rect 20732 7584 20796 7588
rect 20812 7644 20876 7648
rect 20812 7588 20816 7644
rect 20816 7588 20872 7644
rect 20872 7588 20876 7644
rect 20812 7584 20876 7588
rect 20892 7644 20956 7648
rect 20892 7588 20896 7644
rect 20896 7588 20952 7644
rect 20952 7588 20956 7644
rect 20892 7584 20956 7588
rect 20972 7644 21036 7648
rect 20972 7588 20976 7644
rect 20976 7588 21032 7644
rect 21032 7588 21036 7644
rect 20972 7584 21036 7588
rect 26652 7644 26716 7648
rect 26652 7588 26656 7644
rect 26656 7588 26712 7644
rect 26712 7588 26716 7644
rect 26652 7584 26716 7588
rect 26732 7644 26796 7648
rect 26732 7588 26736 7644
rect 26736 7588 26792 7644
rect 26792 7588 26796 7644
rect 26732 7584 26796 7588
rect 26812 7644 26876 7648
rect 26812 7588 26816 7644
rect 26816 7588 26872 7644
rect 26872 7588 26876 7644
rect 26812 7584 26876 7588
rect 26892 7644 26956 7648
rect 26892 7588 26896 7644
rect 26896 7588 26952 7644
rect 26952 7588 26956 7644
rect 26892 7584 26956 7588
rect 26972 7644 27036 7648
rect 26972 7588 26976 7644
rect 26976 7588 27032 7644
rect 27032 7588 27036 7644
rect 26972 7584 27036 7588
rect 32652 7644 32716 7648
rect 32652 7588 32656 7644
rect 32656 7588 32712 7644
rect 32712 7588 32716 7644
rect 32652 7584 32716 7588
rect 32732 7644 32796 7648
rect 32732 7588 32736 7644
rect 32736 7588 32792 7644
rect 32792 7588 32796 7644
rect 32732 7584 32796 7588
rect 32812 7644 32876 7648
rect 32812 7588 32816 7644
rect 32816 7588 32872 7644
rect 32872 7588 32876 7644
rect 32812 7584 32876 7588
rect 32892 7644 32956 7648
rect 32892 7588 32896 7644
rect 32896 7588 32952 7644
rect 32952 7588 32956 7644
rect 32892 7584 32956 7588
rect 32972 7644 33036 7648
rect 32972 7588 32976 7644
rect 32976 7588 33032 7644
rect 33032 7588 33036 7644
rect 32972 7584 33036 7588
rect 38652 7644 38716 7648
rect 38652 7588 38656 7644
rect 38656 7588 38712 7644
rect 38712 7588 38716 7644
rect 38652 7584 38716 7588
rect 38732 7644 38796 7648
rect 38732 7588 38736 7644
rect 38736 7588 38792 7644
rect 38792 7588 38796 7644
rect 38732 7584 38796 7588
rect 38812 7644 38876 7648
rect 38812 7588 38816 7644
rect 38816 7588 38872 7644
rect 38872 7588 38876 7644
rect 38812 7584 38876 7588
rect 38892 7644 38956 7648
rect 38892 7588 38896 7644
rect 38896 7588 38952 7644
rect 38952 7588 38956 7644
rect 38892 7584 38956 7588
rect 38972 7644 39036 7648
rect 38972 7588 38976 7644
rect 38976 7588 39032 7644
rect 39032 7588 39036 7644
rect 38972 7584 39036 7588
rect 20484 7516 20548 7580
rect 26372 7516 26436 7580
rect 21588 7108 21652 7172
rect 21772 7108 21836 7172
rect 26372 7108 26436 7172
rect 32444 7168 32508 7172
rect 32444 7112 32494 7168
rect 32494 7112 32508 7168
rect 32444 7108 32508 7112
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 14152 7100 14216 7104
rect 14152 7044 14156 7100
rect 14156 7044 14212 7100
rect 14212 7044 14216 7100
rect 14152 7040 14216 7044
rect 14232 7100 14296 7104
rect 14232 7044 14236 7100
rect 14236 7044 14292 7100
rect 14292 7044 14296 7100
rect 14232 7040 14296 7044
rect 19912 7100 19976 7104
rect 19912 7044 19916 7100
rect 19916 7044 19972 7100
rect 19972 7044 19976 7100
rect 19912 7040 19976 7044
rect 19992 7100 20056 7104
rect 19992 7044 19996 7100
rect 19996 7044 20052 7100
rect 20052 7044 20056 7100
rect 19992 7040 20056 7044
rect 20072 7100 20136 7104
rect 20072 7044 20076 7100
rect 20076 7044 20132 7100
rect 20132 7044 20136 7100
rect 20072 7040 20136 7044
rect 20152 7100 20216 7104
rect 20152 7044 20156 7100
rect 20156 7044 20212 7100
rect 20212 7044 20216 7100
rect 20152 7040 20216 7044
rect 20232 7100 20296 7104
rect 20232 7044 20236 7100
rect 20236 7044 20292 7100
rect 20292 7044 20296 7100
rect 20232 7040 20296 7044
rect 25912 7100 25976 7104
rect 25912 7044 25916 7100
rect 25916 7044 25972 7100
rect 25972 7044 25976 7100
rect 25912 7040 25976 7044
rect 25992 7100 26056 7104
rect 25992 7044 25996 7100
rect 25996 7044 26052 7100
rect 26052 7044 26056 7100
rect 25992 7040 26056 7044
rect 26072 7100 26136 7104
rect 26072 7044 26076 7100
rect 26076 7044 26132 7100
rect 26132 7044 26136 7100
rect 26072 7040 26136 7044
rect 26152 7100 26216 7104
rect 26152 7044 26156 7100
rect 26156 7044 26212 7100
rect 26212 7044 26216 7100
rect 26152 7040 26216 7044
rect 26232 7100 26296 7104
rect 26232 7044 26236 7100
rect 26236 7044 26292 7100
rect 26292 7044 26296 7100
rect 26232 7040 26296 7044
rect 31912 7100 31976 7104
rect 31912 7044 31916 7100
rect 31916 7044 31972 7100
rect 31972 7044 31976 7100
rect 31912 7040 31976 7044
rect 31992 7100 32056 7104
rect 31992 7044 31996 7100
rect 31996 7044 32052 7100
rect 32052 7044 32056 7100
rect 31992 7040 32056 7044
rect 32072 7100 32136 7104
rect 32072 7044 32076 7100
rect 32076 7044 32132 7100
rect 32132 7044 32136 7100
rect 32072 7040 32136 7044
rect 32152 7100 32216 7104
rect 32152 7044 32156 7100
rect 32156 7044 32212 7100
rect 32212 7044 32216 7100
rect 32152 7040 32216 7044
rect 32232 7100 32296 7104
rect 32232 7044 32236 7100
rect 32236 7044 32292 7100
rect 32292 7044 32296 7100
rect 32232 7040 32296 7044
rect 37912 7100 37976 7104
rect 37912 7044 37916 7100
rect 37916 7044 37972 7100
rect 37972 7044 37976 7100
rect 37912 7040 37976 7044
rect 37992 7100 38056 7104
rect 37992 7044 37996 7100
rect 37996 7044 38052 7100
rect 38052 7044 38056 7100
rect 37992 7040 38056 7044
rect 38072 7100 38136 7104
rect 38072 7044 38076 7100
rect 38076 7044 38132 7100
rect 38132 7044 38136 7100
rect 38072 7040 38136 7044
rect 38152 7100 38216 7104
rect 38152 7044 38156 7100
rect 38156 7044 38212 7100
rect 38212 7044 38216 7100
rect 38152 7040 38216 7044
rect 38232 7100 38296 7104
rect 38232 7044 38236 7100
rect 38236 7044 38292 7100
rect 38292 7044 38296 7100
rect 38232 7040 38296 7044
rect 19196 6972 19260 7036
rect 21220 6972 21284 7036
rect 26372 6972 26436 7036
rect 19012 6836 19076 6900
rect 20484 6564 20548 6628
rect 2652 6556 2716 6560
rect 2652 6500 2656 6556
rect 2656 6500 2712 6556
rect 2712 6500 2716 6556
rect 2652 6496 2716 6500
rect 2732 6556 2796 6560
rect 2732 6500 2736 6556
rect 2736 6500 2792 6556
rect 2792 6500 2796 6556
rect 2732 6496 2796 6500
rect 2812 6556 2876 6560
rect 2812 6500 2816 6556
rect 2816 6500 2872 6556
rect 2872 6500 2876 6556
rect 2812 6496 2876 6500
rect 2892 6556 2956 6560
rect 2892 6500 2896 6556
rect 2896 6500 2952 6556
rect 2952 6500 2956 6556
rect 2892 6496 2956 6500
rect 2972 6556 3036 6560
rect 2972 6500 2976 6556
rect 2976 6500 3032 6556
rect 3032 6500 3036 6556
rect 2972 6496 3036 6500
rect 8652 6556 8716 6560
rect 8652 6500 8656 6556
rect 8656 6500 8712 6556
rect 8712 6500 8716 6556
rect 8652 6496 8716 6500
rect 8732 6556 8796 6560
rect 8732 6500 8736 6556
rect 8736 6500 8792 6556
rect 8792 6500 8796 6556
rect 8732 6496 8796 6500
rect 8812 6556 8876 6560
rect 8812 6500 8816 6556
rect 8816 6500 8872 6556
rect 8872 6500 8876 6556
rect 8812 6496 8876 6500
rect 8892 6556 8956 6560
rect 8892 6500 8896 6556
rect 8896 6500 8952 6556
rect 8952 6500 8956 6556
rect 8892 6496 8956 6500
rect 8972 6556 9036 6560
rect 8972 6500 8976 6556
rect 8976 6500 9032 6556
rect 9032 6500 9036 6556
rect 8972 6496 9036 6500
rect 14652 6556 14716 6560
rect 14652 6500 14656 6556
rect 14656 6500 14712 6556
rect 14712 6500 14716 6556
rect 14652 6496 14716 6500
rect 14732 6556 14796 6560
rect 14732 6500 14736 6556
rect 14736 6500 14792 6556
rect 14792 6500 14796 6556
rect 14732 6496 14796 6500
rect 14812 6556 14876 6560
rect 14812 6500 14816 6556
rect 14816 6500 14872 6556
rect 14872 6500 14876 6556
rect 14812 6496 14876 6500
rect 14892 6556 14956 6560
rect 14892 6500 14896 6556
rect 14896 6500 14952 6556
rect 14952 6500 14956 6556
rect 14892 6496 14956 6500
rect 14972 6556 15036 6560
rect 14972 6500 14976 6556
rect 14976 6500 15032 6556
rect 15032 6500 15036 6556
rect 14972 6496 15036 6500
rect 20652 6556 20716 6560
rect 20652 6500 20656 6556
rect 20656 6500 20712 6556
rect 20712 6500 20716 6556
rect 20652 6496 20716 6500
rect 20732 6556 20796 6560
rect 20732 6500 20736 6556
rect 20736 6500 20792 6556
rect 20792 6500 20796 6556
rect 20732 6496 20796 6500
rect 20812 6556 20876 6560
rect 20812 6500 20816 6556
rect 20816 6500 20872 6556
rect 20872 6500 20876 6556
rect 20812 6496 20876 6500
rect 20892 6556 20956 6560
rect 20892 6500 20896 6556
rect 20896 6500 20952 6556
rect 20952 6500 20956 6556
rect 20892 6496 20956 6500
rect 20972 6556 21036 6560
rect 20972 6500 20976 6556
rect 20976 6500 21032 6556
rect 21032 6500 21036 6556
rect 20972 6496 21036 6500
rect 26652 6556 26716 6560
rect 26652 6500 26656 6556
rect 26656 6500 26712 6556
rect 26712 6500 26716 6556
rect 26652 6496 26716 6500
rect 26732 6556 26796 6560
rect 26732 6500 26736 6556
rect 26736 6500 26792 6556
rect 26792 6500 26796 6556
rect 26732 6496 26796 6500
rect 26812 6556 26876 6560
rect 26812 6500 26816 6556
rect 26816 6500 26872 6556
rect 26872 6500 26876 6556
rect 26812 6496 26876 6500
rect 26892 6556 26956 6560
rect 26892 6500 26896 6556
rect 26896 6500 26952 6556
rect 26952 6500 26956 6556
rect 26892 6496 26956 6500
rect 26972 6556 27036 6560
rect 26972 6500 26976 6556
rect 26976 6500 27032 6556
rect 27032 6500 27036 6556
rect 26972 6496 27036 6500
rect 32652 6556 32716 6560
rect 32652 6500 32656 6556
rect 32656 6500 32712 6556
rect 32712 6500 32716 6556
rect 32652 6496 32716 6500
rect 32732 6556 32796 6560
rect 32732 6500 32736 6556
rect 32736 6500 32792 6556
rect 32792 6500 32796 6556
rect 32732 6496 32796 6500
rect 32812 6556 32876 6560
rect 32812 6500 32816 6556
rect 32816 6500 32872 6556
rect 32872 6500 32876 6556
rect 32812 6496 32876 6500
rect 32892 6556 32956 6560
rect 32892 6500 32896 6556
rect 32896 6500 32952 6556
rect 32952 6500 32956 6556
rect 32892 6496 32956 6500
rect 32972 6556 33036 6560
rect 32972 6500 32976 6556
rect 32976 6500 33032 6556
rect 33032 6500 33036 6556
rect 32972 6496 33036 6500
rect 38652 6556 38716 6560
rect 38652 6500 38656 6556
rect 38656 6500 38712 6556
rect 38712 6500 38716 6556
rect 38652 6496 38716 6500
rect 38732 6556 38796 6560
rect 38732 6500 38736 6556
rect 38736 6500 38792 6556
rect 38792 6500 38796 6556
rect 38732 6496 38796 6500
rect 38812 6556 38876 6560
rect 38812 6500 38816 6556
rect 38816 6500 38872 6556
rect 38872 6500 38876 6556
rect 38812 6496 38876 6500
rect 38892 6556 38956 6560
rect 38892 6500 38896 6556
rect 38896 6500 38952 6556
rect 38952 6500 38956 6556
rect 38892 6496 38956 6500
rect 38972 6556 39036 6560
rect 38972 6500 38976 6556
rect 38976 6500 39032 6556
rect 39032 6500 39036 6556
rect 38972 6496 39036 6500
rect 26372 6428 26436 6492
rect 27108 6428 27172 6492
rect 32444 6292 32508 6356
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 14152 6012 14216 6016
rect 14152 5956 14156 6012
rect 14156 5956 14212 6012
rect 14212 5956 14216 6012
rect 14152 5952 14216 5956
rect 14232 6012 14296 6016
rect 14232 5956 14236 6012
rect 14236 5956 14292 6012
rect 14292 5956 14296 6012
rect 14232 5952 14296 5956
rect 20484 6020 20548 6084
rect 19912 6012 19976 6016
rect 19912 5956 19916 6012
rect 19916 5956 19972 6012
rect 19972 5956 19976 6012
rect 19912 5952 19976 5956
rect 19992 6012 20056 6016
rect 19992 5956 19996 6012
rect 19996 5956 20052 6012
rect 20052 5956 20056 6012
rect 19992 5952 20056 5956
rect 20072 6012 20136 6016
rect 20072 5956 20076 6012
rect 20076 5956 20132 6012
rect 20132 5956 20136 6012
rect 20072 5952 20136 5956
rect 20152 6012 20216 6016
rect 20152 5956 20156 6012
rect 20156 5956 20212 6012
rect 20212 5956 20216 6012
rect 20152 5952 20216 5956
rect 20232 6012 20296 6016
rect 20232 5956 20236 6012
rect 20236 5956 20292 6012
rect 20292 5956 20296 6012
rect 20232 5952 20296 5956
rect 25912 6012 25976 6016
rect 25912 5956 25916 6012
rect 25916 5956 25972 6012
rect 25972 5956 25976 6012
rect 25912 5952 25976 5956
rect 25992 6012 26056 6016
rect 25992 5956 25996 6012
rect 25996 5956 26052 6012
rect 26052 5956 26056 6012
rect 25992 5952 26056 5956
rect 26072 6012 26136 6016
rect 26072 5956 26076 6012
rect 26076 5956 26132 6012
rect 26132 5956 26136 6012
rect 26072 5952 26136 5956
rect 26152 6012 26216 6016
rect 26152 5956 26156 6012
rect 26156 5956 26212 6012
rect 26212 5956 26216 6012
rect 26152 5952 26216 5956
rect 26232 6012 26296 6016
rect 26232 5956 26236 6012
rect 26236 5956 26292 6012
rect 26292 5956 26296 6012
rect 26232 5952 26296 5956
rect 20484 5884 20548 5948
rect 9444 5748 9508 5812
rect 27108 6020 27172 6084
rect 31912 6012 31976 6016
rect 31912 5956 31916 6012
rect 31916 5956 31972 6012
rect 31972 5956 31976 6012
rect 31912 5952 31976 5956
rect 31992 6012 32056 6016
rect 31992 5956 31996 6012
rect 31996 5956 32052 6012
rect 32052 5956 32056 6012
rect 31992 5952 32056 5956
rect 32072 6012 32136 6016
rect 32072 5956 32076 6012
rect 32076 5956 32132 6012
rect 32132 5956 32136 6012
rect 32072 5952 32136 5956
rect 32152 6012 32216 6016
rect 32152 5956 32156 6012
rect 32156 5956 32212 6012
rect 32212 5956 32216 6012
rect 32152 5952 32216 5956
rect 32232 6012 32296 6016
rect 32232 5956 32236 6012
rect 32236 5956 32292 6012
rect 32292 5956 32296 6012
rect 32232 5952 32296 5956
rect 37912 6012 37976 6016
rect 37912 5956 37916 6012
rect 37916 5956 37972 6012
rect 37972 5956 37976 6012
rect 37912 5952 37976 5956
rect 37992 6012 38056 6016
rect 37992 5956 37996 6012
rect 37996 5956 38052 6012
rect 38052 5956 38056 6012
rect 37992 5952 38056 5956
rect 38072 6012 38136 6016
rect 38072 5956 38076 6012
rect 38076 5956 38132 6012
rect 38132 5956 38136 6012
rect 38072 5952 38136 5956
rect 38152 6012 38216 6016
rect 38152 5956 38156 6012
rect 38156 5956 38212 6012
rect 38212 5956 38216 6012
rect 38152 5952 38216 5956
rect 38232 6012 38296 6016
rect 38232 5956 38236 6012
rect 38236 5956 38292 6012
rect 38292 5956 38296 6012
rect 38232 5952 38296 5956
rect 28028 5884 28092 5948
rect 4292 5612 4356 5676
rect 12572 5612 12636 5676
rect 19564 5672 19628 5676
rect 19564 5616 19614 5672
rect 19614 5616 19628 5672
rect 19564 5612 19628 5616
rect 21404 5612 21468 5676
rect 2652 5468 2716 5472
rect 2652 5412 2656 5468
rect 2656 5412 2712 5468
rect 2712 5412 2716 5468
rect 2652 5408 2716 5412
rect 2732 5468 2796 5472
rect 2732 5412 2736 5468
rect 2736 5412 2792 5468
rect 2792 5412 2796 5468
rect 2732 5408 2796 5412
rect 2812 5468 2876 5472
rect 2812 5412 2816 5468
rect 2816 5412 2872 5468
rect 2872 5412 2876 5468
rect 2812 5408 2876 5412
rect 2892 5468 2956 5472
rect 2892 5412 2896 5468
rect 2896 5412 2952 5468
rect 2952 5412 2956 5468
rect 2892 5408 2956 5412
rect 2972 5468 3036 5472
rect 2972 5412 2976 5468
rect 2976 5412 3032 5468
rect 3032 5412 3036 5468
rect 2972 5408 3036 5412
rect 8652 5468 8716 5472
rect 8652 5412 8656 5468
rect 8656 5412 8712 5468
rect 8712 5412 8716 5468
rect 8652 5408 8716 5412
rect 8732 5468 8796 5472
rect 8732 5412 8736 5468
rect 8736 5412 8792 5468
rect 8792 5412 8796 5468
rect 8732 5408 8796 5412
rect 8812 5468 8876 5472
rect 8812 5412 8816 5468
rect 8816 5412 8872 5468
rect 8872 5412 8876 5468
rect 8812 5408 8876 5412
rect 8892 5468 8956 5472
rect 8892 5412 8896 5468
rect 8896 5412 8952 5468
rect 8952 5412 8956 5468
rect 8892 5408 8956 5412
rect 8972 5468 9036 5472
rect 8972 5412 8976 5468
rect 8976 5412 9032 5468
rect 9032 5412 9036 5468
rect 8972 5408 9036 5412
rect 14652 5468 14716 5472
rect 14652 5412 14656 5468
rect 14656 5412 14712 5468
rect 14712 5412 14716 5468
rect 14652 5408 14716 5412
rect 14732 5468 14796 5472
rect 14732 5412 14736 5468
rect 14736 5412 14792 5468
rect 14792 5412 14796 5468
rect 14732 5408 14796 5412
rect 14812 5468 14876 5472
rect 14812 5412 14816 5468
rect 14816 5412 14872 5468
rect 14872 5412 14876 5468
rect 14812 5408 14876 5412
rect 14892 5468 14956 5472
rect 14892 5412 14896 5468
rect 14896 5412 14952 5468
rect 14952 5412 14956 5468
rect 14892 5408 14956 5412
rect 14972 5468 15036 5472
rect 14972 5412 14976 5468
rect 14976 5412 15032 5468
rect 15032 5412 15036 5468
rect 14972 5408 15036 5412
rect 20652 5468 20716 5472
rect 20652 5412 20656 5468
rect 20656 5412 20712 5468
rect 20712 5412 20716 5468
rect 20652 5408 20716 5412
rect 20732 5468 20796 5472
rect 20732 5412 20736 5468
rect 20736 5412 20792 5468
rect 20792 5412 20796 5468
rect 20732 5408 20796 5412
rect 20812 5468 20876 5472
rect 20812 5412 20816 5468
rect 20816 5412 20872 5468
rect 20872 5412 20876 5468
rect 20812 5408 20876 5412
rect 20892 5468 20956 5472
rect 20892 5412 20896 5468
rect 20896 5412 20952 5468
rect 20952 5412 20956 5468
rect 20892 5408 20956 5412
rect 20972 5468 21036 5472
rect 20972 5412 20976 5468
rect 20976 5412 21032 5468
rect 21032 5412 21036 5468
rect 20972 5408 21036 5412
rect 20484 5340 20548 5404
rect 27660 5476 27724 5540
rect 26652 5468 26716 5472
rect 26652 5412 26656 5468
rect 26656 5412 26712 5468
rect 26712 5412 26716 5468
rect 26652 5408 26716 5412
rect 26732 5468 26796 5472
rect 26732 5412 26736 5468
rect 26736 5412 26792 5468
rect 26792 5412 26796 5468
rect 26732 5408 26796 5412
rect 26812 5468 26876 5472
rect 26812 5412 26816 5468
rect 26816 5412 26872 5468
rect 26872 5412 26876 5468
rect 26812 5408 26876 5412
rect 26892 5468 26956 5472
rect 26892 5412 26896 5468
rect 26896 5412 26952 5468
rect 26952 5412 26956 5468
rect 26892 5408 26956 5412
rect 26972 5468 27036 5472
rect 26972 5412 26976 5468
rect 26976 5412 27032 5468
rect 27032 5412 27036 5468
rect 26972 5408 27036 5412
rect 32652 5468 32716 5472
rect 32652 5412 32656 5468
rect 32656 5412 32712 5468
rect 32712 5412 32716 5468
rect 32652 5408 32716 5412
rect 32732 5468 32796 5472
rect 32732 5412 32736 5468
rect 32736 5412 32792 5468
rect 32792 5412 32796 5468
rect 32732 5408 32796 5412
rect 32812 5468 32876 5472
rect 32812 5412 32816 5468
rect 32816 5412 32872 5468
rect 32872 5412 32876 5468
rect 32812 5408 32876 5412
rect 32892 5468 32956 5472
rect 32892 5412 32896 5468
rect 32896 5412 32952 5468
rect 32952 5412 32956 5468
rect 32892 5408 32956 5412
rect 32972 5468 33036 5472
rect 32972 5412 32976 5468
rect 32976 5412 33032 5468
rect 33032 5412 33036 5468
rect 32972 5408 33036 5412
rect 38652 5468 38716 5472
rect 38652 5412 38656 5468
rect 38656 5412 38712 5468
rect 38712 5412 38716 5468
rect 38652 5408 38716 5412
rect 38732 5468 38796 5472
rect 38732 5412 38736 5468
rect 38736 5412 38792 5468
rect 38792 5412 38796 5468
rect 38732 5408 38796 5412
rect 38812 5468 38876 5472
rect 38812 5412 38816 5468
rect 38816 5412 38872 5468
rect 38872 5412 38876 5468
rect 38812 5408 38876 5412
rect 38892 5468 38956 5472
rect 38892 5412 38896 5468
rect 38896 5412 38952 5468
rect 38952 5412 38956 5468
rect 38892 5408 38956 5412
rect 38972 5468 39036 5472
rect 38972 5412 38976 5468
rect 38976 5412 39032 5468
rect 39032 5412 39036 5468
rect 38972 5408 39036 5412
rect 27844 5204 27908 5268
rect 13676 4932 13740 4996
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 14152 4924 14216 4928
rect 14152 4868 14156 4924
rect 14156 4868 14212 4924
rect 14212 4868 14216 4924
rect 14152 4864 14216 4868
rect 14232 4924 14296 4928
rect 14232 4868 14236 4924
rect 14236 4868 14292 4924
rect 14292 4868 14296 4924
rect 14232 4864 14296 4868
rect 19912 4924 19976 4928
rect 19912 4868 19916 4924
rect 19916 4868 19972 4924
rect 19972 4868 19976 4924
rect 19912 4864 19976 4868
rect 19992 4924 20056 4928
rect 19992 4868 19996 4924
rect 19996 4868 20052 4924
rect 20052 4868 20056 4924
rect 19992 4864 20056 4868
rect 20072 4924 20136 4928
rect 20072 4868 20076 4924
rect 20076 4868 20132 4924
rect 20132 4868 20136 4924
rect 20072 4864 20136 4868
rect 20152 4924 20216 4928
rect 20152 4868 20156 4924
rect 20156 4868 20212 4924
rect 20212 4868 20216 4924
rect 20152 4864 20216 4868
rect 20232 4924 20296 4928
rect 20232 4868 20236 4924
rect 20236 4868 20292 4924
rect 20292 4868 20296 4924
rect 20232 4864 20296 4868
rect 15148 4796 15212 4860
rect 26372 4932 26436 4996
rect 25912 4924 25976 4928
rect 25912 4868 25916 4924
rect 25916 4868 25972 4924
rect 25972 4868 25976 4924
rect 25912 4864 25976 4868
rect 25992 4924 26056 4928
rect 25992 4868 25996 4924
rect 25996 4868 26052 4924
rect 26052 4868 26056 4924
rect 25992 4864 26056 4868
rect 26072 4924 26136 4928
rect 26072 4868 26076 4924
rect 26076 4868 26132 4924
rect 26132 4868 26136 4924
rect 26072 4864 26136 4868
rect 26152 4924 26216 4928
rect 26152 4868 26156 4924
rect 26156 4868 26212 4924
rect 26212 4868 26216 4924
rect 26152 4864 26216 4868
rect 26232 4924 26296 4928
rect 26232 4868 26236 4924
rect 26236 4868 26292 4924
rect 26292 4868 26296 4924
rect 26232 4864 26296 4868
rect 31912 4924 31976 4928
rect 31912 4868 31916 4924
rect 31916 4868 31972 4924
rect 31972 4868 31976 4924
rect 31912 4864 31976 4868
rect 31992 4924 32056 4928
rect 31992 4868 31996 4924
rect 31996 4868 32052 4924
rect 32052 4868 32056 4924
rect 31992 4864 32056 4868
rect 32072 4924 32136 4928
rect 32072 4868 32076 4924
rect 32076 4868 32132 4924
rect 32132 4868 32136 4924
rect 32072 4864 32136 4868
rect 32152 4924 32216 4928
rect 32152 4868 32156 4924
rect 32156 4868 32212 4924
rect 32212 4868 32216 4924
rect 32152 4864 32216 4868
rect 32232 4924 32296 4928
rect 32232 4868 32236 4924
rect 32236 4868 32292 4924
rect 32292 4868 32296 4924
rect 32232 4864 32296 4868
rect 37912 4924 37976 4928
rect 37912 4868 37916 4924
rect 37916 4868 37972 4924
rect 37972 4868 37976 4924
rect 37912 4864 37976 4868
rect 37992 4924 38056 4928
rect 37992 4868 37996 4924
rect 37996 4868 38052 4924
rect 38052 4868 38056 4924
rect 37992 4864 38056 4868
rect 38072 4924 38136 4928
rect 38072 4868 38076 4924
rect 38076 4868 38132 4924
rect 38132 4868 38136 4924
rect 38072 4864 38136 4868
rect 38152 4924 38216 4928
rect 38152 4868 38156 4924
rect 38156 4868 38212 4924
rect 38212 4868 38216 4924
rect 38152 4864 38216 4868
rect 38232 4924 38296 4928
rect 38232 4868 38236 4924
rect 38236 4868 38292 4924
rect 38292 4868 38296 4924
rect 38232 4864 38296 4868
rect 35020 4856 35084 4860
rect 35020 4800 35070 4856
rect 35070 4800 35084 4856
rect 35020 4796 35084 4800
rect 28028 4660 28092 4724
rect 13492 4388 13556 4452
rect 26372 4388 26436 4452
rect 2652 4380 2716 4384
rect 2652 4324 2656 4380
rect 2656 4324 2712 4380
rect 2712 4324 2716 4380
rect 2652 4320 2716 4324
rect 2732 4380 2796 4384
rect 2732 4324 2736 4380
rect 2736 4324 2792 4380
rect 2792 4324 2796 4380
rect 2732 4320 2796 4324
rect 2812 4380 2876 4384
rect 2812 4324 2816 4380
rect 2816 4324 2872 4380
rect 2872 4324 2876 4380
rect 2812 4320 2876 4324
rect 2892 4380 2956 4384
rect 2892 4324 2896 4380
rect 2896 4324 2952 4380
rect 2952 4324 2956 4380
rect 2892 4320 2956 4324
rect 2972 4380 3036 4384
rect 2972 4324 2976 4380
rect 2976 4324 3032 4380
rect 3032 4324 3036 4380
rect 2972 4320 3036 4324
rect 8652 4380 8716 4384
rect 8652 4324 8656 4380
rect 8656 4324 8712 4380
rect 8712 4324 8716 4380
rect 8652 4320 8716 4324
rect 8732 4380 8796 4384
rect 8732 4324 8736 4380
rect 8736 4324 8792 4380
rect 8792 4324 8796 4380
rect 8732 4320 8796 4324
rect 8812 4380 8876 4384
rect 8812 4324 8816 4380
rect 8816 4324 8872 4380
rect 8872 4324 8876 4380
rect 8812 4320 8876 4324
rect 8892 4380 8956 4384
rect 8892 4324 8896 4380
rect 8896 4324 8952 4380
rect 8952 4324 8956 4380
rect 8892 4320 8956 4324
rect 8972 4380 9036 4384
rect 8972 4324 8976 4380
rect 8976 4324 9032 4380
rect 9032 4324 9036 4380
rect 8972 4320 9036 4324
rect 14652 4380 14716 4384
rect 14652 4324 14656 4380
rect 14656 4324 14712 4380
rect 14712 4324 14716 4380
rect 14652 4320 14716 4324
rect 14732 4380 14796 4384
rect 14732 4324 14736 4380
rect 14736 4324 14792 4380
rect 14792 4324 14796 4380
rect 14732 4320 14796 4324
rect 14812 4380 14876 4384
rect 14812 4324 14816 4380
rect 14816 4324 14872 4380
rect 14872 4324 14876 4380
rect 14812 4320 14876 4324
rect 14892 4380 14956 4384
rect 14892 4324 14896 4380
rect 14896 4324 14952 4380
rect 14952 4324 14956 4380
rect 14892 4320 14956 4324
rect 14972 4380 15036 4384
rect 14972 4324 14976 4380
rect 14976 4324 15032 4380
rect 15032 4324 15036 4380
rect 14972 4320 15036 4324
rect 20652 4380 20716 4384
rect 20652 4324 20656 4380
rect 20656 4324 20712 4380
rect 20712 4324 20716 4380
rect 20652 4320 20716 4324
rect 20732 4380 20796 4384
rect 20732 4324 20736 4380
rect 20736 4324 20792 4380
rect 20792 4324 20796 4380
rect 20732 4320 20796 4324
rect 20812 4380 20876 4384
rect 20812 4324 20816 4380
rect 20816 4324 20872 4380
rect 20872 4324 20876 4380
rect 20812 4320 20876 4324
rect 20892 4380 20956 4384
rect 20892 4324 20896 4380
rect 20896 4324 20952 4380
rect 20952 4324 20956 4380
rect 20892 4320 20956 4324
rect 20972 4380 21036 4384
rect 20972 4324 20976 4380
rect 20976 4324 21032 4380
rect 21032 4324 21036 4380
rect 20972 4320 21036 4324
rect 26652 4380 26716 4384
rect 26652 4324 26656 4380
rect 26656 4324 26712 4380
rect 26712 4324 26716 4380
rect 26652 4320 26716 4324
rect 26732 4380 26796 4384
rect 26732 4324 26736 4380
rect 26736 4324 26792 4380
rect 26792 4324 26796 4380
rect 26732 4320 26796 4324
rect 26812 4380 26876 4384
rect 26812 4324 26816 4380
rect 26816 4324 26872 4380
rect 26872 4324 26876 4380
rect 26812 4320 26876 4324
rect 26892 4380 26956 4384
rect 26892 4324 26896 4380
rect 26896 4324 26952 4380
rect 26952 4324 26956 4380
rect 26892 4320 26956 4324
rect 26972 4380 27036 4384
rect 26972 4324 26976 4380
rect 26976 4324 27032 4380
rect 27032 4324 27036 4380
rect 26972 4320 27036 4324
rect 17908 4252 17972 4316
rect 21220 4312 21284 4316
rect 32652 4380 32716 4384
rect 32652 4324 32656 4380
rect 32656 4324 32712 4380
rect 32712 4324 32716 4380
rect 32652 4320 32716 4324
rect 32732 4380 32796 4384
rect 32732 4324 32736 4380
rect 32736 4324 32792 4380
rect 32792 4324 32796 4380
rect 32732 4320 32796 4324
rect 32812 4380 32876 4384
rect 32812 4324 32816 4380
rect 32816 4324 32872 4380
rect 32872 4324 32876 4380
rect 32812 4320 32876 4324
rect 32892 4380 32956 4384
rect 32892 4324 32896 4380
rect 32896 4324 32952 4380
rect 32952 4324 32956 4380
rect 32892 4320 32956 4324
rect 32972 4380 33036 4384
rect 32972 4324 32976 4380
rect 32976 4324 33032 4380
rect 33032 4324 33036 4380
rect 32972 4320 33036 4324
rect 38652 4380 38716 4384
rect 38652 4324 38656 4380
rect 38656 4324 38712 4380
rect 38712 4324 38716 4380
rect 38652 4320 38716 4324
rect 38732 4380 38796 4384
rect 38732 4324 38736 4380
rect 38736 4324 38792 4380
rect 38792 4324 38796 4380
rect 38732 4320 38796 4324
rect 38812 4380 38876 4384
rect 38812 4324 38816 4380
rect 38816 4324 38872 4380
rect 38872 4324 38876 4380
rect 38812 4320 38876 4324
rect 38892 4380 38956 4384
rect 38892 4324 38896 4380
rect 38896 4324 38952 4380
rect 38952 4324 38956 4380
rect 38892 4320 38956 4324
rect 38972 4380 39036 4384
rect 38972 4324 38976 4380
rect 38976 4324 39032 4380
rect 39032 4324 39036 4380
rect 38972 4320 39036 4324
rect 21220 4256 21234 4312
rect 21234 4256 21284 4312
rect 21220 4252 21284 4256
rect 21772 4116 21836 4180
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 14152 3836 14216 3840
rect 14152 3780 14156 3836
rect 14156 3780 14212 3836
rect 14212 3780 14216 3836
rect 14152 3776 14216 3780
rect 14232 3836 14296 3840
rect 14232 3780 14236 3836
rect 14236 3780 14292 3836
rect 14292 3780 14296 3836
rect 14232 3776 14296 3780
rect 33916 3904 33980 3908
rect 33916 3848 33966 3904
rect 33966 3848 33980 3904
rect 33916 3844 33980 3848
rect 19912 3836 19976 3840
rect 19912 3780 19916 3836
rect 19916 3780 19972 3836
rect 19972 3780 19976 3836
rect 19912 3776 19976 3780
rect 19992 3836 20056 3840
rect 19992 3780 19996 3836
rect 19996 3780 20052 3836
rect 20052 3780 20056 3836
rect 19992 3776 20056 3780
rect 20072 3836 20136 3840
rect 20072 3780 20076 3836
rect 20076 3780 20132 3836
rect 20132 3780 20136 3836
rect 20072 3776 20136 3780
rect 20152 3836 20216 3840
rect 20152 3780 20156 3836
rect 20156 3780 20212 3836
rect 20212 3780 20216 3836
rect 20152 3776 20216 3780
rect 20232 3836 20296 3840
rect 20232 3780 20236 3836
rect 20236 3780 20292 3836
rect 20292 3780 20296 3836
rect 20232 3776 20296 3780
rect 25912 3836 25976 3840
rect 25912 3780 25916 3836
rect 25916 3780 25972 3836
rect 25972 3780 25976 3836
rect 25912 3776 25976 3780
rect 25992 3836 26056 3840
rect 25992 3780 25996 3836
rect 25996 3780 26052 3836
rect 26052 3780 26056 3836
rect 25992 3776 26056 3780
rect 26072 3836 26136 3840
rect 26072 3780 26076 3836
rect 26076 3780 26132 3836
rect 26132 3780 26136 3836
rect 26072 3776 26136 3780
rect 26152 3836 26216 3840
rect 26152 3780 26156 3836
rect 26156 3780 26212 3836
rect 26212 3780 26216 3836
rect 26152 3776 26216 3780
rect 26232 3836 26296 3840
rect 26232 3780 26236 3836
rect 26236 3780 26292 3836
rect 26292 3780 26296 3836
rect 26232 3776 26296 3780
rect 31912 3836 31976 3840
rect 31912 3780 31916 3836
rect 31916 3780 31972 3836
rect 31972 3780 31976 3836
rect 31912 3776 31976 3780
rect 31992 3836 32056 3840
rect 31992 3780 31996 3836
rect 31996 3780 32052 3836
rect 32052 3780 32056 3836
rect 31992 3776 32056 3780
rect 32072 3836 32136 3840
rect 32072 3780 32076 3836
rect 32076 3780 32132 3836
rect 32132 3780 32136 3836
rect 32072 3776 32136 3780
rect 32152 3836 32216 3840
rect 32152 3780 32156 3836
rect 32156 3780 32212 3836
rect 32212 3780 32216 3836
rect 32152 3776 32216 3780
rect 32232 3836 32296 3840
rect 32232 3780 32236 3836
rect 32236 3780 32292 3836
rect 32292 3780 32296 3836
rect 32232 3776 32296 3780
rect 37912 3836 37976 3840
rect 37912 3780 37916 3836
rect 37916 3780 37972 3836
rect 37972 3780 37976 3836
rect 37912 3776 37976 3780
rect 37992 3836 38056 3840
rect 37992 3780 37996 3836
rect 37996 3780 38052 3836
rect 38052 3780 38056 3836
rect 37992 3776 38056 3780
rect 38072 3836 38136 3840
rect 38072 3780 38076 3836
rect 38076 3780 38132 3836
rect 38132 3780 38136 3836
rect 38072 3776 38136 3780
rect 38152 3836 38216 3840
rect 38152 3780 38156 3836
rect 38156 3780 38212 3836
rect 38212 3780 38216 3836
rect 38152 3776 38216 3780
rect 38232 3836 38296 3840
rect 38232 3780 38236 3836
rect 38236 3780 38292 3836
rect 38292 3780 38296 3836
rect 38232 3776 38296 3780
rect 15332 3708 15396 3772
rect 15516 3708 15580 3772
rect 21588 3436 21652 3500
rect 2652 3292 2716 3296
rect 2652 3236 2656 3292
rect 2656 3236 2712 3292
rect 2712 3236 2716 3292
rect 2652 3232 2716 3236
rect 2732 3292 2796 3296
rect 2732 3236 2736 3292
rect 2736 3236 2792 3292
rect 2792 3236 2796 3292
rect 2732 3232 2796 3236
rect 2812 3292 2876 3296
rect 2812 3236 2816 3292
rect 2816 3236 2872 3292
rect 2872 3236 2876 3292
rect 2812 3232 2876 3236
rect 2892 3292 2956 3296
rect 2892 3236 2896 3292
rect 2896 3236 2952 3292
rect 2952 3236 2956 3292
rect 2892 3232 2956 3236
rect 2972 3292 3036 3296
rect 2972 3236 2976 3292
rect 2976 3236 3032 3292
rect 3032 3236 3036 3292
rect 2972 3232 3036 3236
rect 8652 3292 8716 3296
rect 8652 3236 8656 3292
rect 8656 3236 8712 3292
rect 8712 3236 8716 3292
rect 8652 3232 8716 3236
rect 8732 3292 8796 3296
rect 8732 3236 8736 3292
rect 8736 3236 8792 3292
rect 8792 3236 8796 3292
rect 8732 3232 8796 3236
rect 8812 3292 8876 3296
rect 8812 3236 8816 3292
rect 8816 3236 8872 3292
rect 8872 3236 8876 3292
rect 8812 3232 8876 3236
rect 8892 3292 8956 3296
rect 8892 3236 8896 3292
rect 8896 3236 8952 3292
rect 8952 3236 8956 3292
rect 8892 3232 8956 3236
rect 8972 3292 9036 3296
rect 8972 3236 8976 3292
rect 8976 3236 9032 3292
rect 9032 3236 9036 3292
rect 8972 3232 9036 3236
rect 14652 3292 14716 3296
rect 14652 3236 14656 3292
rect 14656 3236 14712 3292
rect 14712 3236 14716 3292
rect 14652 3232 14716 3236
rect 14732 3292 14796 3296
rect 14732 3236 14736 3292
rect 14736 3236 14792 3292
rect 14792 3236 14796 3292
rect 14732 3232 14796 3236
rect 14812 3292 14876 3296
rect 14812 3236 14816 3292
rect 14816 3236 14872 3292
rect 14872 3236 14876 3292
rect 14812 3232 14876 3236
rect 14892 3292 14956 3296
rect 14892 3236 14896 3292
rect 14896 3236 14952 3292
rect 14952 3236 14956 3292
rect 14892 3232 14956 3236
rect 14972 3292 15036 3296
rect 14972 3236 14976 3292
rect 14976 3236 15032 3292
rect 15032 3236 15036 3292
rect 14972 3232 15036 3236
rect 20652 3292 20716 3296
rect 20652 3236 20656 3292
rect 20656 3236 20712 3292
rect 20712 3236 20716 3292
rect 20652 3232 20716 3236
rect 20732 3292 20796 3296
rect 20732 3236 20736 3292
rect 20736 3236 20792 3292
rect 20792 3236 20796 3292
rect 20732 3232 20796 3236
rect 20812 3292 20876 3296
rect 20812 3236 20816 3292
rect 20816 3236 20872 3292
rect 20872 3236 20876 3292
rect 20812 3232 20876 3236
rect 20892 3292 20956 3296
rect 20892 3236 20896 3292
rect 20896 3236 20952 3292
rect 20952 3236 20956 3292
rect 20892 3232 20956 3236
rect 20972 3292 21036 3296
rect 20972 3236 20976 3292
rect 20976 3236 21032 3292
rect 21032 3236 21036 3292
rect 20972 3232 21036 3236
rect 16988 3164 17052 3228
rect 17356 3164 17420 3228
rect 19012 3164 19076 3228
rect 26652 3292 26716 3296
rect 26652 3236 26656 3292
rect 26656 3236 26712 3292
rect 26712 3236 26716 3292
rect 26652 3232 26716 3236
rect 26732 3292 26796 3296
rect 26732 3236 26736 3292
rect 26736 3236 26792 3292
rect 26792 3236 26796 3292
rect 26732 3232 26796 3236
rect 26812 3292 26876 3296
rect 26812 3236 26816 3292
rect 26816 3236 26872 3292
rect 26872 3236 26876 3292
rect 26812 3232 26876 3236
rect 26892 3292 26956 3296
rect 26892 3236 26896 3292
rect 26896 3236 26952 3292
rect 26952 3236 26956 3292
rect 26892 3232 26956 3236
rect 26972 3292 27036 3296
rect 26972 3236 26976 3292
rect 26976 3236 27032 3292
rect 27032 3236 27036 3292
rect 26972 3232 27036 3236
rect 32652 3292 32716 3296
rect 32652 3236 32656 3292
rect 32656 3236 32712 3292
rect 32712 3236 32716 3292
rect 32652 3232 32716 3236
rect 32732 3292 32796 3296
rect 32732 3236 32736 3292
rect 32736 3236 32792 3292
rect 32792 3236 32796 3292
rect 32732 3232 32796 3236
rect 32812 3292 32876 3296
rect 32812 3236 32816 3292
rect 32816 3236 32872 3292
rect 32872 3236 32876 3292
rect 32812 3232 32876 3236
rect 32892 3292 32956 3296
rect 32892 3236 32896 3292
rect 32896 3236 32952 3292
rect 32952 3236 32956 3292
rect 32892 3232 32956 3236
rect 32972 3292 33036 3296
rect 32972 3236 32976 3292
rect 32976 3236 33032 3292
rect 33032 3236 33036 3292
rect 32972 3232 33036 3236
rect 38652 3292 38716 3296
rect 38652 3236 38656 3292
rect 38656 3236 38712 3292
rect 38712 3236 38716 3292
rect 38652 3232 38716 3236
rect 38732 3292 38796 3296
rect 38732 3236 38736 3292
rect 38736 3236 38792 3292
rect 38792 3236 38796 3292
rect 38732 3232 38796 3236
rect 38812 3292 38876 3296
rect 38812 3236 38816 3292
rect 38816 3236 38872 3292
rect 38872 3236 38876 3292
rect 38812 3232 38876 3236
rect 38892 3292 38956 3296
rect 38892 3236 38896 3292
rect 38896 3236 38952 3292
rect 38952 3236 38956 3292
rect 38892 3232 38956 3236
rect 38972 3292 39036 3296
rect 38972 3236 38976 3292
rect 38976 3236 39032 3292
rect 39032 3236 39036 3292
rect 38972 3232 39036 3236
rect 32444 3224 32508 3228
rect 32444 3168 32458 3224
rect 32458 3168 32508 3224
rect 32444 3164 32508 3168
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 9444 2892 9508 2956
rect 10916 2892 10980 2956
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 14152 2748 14216 2752
rect 14152 2692 14156 2748
rect 14156 2692 14212 2748
rect 14212 2692 14216 2748
rect 14152 2688 14216 2692
rect 14232 2748 14296 2752
rect 14232 2692 14236 2748
rect 14236 2692 14292 2748
rect 14292 2692 14296 2748
rect 14232 2688 14296 2692
rect 19912 2748 19976 2752
rect 19912 2692 19916 2748
rect 19916 2692 19972 2748
rect 19972 2692 19976 2748
rect 19912 2688 19976 2692
rect 19992 2748 20056 2752
rect 19992 2692 19996 2748
rect 19996 2692 20052 2748
rect 20052 2692 20056 2748
rect 19992 2688 20056 2692
rect 20072 2748 20136 2752
rect 20072 2692 20076 2748
rect 20076 2692 20132 2748
rect 20132 2692 20136 2748
rect 20072 2688 20136 2692
rect 20152 2748 20216 2752
rect 20152 2692 20156 2748
rect 20156 2692 20212 2748
rect 20212 2692 20216 2748
rect 20152 2688 20216 2692
rect 20232 2748 20296 2752
rect 20232 2692 20236 2748
rect 20236 2692 20292 2748
rect 20292 2692 20296 2748
rect 20232 2688 20296 2692
rect 25912 2748 25976 2752
rect 25912 2692 25916 2748
rect 25916 2692 25972 2748
rect 25972 2692 25976 2748
rect 25912 2688 25976 2692
rect 25992 2748 26056 2752
rect 25992 2692 25996 2748
rect 25996 2692 26052 2748
rect 26052 2692 26056 2748
rect 25992 2688 26056 2692
rect 26072 2748 26136 2752
rect 26072 2692 26076 2748
rect 26076 2692 26132 2748
rect 26132 2692 26136 2748
rect 26072 2688 26136 2692
rect 26152 2748 26216 2752
rect 26152 2692 26156 2748
rect 26156 2692 26212 2748
rect 26212 2692 26216 2748
rect 26152 2688 26216 2692
rect 26232 2748 26296 2752
rect 26232 2692 26236 2748
rect 26236 2692 26292 2748
rect 26292 2692 26296 2748
rect 26232 2688 26296 2692
rect 31912 2748 31976 2752
rect 31912 2692 31916 2748
rect 31916 2692 31972 2748
rect 31972 2692 31976 2748
rect 31912 2688 31976 2692
rect 31992 2748 32056 2752
rect 31992 2692 31996 2748
rect 31996 2692 32052 2748
rect 32052 2692 32056 2748
rect 31992 2688 32056 2692
rect 32072 2748 32136 2752
rect 32072 2692 32076 2748
rect 32076 2692 32132 2748
rect 32132 2692 32136 2748
rect 32072 2688 32136 2692
rect 32152 2748 32216 2752
rect 32152 2692 32156 2748
rect 32156 2692 32212 2748
rect 32212 2692 32216 2748
rect 32152 2688 32216 2692
rect 32232 2748 32296 2752
rect 32232 2692 32236 2748
rect 32236 2692 32292 2748
rect 32292 2692 32296 2748
rect 32232 2688 32296 2692
rect 37912 2748 37976 2752
rect 37912 2692 37916 2748
rect 37916 2692 37972 2748
rect 37972 2692 37976 2748
rect 37912 2688 37976 2692
rect 37992 2748 38056 2752
rect 37992 2692 37996 2748
rect 37996 2692 38052 2748
rect 38052 2692 38056 2748
rect 37992 2688 38056 2692
rect 38072 2748 38136 2752
rect 38072 2692 38076 2748
rect 38076 2692 38132 2748
rect 38132 2692 38136 2748
rect 38072 2688 38136 2692
rect 38152 2748 38216 2752
rect 38152 2692 38156 2748
rect 38156 2692 38212 2748
rect 38212 2692 38216 2748
rect 38152 2688 38216 2692
rect 38232 2748 38296 2752
rect 38232 2692 38236 2748
rect 38236 2692 38292 2748
rect 38292 2692 38296 2748
rect 38232 2688 38296 2692
rect 10732 2484 10796 2548
rect 2652 2204 2716 2208
rect 2652 2148 2656 2204
rect 2656 2148 2712 2204
rect 2712 2148 2716 2204
rect 2652 2144 2716 2148
rect 2732 2204 2796 2208
rect 2732 2148 2736 2204
rect 2736 2148 2792 2204
rect 2792 2148 2796 2204
rect 2732 2144 2796 2148
rect 2812 2204 2876 2208
rect 2812 2148 2816 2204
rect 2816 2148 2872 2204
rect 2872 2148 2876 2204
rect 2812 2144 2876 2148
rect 2892 2204 2956 2208
rect 2892 2148 2896 2204
rect 2896 2148 2952 2204
rect 2952 2148 2956 2204
rect 2892 2144 2956 2148
rect 2972 2204 3036 2208
rect 2972 2148 2976 2204
rect 2976 2148 3032 2204
rect 3032 2148 3036 2204
rect 2972 2144 3036 2148
rect 8652 2204 8716 2208
rect 8652 2148 8656 2204
rect 8656 2148 8712 2204
rect 8712 2148 8716 2204
rect 8652 2144 8716 2148
rect 8732 2204 8796 2208
rect 8732 2148 8736 2204
rect 8736 2148 8792 2204
rect 8792 2148 8796 2204
rect 8732 2144 8796 2148
rect 8812 2204 8876 2208
rect 8812 2148 8816 2204
rect 8816 2148 8872 2204
rect 8872 2148 8876 2204
rect 8812 2144 8876 2148
rect 8892 2204 8956 2208
rect 8892 2148 8896 2204
rect 8896 2148 8952 2204
rect 8952 2148 8956 2204
rect 8892 2144 8956 2148
rect 8972 2204 9036 2208
rect 8972 2148 8976 2204
rect 8976 2148 9032 2204
rect 9032 2148 9036 2204
rect 8972 2144 9036 2148
rect 14652 2204 14716 2208
rect 14652 2148 14656 2204
rect 14656 2148 14712 2204
rect 14712 2148 14716 2204
rect 14652 2144 14716 2148
rect 14732 2204 14796 2208
rect 14732 2148 14736 2204
rect 14736 2148 14792 2204
rect 14792 2148 14796 2204
rect 14732 2144 14796 2148
rect 14812 2204 14876 2208
rect 14812 2148 14816 2204
rect 14816 2148 14872 2204
rect 14872 2148 14876 2204
rect 14812 2144 14876 2148
rect 14892 2204 14956 2208
rect 14892 2148 14896 2204
rect 14896 2148 14952 2204
rect 14952 2148 14956 2204
rect 14892 2144 14956 2148
rect 14972 2204 15036 2208
rect 14972 2148 14976 2204
rect 14976 2148 15032 2204
rect 15032 2148 15036 2204
rect 14972 2144 15036 2148
rect 20652 2204 20716 2208
rect 20652 2148 20656 2204
rect 20656 2148 20712 2204
rect 20712 2148 20716 2204
rect 20652 2144 20716 2148
rect 20732 2204 20796 2208
rect 20732 2148 20736 2204
rect 20736 2148 20792 2204
rect 20792 2148 20796 2204
rect 20732 2144 20796 2148
rect 20812 2204 20876 2208
rect 20812 2148 20816 2204
rect 20816 2148 20872 2204
rect 20872 2148 20876 2204
rect 20812 2144 20876 2148
rect 20892 2204 20956 2208
rect 20892 2148 20896 2204
rect 20896 2148 20952 2204
rect 20952 2148 20956 2204
rect 20892 2144 20956 2148
rect 20972 2204 21036 2208
rect 20972 2148 20976 2204
rect 20976 2148 21032 2204
rect 21032 2148 21036 2204
rect 20972 2144 21036 2148
rect 26652 2204 26716 2208
rect 26652 2148 26656 2204
rect 26656 2148 26712 2204
rect 26712 2148 26716 2204
rect 26652 2144 26716 2148
rect 26732 2204 26796 2208
rect 26732 2148 26736 2204
rect 26736 2148 26792 2204
rect 26792 2148 26796 2204
rect 26732 2144 26796 2148
rect 26812 2204 26876 2208
rect 26812 2148 26816 2204
rect 26816 2148 26872 2204
rect 26872 2148 26876 2204
rect 26812 2144 26876 2148
rect 26892 2204 26956 2208
rect 26892 2148 26896 2204
rect 26896 2148 26952 2204
rect 26952 2148 26956 2204
rect 26892 2144 26956 2148
rect 26972 2204 27036 2208
rect 26972 2148 26976 2204
rect 26976 2148 27032 2204
rect 27032 2148 27036 2204
rect 26972 2144 27036 2148
rect 32652 2204 32716 2208
rect 32652 2148 32656 2204
rect 32656 2148 32712 2204
rect 32712 2148 32716 2204
rect 32652 2144 32716 2148
rect 32732 2204 32796 2208
rect 32732 2148 32736 2204
rect 32736 2148 32792 2204
rect 32792 2148 32796 2204
rect 32732 2144 32796 2148
rect 32812 2204 32876 2208
rect 32812 2148 32816 2204
rect 32816 2148 32872 2204
rect 32872 2148 32876 2204
rect 32812 2144 32876 2148
rect 32892 2204 32956 2208
rect 32892 2148 32896 2204
rect 32896 2148 32952 2204
rect 32952 2148 32956 2204
rect 32892 2144 32956 2148
rect 32972 2204 33036 2208
rect 32972 2148 32976 2204
rect 32976 2148 33032 2204
rect 33032 2148 33036 2204
rect 32972 2144 33036 2148
rect 38652 2204 38716 2208
rect 38652 2148 38656 2204
rect 38656 2148 38712 2204
rect 38712 2148 38716 2204
rect 38652 2144 38716 2148
rect 38732 2204 38796 2208
rect 38732 2148 38736 2204
rect 38736 2148 38792 2204
rect 38792 2148 38796 2204
rect 38732 2144 38796 2148
rect 38812 2204 38876 2208
rect 38812 2148 38816 2204
rect 38816 2148 38872 2204
rect 38872 2148 38876 2204
rect 38812 2144 38876 2148
rect 38892 2204 38956 2208
rect 38892 2148 38896 2204
rect 38896 2148 38952 2204
rect 38952 2148 38956 2204
rect 38892 2144 38956 2148
rect 38972 2204 39036 2208
rect 38972 2148 38976 2204
rect 38976 2148 39032 2204
rect 39032 2148 39036 2204
rect 38972 2144 39036 2148
rect 19196 1804 19260 1868
rect 27844 1804 27908 1868
rect 10364 1260 10428 1324
<< metal4 >>
rect 1904 8192 2304 11250
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 2752 2304 3776
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 0 2304 2688
rect 2644 8736 3044 11250
rect 6315 10572 6381 10573
rect 6315 10508 6316 10572
rect 6380 10508 6381 10572
rect 6315 10507 6381 10508
rect 5947 10164 6013 10165
rect 5947 10100 5948 10164
rect 6012 10100 6013 10164
rect 5947 10099 6013 10100
rect 2644 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3044 8736
rect 2644 7648 3044 8672
rect 5950 7717 6010 10099
rect 6318 7717 6378 10507
rect 7904 8192 8304 11250
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 4291 7716 4357 7717
rect 4291 7652 4292 7716
rect 4356 7652 4357 7716
rect 4291 7651 4357 7652
rect 5947 7716 6013 7717
rect 5947 7652 5948 7716
rect 6012 7652 6013 7716
rect 5947 7651 6013 7652
rect 6315 7716 6381 7717
rect 6315 7652 6316 7716
rect 6380 7652 6381 7716
rect 6315 7651 6381 7652
rect 2644 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3044 7648
rect 2644 6560 3044 7584
rect 2644 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3044 6560
rect 2644 5472 3044 6496
rect 4294 5677 4354 7651
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 4291 5676 4357 5677
rect 4291 5612 4292 5676
rect 4356 5612 4357 5676
rect 4291 5611 4357 5612
rect 2644 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3044 5472
rect 2644 4384 3044 5408
rect 2644 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3044 4384
rect 2644 3296 3044 4320
rect 2644 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3044 3296
rect 2644 2208 3044 3232
rect 2644 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3044 2208
rect 2644 0 3044 2144
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 2752 8304 3776
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 0 8304 2688
rect 8644 8736 9044 11250
rect 10363 10436 10429 10437
rect 10363 10372 10364 10436
rect 10428 10372 10429 10436
rect 10363 10371 10429 10372
rect 8644 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9044 8736
rect 8644 7648 9044 8672
rect 8644 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9044 7648
rect 8644 6560 9044 7584
rect 8644 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9044 6560
rect 8644 5472 9044 6496
rect 9443 5812 9509 5813
rect 9443 5748 9444 5812
rect 9508 5748 9509 5812
rect 9443 5747 9509 5748
rect 8644 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9044 5472
rect 8644 4384 9044 5408
rect 8644 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9044 4384
rect 8644 3296 9044 4320
rect 8644 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9044 3296
rect 8644 2208 9044 3232
rect 9446 2957 9506 5747
rect 9443 2956 9509 2957
rect 9443 2892 9444 2956
rect 9508 2892 9509 2956
rect 9443 2891 9509 2892
rect 8644 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9044 2208
rect 8644 0 9044 2144
rect 10366 1325 10426 10371
rect 10731 8396 10797 8397
rect 10731 8332 10732 8396
rect 10796 8332 10797 8396
rect 10731 8331 10797 8332
rect 10734 2954 10794 8331
rect 13491 8260 13557 8261
rect 13491 8196 13492 8260
rect 13556 8196 13557 8260
rect 13491 8195 13557 8196
rect 12571 7580 12637 7581
rect 12571 7516 12572 7580
rect 12636 7516 12637 7580
rect 12571 7515 12637 7516
rect 12574 5677 12634 7515
rect 12571 5676 12637 5677
rect 12571 5612 12572 5676
rect 12636 5612 12637 5676
rect 12571 5611 12637 5612
rect 13494 4453 13554 8195
rect 13904 8192 14304 11250
rect 13904 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14304 8192
rect 13675 7852 13741 7853
rect 13675 7788 13676 7852
rect 13740 7788 13741 7852
rect 13675 7787 13741 7788
rect 13678 4997 13738 7787
rect 13904 7104 14304 8128
rect 13904 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14304 7104
rect 13904 6016 14304 7040
rect 13904 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14304 6016
rect 13675 4996 13741 4997
rect 13675 4932 13676 4996
rect 13740 4932 13741 4996
rect 13675 4931 13741 4932
rect 13904 4928 14304 5952
rect 13904 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14304 4928
rect 13491 4452 13557 4453
rect 13491 4388 13492 4452
rect 13556 4388 13557 4452
rect 13491 4387 13557 4388
rect 13904 3840 14304 4864
rect 13904 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14304 3840
rect 10915 2956 10981 2957
rect 10915 2954 10916 2956
rect 10734 2894 10916 2954
rect 10734 2549 10794 2894
rect 10915 2892 10916 2894
rect 10980 2892 10981 2956
rect 10915 2891 10981 2892
rect 13904 2752 14304 3776
rect 13904 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14304 2752
rect 10731 2548 10797 2549
rect 10731 2484 10732 2548
rect 10796 2484 10797 2548
rect 10731 2483 10797 2484
rect 10363 1324 10429 1325
rect 10363 1260 10364 1324
rect 10428 1260 10429 1324
rect 10363 1259 10429 1260
rect 13904 0 14304 2688
rect 14644 8736 15044 11250
rect 17355 9892 17421 9893
rect 17355 9828 17356 9892
rect 17420 9828 17421 9892
rect 17355 9827 17421 9828
rect 16987 9756 17053 9757
rect 16987 9692 16988 9756
rect 17052 9692 17053 9756
rect 16987 9691 17053 9692
rect 15147 9484 15213 9485
rect 15147 9420 15148 9484
rect 15212 9420 15213 9484
rect 15147 9419 15213 9420
rect 14644 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15044 8736
rect 14644 7648 15044 8672
rect 14644 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15044 7648
rect 14644 6560 15044 7584
rect 14644 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15044 6560
rect 14644 5472 15044 6496
rect 14644 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15044 5472
rect 14644 4384 15044 5408
rect 15150 4861 15210 9419
rect 15331 8668 15397 8669
rect 15331 8604 15332 8668
rect 15396 8604 15397 8668
rect 15331 8603 15397 8604
rect 15147 4860 15213 4861
rect 15147 4796 15148 4860
rect 15212 4796 15213 4860
rect 15147 4795 15213 4796
rect 14644 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15044 4384
rect 14644 3296 15044 4320
rect 15334 3773 15394 8603
rect 15515 8396 15581 8397
rect 15515 8332 15516 8396
rect 15580 8332 15581 8396
rect 15515 8331 15581 8332
rect 15518 3773 15578 8331
rect 15331 3772 15397 3773
rect 15331 3708 15332 3772
rect 15396 3708 15397 3772
rect 15331 3707 15397 3708
rect 15515 3772 15581 3773
rect 15515 3708 15516 3772
rect 15580 3708 15581 3772
rect 15515 3707 15581 3708
rect 14644 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15044 3296
rect 14644 2208 15044 3232
rect 16990 3229 17050 9691
rect 17358 3229 17418 9827
rect 17726 9150 17970 9210
rect 17726 9077 17786 9150
rect 17723 9076 17789 9077
rect 17723 9012 17724 9076
rect 17788 9012 17789 9076
rect 17723 9011 17789 9012
rect 17910 4317 17970 9150
rect 19563 8804 19629 8805
rect 19563 8740 19564 8804
rect 19628 8740 19629 8804
rect 19563 8739 19629 8740
rect 19195 7036 19261 7037
rect 19195 6972 19196 7036
rect 19260 6972 19261 7036
rect 19195 6971 19261 6972
rect 19011 6900 19077 6901
rect 19011 6836 19012 6900
rect 19076 6836 19077 6900
rect 19011 6835 19077 6836
rect 17907 4316 17973 4317
rect 17907 4252 17908 4316
rect 17972 4252 17973 4316
rect 17907 4251 17973 4252
rect 19014 3229 19074 6835
rect 16987 3228 17053 3229
rect 16987 3164 16988 3228
rect 17052 3164 17053 3228
rect 16987 3163 17053 3164
rect 17355 3228 17421 3229
rect 17355 3164 17356 3228
rect 17420 3164 17421 3228
rect 17355 3163 17421 3164
rect 19011 3228 19077 3229
rect 19011 3164 19012 3228
rect 19076 3164 19077 3228
rect 19011 3163 19077 3164
rect 14644 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15044 2208
rect 14644 0 15044 2144
rect 19198 1869 19258 6971
rect 19566 5677 19626 8739
rect 19904 8192 20304 11250
rect 19904 8128 19912 8192
rect 19976 8128 19992 8192
rect 20056 8128 20072 8192
rect 20136 8128 20152 8192
rect 20216 8128 20232 8192
rect 20296 8128 20304 8192
rect 19904 7104 20304 8128
rect 20644 8736 21044 11250
rect 21219 10300 21285 10301
rect 21219 10236 21220 10300
rect 21284 10236 21285 10300
rect 21219 10235 21285 10236
rect 21222 9485 21282 10235
rect 21219 9484 21285 9485
rect 21219 9420 21220 9484
rect 21284 9420 21285 9484
rect 21219 9419 21285 9420
rect 20644 8672 20652 8736
rect 20716 8672 20732 8736
rect 20796 8672 20812 8736
rect 20876 8672 20892 8736
rect 20956 8672 20972 8736
rect 21036 8672 21044 8736
rect 20483 8124 20549 8125
rect 20483 8060 20484 8124
rect 20548 8060 20549 8124
rect 20483 8059 20549 8060
rect 20486 7581 20546 8059
rect 20644 7648 21044 8672
rect 25904 8192 26304 11250
rect 25904 8128 25912 8192
rect 25976 8128 25992 8192
rect 26056 8128 26072 8192
rect 26136 8128 26152 8192
rect 26216 8128 26232 8192
rect 26296 8128 26304 8192
rect 21403 7716 21469 7717
rect 21403 7652 21404 7716
rect 21468 7652 21469 7716
rect 21403 7651 21469 7652
rect 20644 7584 20652 7648
rect 20716 7584 20732 7648
rect 20796 7584 20812 7648
rect 20876 7584 20892 7648
rect 20956 7584 20972 7648
rect 21036 7584 21044 7648
rect 20483 7580 20549 7581
rect 20483 7516 20484 7580
rect 20548 7516 20549 7580
rect 20483 7515 20549 7516
rect 19904 7040 19912 7104
rect 19976 7040 19992 7104
rect 20056 7040 20072 7104
rect 20136 7040 20152 7104
rect 20216 7040 20232 7104
rect 20296 7040 20304 7104
rect 19904 6016 20304 7040
rect 20483 6628 20549 6629
rect 20483 6564 20484 6628
rect 20548 6564 20549 6628
rect 20483 6563 20549 6564
rect 20486 6085 20546 6563
rect 20644 6560 21044 7584
rect 21219 7036 21285 7037
rect 21219 6972 21220 7036
rect 21284 6972 21285 7036
rect 21219 6971 21285 6972
rect 20644 6496 20652 6560
rect 20716 6496 20732 6560
rect 20796 6496 20812 6560
rect 20876 6496 20892 6560
rect 20956 6496 20972 6560
rect 21036 6496 21044 6560
rect 20483 6084 20549 6085
rect 20483 6020 20484 6084
rect 20548 6020 20549 6084
rect 20483 6019 20549 6020
rect 19904 5952 19912 6016
rect 19976 5952 19992 6016
rect 20056 5952 20072 6016
rect 20136 5952 20152 6016
rect 20216 5952 20232 6016
rect 20296 5952 20304 6016
rect 19563 5676 19629 5677
rect 19563 5612 19564 5676
rect 19628 5612 19629 5676
rect 19563 5611 19629 5612
rect 19904 4928 20304 5952
rect 20483 5948 20549 5949
rect 20483 5884 20484 5948
rect 20548 5884 20549 5948
rect 20483 5883 20549 5884
rect 20486 5405 20546 5883
rect 20644 5472 21044 6496
rect 20644 5408 20652 5472
rect 20716 5408 20732 5472
rect 20796 5408 20812 5472
rect 20876 5408 20892 5472
rect 20956 5408 20972 5472
rect 21036 5408 21044 5472
rect 20483 5404 20549 5405
rect 20483 5340 20484 5404
rect 20548 5340 20549 5404
rect 20483 5339 20549 5340
rect 19904 4864 19912 4928
rect 19976 4864 19992 4928
rect 20056 4864 20072 4928
rect 20136 4864 20152 4928
rect 20216 4864 20232 4928
rect 20296 4864 20304 4928
rect 19904 3840 20304 4864
rect 19904 3776 19912 3840
rect 19976 3776 19992 3840
rect 20056 3776 20072 3840
rect 20136 3776 20152 3840
rect 20216 3776 20232 3840
rect 20296 3776 20304 3840
rect 19904 2752 20304 3776
rect 19904 2688 19912 2752
rect 19976 2688 19992 2752
rect 20056 2688 20072 2752
rect 20136 2688 20152 2752
rect 20216 2688 20232 2752
rect 20296 2688 20304 2752
rect 19195 1868 19261 1869
rect 19195 1804 19196 1868
rect 19260 1804 19261 1868
rect 19195 1803 19261 1804
rect 19904 0 20304 2688
rect 20644 4384 21044 5408
rect 20644 4320 20652 4384
rect 20716 4320 20732 4384
rect 20796 4320 20812 4384
rect 20876 4320 20892 4384
rect 20956 4320 20972 4384
rect 21036 4320 21044 4384
rect 20644 3296 21044 4320
rect 21222 4317 21282 6971
rect 21406 5677 21466 7651
rect 21587 7172 21653 7173
rect 21587 7108 21588 7172
rect 21652 7108 21653 7172
rect 21587 7107 21653 7108
rect 21771 7172 21837 7173
rect 21771 7108 21772 7172
rect 21836 7108 21837 7172
rect 21771 7107 21837 7108
rect 21403 5676 21469 5677
rect 21403 5612 21404 5676
rect 21468 5612 21469 5676
rect 21403 5611 21469 5612
rect 21219 4316 21285 4317
rect 21219 4252 21220 4316
rect 21284 4252 21285 4316
rect 21219 4251 21285 4252
rect 21590 3501 21650 7107
rect 21774 4181 21834 7107
rect 25904 7104 26304 8128
rect 26644 8736 27044 11250
rect 27659 8940 27725 8941
rect 27659 8876 27660 8940
rect 27724 8876 27725 8940
rect 27659 8875 27725 8876
rect 26644 8672 26652 8736
rect 26716 8672 26732 8736
rect 26796 8672 26812 8736
rect 26876 8672 26892 8736
rect 26956 8672 26972 8736
rect 27036 8672 27044 8736
rect 26371 8124 26437 8125
rect 26371 8060 26372 8124
rect 26436 8060 26437 8124
rect 26371 8059 26437 8060
rect 26374 7853 26434 8059
rect 26371 7852 26437 7853
rect 26371 7788 26372 7852
rect 26436 7788 26437 7852
rect 26371 7787 26437 7788
rect 26644 7648 27044 8672
rect 26644 7584 26652 7648
rect 26716 7584 26732 7648
rect 26796 7584 26812 7648
rect 26876 7584 26892 7648
rect 26956 7584 26972 7648
rect 27036 7584 27044 7648
rect 26371 7580 26437 7581
rect 26371 7516 26372 7580
rect 26436 7516 26437 7580
rect 26371 7515 26437 7516
rect 26374 7173 26434 7515
rect 26371 7172 26437 7173
rect 26371 7108 26372 7172
rect 26436 7108 26437 7172
rect 26371 7107 26437 7108
rect 25904 7040 25912 7104
rect 25976 7040 25992 7104
rect 26056 7040 26072 7104
rect 26136 7040 26152 7104
rect 26216 7040 26232 7104
rect 26296 7040 26304 7104
rect 25904 6016 26304 7040
rect 26371 7036 26437 7037
rect 26371 6972 26372 7036
rect 26436 6972 26437 7036
rect 26371 6971 26437 6972
rect 26374 6493 26434 6971
rect 26644 6560 27044 7584
rect 26644 6496 26652 6560
rect 26716 6496 26732 6560
rect 26796 6496 26812 6560
rect 26876 6496 26892 6560
rect 26956 6496 26972 6560
rect 27036 6496 27044 6560
rect 26371 6492 26437 6493
rect 26371 6428 26372 6492
rect 26436 6428 26437 6492
rect 26371 6427 26437 6428
rect 25904 5952 25912 6016
rect 25976 5952 25992 6016
rect 26056 5952 26072 6016
rect 26136 5952 26152 6016
rect 26216 5952 26232 6016
rect 26296 5952 26304 6016
rect 25904 4928 26304 5952
rect 26644 5472 27044 6496
rect 27107 6492 27173 6493
rect 27107 6428 27108 6492
rect 27172 6428 27173 6492
rect 27107 6427 27173 6428
rect 27110 6085 27170 6427
rect 27107 6084 27173 6085
rect 27107 6020 27108 6084
rect 27172 6020 27173 6084
rect 27107 6019 27173 6020
rect 27662 5541 27722 8875
rect 31904 8192 32304 11250
rect 32644 8736 33044 11250
rect 35019 9076 35085 9077
rect 35019 9012 35020 9076
rect 35084 9012 35085 9076
rect 35019 9011 35085 9012
rect 32644 8672 32652 8736
rect 32716 8672 32732 8736
rect 32796 8672 32812 8736
rect 32876 8672 32892 8736
rect 32956 8672 32972 8736
rect 33036 8672 33044 8736
rect 32443 8668 32509 8669
rect 32443 8604 32444 8668
rect 32508 8604 32509 8668
rect 32443 8603 32509 8604
rect 31904 8128 31912 8192
rect 31976 8128 31992 8192
rect 32056 8128 32072 8192
rect 32136 8128 32152 8192
rect 32216 8128 32232 8192
rect 32296 8128 32304 8192
rect 31904 7104 32304 8128
rect 32446 7173 32506 8603
rect 32644 7648 33044 8672
rect 33915 8260 33981 8261
rect 33915 8196 33916 8260
rect 33980 8196 33981 8260
rect 33915 8195 33981 8196
rect 32644 7584 32652 7648
rect 32716 7584 32732 7648
rect 32796 7584 32812 7648
rect 32876 7584 32892 7648
rect 32956 7584 32972 7648
rect 33036 7584 33044 7648
rect 32443 7172 32509 7173
rect 32443 7108 32444 7172
rect 32508 7108 32509 7172
rect 32443 7107 32509 7108
rect 31904 7040 31912 7104
rect 31976 7040 31992 7104
rect 32056 7040 32072 7104
rect 32136 7040 32152 7104
rect 32216 7040 32232 7104
rect 32296 7040 32304 7104
rect 31904 6016 32304 7040
rect 32644 6560 33044 7584
rect 32644 6496 32652 6560
rect 32716 6496 32732 6560
rect 32796 6496 32812 6560
rect 32876 6496 32892 6560
rect 32956 6496 32972 6560
rect 33036 6496 33044 6560
rect 32443 6356 32509 6357
rect 32443 6292 32444 6356
rect 32508 6292 32509 6356
rect 32443 6291 32509 6292
rect 31904 5952 31912 6016
rect 31976 5952 31992 6016
rect 32056 5952 32072 6016
rect 32136 5952 32152 6016
rect 32216 5952 32232 6016
rect 32296 5952 32304 6016
rect 28027 5948 28093 5949
rect 28027 5884 28028 5948
rect 28092 5884 28093 5948
rect 28027 5883 28093 5884
rect 27659 5540 27725 5541
rect 27659 5476 27660 5540
rect 27724 5476 27725 5540
rect 27659 5475 27725 5476
rect 26644 5408 26652 5472
rect 26716 5408 26732 5472
rect 26796 5408 26812 5472
rect 26876 5408 26892 5472
rect 26956 5408 26972 5472
rect 27036 5408 27044 5472
rect 26371 4996 26437 4997
rect 26371 4932 26372 4996
rect 26436 4932 26437 4996
rect 26371 4931 26437 4932
rect 25904 4864 25912 4928
rect 25976 4864 25992 4928
rect 26056 4864 26072 4928
rect 26136 4864 26152 4928
rect 26216 4864 26232 4928
rect 26296 4864 26304 4928
rect 21771 4180 21837 4181
rect 21771 4116 21772 4180
rect 21836 4116 21837 4180
rect 21771 4115 21837 4116
rect 25904 3840 26304 4864
rect 26374 4453 26434 4931
rect 26371 4452 26437 4453
rect 26371 4388 26372 4452
rect 26436 4388 26437 4452
rect 26371 4387 26437 4388
rect 25904 3776 25912 3840
rect 25976 3776 25992 3840
rect 26056 3776 26072 3840
rect 26136 3776 26152 3840
rect 26216 3776 26232 3840
rect 26296 3776 26304 3840
rect 21587 3500 21653 3501
rect 21587 3436 21588 3500
rect 21652 3436 21653 3500
rect 21587 3435 21653 3436
rect 20644 3232 20652 3296
rect 20716 3232 20732 3296
rect 20796 3232 20812 3296
rect 20876 3232 20892 3296
rect 20956 3232 20972 3296
rect 21036 3232 21044 3296
rect 20644 2208 21044 3232
rect 20644 2144 20652 2208
rect 20716 2144 20732 2208
rect 20796 2144 20812 2208
rect 20876 2144 20892 2208
rect 20956 2144 20972 2208
rect 21036 2144 21044 2208
rect 20644 0 21044 2144
rect 25904 2752 26304 3776
rect 25904 2688 25912 2752
rect 25976 2688 25992 2752
rect 26056 2688 26072 2752
rect 26136 2688 26152 2752
rect 26216 2688 26232 2752
rect 26296 2688 26304 2752
rect 25904 0 26304 2688
rect 26644 4384 27044 5408
rect 27843 5268 27909 5269
rect 27843 5204 27844 5268
rect 27908 5204 27909 5268
rect 27843 5203 27909 5204
rect 26644 4320 26652 4384
rect 26716 4320 26732 4384
rect 26796 4320 26812 4384
rect 26876 4320 26892 4384
rect 26956 4320 26972 4384
rect 27036 4320 27044 4384
rect 26644 3296 27044 4320
rect 26644 3232 26652 3296
rect 26716 3232 26732 3296
rect 26796 3232 26812 3296
rect 26876 3232 26892 3296
rect 26956 3232 26972 3296
rect 27036 3232 27044 3296
rect 26644 2208 27044 3232
rect 26644 2144 26652 2208
rect 26716 2144 26732 2208
rect 26796 2144 26812 2208
rect 26876 2144 26892 2208
rect 26956 2144 26972 2208
rect 27036 2144 27044 2208
rect 26644 0 27044 2144
rect 27846 1869 27906 5203
rect 28030 4725 28090 5883
rect 31904 4928 32304 5952
rect 31904 4864 31912 4928
rect 31976 4864 31992 4928
rect 32056 4864 32072 4928
rect 32136 4864 32152 4928
rect 32216 4864 32232 4928
rect 32296 4864 32304 4928
rect 28027 4724 28093 4725
rect 28027 4660 28028 4724
rect 28092 4660 28093 4724
rect 28027 4659 28093 4660
rect 31904 3840 32304 4864
rect 31904 3776 31912 3840
rect 31976 3776 31992 3840
rect 32056 3776 32072 3840
rect 32136 3776 32152 3840
rect 32216 3776 32232 3840
rect 32296 3776 32304 3840
rect 31904 2752 32304 3776
rect 32446 3229 32506 6291
rect 32644 5472 33044 6496
rect 32644 5408 32652 5472
rect 32716 5408 32732 5472
rect 32796 5408 32812 5472
rect 32876 5408 32892 5472
rect 32956 5408 32972 5472
rect 33036 5408 33044 5472
rect 32644 4384 33044 5408
rect 32644 4320 32652 4384
rect 32716 4320 32732 4384
rect 32796 4320 32812 4384
rect 32876 4320 32892 4384
rect 32956 4320 32972 4384
rect 33036 4320 33044 4384
rect 32644 3296 33044 4320
rect 33918 3909 33978 8195
rect 35022 4861 35082 9011
rect 37904 8192 38304 11250
rect 37904 8128 37912 8192
rect 37976 8128 37992 8192
rect 38056 8128 38072 8192
rect 38136 8128 38152 8192
rect 38216 8128 38232 8192
rect 38296 8128 38304 8192
rect 37904 7104 38304 8128
rect 37904 7040 37912 7104
rect 37976 7040 37992 7104
rect 38056 7040 38072 7104
rect 38136 7040 38152 7104
rect 38216 7040 38232 7104
rect 38296 7040 38304 7104
rect 37904 6016 38304 7040
rect 37904 5952 37912 6016
rect 37976 5952 37992 6016
rect 38056 5952 38072 6016
rect 38136 5952 38152 6016
rect 38216 5952 38232 6016
rect 38296 5952 38304 6016
rect 37904 4928 38304 5952
rect 37904 4864 37912 4928
rect 37976 4864 37992 4928
rect 38056 4864 38072 4928
rect 38136 4864 38152 4928
rect 38216 4864 38232 4928
rect 38296 4864 38304 4928
rect 35019 4860 35085 4861
rect 35019 4796 35020 4860
rect 35084 4796 35085 4860
rect 35019 4795 35085 4796
rect 33915 3908 33981 3909
rect 33915 3844 33916 3908
rect 33980 3844 33981 3908
rect 33915 3843 33981 3844
rect 32644 3232 32652 3296
rect 32716 3232 32732 3296
rect 32796 3232 32812 3296
rect 32876 3232 32892 3296
rect 32956 3232 32972 3296
rect 33036 3232 33044 3296
rect 32443 3228 32509 3229
rect 32443 3164 32444 3228
rect 32508 3164 32509 3228
rect 32443 3163 32509 3164
rect 31904 2688 31912 2752
rect 31976 2688 31992 2752
rect 32056 2688 32072 2752
rect 32136 2688 32152 2752
rect 32216 2688 32232 2752
rect 32296 2688 32304 2752
rect 27843 1868 27909 1869
rect 27843 1804 27844 1868
rect 27908 1804 27909 1868
rect 27843 1803 27909 1804
rect 31904 0 32304 2688
rect 32644 2208 33044 3232
rect 32644 2144 32652 2208
rect 32716 2144 32732 2208
rect 32796 2144 32812 2208
rect 32876 2144 32892 2208
rect 32956 2144 32972 2208
rect 33036 2144 33044 2208
rect 32644 0 33044 2144
rect 37904 3840 38304 4864
rect 37904 3776 37912 3840
rect 37976 3776 37992 3840
rect 38056 3776 38072 3840
rect 38136 3776 38152 3840
rect 38216 3776 38232 3840
rect 38296 3776 38304 3840
rect 37904 2752 38304 3776
rect 37904 2688 37912 2752
rect 37976 2688 37992 2752
rect 38056 2688 38072 2752
rect 38136 2688 38152 2752
rect 38216 2688 38232 2752
rect 38296 2688 38304 2752
rect 37904 0 38304 2688
rect 38644 8736 39044 11250
rect 38644 8672 38652 8736
rect 38716 8672 38732 8736
rect 38796 8672 38812 8736
rect 38876 8672 38892 8736
rect 38956 8672 38972 8736
rect 39036 8672 39044 8736
rect 38644 7648 39044 8672
rect 38644 7584 38652 7648
rect 38716 7584 38732 7648
rect 38796 7584 38812 7648
rect 38876 7584 38892 7648
rect 38956 7584 38972 7648
rect 39036 7584 39044 7648
rect 38644 6560 39044 7584
rect 38644 6496 38652 6560
rect 38716 6496 38732 6560
rect 38796 6496 38812 6560
rect 38876 6496 38892 6560
rect 38956 6496 38972 6560
rect 39036 6496 39044 6560
rect 38644 5472 39044 6496
rect 38644 5408 38652 5472
rect 38716 5408 38732 5472
rect 38796 5408 38812 5472
rect 38876 5408 38892 5472
rect 38956 5408 38972 5472
rect 39036 5408 39044 5472
rect 38644 4384 39044 5408
rect 38644 4320 38652 4384
rect 38716 4320 38732 4384
rect 38796 4320 38812 4384
rect 38876 4320 38892 4384
rect 38956 4320 38972 4384
rect 39036 4320 39044 4384
rect 38644 3296 39044 4320
rect 38644 3232 38652 3296
rect 38716 3232 38732 3296
rect 38796 3232 38812 3296
rect 38876 3232 38892 3296
rect 38956 3232 38972 3296
rect 39036 3232 39044 3296
rect 38644 2208 39044 3232
rect 38644 2144 38652 2208
rect 38716 2144 38732 2208
rect 38796 2144 38812 2208
rect 38876 2144 38892 2208
rect 38956 2144 38972 2208
rect 39036 2144 39044 2208
rect 38644 0 39044 2144
use sky130_fd_sc_hd__mux4_1  _032_
timestamp -3599
transform 1 0 31464 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _033_
timestamp -3599
transform 1 0 12696 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _034_
timestamp -3599
transform 1 0 35512 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _035_
timestamp -3599
transform -1 0 12788 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _036_
timestamp -3599
transform 1 0 27508 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _037_
timestamp -3599
transform 1 0 14536 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _038_
timestamp -3599
transform -1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _039_
timestamp -3599
transform -1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _040_
timestamp -3599
transform -1 0 11316 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _041_
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _042_
timestamp -3599
transform -1 0 26404 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _043_
timestamp -3599
transform -1 0 25760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _044_
timestamp -3599
transform 1 0 24656 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _045_
timestamp -3599
transform -1 0 26772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _046_
timestamp -3599
transform -1 0 25484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _047_
timestamp -3599
transform 1 0 25576 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _048_
timestamp -3599
transform 1 0 18216 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _049_
timestamp -3599
transform 1 0 18492 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _050_
timestamp -3599
transform 1 0 18492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _051_
timestamp -3599
transform -1 0 19872 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _052_
timestamp -3599
transform -1 0 19412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _053_
timestamp -3599
transform -1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _054_
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp -3599
transform 1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp -3599
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _057_
timestamp -3599
transform -1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp -3599
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _059_
timestamp -3599
transform -1 0 26772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _060_
timestamp -3599
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _061_
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _062_
timestamp -3599
transform -1 0 24840 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _063_
timestamp -3599
transform 1 0 19780 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _064_
timestamp -3599
transform -1 0 24012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _065_
timestamp -3599
transform 1 0 19780 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _066_
timestamp -3599
transform 1 0 22908 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _068_
timestamp -3599
transform -1 0 24380 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _069_
timestamp -3599
transform 1 0 19780 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _070_
timestamp -3599
transform 1 0 21804 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _071_
timestamp -3599
transform 1 0 19780 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _072_
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _073_
timestamp -3599
transform -1 0 24288 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _074_
timestamp -3599
transform 1 0 19872 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _075_
timestamp -3599
transform -1 0 22632 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _076_
timestamp -3599
transform -1 0 22448 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _077_
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _078_
timestamp -3599
transform -1 0 17020 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _079_
timestamp -3599
transform 1 0 25668 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _080_
timestamp -3599
transform 1 0 38548 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _081_
timestamp -3599
transform 1 0 2760 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _082_
timestamp -3599
transform 1 0 32844 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _083_
timestamp -3599
transform 1 0 28152 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _084_
timestamp -3599
transform 1 0 4416 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _085_
timestamp -3599
transform 1 0 28796 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _086_
timestamp -3599
transform 1 0 14628 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _087_
timestamp -3599
transform -1 0 21620 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _088_
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _089_
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _090_
timestamp -3599
transform 1 0 38364 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _091_
timestamp -3599
transform 1 0 2576 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _092_
timestamp -3599
transform 1 0 32384 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _093_
timestamp -3599
transform 1 0 34316 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _094_
timestamp -3599
transform 1 0 25024 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _095_
timestamp -3599
transform 1 0 7912 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _096_
timestamp -3599
transform 1 0 35880 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _097_
timestamp -3599
transform 1 0 5244 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _098_
timestamp -3599
transform 1 0 29992 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _099_
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _100_
timestamp -3599
transform -1 0 18584 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _101_
timestamp -3599
transform 1 0 7912 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _102_
timestamp -3599
transform 1 0 30728 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _103_
timestamp -3599
transform -1 0 10948 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _104_
timestamp -3599
transform -1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _105_
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _106_
timestamp -3599
transform 1 0 33672 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _107_
timestamp -3599
transform -1 0 8924 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _108_
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _109_
timestamp -3599
transform 1 0 34316 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _110_
timestamp -3599
transform 1 0 25484 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _111_
timestamp -3599
transform 1 0 8648 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _112_
timestamp -3599
transform 1 0 36156 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _113_
timestamp -3599
transform -1 0 7820 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _114_
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _115_
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _116_
timestamp -3599
transform -1 0 21160 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _117_
timestamp -3599
transform 1 0 32384 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _118_
timestamp -3599
transform 1 0 28336 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _119_
timestamp -3599
transform -1 0 10856 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  _120_
timestamp -3599
transform -1 0 33764 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _121_
timestamp -3599
transform -1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _122_
timestamp -3599
transform 1 0 3128 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _123_
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _124_
timestamp -3599
transform -1 0 39560 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _125_
timestamp -3599
transform 1 0 38456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _126_
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _127_
timestamp -3599
transform 1 0 11592 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _128_
timestamp -3599
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _129_
timestamp -3599
transform -1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _130_
timestamp -3599
transform -1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _131_
timestamp -3599
transform 1 0 13432 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _132_
timestamp -3599
transform -1 0 29256 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _133_
timestamp -3599
transform 1 0 27048 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _134_
timestamp -3599
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _135_
timestamp -3599
transform 1 0 10304 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _136_
timestamp -3599
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _137_
timestamp -3599
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _138_
timestamp -3599
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _139_
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _140_
timestamp -3599
transform 1 0 30360 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _141_
timestamp -3599
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _142_
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _143_
timestamp -3599
transform 1 0 6716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _144_
timestamp -3599
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _145_
timestamp -3599
transform 1 0 27876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _146_
timestamp -3599
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _147_
timestamp -3599
transform 1 0 31556 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _148_
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _149_
timestamp -3599
transform 1 0 17756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _150_
timestamp -3599
transform 1 0 10488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _151_
timestamp -3599
transform 1 0 10396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _152_
timestamp -3599
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _153_
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _154_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _155_
timestamp -3599
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _156_
timestamp -3599
transform 1 0 36064 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _157_
timestamp -3599
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _158_
timestamp -3599
transform -1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _159_
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _160_
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _161_
timestamp -3599
transform 1 0 25208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _162_
timestamp -3599
transform -1 0 36340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _163_
timestamp -3599
transform 1 0 37260 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _164_
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _165_
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _166_
timestamp -3599
transform 1 0 6440 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _167_
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _168_
timestamp -3599
transform -1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _169_
timestamp -3599
transform -1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _170_
timestamp -3599
transform 1 0 4600 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _171_
timestamp -3599
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _172_
timestamp -3599
transform 1 0 17480 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _173_
timestamp -3599
transform 1 0 17572 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _174_
timestamp -3599
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _175_
timestamp -3599
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _176_
timestamp -3599
transform 1 0 30084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _177_
timestamp -3599
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _178_
timestamp -3599
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _179_
timestamp -3599
transform -1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _180_
timestamp -3599
transform 1 0 15548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _181_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _182_
timestamp -3599
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _183_
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _184_
timestamp -3599
transform -1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _185_
timestamp -3599
transform 1 0 29716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _186_
timestamp -3599
transform 1 0 4784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _187_
timestamp -3599
transform 1 0 4784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _188_
timestamp -3599
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _189_
timestamp -3599
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _190_
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _191_
timestamp -3599
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _192_
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _193_
timestamp -3599
transform 1 0 24104 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _194_
timestamp -3599
transform -1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _195_
timestamp -3599
transform -1 0 36892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _196_
timestamp -3599
transform 1 0 32660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _197_
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _198_
timestamp -3599
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _199_
timestamp -3599
transform 1 0 1472 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _200_
timestamp -3599
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _201_
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _202_
timestamp -3599
transform -1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _203_
timestamp -3599
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _204_
timestamp -3599
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _205_
timestamp -3599
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _206_
timestamp -3599
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _207_
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _208_
timestamp -3599
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _209_
timestamp -3599
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _210_
timestamp -3599
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _211_
timestamp -3599
transform 1 0 28244 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _212_
timestamp -3599
transform 1 0 4140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _213_
timestamp -3599
transform 1 0 4232 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _214_
timestamp -3599
transform 1 0 22632 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _215_
timestamp -3599
transform 1 0 27508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _216_
timestamp -3599
transform 1 0 32568 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _217_
timestamp -3599
transform 1 0 32660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _218_
timestamp -3599
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _219_
timestamp -3599
transform -1 0 2760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _220_
timestamp -3599
transform 1 0 38180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _221_
timestamp -3599
transform 1 0 37444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _222_
timestamp -3599
transform 1 0 24932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _223_
timestamp -3599
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _224_
timestamp -3599
transform -1 0 16836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _225_
timestamp -3599
transform -1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _226_
timestamp -3599
transform 1 0 28244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _227_
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _228_
timestamp -3599
transform -1 0 23276 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _229_
timestamp -3599
transform 1 0 19596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _230_
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _231_
timestamp -3599
transform 1 0 16468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _232_
timestamp -3599
transform -1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _233_
timestamp -3599
transform -1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _234_
timestamp -3599
transform -1 0 26404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _235_
timestamp -3599
transform -1 0 23276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _236_
timestamp -3599
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _237_
timestamp -3599
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _238_
timestamp -3599
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _239_
timestamp -3599
transform 1 0 14628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _240_
timestamp -3599
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _241_
timestamp -3599
transform 1 0 17572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _242_
timestamp -3599
transform 1 0 11960 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _243_
timestamp -3599
transform -1 0 11408 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _245_
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _246_
timestamp -3599
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _247_
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _248_
timestamp -3599
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _249_
timestamp -3599
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _250_
timestamp -3599
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _251_
timestamp -3599
transform 1 0 35144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _252_
timestamp -3599
transform 1 0 33764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _253_
timestamp -3599
transform 1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _254_
timestamp -3599
transform 1 0 3128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp -3599
transform -1 0 39560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp -3599
transform -1 0 38180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _257_
timestamp -3599
transform 1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _258_
timestamp -3599
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _259_
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _260_
timestamp -3599
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _261_
timestamp -3599
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _262_
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _263_
timestamp -3599
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _264_
timestamp -3599
transform 1 0 30084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _265_
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _266_
timestamp -3599
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _267_
timestamp -3599
transform -1 0 39744 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp -3599
transform -1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _269_
timestamp -3599
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _270_
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _271_
timestamp -3599
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _272_
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _273_
timestamp -3599
transform 1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _274_
timestamp -3599
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _275_
timestamp -3599
transform 1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _276_
timestamp -3599
transform 1 0 31464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp -3599
transform 1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp -3599
transform 1 0 38916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp -3599
transform 1 0 36708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _280_
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _281_
timestamp -3599
transform -1 0 42320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _282_
timestamp -3599
transform -1 0 42596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _283_
timestamp -3599
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp -3599
transform 1 0 41768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp -3599
transform -1 0 38640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp -3599
transform 1 0 42044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp -3599
transform 1 0 42596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp -3599
transform -1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp -3599
transform 1 0 40388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp -3599
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp -3599
transform 1 0 41492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp -3599
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp -3599
transform 1 0 42596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp -3599
transform -1 0 41676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp -3599
transform 1 0 42320 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp -3599
transform 1 0 42044 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp -3599
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _298_
timestamp -3599
transform -1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp -3599
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _300_
timestamp -3599
transform -1 0 13800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _301_
timestamp -3599
transform -1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp -3599
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _303_
timestamp -3599
transform -1 0 38548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp -3599
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _305_
timestamp -3599
transform -1 0 33488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _307_
timestamp -3599
transform -1 0 30636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _308_
timestamp -3599
transform -1 0 34408 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _309_
timestamp -3599
transform -1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp -3599
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp -3599
transform -1 0 37168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp -3599
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _313_
timestamp -3599
transform -1 0 38456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp -3599
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp -3599
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _316_
timestamp -3599
transform -1 0 35328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _317_
timestamp -3599
transform -1 0 21620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _319_
timestamp -3599
transform -1 0 35880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp -3599
transform -1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp -3599
transform -1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp -3599
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp -3599
transform -1 0 32016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp -3599
transform 1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp -3599
transform 1 0 17204 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _327_
timestamp -3599
transform -1 0 32292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp -3599
transform -1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _329_
timestamp -3599
transform -1 0 37628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp -3599
transform -1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _331_
timestamp -3599
transform -1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _332_
timestamp -3599
transform -1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp -3599
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _334_
timestamp -3599
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _335_
timestamp -3599
transform -1 0 40940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _336_
timestamp -3599
transform -1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _337_
timestamp -3599
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _338_
timestamp -3599
transform 1 0 19596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp -3599
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _340_
timestamp -3599
transform -1 0 31004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _341_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _342_
timestamp -3599
transform -1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _343_
timestamp -3599
transform -1 0 34592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _344_
timestamp -3599
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp -3599
transform 1 0 40480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _346_
timestamp -3599
transform -1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp -3599
transform -1 0 14352 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _348_
timestamp -3599
transform -1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _349_
timestamp -3599
transform -1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 43240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform 1 0 42688 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 38272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 17112 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp -3599
transform 1 0 12144 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK
timestamp -3599
transform -1 0 13340 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp -3599
transform -1 0 11960 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp -3599
transform -1 0 13340 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp -3599
transform 1 0 14260 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp -3599
transform -1 0 8648 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp -3599
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp -3599
transform -1 0 38916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp -3599
transform 1 0 38456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout51
timestamp -3599
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp -3599
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout54
timestamp -3599
transform -1 0 19136 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp -3599
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp -3599
transform -1 0 36892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp -3599
transform -1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp -3599
transform -1 0 13892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp -3599
transform -1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp -3599
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp -3599
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp -3599
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42
timestamp -3599
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp -3599
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp -3599
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp -3599
transform 1 0 14812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp -3599
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp -3599
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp -3599
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp -3599
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp -3599
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_243
timestamp -3599
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp -3599
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_253
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp -3599
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp -3599
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp -3599
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_317
timestamp -3599
transform 1 0 30268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp -3599
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp -3599
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636964856
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636964856
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp -3599
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636964856
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_433
timestamp -3599
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_441
timestamp -3599
transform 1 0 41676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_449
timestamp -3599
transform 1 0 42412 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_21
timestamp 1636964856
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1636964856
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_45
timestamp -3599
transform 1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp -3599
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp -3599
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_95
timestamp -3599
transform 1 0 9844 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp -3599
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp -3599
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp -3599
transform 1 0 23644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp -3599
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_286
timestamp -3599
transform 1 0 27416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp -3599
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_318
timestamp -3599
transform 1 0 30360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp -3599
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp -3599
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp -3599
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636964856
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_408
timestamp -3599
transform 1 0 38640 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_412
timestamp 1636964856
transform 1 0 39008 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_424
timestamp -3599
transform 1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_430
timestamp -3599
transform 1 0 40664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_434
timestamp -3599
transform 1 0 41032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_441
timestamp -3599
transform 1 0 41676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_449
timestamp -3599
transform 1 0 42412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_19
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp -3599
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp -3599
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_76
timestamp -3599
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_101
timestamp -3599
transform 1 0 10396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_130
timestamp -3599
transform 1 0 13064 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp -3599
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_150
timestamp -3599
transform 1 0 14904 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_168
timestamp -3599
transform 1 0 16560 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp -3599
transform 1 0 17296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp -3599
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_213
timestamp 1636964856
transform 1 0 20700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_228
timestamp -3599
transform 1 0 22080 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp -3599
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_262
timestamp -3599
transform 1 0 25208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_266
timestamp -3599
transform 1 0 25576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_288
timestamp -3599
transform 1 0 27600 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_294
timestamp -3599
transform 1 0 28152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp -3599
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp -3599
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_329
timestamp -3599
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp -3599
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp -3599
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_368
timestamp -3599
transform 1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_383
timestamp -3599
transform 1 0 36340 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_391
timestamp -3599
transform 1 0 37076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_414
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636964856
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636964856
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_37
timestamp -3599
transform 1 0 4508 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp -3599
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp -3599
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp -3599
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp -3599
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp -3599
transform 1 0 12328 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_147
timestamp 1636964856
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp -3599
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_193
timestamp -3599
transform 1 0 18860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp -3599
transform 1 0 19596 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_234
timestamp -3599
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp -3599
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_265
timestamp -3599
transform 1 0 25484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_274
timestamp -3599
transform 1 0 26312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_290
timestamp -3599
transform 1 0 27784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_294
timestamp -3599
transform 1 0 28152 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_307
timestamp 1636964856
transform 1 0 29348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_322
timestamp 1636964856
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp -3599
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_337
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_382
timestamp -3599
transform 1 0 36248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_386
timestamp -3599
transform 1 0 36616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp -3599
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp -3599
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_401
timestamp -3599
transform 1 0 37996 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_413
timestamp 1636964856
transform 1 0 39100 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_425
timestamp 1636964856
transform 1 0 40204 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_437
timestamp -3599
transform 1 0 41308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_452
timestamp -3599
transform 1 0 42688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp -3599
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp -3599
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp -3599
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_113
timestamp -3599
transform 1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_159
timestamp -3599
transform 1 0 15732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_164
timestamp -3599
transform 1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_179
timestamp -3599
transform 1 0 17572 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp -3599
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_230
timestamp -3599
transform 1 0 22264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_291
timestamp -3599
transform 1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_351
timestamp -3599
transform 1 0 33396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_357
timestamp -3599
transform 1 0 33948 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp -3599
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_372
timestamp -3599
transform 1 0 35328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_380
timestamp -3599
transform 1 0 36064 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp -3599
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636964856
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636964856
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_445
timestamp -3599
transform 1 0 42044 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_453
timestamp -3599
transform 1 0 42780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_39
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp -3599
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp -3599
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp -3599
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_134
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp -3599
transform 1 0 14444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp -3599
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_235
timestamp -3599
transform 1 0 22724 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp -3599
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_296
timestamp -3599
transform 1 0 28336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_300
timestamp -3599
transform 1 0 28704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_325
timestamp -3599
transform 1 0 31004 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_352
timestamp -3599
transform 1 0 33488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_378
timestamp -3599
transform 1 0 35880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_418
timestamp 1636964856
transform 1 0 39560 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_430
timestamp 1636964856
transform 1 0 40664 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_442
timestamp -3599
transform 1 0 41768 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp -3599
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_453
timestamp -3599
transform 1 0 42780 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_7
timestamp -3599
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp -3599
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp -3599
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_150
timestamp -3599
transform 1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp -3599
transform 1 0 17020 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_230
timestamp 1636964856
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_242
timestamp -3599
transform 1 0 23368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp -3599
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_265
timestamp -3599
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp -3599
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_312
timestamp -3599
transform 1 0 29808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_320
timestamp -3599
transform 1 0 30544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_358
timestamp -3599
transform 1 0 34040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_389
timestamp -3599
transform 1 0 36892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_393
timestamp -3599
transform 1 0 37260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_397
timestamp -3599
transform 1 0 37628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp -3599
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636964856
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636964856
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_445
timestamp -3599
transform 1 0 42044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_453
timestamp -3599
transform 1 0 42780 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_40
timestamp -3599
transform 1 0 4784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp -3599
transform 1 0 14076 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp -3599
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_177
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp -3599
transform 1 0 19044 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_231
timestamp 1636964856
transform 1 0 22356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_258
timestamp -3599
transform 1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_344
timestamp -3599
transform 1 0 32752 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp -3599
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_431
timestamp 1636964856
transform 1 0 40756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_443
timestamp -3599
transform 1 0 41860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp -3599
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp -3599
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp -3599
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_33
timestamp -3599
transform 1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp -3599
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp -3599
transform 1 0 7544 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_119
timestamp -3599
transform 1 0 12052 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_171
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_230
timestamp -3599
transform 1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp -3599
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_286
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636964856
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636964856
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_445
timestamp -3599
transform 1 0 42044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_451
timestamp -3599
transform 1 0 42596 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_25
timestamp -3599
transform 1 0 3404 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp -3599
transform 1 0 4140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp -3599
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_92
timestamp -3599
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_149
timestamp -3599
transform 1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp -3599
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_274
timestamp -3599
transform 1 0 26312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_295
timestamp -3599
transform 1 0 28244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp -3599
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_433
timestamp 1636964856
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_449
timestamp -3599
transform 1 0 42412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_23
timestamp -3599
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_73
timestamp -3599
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_135
timestamp -3599
transform 1 0 13524 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_190
timestamp -3599
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp -3599
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp -3599
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_359
timestamp -3599
transform 1 0 34132 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_373
timestamp -3599
transform 1 0 35420 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp -3599
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_437
timestamp -3599
transform 1 0 41308 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_13
timestamp -3599
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_125
timestamp -3599
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp -3599
transform 1 0 19688 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -3599
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_309
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_341
timestamp -3599
transform 1 0 32476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp -3599
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_419
timestamp -3599
transform 1 0 39652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_441
timestamp -3599
transform 1 0 41676 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_449
timestamp -3599
transform 1 0 42412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input1
timestamp -3599
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp -3599
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp -3599
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp -3599
transform 1 0 3128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp -3599
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input17
timestamp -3599
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp -3599
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -3599
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp -3599
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp -3599
transform 1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp -3599
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp -3599
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp -3599
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp -3599
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp -3599
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp -3599
transform -1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp -3599
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp -3599
transform 1 0 19872 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -3599
transform -1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp -3599
transform -1 0 19136 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp -3599
transform -1 0 22448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input41
timestamp -3599
transform 1 0 23552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp -3599
transform 1 0 23368 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp -3599
transform 1 0 25484 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input45
timestamp -3599
transform 1 0 24748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input47
timestamp -3599
transform -1 0 24104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp -3599
transform 1 0 20976 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input49
timestamp -3599
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp -3599
transform -1 0 21712 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input51
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp -3599
transform -1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp -3599
transform 1 0 22356 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp -3599
transform 1 0 23276 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp -3599
transform 1 0 22448 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input56
timestamp -3599
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp -3599
transform -1 0 29348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input58
timestamp -3599
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp -3599
transform -1 0 29808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp -3599
transform -1 0 30084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp -3599
transform -1 0 32016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp -3599
transform -1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp -3599
transform 1 0 26956 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp -3599
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp -3599
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp -3599
transform 1 0 30820 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp -3599
transform -1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp -3599
transform 1 0 27968 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp -3599
transform -1 0 29348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input71
timestamp -3599
transform 1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp -3599
transform 1 0 31556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp -3599
transform 1 0 33672 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input74
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp -3599
transform 1 0 33764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp -3599
transform -1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input79
timestamp -3599
transform -1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp -3599
transform 1 0 30360 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input81
timestamp -3599
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input83
timestamp -3599
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp -3599
transform 1 0 35604 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input85
timestamp -3599
transform -1 0 32568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp -3599
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input87
timestamp -3599
transform -1 0 32752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 42504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 43240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 42872 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 43240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 42872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 43240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 42872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 43240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 42872 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 43240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform 1 0 42688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform 1 0 43240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform 1 0 43240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform 1 0 42872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform 1 0 43240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform 1 0 42504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform 1 0 43240 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform 1 0 41952 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 42504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform 1 0 42872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform 1 0 42504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform 1 0 42136 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform 1 0 41768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform 1 0 43240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform 1 0 43240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 43240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform 1 0 42872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform -1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform -1 0 39652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform 1 0 38916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 39652 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 40572 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform -1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform -1 0 41308 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform -1 0 41676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform -1 0 40664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform -1 0 41308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform -1 0 35420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform -1 0 36892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 34592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform -1 0 38548 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform -1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 38916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform 1 0 38916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform -1 0 38916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform -1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform -1 0 2944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform -1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform -1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform -1 0 6992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform -1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp -3599
transform -1 0 5520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp -3599
transform -1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp -3599
transform -1 0 7728 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp -3599
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp -3599
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp -3599
transform -1 0 6992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp -3599
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp -3599
transform -1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp -3599
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp -3599
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp -3599
transform -1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp -3599
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp -3599
transform -1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp -3599
transform -1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp -3599
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp -3599
transform -1 0 8832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp -3599
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp -3599
transform -1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp -3599
transform -1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp -3599
transform -1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp -3599
transform -1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp -3599
transform -1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp -3599
transform -1 0 13708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp -3599
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp -3599
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp -3599
transform -1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp -3599
transform -1 0 19136 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp -3599
transform -1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp -3599
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp -3599
transform -1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp -3599
transform -1 0 16560 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp -3599
transform -1 0 13984 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp -3599
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output204
timestamp -3599
transform -1 0 35880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 43884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 43884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 43884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 43884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 43884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 43884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 43884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 43884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 43884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_IO_205
timestamp -3599
transform 1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp -3599
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp -3599
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_45
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp -3599
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_54
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_55
timestamp -3599
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_59
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp -3599
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_70
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp -3599
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_73
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_86
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -3599
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_91
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_92
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_93
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_94
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_95
timestamp -3599
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_96
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_97
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_98
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp -3599
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_106
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_110
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp -3599
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_118
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_119
timestamp -3599
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_122
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_123
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_124
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_125
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_126
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_127
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_128
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_129
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_130
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_131
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp -3599
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp -3599
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 B_I_top
port 7 nsew signal output
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 B_O_top
port 8 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 B_T_top
port 9 nsew signal output
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal2 s 19522 10450 19578 11250 0 FreeSans 224 90 0 0 Co
port 14 nsew signal output
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 15 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 16 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 17 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 18 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 19 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 20 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 21 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 22 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 23 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 24 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 25 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 26 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 27 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 28 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 29 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 30 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 31 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 32 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 33 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 34 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 35 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 36 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 37 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 38 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 39 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 40 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 41 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 42 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 43 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 44 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 45 nsew signal input
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 46 nsew signal input
flabel metal3 s 44200 1368 45000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 47 nsew signal output
flabel metal3 s 44200 4088 45000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 48 nsew signal output
flabel metal3 s 44200 4360 45000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 49 nsew signal output
flabel metal3 s 44200 4632 45000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 50 nsew signal output
flabel metal3 s 44200 4904 45000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 51 nsew signal output
flabel metal3 s 44200 5176 45000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 52 nsew signal output
flabel metal3 s 44200 5448 45000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 53 nsew signal output
flabel metal3 s 44200 5720 45000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 54 nsew signal output
flabel metal3 s 44200 5992 45000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 55 nsew signal output
flabel metal3 s 44200 6264 45000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 56 nsew signal output
flabel metal3 s 44200 6536 45000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 57 nsew signal output
flabel metal3 s 44200 1640 45000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 58 nsew signal output
flabel metal3 s 44200 6808 45000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 59 nsew signal output
flabel metal3 s 44200 7080 45000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 60 nsew signal output
flabel metal3 s 44200 7352 45000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 61 nsew signal output
flabel metal3 s 44200 7624 45000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 62 nsew signal output
flabel metal3 s 44200 7896 45000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 63 nsew signal output
flabel metal3 s 44200 8168 45000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 64 nsew signal output
flabel metal3 s 44200 8440 45000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 65 nsew signal output
flabel metal3 s 44200 8712 45000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 66 nsew signal output
flabel metal3 s 44200 8984 45000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 67 nsew signal output
flabel metal3 s 44200 9256 45000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 68 nsew signal output
flabel metal3 s 44200 1912 45000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 69 nsew signal output
flabel metal3 s 44200 9528 45000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 70 nsew signal output
flabel metal3 s 44200 9800 45000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 71 nsew signal output
flabel metal3 s 44200 2184 45000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 72 nsew signal output
flabel metal3 s 44200 2456 45000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 73 nsew signal output
flabel metal3 s 44200 2728 45000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 74 nsew signal output
flabel metal3 s 44200 3000 45000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 75 nsew signal output
flabel metal3 s 44200 3272 45000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 76 nsew signal output
flabel metal3 s 44200 3544 45000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 77 nsew signal output
flabel metal3 s 44200 3816 45000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 78 nsew signal output
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 79 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 80 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 81 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 82 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 83 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 84 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 85 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 86 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 87 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 88 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 89 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 90 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 91 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 92 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 93 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 94 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 95 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 96 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 97 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 98 nsew signal input
flabel metal2 s 34426 10450 34482 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 99 nsew signal output
flabel metal2 s 37186 10450 37242 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 100 nsew signal output
flabel metal2 s 37462 10450 37518 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 101 nsew signal output
flabel metal2 s 37738 10450 37794 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 102 nsew signal output
flabel metal2 s 38014 10450 38070 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 103 nsew signal output
flabel metal2 s 38290 10450 38346 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 104 nsew signal output
flabel metal2 s 38566 10450 38622 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 105 nsew signal output
flabel metal2 s 38842 10450 38898 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 106 nsew signal output
flabel metal2 s 39118 10450 39174 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 107 nsew signal output
flabel metal2 s 39394 10450 39450 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 108 nsew signal output
flabel metal2 s 39670 10450 39726 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 109 nsew signal output
flabel metal2 s 34702 10450 34758 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 110 nsew signal output
flabel metal2 s 34978 10450 35034 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 111 nsew signal output
flabel metal2 s 35254 10450 35310 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 112 nsew signal output
flabel metal2 s 35530 10450 35586 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 113 nsew signal output
flabel metal2 s 35806 10450 35862 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 114 nsew signal output
flabel metal2 s 36082 10450 36138 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 115 nsew signal output
flabel metal2 s 36358 10450 36414 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 116 nsew signal output
flabel metal2 s 36634 10450 36690 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 117 nsew signal output
flabel metal2 s 36910 10450 36966 11250 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 118 nsew signal output
flabel metal2 s 5170 10450 5226 11250 0 FreeSans 224 90 0 0 N1BEG[0]
port 119 nsew signal output
flabel metal2 s 5446 10450 5502 11250 0 FreeSans 224 90 0 0 N1BEG[1]
port 120 nsew signal output
flabel metal2 s 5722 10450 5778 11250 0 FreeSans 224 90 0 0 N1BEG[2]
port 121 nsew signal output
flabel metal2 s 5998 10450 6054 11250 0 FreeSans 224 90 0 0 N1BEG[3]
port 122 nsew signal output
flabel metal2 s 6274 10450 6330 11250 0 FreeSans 224 90 0 0 N2BEG[0]
port 123 nsew signal output
flabel metal2 s 6550 10450 6606 11250 0 FreeSans 224 90 0 0 N2BEG[1]
port 124 nsew signal output
flabel metal2 s 6826 10450 6882 11250 0 FreeSans 224 90 0 0 N2BEG[2]
port 125 nsew signal output
flabel metal2 s 7102 10450 7158 11250 0 FreeSans 224 90 0 0 N2BEG[3]
port 126 nsew signal output
flabel metal2 s 7378 10450 7434 11250 0 FreeSans 224 90 0 0 N2BEG[4]
port 127 nsew signal output
flabel metal2 s 7654 10450 7710 11250 0 FreeSans 224 90 0 0 N2BEG[5]
port 128 nsew signal output
flabel metal2 s 7930 10450 7986 11250 0 FreeSans 224 90 0 0 N2BEG[6]
port 129 nsew signal output
flabel metal2 s 8206 10450 8262 11250 0 FreeSans 224 90 0 0 N2BEG[7]
port 130 nsew signal output
flabel metal2 s 8482 10450 8538 11250 0 FreeSans 224 90 0 0 N2BEGb[0]
port 131 nsew signal output
flabel metal2 s 8758 10450 8814 11250 0 FreeSans 224 90 0 0 N2BEGb[1]
port 132 nsew signal output
flabel metal2 s 9034 10450 9090 11250 0 FreeSans 224 90 0 0 N2BEGb[2]
port 133 nsew signal output
flabel metal2 s 9310 10450 9366 11250 0 FreeSans 224 90 0 0 N2BEGb[3]
port 134 nsew signal output
flabel metal2 s 9586 10450 9642 11250 0 FreeSans 224 90 0 0 N2BEGb[4]
port 135 nsew signal output
flabel metal2 s 9862 10450 9918 11250 0 FreeSans 224 90 0 0 N2BEGb[5]
port 136 nsew signal output
flabel metal2 s 10138 10450 10194 11250 0 FreeSans 224 90 0 0 N2BEGb[6]
port 137 nsew signal output
flabel metal2 s 10414 10450 10470 11250 0 FreeSans 224 90 0 0 N2BEGb[7]
port 138 nsew signal output
flabel metal2 s 10690 10450 10746 11250 0 FreeSans 224 90 0 0 N4BEG[0]
port 139 nsew signal output
flabel metal2 s 13450 10450 13506 11250 0 FreeSans 224 90 0 0 N4BEG[10]
port 140 nsew signal output
flabel metal2 s 13726 10450 13782 11250 0 FreeSans 224 90 0 0 N4BEG[11]
port 141 nsew signal output
flabel metal2 s 14002 10450 14058 11250 0 FreeSans 224 90 0 0 N4BEG[12]
port 142 nsew signal output
flabel metal2 s 14278 10450 14334 11250 0 FreeSans 224 90 0 0 N4BEG[13]
port 143 nsew signal output
flabel metal2 s 14554 10450 14610 11250 0 FreeSans 224 90 0 0 N4BEG[14]
port 144 nsew signal output
flabel metal2 s 14830 10450 14886 11250 0 FreeSans 224 90 0 0 N4BEG[15]
port 145 nsew signal output
flabel metal2 s 10966 10450 11022 11250 0 FreeSans 224 90 0 0 N4BEG[1]
port 146 nsew signal output
flabel metal2 s 11242 10450 11298 11250 0 FreeSans 224 90 0 0 N4BEG[2]
port 147 nsew signal output
flabel metal2 s 11518 10450 11574 11250 0 FreeSans 224 90 0 0 N4BEG[3]
port 148 nsew signal output
flabel metal2 s 11794 10450 11850 11250 0 FreeSans 224 90 0 0 N4BEG[4]
port 149 nsew signal output
flabel metal2 s 12070 10450 12126 11250 0 FreeSans 224 90 0 0 N4BEG[5]
port 150 nsew signal output
flabel metal2 s 12346 10450 12402 11250 0 FreeSans 224 90 0 0 N4BEG[6]
port 151 nsew signal output
flabel metal2 s 12622 10450 12678 11250 0 FreeSans 224 90 0 0 N4BEG[7]
port 152 nsew signal output
flabel metal2 s 12898 10450 12954 11250 0 FreeSans 224 90 0 0 N4BEG[8]
port 153 nsew signal output
flabel metal2 s 13174 10450 13230 11250 0 FreeSans 224 90 0 0 N4BEG[9]
port 154 nsew signal output
flabel metal2 s 15106 10450 15162 11250 0 FreeSans 224 90 0 0 NN4BEG[0]
port 155 nsew signal output
flabel metal2 s 17866 10450 17922 11250 0 FreeSans 224 90 0 0 NN4BEG[10]
port 156 nsew signal output
flabel metal2 s 18142 10450 18198 11250 0 FreeSans 224 90 0 0 NN4BEG[11]
port 157 nsew signal output
flabel metal2 s 18418 10450 18474 11250 0 FreeSans 224 90 0 0 NN4BEG[12]
port 158 nsew signal output
flabel metal2 s 18694 10450 18750 11250 0 FreeSans 224 90 0 0 NN4BEG[13]
port 159 nsew signal output
flabel metal2 s 18970 10450 19026 11250 0 FreeSans 224 90 0 0 NN4BEG[14]
port 160 nsew signal output
flabel metal2 s 19246 10450 19302 11250 0 FreeSans 224 90 0 0 NN4BEG[15]
port 161 nsew signal output
flabel metal2 s 15382 10450 15438 11250 0 FreeSans 224 90 0 0 NN4BEG[1]
port 162 nsew signal output
flabel metal2 s 15658 10450 15714 11250 0 FreeSans 224 90 0 0 NN4BEG[2]
port 163 nsew signal output
flabel metal2 s 15934 10450 15990 11250 0 FreeSans 224 90 0 0 NN4BEG[3]
port 164 nsew signal output
flabel metal2 s 16210 10450 16266 11250 0 FreeSans 224 90 0 0 NN4BEG[4]
port 165 nsew signal output
flabel metal2 s 16486 10450 16542 11250 0 FreeSans 224 90 0 0 NN4BEG[5]
port 166 nsew signal output
flabel metal2 s 16762 10450 16818 11250 0 FreeSans 224 90 0 0 NN4BEG[6]
port 167 nsew signal output
flabel metal2 s 17038 10450 17094 11250 0 FreeSans 224 90 0 0 NN4BEG[7]
port 168 nsew signal output
flabel metal2 s 17314 10450 17370 11250 0 FreeSans 224 90 0 0 NN4BEG[8]
port 169 nsew signal output
flabel metal2 s 17590 10450 17646 11250 0 FreeSans 224 90 0 0 NN4BEG[9]
port 170 nsew signal output
flabel metal2 s 19798 10450 19854 11250 0 FreeSans 224 90 0 0 S1END[0]
port 171 nsew signal input
flabel metal2 s 20074 10450 20130 11250 0 FreeSans 224 90 0 0 S1END[1]
port 172 nsew signal input
flabel metal2 s 20350 10450 20406 11250 0 FreeSans 224 90 0 0 S1END[2]
port 173 nsew signal input
flabel metal2 s 20626 10450 20682 11250 0 FreeSans 224 90 0 0 S1END[3]
port 174 nsew signal input
flabel metal2 s 23110 10450 23166 11250 0 FreeSans 224 90 0 0 S2END[0]
port 175 nsew signal input
flabel metal2 s 23386 10450 23442 11250 0 FreeSans 224 90 0 0 S2END[1]
port 176 nsew signal input
flabel metal2 s 23662 10450 23718 11250 0 FreeSans 224 90 0 0 S2END[2]
port 177 nsew signal input
flabel metal2 s 23938 10450 23994 11250 0 FreeSans 224 90 0 0 S2END[3]
port 178 nsew signal input
flabel metal2 s 24214 10450 24270 11250 0 FreeSans 224 90 0 0 S2END[4]
port 179 nsew signal input
flabel metal2 s 24490 10450 24546 11250 0 FreeSans 224 90 0 0 S2END[5]
port 180 nsew signal input
flabel metal2 s 24766 10450 24822 11250 0 FreeSans 224 90 0 0 S2END[6]
port 181 nsew signal input
flabel metal2 s 25042 10450 25098 11250 0 FreeSans 224 90 0 0 S2END[7]
port 182 nsew signal input
flabel metal2 s 20902 10450 20958 11250 0 FreeSans 224 90 0 0 S2MID[0]
port 183 nsew signal input
flabel metal2 s 21178 10450 21234 11250 0 FreeSans 224 90 0 0 S2MID[1]
port 184 nsew signal input
flabel metal2 s 21454 10450 21510 11250 0 FreeSans 224 90 0 0 S2MID[2]
port 185 nsew signal input
flabel metal2 s 21730 10450 21786 11250 0 FreeSans 224 90 0 0 S2MID[3]
port 186 nsew signal input
flabel metal2 s 22006 10450 22062 11250 0 FreeSans 224 90 0 0 S2MID[4]
port 187 nsew signal input
flabel metal2 s 22282 10450 22338 11250 0 FreeSans 224 90 0 0 S2MID[5]
port 188 nsew signal input
flabel metal2 s 22558 10450 22614 11250 0 FreeSans 224 90 0 0 S2MID[6]
port 189 nsew signal input
flabel metal2 s 22834 10450 22890 11250 0 FreeSans 224 90 0 0 S2MID[7]
port 190 nsew signal input
flabel metal2 s 25318 10450 25374 11250 0 FreeSans 224 90 0 0 S4END[0]
port 191 nsew signal input
flabel metal2 s 28078 10450 28134 11250 0 FreeSans 224 90 0 0 S4END[10]
port 192 nsew signal input
flabel metal2 s 28354 10450 28410 11250 0 FreeSans 224 90 0 0 S4END[11]
port 193 nsew signal input
flabel metal2 s 28630 10450 28686 11250 0 FreeSans 224 90 0 0 S4END[12]
port 194 nsew signal input
flabel metal2 s 28906 10450 28962 11250 0 FreeSans 224 90 0 0 S4END[13]
port 195 nsew signal input
flabel metal2 s 29182 10450 29238 11250 0 FreeSans 224 90 0 0 S4END[14]
port 196 nsew signal input
flabel metal2 s 29458 10450 29514 11250 0 FreeSans 224 90 0 0 S4END[15]
port 197 nsew signal input
flabel metal2 s 25594 10450 25650 11250 0 FreeSans 224 90 0 0 S4END[1]
port 198 nsew signal input
flabel metal2 s 25870 10450 25926 11250 0 FreeSans 224 90 0 0 S4END[2]
port 199 nsew signal input
flabel metal2 s 26146 10450 26202 11250 0 FreeSans 224 90 0 0 S4END[3]
port 200 nsew signal input
flabel metal2 s 26422 10450 26478 11250 0 FreeSans 224 90 0 0 S4END[4]
port 201 nsew signal input
flabel metal2 s 26698 10450 26754 11250 0 FreeSans 224 90 0 0 S4END[5]
port 202 nsew signal input
flabel metal2 s 26974 10450 27030 11250 0 FreeSans 224 90 0 0 S4END[6]
port 203 nsew signal input
flabel metal2 s 27250 10450 27306 11250 0 FreeSans 224 90 0 0 S4END[7]
port 204 nsew signal input
flabel metal2 s 27526 10450 27582 11250 0 FreeSans 224 90 0 0 S4END[8]
port 205 nsew signal input
flabel metal2 s 27802 10450 27858 11250 0 FreeSans 224 90 0 0 S4END[9]
port 206 nsew signal input
flabel metal2 s 29734 10450 29790 11250 0 FreeSans 224 90 0 0 SS4END[0]
port 207 nsew signal input
flabel metal2 s 32494 10450 32550 11250 0 FreeSans 224 90 0 0 SS4END[10]
port 208 nsew signal input
flabel metal2 s 32770 10450 32826 11250 0 FreeSans 224 90 0 0 SS4END[11]
port 209 nsew signal input
flabel metal2 s 33046 10450 33102 11250 0 FreeSans 224 90 0 0 SS4END[12]
port 210 nsew signal input
flabel metal2 s 33322 10450 33378 11250 0 FreeSans 224 90 0 0 SS4END[13]
port 211 nsew signal input
flabel metal2 s 33598 10450 33654 11250 0 FreeSans 224 90 0 0 SS4END[14]
port 212 nsew signal input
flabel metal2 s 33874 10450 33930 11250 0 FreeSans 224 90 0 0 SS4END[15]
port 213 nsew signal input
flabel metal2 s 30010 10450 30066 11250 0 FreeSans 224 90 0 0 SS4END[1]
port 214 nsew signal input
flabel metal2 s 30286 10450 30342 11250 0 FreeSans 224 90 0 0 SS4END[2]
port 215 nsew signal input
flabel metal2 s 30562 10450 30618 11250 0 FreeSans 224 90 0 0 SS4END[3]
port 216 nsew signal input
flabel metal2 s 30838 10450 30894 11250 0 FreeSans 224 90 0 0 SS4END[4]
port 217 nsew signal input
flabel metal2 s 31114 10450 31170 11250 0 FreeSans 224 90 0 0 SS4END[5]
port 218 nsew signal input
flabel metal2 s 31390 10450 31446 11250 0 FreeSans 224 90 0 0 SS4END[6]
port 219 nsew signal input
flabel metal2 s 31666 10450 31722 11250 0 FreeSans 224 90 0 0 SS4END[7]
port 220 nsew signal input
flabel metal2 s 31942 10450 31998 11250 0 FreeSans 224 90 0 0 SS4END[8]
port 221 nsew signal input
flabel metal2 s 32218 10450 32274 11250 0 FreeSans 224 90 0 0 SS4END[9]
port 222 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 UserCLK
port 223 nsew signal input
flabel metal2 s 34150 10450 34206 11250 0 FreeSans 224 90 0 0 UserCLKo
port 224 nsew signal output
flabel metal4 s 2644 0 3044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 2644 0 3044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 2644 11190 3044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 8644 0 9044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 8644 0 9044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 8644 11190 9044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 14644 0 15044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 14644 0 15044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 14644 11190 15044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 20644 0 21044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 20644 0 21044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 20644 11190 21044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 26644 0 27044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 26644 0 27044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 26644 11190 27044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 32644 0 33044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 32644 0 33044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 32644 11190 33044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 38644 0 39044 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 38644 0 39044 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 38644 11190 39044 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 1904 0 2304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 1904 0 2304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 1904 11190 2304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 7904 0 8304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 7904 0 8304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 7904 11190 8304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 13904 0 14304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 13904 0 14304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 13904 11190 14304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 19904 0 20304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 19904 0 20304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 19904 11190 20304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 25904 0 26304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 25904 0 26304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 25904 11190 26304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 31904 0 32304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 31904 0 32304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 31904 11190 32304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 37904 0 38304 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 37904 0 38304 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 37904 11190 38304 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
rlabel metal1 22494 8704 22494 8704 0 VGND
rlabel metal1 22494 8160 22494 8160 0 VPWR
rlabel metal2 3358 959 3358 959 0 A_I_top
rlabel metal2 2162 1163 2162 1163 0 A_O_top
rlabel metal2 4554 1520 4554 1520 0 A_T_top
rlabel metal2 9338 823 9338 823 0 A_config_C_bit0
rlabel metal2 10534 823 10534 823 0 A_config_C_bit1
rlabel metal2 12834 1734 12834 1734 0 A_config_C_bit2
rlabel metal2 12926 1520 12926 1520 0 A_config_C_bit3
rlabel metal2 6946 1520 6946 1520 0 B_I_top
rlabel metal2 5750 1554 5750 1554 0 B_O_top
rlabel metal2 8142 823 8142 823 0 B_T_top
rlabel metal2 14122 1656 14122 1656 0 B_config_C_bit0
rlabel metal2 15318 1520 15318 1520 0 B_config_C_bit1
rlabel metal2 16606 1717 16606 1717 0 B_config_C_bit2
rlabel metal2 17710 1520 17710 1520 0 B_config_C_bit3
rlabel metal3 1556 1428 1556 1428 0 FrameData[0]
rlabel metal3 1464 4148 1464 4148 0 FrameData[10]
rlabel metal3 1050 4420 1050 4420 0 FrameData[11]
rlabel metal3 1280 4692 1280 4692 0 FrameData[12]
rlabel metal3 1096 4964 1096 4964 0 FrameData[13]
rlabel metal3 2062 5236 2062 5236 0 FrameData[14]
rlabel metal3 1602 5508 1602 5508 0 FrameData[15]
rlabel metal3 1188 5780 1188 5780 0 FrameData[16]
rlabel metal3 1050 6052 1050 6052 0 FrameData[17]
rlabel metal3 1510 6324 1510 6324 0 FrameData[18]
rlabel metal3 1096 6596 1096 6596 0 FrameData[19]
rlabel metal2 3358 2023 3358 2023 0 FrameData[1]
rlabel metal3 1050 6868 1050 6868 0 FrameData[20]
rlabel metal3 1050 7140 1050 7140 0 FrameData[21]
rlabel metal3 1510 7412 1510 7412 0 FrameData[22]
rlabel metal3 1579 7684 1579 7684 0 FrameData[23]
rlabel metal3 1096 7956 1096 7956 0 FrameData[24]
rlabel metal3 1211 8228 1211 8228 0 FrameData[25]
rlabel metal3 1188 8500 1188 8500 0 FrameData[26]
rlabel metal3 1510 8772 1510 8772 0 FrameData[27]
rlabel metal2 3174 8245 3174 8245 0 FrameData[28]
rlabel metal3 1050 9316 1050 9316 0 FrameData[29]
rlabel metal3 1234 1972 1234 1972 0 FrameData[2]
rlabel metal2 3082 9044 3082 9044 0 FrameData[30]
rlabel metal2 3450 8823 3450 8823 0 FrameData[31]
rlabel metal3 1050 2244 1050 2244 0 FrameData[3]
rlabel metal3 1050 2516 1050 2516 0 FrameData[4]
rlabel metal3 1050 2788 1050 2788 0 FrameData[5]
rlabel metal3 935 3060 935 3060 0 FrameData[6]
rlabel metal3 1280 3332 1280 3332 0 FrameData[7]
rlabel metal3 1142 3604 1142 3604 0 FrameData[8]
rlabel metal3 1096 3876 1096 3876 0 FrameData[9]
rlabel metal1 42826 2278 42826 2278 0 FrameData_O[0]
rlabel metal2 43470 4063 43470 4063 0 FrameData_O[10]
rlabel via2 43102 4437 43102 4437 0 FrameData_O[11]
rlabel via2 43470 4709 43470 4709 0 FrameData_O[12]
rlabel via2 43102 4981 43102 4981 0 FrameData_O[13]
rlabel metal2 43470 5287 43470 5287 0 FrameData_O[14]
rlabel via2 43102 5525 43102 5525 0 FrameData_O[15]
rlabel via2 43470 5797 43470 5797 0 FrameData_O[16]
rlabel via2 43102 6069 43102 6069 0 FrameData_O[17]
rlabel metal2 43470 6375 43470 6375 0 FrameData_O[18]
rlabel via2 42918 6613 42918 6613 0 FrameData_O[19]
rlabel metal1 42504 2550 42504 2550 0 FrameData_O[1]
rlabel metal2 43470 6749 43470 6749 0 FrameData_O[20]
rlabel via2 43470 7157 43470 7157 0 FrameData_O[21]
rlabel metal2 43102 7565 43102 7565 0 FrameData_O[22]
rlabel via2 43470 7701 43470 7701 0 FrameData_O[23]
rlabel metal1 42826 7514 42826 7514 0 FrameData_O[24]
rlabel metal2 43102 8279 43102 8279 0 FrameData_O[25]
rlabel metal2 43470 8551 43470 8551 0 FrameData_O[26]
rlabel metal1 42504 8602 42504 8602 0 FrameData_O[27]
rlabel metal1 42964 8058 42964 8058 0 FrameData_O[28]
rlabel metal1 43194 7514 43194 7514 0 FrameData_O[29]
rlabel metal1 42826 2890 42826 2890 0 FrameData_O[2]
rlabel metal1 42872 7990 42872 7990 0 FrameData_O[30]
rlabel metal1 41998 7956 41998 7956 0 FrameData_O[31]
rlabel via2 43102 2261 43102 2261 0 FrameData_O[3]
rlabel via2 43470 2533 43470 2533 0 FrameData_O[4]
rlabel via2 43102 2805 43102 2805 0 FrameData_O[5]
rlabel metal2 43470 3111 43470 3111 0 FrameData_O[6]
rlabel via2 43102 3349 43102 3349 0 FrameData_O[7]
rlabel via2 43470 3621 43470 3621 0 FrameData_O[8]
rlabel via2 43102 3893 43102 3893 0 FrameData_O[9]
rlabel metal2 20102 1010 20102 1010 0 FrameStrobe[0]
rlabel metal2 42734 5474 42734 5474 0 FrameStrobe[10]
rlabel metal2 33258 823 33258 823 0 FrameStrobe[11]
rlabel metal2 34454 1044 34454 1044 0 FrameStrobe[12]
rlabel metal2 42642 2312 42642 2312 0 FrameStrobe[13]
rlabel metal1 42182 7752 42182 7752 0 FrameStrobe[14]
rlabel metal2 42182 2193 42182 2193 0 FrameStrobe[15]
rlabel metal2 43286 2312 43286 2312 0 FrameStrobe[16]
rlabel metal2 41446 2176 41446 2176 0 FrameStrobe[17]
rlabel metal2 41630 1911 41630 1911 0 FrameStrobe[18]
rlabel metal2 42826 1027 42826 1027 0 FrameStrobe[19]
rlabel metal2 21206 476 21206 476 0 FrameStrobe[1]
rlabel metal2 22494 1554 22494 1554 0 FrameStrobe[2]
rlabel metal1 32982 1972 32982 1972 0 FrameStrobe[3]
rlabel metal2 42274 2244 42274 2244 0 FrameStrobe[4]
rlabel metal2 42550 1802 42550 1802 0 FrameStrobe[5]
rlabel metal2 41354 1598 41354 1598 0 FrameStrobe[6]
rlabel metal2 41998 2346 41998 2346 0 FrameStrobe[7]
rlabel metal2 38410 2040 38410 2040 0 FrameStrobe[8]
rlabel metal2 42090 2244 42090 2244 0 FrameStrobe[9]
rlabel metal1 34684 8058 34684 8058 0 FrameStrobe_O[0]
rlabel metal1 39376 8330 39376 8330 0 FrameStrobe_O[10]
rlabel metal1 39330 7990 39330 7990 0 FrameStrobe_O[11]
rlabel metal1 39606 8058 39606 8058 0 FrameStrobe_O[12]
rlabel metal2 39974 9112 39974 9112 0 FrameStrobe_O[13]
rlabel metal1 40204 8262 40204 8262 0 FrameStrobe_O[14]
rlabel metal2 40710 9112 40710 9112 0 FrameStrobe_O[15]
rlabel metal2 41078 9146 41078 9146 0 FrameStrobe_O[16]
rlabel metal1 41584 8330 41584 8330 0 FrameStrobe_O[17]
rlabel metal1 40388 7514 40388 7514 0 FrameStrobe_O[18]
rlabel metal1 40618 8058 40618 8058 0 FrameStrobe_O[19]
rlabel metal1 34960 7990 34960 7990 0 FrameStrobe_O[1]
rlabel metal2 36662 9112 36662 9112 0 FrameStrobe_O[2]
rlabel metal2 34362 8942 34362 8942 0 FrameStrobe_O[3]
rlabel metal1 38272 8330 38272 8330 0 FrameStrobe_O[4]
rlabel metal2 37582 9010 37582 9010 0 FrameStrobe_O[5]
rlabel metal1 37904 8058 37904 8058 0 FrameStrobe_O[6]
rlabel metal2 38686 8432 38686 8432 0 FrameStrobe_O[7]
rlabel metal2 39146 8891 39146 8891 0 FrameStrobe_O[8]
rlabel metal1 38962 8058 38962 8058 0 FrameStrobe_O[9]
rlabel metal1 39100 6222 39100 6222 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal1 15134 3026 15134 3026 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal1 29670 4794 29670 4794 0 Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal1 29394 4250 29394 4250 0 Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 39238 6018 39238 6018 0 Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 39790 6154 39790 6154 0 Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal1 26174 2618 26174 2618 0 Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal1 26220 3162 26220 3162 0 Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 15778 6154 15778 6154 0 Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 16330 5848 16330 5848 0 Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal1 29762 3706 29762 3706 0 Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 30590 4250 30590 4250 0 Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal1 22264 2890 22264 2890 0 Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 21022 3842 21022 3842 0 Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 5658 7412 5658 7412 0 Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal1 21850 4590 21850 4590 0 Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel via2 17526 4811 17526 4811 0 Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 25898 4080 25898 4080 0 Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal1 27232 4794 27232 4794 0 Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal1 25714 4794 25714 4794 0 Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal1 23644 5066 23644 5066 0 Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal1 21114 5134 21114 5134 0 Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal1 25254 5644 25254 5644 0 Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 23506 6460 23506 6460 0 Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal1 18078 5236 18078 5236 0 Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 5106 7038 5106 7038 0 Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 18814 4590 18814 4590 0 Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 19090 4862 19090 4862 0 Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal1 23690 3400 23690 3400 0 Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 29394 6562 29394 6562 0 Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 33534 6426 33534 6426 0 Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal1 33902 5882 33902 5882 0 Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 3450 4930 3450 4930 0 Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal1 4186 5134 4186 5134 0 Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal1 8694 4794 8694 4794 0 Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal1 9062 4794 9062 4794 0 Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal1 37030 6426 37030 6426 0 Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal1 36708 5882 36708 5882 0 Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal1 7820 2618 7820 2618 0 Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal1 8556 2618 8556 2618 0 Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal1 25576 7990 25576 7990 0 Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal1 25714 7514 25714 7514 0 Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal1 34868 2890 34868 2890 0 Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal1 35742 2618 35742 2618 0 Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 33074 3162 33074 3162 0 Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal1 33350 2618 33350 2618 0 Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 17894 8228 17894 8228 0 Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 3082 6018 3082 6018 0 Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 3818 6375 3818 6375 0 Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal1 38962 6970 38962 6970 0 Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal1 39790 7310 39790 7310 0 Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal1 26542 5746 26542 5746 0 Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 27232 5678 27232 5678 0 Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 16514 3570 16514 3570 0 Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal1 17204 3706 17204 3706 0 Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal1 20930 7208 20930 7208 0 Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal1 19780 7310 19780 7310 0 Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal1 17526 7514 17526 7514 0 Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 15870 6188 15870 6188 0 Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal1 14214 4726 14214 4726 0 Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal1 11776 2890 11776 2890 0 Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal1 12650 2618 12650 2618 0 Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal1 31970 7956 31970 7956 0 Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal1 30728 7990 30728 7990 0 Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 6486 4828 6486 4828 0 Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal1 5612 4250 5612 4250 0 Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 33074 4522 33074 4522 0 Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal1 33120 3706 33120 3706 0 Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 36846 4862 36846 4862 0 Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 37398 4828 37398 4828 0 Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal1 9154 2618 9154 2618 0 Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal1 9936 3706 9936 3706 0 Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal1 25806 6834 25806 6834 0 Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 26680 6766 26680 6766 0 Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal1 35144 3706 35144 3706 0 Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal1 36938 3706 36938 3706 0 Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal1 20332 2618 20332 2618 0 Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal1 21022 2958 21022 2958 0 Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 20470 7004 20470 7004 0 Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 8234 6426 8234 6426 0 Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal1 7544 5338 7544 5338 0 Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 34914 5644 34914 5644 0 Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal1 34362 5100 34362 5100 0 Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 6900 5678 6900 5678 0 Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 6394 5950 6394 5950 0 Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 18170 3196 18170 3196 0 Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal1 18676 2618 18676 2618 0 Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 9706 6970 9706 6970 0 Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 10258 6732 10258 6732 0 Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 19918 6698 19918 6698 0 Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal1 31372 5814 31372 5814 0 Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal1 31740 5746 31740 5746 0 Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 11546 3808 11546 3808 0 Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal1 12098 4794 12098 4794 0 Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 33902 7514 33902 7514 0 Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 34454 7242 34454 7242 0 Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 7406 3366 7406 3366 0 Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal1 6210 3570 6210 3570 0 Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal1 10718 8364 10718 8364 0 Inst_S_IO_ConfigMem.Inst_frame3_bit14.Q
rlabel metal1 19090 7378 19090 7378 0 Inst_S_IO_ConfigMem.Inst_frame3_bit15.Q
rlabel metal1 14260 4794 14260 4794 0 Inst_S_IO_ConfigMem.Inst_frame3_bit16.Q
rlabel metal1 15134 2924 15134 2924 0 Inst_S_IO_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 28198 2754 28198 2754 0 Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q
rlabel metal1 28244 2550 28244 2550 0 Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 12098 6222 12098 6222 0 Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q
rlabel metal1 11454 5338 11454 5338 0 Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q
rlabel metal1 37858 7922 37858 7922 0 Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal1 36616 7514 36616 7514 0 Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 13386 4250 13386 4250 0 Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 13984 4046 13984 4046 0 Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal1 31556 2618 31556 2618 0 Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal1 32016 3162 32016 3162 0 Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 10166 6766 10166 6766 0 Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal1 8648 5746 8648 5746 0 Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 29026 7514 29026 7514 0 Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 29578 7854 29578 7854 0 Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 11362 7820 11362 7820 0 Inst_S_IO_switch_matrix.N1BEG0
rlabel metal2 19734 6732 19734 6732 0 Inst_S_IO_switch_matrix.N1BEG1
rlabel metal1 15364 4590 15364 4590 0 Inst_S_IO_switch_matrix.N1BEG2
rlabel metal1 14168 2414 14168 2414 0 Inst_S_IO_switch_matrix.N1BEG3
rlabel metal1 29532 3026 29532 3026 0 Inst_S_IO_switch_matrix.N2BEG0
rlabel metal1 12282 4148 12282 4148 0 Inst_S_IO_switch_matrix.N2BEG1
rlabel metal1 37904 7786 37904 7786 0 Inst_S_IO_switch_matrix.N2BEG2
rlabel metal1 15134 4114 15134 4114 0 Inst_S_IO_switch_matrix.N2BEG3
rlabel metal2 33350 4998 33350 4998 0 Inst_S_IO_switch_matrix.N2BEG4
rlabel metal1 8694 5678 8694 5678 0 Inst_S_IO_switch_matrix.N2BEG5
rlabel metal2 30590 6970 30590 6970 0 Inst_S_IO_switch_matrix.N2BEG6
rlabel metal2 34270 4386 34270 4386 0 Inst_S_IO_switch_matrix.N2BEG7
rlabel metal2 19366 6154 19366 6154 0 Inst_S_IO_switch_matrix.N2BEGb0
rlabel metal1 13708 3502 13708 3502 0 Inst_S_IO_switch_matrix.N2BEGb1
rlabel metal1 37122 7412 37122 7412 0 Inst_S_IO_switch_matrix.N2BEGb2
rlabel metal1 8050 3468 8050 3468 0 Inst_S_IO_switch_matrix.N2BEGb3
rlabel metal1 38180 4522 38180 4522 0 Inst_S_IO_switch_matrix.N2BEGb4
rlabel metal1 11086 4080 11086 4080 0 Inst_S_IO_switch_matrix.N2BEGb5
rlabel metal1 28842 6732 28842 6732 0 Inst_S_IO_switch_matrix.N2BEGb6
rlabel metal1 36156 4046 36156 4046 0 Inst_S_IO_switch_matrix.N2BEGb7
rlabel metal1 21436 3026 21436 3026 0 Inst_S_IO_switch_matrix.N4BEG0
rlabel metal1 8050 5678 8050 5678 0 Inst_S_IO_switch_matrix.N4BEG1
rlabel metal1 32292 6766 32292 6766 0 Inst_S_IO_switch_matrix.N4BEG10
rlabel metal2 7130 4998 7130 4998 0 Inst_S_IO_switch_matrix.N4BEG11
rlabel metal2 37582 6290 37582 6290 0 Inst_S_IO_switch_matrix.N4BEG12
rlabel via1 10074 2409 10074 2409 0 Inst_S_IO_switch_matrix.N4BEG13
rlabel metal1 29072 7854 29072 7854 0 Inst_S_IO_switch_matrix.N4BEG14
rlabel metal1 35558 3162 35558 3162 0 Inst_S_IO_switch_matrix.N4BEG15
rlabel metal1 35696 5202 35696 5202 0 Inst_S_IO_switch_matrix.N4BEG2
rlabel metal1 7636 5678 7636 5678 0 Inst_S_IO_switch_matrix.N4BEG3
rlabel metal1 18538 3162 18538 3162 0 Inst_S_IO_switch_matrix.N4BEG4
rlabel metal2 10258 5780 10258 5780 0 Inst_S_IO_switch_matrix.N4BEG5
rlabel metal2 31970 5372 31970 5372 0 Inst_S_IO_switch_matrix.N4BEG6
rlabel metal2 10810 4556 10810 4556 0 Inst_S_IO_switch_matrix.N4BEG7
rlabel metal2 17434 7242 17434 7242 0 Inst_S_IO_switch_matrix.N4BEG8
rlabel metal1 13846 3162 13846 3162 0 Inst_S_IO_switch_matrix.N4BEG9
rlabel metal1 34224 2822 34224 2822 0 Inst_S_IO_switch_matrix.NN4BEG0
rlabel metal1 4508 6290 4508 6290 0 Inst_S_IO_switch_matrix.NN4BEG1
rlabel metal2 34546 5882 34546 5882 0 Inst_S_IO_switch_matrix.NN4BEG10
rlabel metal1 4462 4114 4462 4114 0 Inst_S_IO_switch_matrix.NN4BEG11
rlabel metal1 40572 6290 40572 6290 0 Inst_S_IO_switch_matrix.NN4BEG12
rlabel metal2 27370 3196 27370 3196 0 Inst_S_IO_switch_matrix.NN4BEG13
rlabel metal1 14766 5882 14766 5882 0 Inst_S_IO_switch_matrix.NN4BEG14
rlabel metal2 30682 4284 30682 4284 0 Inst_S_IO_switch_matrix.NN4BEG15
rlabel metal1 40894 7412 40894 7412 0 Inst_S_IO_switch_matrix.NN4BEG2
rlabel metal2 28290 5372 28290 5372 0 Inst_S_IO_switch_matrix.NN4BEG3
rlabel metal1 18676 4114 18676 4114 0 Inst_S_IO_switch_matrix.NN4BEG4
rlabel metal2 19734 7684 19734 7684 0 Inst_S_IO_switch_matrix.NN4BEG5
rlabel metal1 16192 4590 16192 4590 0 Inst_S_IO_switch_matrix.NN4BEG6
rlabel metal1 30820 5202 30820 5202 0 Inst_S_IO_switch_matrix.NN4BEG7
rlabel metal2 6394 6460 6394 6460 0 Inst_S_IO_switch_matrix.NN4BEG8
rlabel metal2 29762 5882 29762 5882 0 Inst_S_IO_switch_matrix.NN4BEG9
rlabel metal2 5198 9122 5198 9122 0 N1BEG[0]
rlabel metal1 4692 8058 4692 8058 0 N1BEG[1]
rlabel metal2 3542 8704 3542 8704 0 N1BEG[2]
rlabel metal1 3082 8568 3082 8568 0 N1BEG[3]
rlabel metal1 4876 8602 4876 8602 0 N2BEG[0]
rlabel metal1 6716 6426 6716 6426 0 N2BEG[1]
rlabel metal2 6118 8160 6118 8160 0 N2BEG[2]
rlabel metal2 4186 9010 4186 9010 0 N2BEG[3]
rlabel metal2 6762 8602 6762 8602 0 N2BEG[4]
rlabel metal1 4554 8364 4554 8364 0 N2BEG[5]
rlabel metal1 7498 7514 7498 7514 0 N2BEG[6]
rlabel metal2 4922 8568 4922 8568 0 N2BEG[7]
rlabel metal2 5290 8908 5290 8908 0 N2BEGb[0]
rlabel metal2 6486 8976 6486 8976 0 N2BEGb[1]
rlabel metal1 5750 8262 5750 8262 0 N2BEGb[2]
rlabel metal1 7406 7242 7406 7242 0 N2BEGb[3]
rlabel metal1 9292 6426 9292 6426 0 N2BEGb[4]
rlabel metal1 6532 8330 6532 8330 0 N2BEGb[5]
rlabel metal1 6716 8602 6716 8602 0 N2BEGb[6]
rlabel metal1 7176 8330 7176 8330 0 N2BEGb[7]
rlabel metal1 8004 8058 8004 8058 0 N4BEG[0]
rlabel metal2 13478 10142 13478 10142 0 N4BEG[10]
rlabel metal2 13754 10244 13754 10244 0 N4BEG[11]
rlabel metal2 14030 10278 14030 10278 0 N4BEG[12]
rlabel metal2 13386 7854 13386 7854 0 N4BEG[13]
rlabel metal1 14122 9758 14122 9758 0 N4BEG[14]
rlabel metal1 14582 6630 14582 6630 0 N4BEG[15]
rlabel metal1 7452 8330 7452 8330 0 N4BEG[1]
rlabel metal1 9936 9690 9936 9690 0 N4BEG[2]
rlabel metal1 10396 10438 10396 10438 0 N4BEG[3]
rlabel metal1 7866 8330 7866 8330 0 N4BEG[4]
rlabel metal2 9798 8670 9798 8670 0 N4BEG[5]
rlabel metal1 8188 8330 8188 8330 0 N4BEG[6]
rlabel metal2 12650 10380 12650 10380 0 N4BEG[7]
rlabel metal1 13432 5338 13432 5338 0 N4BEG[8]
rlabel metal2 13846 8058 13846 8058 0 N4BEG[9]
rlabel metal1 13524 7174 13524 7174 0 NN4BEG[0]
rlabel metal1 17572 8330 17572 8330 0 NN4BEG[10]
rlabel metal1 17802 8602 17802 8602 0 NN4BEG[11]
rlabel metal1 18216 8602 18216 8602 0 NN4BEG[12]
rlabel metal1 18814 8058 18814 8058 0 NN4BEG[13]
rlabel metal1 19228 8058 19228 8058 0 NN4BEG[14]
rlabel metal1 19366 8330 19366 8330 0 NN4BEG[15]
rlabel metal1 15364 8602 15364 8602 0 NN4BEG[1]
rlabel metal1 15502 8058 15502 8058 0 NN4BEG[2]
rlabel metal1 16146 7514 16146 7514 0 NN4BEG[3]
rlabel metal1 14766 10234 14766 10234 0 NN4BEG[4]
rlabel metal2 14490 9248 14490 9248 0 NN4BEG[5]
rlabel metal1 14996 8602 14996 8602 0 NN4BEG[6]
rlabel metal1 16330 8330 16330 8330 0 NN4BEG[7]
rlabel metal2 16054 9146 16054 9146 0 NN4BEG[8]
rlabel metal2 16330 9180 16330 9180 0 NN4BEG[9]
rlabel metal3 19711 8772 19711 8772 0 S1END[0]
rlabel metal1 20010 8466 20010 8466 0 S1END[1]
rlabel metal1 19458 6358 19458 6358 0 S1END[2]
rlabel metal1 19136 6766 19136 6766 0 S1END[3]
rlabel metal1 22724 8534 22724 8534 0 S2END[0]
rlabel metal2 23598 8959 23598 8959 0 S2END[1]
rlabel metal2 23414 9078 23414 9078 0 S2END[2]
rlabel metal2 25530 9078 25530 9078 0 S2END[3]
rlabel metal1 24380 7786 24380 7786 0 S2END[4]
rlabel metal1 24656 7854 24656 7854 0 S2END[5]
rlabel metal1 26496 8466 26496 8466 0 S2END[6]
rlabel metal2 24840 9690 24840 9690 0 S2END[7]
rlabel metal1 21068 7922 21068 7922 0 S2MID[0]
rlabel metal2 21206 10108 21206 10108 0 S2MID[1]
rlabel metal2 21666 9503 21666 9503 0 S2MID[2]
rlabel metal2 21811 10540 21811 10540 0 S2MID[3]
rlabel metal2 22034 9496 22034 9496 0 S2MID[4]
rlabel metal2 22356 7378 22356 7378 0 S2MID[5]
rlabel metal1 23276 7922 23276 7922 0 S2MID[6]
rlabel metal1 22678 8466 22678 8466 0 S2MID[7]
rlabel metal1 26266 9894 26266 9894 0 S4END[0]
rlabel metal2 29164 7786 29164 7786 0 S4END[10]
rlabel metal1 29256 6766 29256 6766 0 S4END[11]
rlabel metal1 29716 6766 29716 6766 0 S4END[12]
rlabel metal2 30038 8398 30038 8398 0 S4END[13]
rlabel metal1 31924 8466 31924 8466 0 S4END[14]
rlabel metal2 31510 8602 31510 8602 0 S4END[15]
rlabel metal1 26910 7922 26910 7922 0 S4END[1]
rlabel metal1 26404 8534 26404 8534 0 S4END[2]
rlabel metal1 26680 7378 26680 7378 0 S4END[3]
rlabel metal1 26542 7446 26542 7446 0 S4END[4]
rlabel metal1 30820 8466 30820 8466 0 S4END[5]
rlabel metal1 28060 7446 28060 7446 0 S4END[6]
rlabel metal1 27968 5746 27968 5746 0 S4END[7]
rlabel metal2 29210 9112 29210 9112 0 S4END[8]
rlabel metal1 28934 6698 28934 6698 0 S4END[9]
rlabel metal2 31602 8806 31602 8806 0 SS4END[0]
rlabel metal2 33718 8262 33718 8262 0 SS4END[10]
rlabel metal2 36938 9350 36938 9350 0 SS4END[11]
rlabel metal1 33718 8466 33718 8466 0 SS4END[12]
rlabel metal1 34684 6834 34684 6834 0 SS4END[13]
rlabel metal1 33994 8534 33994 8534 0 SS4END[14]
rlabel metal2 37306 9452 37306 9452 0 SS4END[15]
rlabel metal2 30038 10448 30038 10448 0 SS4END[1]
rlabel metal2 30406 8959 30406 8959 0 SS4END[2]
rlabel metal1 30958 6290 30958 6290 0 SS4END[3]
rlabel metal2 34822 9248 34822 9248 0 SS4END[4]
rlabel metal1 31924 8942 31924 8942 0 SS4END[5]
rlabel metal2 34914 9282 34914 9282 0 SS4END[6]
rlabel metal3 32407 8636 32407 8636 0 SS4END[7]
rlabel metal1 32154 8534 32154 8534 0 SS4END[8]
rlabel metal2 32338 9962 32338 9962 0 SS4END[9]
rlabel metal2 13938 4199 13938 4199 0 UserCLK
rlabel metal1 10534 3944 10534 3944 0 UserCLK_regs
rlabel metal2 35650 8160 35650 8160 0 UserCLKo
rlabel metal1 24242 5746 24242 5746 0 _000_
rlabel metal1 24334 6256 24334 6256 0 _001_
rlabel metal1 22379 5338 22379 5338 0 _002_
rlabel metal1 20562 5338 20562 5338 0 _003_
rlabel metal1 26427 3910 26427 3910 0 _004_
rlabel metal1 18088 4658 18088 4658 0 _005_
rlabel metal1 24748 4046 24748 4046 0 _006_
rlabel metal1 24242 6358 24242 6358 0 _007_
rlabel metal2 21666 5984 21666 5984 0 _008_
rlabel metal2 23966 6086 23966 6086 0 _009_
rlabel metal1 21896 5338 21896 5338 0 _010_
rlabel metal2 24794 5508 24794 5508 0 _011_
rlabel metal1 24288 5882 24288 5882 0 _012_
rlabel metal1 21758 4250 21758 4250 0 _013_
rlabel metal1 22172 4794 22172 4794 0 _014_
rlabel metal1 21896 5746 21896 5746 0 _015_
rlabel metal2 22034 5372 22034 5372 0 _016_
rlabel metal1 22310 4250 22310 4250 0 _017_
rlabel metal2 22126 4284 22126 4284 0 _018_
rlabel metal1 22540 4250 22540 4250 0 _019_
rlabel metal1 27186 3910 27186 3910 0 _020_
rlabel metal1 25622 4998 25622 4998 0 _021_
rlabel metal1 25810 4148 25810 4148 0 _022_
rlabel metal1 25622 4250 25622 4250 0 _023_
rlabel metal1 26266 4250 26266 4250 0 _024_
rlabel metal1 26266 4012 26266 4012 0 _025_
rlabel metal1 18354 4726 18354 4726 0 _026_
rlabel metal1 18906 5202 18906 5202 0 _027_
rlabel metal1 17986 5100 17986 5100 0 _028_
rlabel metal2 19274 5032 19274 5032 0 _029_
rlabel metal1 18722 5270 18722 5270 0 _030_
rlabel metal1 18308 5202 18308 5202 0 _031_
rlabel metal2 12006 6902 12006 6902 0 clknet_0_UserCLK
rlabel metal2 13478 7344 13478 7344 0 clknet_0_UserCLK_regs
rlabel metal1 10258 6290 10258 6290 0 clknet_1_0__leaf_UserCLK
rlabel metal1 11316 7922 11316 7922 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal1 11362 6188 11362 6188 0 clknet_1_1__leaf_UserCLK_regs
rlabel via2 2530 2907 2530 2907 0 net1
rlabel via2 2070 4539 2070 4539 0 net10
rlabel metal1 19366 2924 19366 2924 0 net100
rlabel metal1 28198 3910 28198 3910 0 net101
rlabel metal2 26542 7123 26542 7123 0 net102
rlabel metal2 21482 4811 21482 4811 0 net103
rlabel metal2 19090 2023 19090 2023 0 net104
rlabel metal2 30130 9690 30130 9690 0 net105
rlabel metal1 10396 3026 10396 3026 0 net106
rlabel metal1 6256 4114 6256 4114 0 net107
rlabel metal2 4830 3230 4830 3230 0 net108
rlabel metal2 14214 2448 14214 2448 0 net109
rlabel metal2 2530 4029 2530 4029 0 net11
rlabel metal3 13524 4216 13524 4216 0 net110
rlabel metal2 17526 2210 17526 2210 0 net111
rlabel metal2 15686 2210 15686 2210 0 net112
rlabel metal1 16629 2414 16629 2414 0 net113
rlabel metal1 17250 2516 17250 2516 0 net114
rlabel metal1 42550 2346 42550 2346 0 net115
rlabel metal1 43148 4114 43148 4114 0 net116
rlabel metal1 42872 4590 42872 4590 0 net117
rlabel metal2 43194 4964 43194 4964 0 net118
rlabel metal2 42918 4998 42918 4998 0 net119
rlabel metal2 32982 3553 32982 3553 0 net12
rlabel via2 43286 5219 43286 5219 0 net120
rlabel metal1 43378 5746 43378 5746 0 net121
rlabel metal1 19366 1326 19366 1326 0 net122
rlabel metal1 42918 6256 42918 6256 0 net123
rlabel metal2 43332 4692 43332 4692 0 net124
rlabel metal2 42734 6273 42734 6273 0 net125
rlabel metal1 41998 2380 41998 2380 0 net126
rlabel via2 43102 6715 43102 6715 0 net127
rlabel metal2 42090 7106 42090 7106 0 net128
rlabel metal1 42964 7854 42964 7854 0 net129
rlabel metal1 32430 2380 32430 2380 0 net13
rlabel metal1 43056 7786 43056 7786 0 net130
rlabel metal2 42458 7820 42458 7820 0 net131
rlabel metal1 42780 8466 42780 8466 0 net132
rlabel metal2 43010 8670 43010 8670 0 net133
rlabel metal1 41998 8534 41998 8534 0 net134
rlabel metal2 42550 9112 42550 9112 0 net135
rlabel via2 42918 7395 42918 7395 0 net136
rlabel metal1 42550 3060 42550 3060 0 net137
rlabel metal2 42182 7905 42182 7905 0 net138
rlabel metal1 41860 7854 41860 7854 0 net139
rlabel metal1 26864 9962 26864 9962 0 net14
rlabel metal1 42918 2448 42918 2448 0 net140
rlabel metal1 43930 2006 43930 2006 0 net141
rlabel metal1 42918 2992 42918 2992 0 net142
rlabel metal2 41998 3298 41998 3298 0 net143
rlabel metal1 42918 3536 42918 3536 0 net144
rlabel metal2 37030 2023 37030 2023 0 net145
rlabel metal1 42918 4080 42918 4080 0 net146
rlabel metal1 37076 3366 37076 3366 0 net147
rlabel metal2 42642 7684 42642 7684 0 net148
rlabel metal1 39054 3162 39054 3162 0 net149
rlabel metal1 6762 6732 6762 6732 0 net15
rlabel metal2 40434 5474 40434 5474 0 net150
rlabel metal1 42136 3910 42136 3910 0 net151
rlabel metal2 41538 8228 41538 8228 0 net152
rlabel metal1 41952 7514 41952 7514 0 net153
rlabel metal1 42044 3638 42044 3638 0 net154
rlabel metal2 41630 5814 41630 5814 0 net155
rlabel metal2 42366 7140 42366 7140 0 net156
rlabel metal1 41814 3706 41814 3706 0 net157
rlabel metal1 38962 6664 38962 6664 0 net158
rlabel metal2 36754 5083 36754 5083 0 net159
rlabel metal1 1748 7310 1748 7310 0 net16
rlabel metal1 37858 3978 37858 3978 0 net160
rlabel metal2 38594 4029 38594 4029 0 net161
rlabel metal1 39054 3434 39054 3434 0 net162
rlabel metal2 41170 5066 41170 5066 0 net163
rlabel metal1 41860 3162 41860 3162 0 net164
rlabel metal1 38594 3128 38594 3128 0 net165
rlabel metal1 42044 3978 42044 3978 0 net166
rlabel metal2 2070 7684 2070 7684 0 net167
rlabel metal2 3864 5746 3864 5746 0 net168
rlabel metal1 15318 4726 15318 4726 0 net169
rlabel metal2 2530 6477 2530 6477 0 net17
rlabel metal2 5244 2924 5244 2924 0 net170
rlabel metal2 29486 2125 29486 2125 0 net171
rlabel metal1 12052 3910 12052 3910 0 net172
rlabel metal1 37720 7990 37720 7990 0 net173
rlabel metal2 4370 8874 4370 8874 0 net174
rlabel metal1 6992 7378 6992 7378 0 net175
rlabel metal1 5842 9214 5842 9214 0 net176
rlabel metal2 15594 714 15594 714 0 net177
rlabel metal1 34132 4590 34132 4590 0 net178
rlabel metal2 5658 8806 5658 8806 0 net179
rlabel metal1 39238 6800 39238 6800 0 net18
rlabel metal1 6624 7854 6624 7854 0 net180
rlabel metal1 36984 7514 36984 7514 0 net181
rlabel metal1 7682 3706 7682 3706 0 net182
rlabel metal1 37766 4454 37766 4454 0 net183
rlabel metal1 10948 3910 10948 3910 0 net184
rlabel metal2 14398 9486 14398 9486 0 net185
rlabel metal2 17986 9197 17986 9197 0 net186
rlabel metal2 15502 1496 15502 1496 0 net187
rlabel metal1 31878 6732 31878 6732 0 net188
rlabel metal1 7636 5066 7636 5066 0 net189
rlabel metal1 5244 5678 5244 5678 0 net19
rlabel metal2 37398 7191 37398 7191 0 net190
rlabel metal2 13202 3876 13202 3876 0 net191
rlabel metal2 26266 1343 26266 1343 0 net192
rlabel metal3 33534 3060 33534 3060 0 net193
rlabel metal1 7774 5882 7774 5882 0 net194
rlabel metal1 35466 4998 35466 4998 0 net195
rlabel metal1 7820 5814 7820 5814 0 net196
rlabel metal2 19366 3961 19366 3961 0 net197
rlabel metal1 10028 5338 10028 5338 0 net198
rlabel via2 31786 5355 31786 5355 0 net199
rlabel metal2 6670 4964 6670 4964 0 net2
rlabel metal2 12742 7582 12742 7582 0 net20
rlabel metal2 10626 6154 10626 6154 0 net200
rlabel metal1 14076 5202 14076 5202 0 net201
rlabel metal1 13984 3706 13984 3706 0 net202
rlabel metal2 12972 2414 12972 2414 0 net203
rlabel metal1 17940 8398 17940 8398 0 net204
rlabel metal2 17526 8670 17526 8670 0 net205
rlabel metal2 18170 8874 18170 8874 0 net206
rlabel metal3 19159 7004 19159 7004 0 net207
rlabel metal1 19274 7888 19274 7888 0 net208
rlabel metal2 19642 8772 19642 8772 0 net209
rlabel via2 2438 7803 2438 7803 0 net21
rlabel metal2 13754 9010 13754 9010 0 net210
rlabel metal1 19182 9826 19182 9826 0 net211
rlabel metal1 19366 510 19366 510 0 net212
rlabel metal1 17664 4250 17664 4250 0 net213
rlabel metal1 19596 8058 19596 8058 0 net214
rlabel metal1 15548 4794 15548 4794 0 net215
rlabel metal2 15778 9010 15778 9010 0 net216
rlabel metal2 15870 9044 15870 9044 0 net217
rlabel metal2 16514 9044 16514 9044 0 net218
rlabel metal2 32798 1683 32798 1683 0 net219
rlabel metal3 19780 2856 19780 2856 0 net22
rlabel metal2 17710 8296 17710 8296 0 net220
rlabel metal1 13340 8466 13340 8466 0 net23
rlabel metal1 14030 7412 14030 7412 0 net24
rlabel metal1 4416 7854 4416 7854 0 net25
rlabel metal1 17756 5678 17756 5678 0 net26
rlabel metal1 17802 6290 17802 6290 0 net27
rlabel via2 16974 7395 16974 7395 0 net28
rlabel metal1 21850 3570 21850 3570 0 net29
rlabel metal1 7544 4590 7544 4590 0 net3
rlabel metal2 6210 3927 6210 3927 0 net30
rlabel metal2 23506 850 23506 850 0 net31
rlabel metal2 1702 2448 1702 2448 0 net32
rlabel metal1 5152 5202 5152 5202 0 net33
rlabel metal1 2576 4250 2576 4250 0 net34
rlabel metal1 18446 6358 18446 6358 0 net35
rlabel metal1 8142 3094 8142 3094 0 net36
rlabel metal2 18354 7769 18354 7769 0 net37
rlabel metal2 19274 6902 19274 6902 0 net38
rlabel metal1 14030 6392 14030 6392 0 net39
rlabel metal2 2530 1462 2530 1462 0 net4
rlabel metal1 24748 4590 24748 4590 0 net40
rlabel metal1 25668 6766 25668 6766 0 net41
rlabel metal2 20930 3876 20930 3876 0 net42
rlabel metal2 23874 3774 23874 3774 0 net43
rlabel metal1 9062 3672 9062 3672 0 net44
rlabel metal1 32246 7208 32246 7208 0 net45
rlabel via1 20907 6222 20907 6222 0 net46
rlabel metal1 20976 7310 20976 7310 0 net47
rlabel metal2 9246 7633 9246 7633 0 net48
rlabel metal1 39514 5066 39514 5066 0 net49
rlabel metal2 1610 2040 1610 2040 0 net5
rlabel metal2 38778 3536 38778 3536 0 net50
rlabel metal2 10442 4114 10442 4114 0 net51
rlabel metal1 8740 5610 8740 5610 0 net52
rlabel metal1 32108 6086 32108 6086 0 net53
rlabel metal1 18814 8500 18814 8500 0 net54
rlabel metal1 1932 5746 1932 5746 0 net55
rlabel metal2 13110 4760 13110 4760 0 net56
rlabel metal2 9430 4165 9430 4165 0 net57
rlabel metal2 13754 7820 13754 7820 0 net58
rlabel metal1 17066 6766 17066 6766 0 net59
rlabel metal1 7084 2414 7084 2414 0 net6
rlabel via2 17618 6307 17618 6307 0 net60
rlabel metal1 39330 5576 39330 5576 0 net61
rlabel metal1 22310 7412 22310 7412 0 net62
rlabel via2 32614 4131 32614 4131 0 net63
rlabel metal1 29762 4624 29762 4624 0 net64
rlabel metal1 21068 8398 21068 8398 0 net65
rlabel metal1 29498 5134 29498 5134 0 net66
rlabel metal1 20746 8330 20746 8330 0 net67
rlabel metal1 28750 5134 28750 5134 0 net68
rlabel via1 20942 4590 20942 4590 0 net69
rlabel metal2 1794 3808 1794 3808 0 net7
rlabel metal2 29762 4964 29762 4964 0 net70
rlabel metal1 27278 6120 27278 6120 0 net71
rlabel metal1 29256 7718 29256 7718 0 net72
rlabel metal2 28014 4794 28014 4794 0 net73
rlabel metal1 20562 918 20562 918 0 net74
rlabel metal2 28980 6188 28980 6188 0 net75
rlabel metal2 31786 8721 31786 8721 0 net76
rlabel metal2 19458 2516 19458 2516 0 net77
rlabel metal1 38732 6290 38732 6290 0 net78
rlabel metal1 8142 5270 8142 5270 0 net79
rlabel metal1 20378 6188 20378 6188 0 net8
rlabel metal1 28198 6324 28198 6324 0 net80
rlabel metal1 12926 4114 12926 4114 0 net81
rlabel metal2 38778 6681 38778 6681 0 net82
rlabel metal1 19458 7956 19458 7956 0 net83
rlabel metal2 18354 3366 18354 3366 0 net84
rlabel metal2 29026 8806 29026 8806 0 net85
rlabel metal1 29164 6630 29164 6630 0 net86
rlabel via1 33454 4114 33454 4114 0 net87
rlabel metal2 33258 8602 33258 8602 0 net88
rlabel metal2 37030 4590 37030 4590 0 net89
rlabel metal3 17388 6324 17388 6324 0 net9
rlabel metal3 15180 3400 15180 3400 0 net90
rlabel metal1 25450 7922 25450 7922 0 net91
rlabel metal2 34178 8840 34178 8840 0 net92
rlabel metal2 28750 3774 28750 3774 0 net93
rlabel via1 26554 6766 26554 6766 0 net94
rlabel metal2 19458 9554 19458 9554 0 net95
rlabel metal2 31418 5440 31418 5440 0 net96
rlabel metal1 13628 4046 13628 4046 0 net97
rlabel via1 34282 7310 34282 7310 0 net98
rlabel metal2 35926 8806 35926 8806 0 net99
<< properties >>
string FIXED_BBOX 0 0 45000 11250
<< end >>
