module N_term_EF_SRAM (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;

 sky130_fd_sc_hd__buf_1 _00_ (.A(FrameData[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 _01_ (.A(FrameData[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 _02_ (.A(FrameData[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 _03_ (.A(FrameData[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 _04_ (.A(FrameData[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 _05_ (.A(FrameData[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(FrameData[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 _07_ (.A(FrameData[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 _08_ (.A(FrameData[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 _09_ (.A(FrameData[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 _10_ (.A(FrameData[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 _11_ (.A(FrameData[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 _12_ (.A(FrameData[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 _13_ (.A(FrameData[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 _14_ (.A(FrameData[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 _15_ (.A(FrameData[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 _16_ (.A(FrameData[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 _17_ (.A(FrameData[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 _18_ (.A(FrameData[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 _19_ (.A(FrameData[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 _20_ (.A(FrameData[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 _21_ (.A(FrameData[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 _22_ (.A(FrameData[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _23_ (.A(FrameData[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 _24_ (.A(FrameData[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 _25_ (.A(FrameData[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 _26_ (.A(FrameData[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _27_ (.A(FrameData[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _28_ (.A(FrameData[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 _29_ (.A(FrameData[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 _30_ (.A(FrameData[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 _31_ (.A(FrameData[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 _32_ (.A(FrameStrobe[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 _33_ (.A(FrameStrobe[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 _34_ (.A(FrameStrobe[2]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _35_ (.A(FrameStrobe[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 _36_ (.A(FrameStrobe[4]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 _37_ (.A(FrameStrobe[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 _38_ (.A(FrameStrobe[6]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 _39_ (.A(FrameStrobe[7]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _40_ (.A(FrameStrobe[8]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _41_ (.A(FrameStrobe[9]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _42_ (.A(FrameStrobe[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 _43_ (.A(FrameStrobe[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 _44_ (.A(FrameStrobe[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _45_ (.A(FrameStrobe[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _46_ (.A(FrameStrobe[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 _47_ (.A(FrameStrobe[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _48_ (.A(FrameStrobe[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _49_ (.A(FrameStrobe[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _50_ (.A(FrameStrobe[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _51_ (.A(FrameStrobe[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _52_ (.A(N1END[3]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _53_ (.A(N1END[2]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _54_ (.A(N1END[1]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 _55_ (.A(N1END[0]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _56_ (.A(N2MID[7]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _57_ (.A(N2MID[6]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _58_ (.A(N2MID[5]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _59_ (.A(N2MID[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 _60_ (.A(N2MID[3]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 _61_ (.A(N2MID[2]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 _62_ (.A(N2MID[1]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 _63_ (.A(N2MID[0]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _64_ (.A(N2END[7]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _65_ (.A(N2END[6]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _66_ (.A(N2END[5]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 _67_ (.A(N2END[4]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 _68_ (.A(N2END[3]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _69_ (.A(N2END[2]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 _70_ (.A(N2END[1]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 _71_ (.A(N2END[0]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _72_ (.A(N4END[15]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _73_ (.A(N4END[14]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _74_ (.A(N4END[13]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _75_ (.A(N4END[12]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _76_ (.A(N4END[11]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _77_ (.A(N4END[10]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _78_ (.A(N4END[9]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _79_ (.A(N4END[8]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _80_ (.A(N4END[7]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _81_ (.A(N4END[6]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _82_ (.A(N4END[5]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _83_ (.A(N4END[4]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _84_ (.A(N4END[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _85_ (.A(N4END[2]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _86_ (.A(N4END[1]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _87_ (.A(N4END[0]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 _88_ (.A(UserCLK),
    .X(net89));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_107 ();
 sky130_fd_sc_hd__buf_2 output1 (.A(net1),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(UserCLKo));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(FrameData[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(FrameData[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(FrameData[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(FrameData[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(FrameData[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(FrameData[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(FrameData[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(FrameData[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(FrameData[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(FrameData[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(FrameData[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(FrameData[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(FrameData[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(FrameData[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(FrameData[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(FrameData[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(FrameData[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(FrameData[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(FrameData[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(FrameData[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(FrameData[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(FrameData[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(FrameData[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(FrameStrobe[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(N4END[2]));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
endmodule
