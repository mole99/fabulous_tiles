* NGSPICE file created from S_term_single.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

.subckt S_term_single Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_10_306 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_5_387 VPWR VGND sg13g2_decap_8
XFILLER_5_310 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_6_129 VPWR VGND sg13g2_fill_1
X_062_ S2MID[2] net62 VPWR VGND sg13g2_buf_1
XFILLER_9_77 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_7_246 VPWR VGND sg13g2_decap_8
X_045_ FrameStrobe[12] net36 VPWR VGND sg13g2_buf_1
XFILLER_3_441 VPWR VGND sg13g2_decap_8
XFILLER_4_216 VPWR VGND sg13g2_decap_8
X_028_ FrameData[27] net20 VPWR VGND sg13g2_buf_1
XANTENNA_5 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XFILLER_3_260 VPWR VGND sg13g2_decap_8
Xoutput20 net20 FrameData_O[27] VPWR VGND sg13g2_buf_1
Xoutput42 net42 FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
Xoutput97 net97 NN4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput75 net75 N4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput86 net86 N4BEG[7] VPWR VGND sg13g2_buf_1
Xoutput64 net64 N2BEG[7] VPWR VGND sg13g2_buf_1
Xoutput53 net53 N1BEG[0] VPWR VGND sg13g2_buf_1
Xoutput7 net7 FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_0_252 VPWR VGND sg13g2_decap_8
Xoutput31 net31 FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_5_366 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_8_182 VPWR VGND sg13g2_decap_8
XFILLER_6_108 VPWR VGND sg13g2_decap_8
XFILLER_2_314 VPWR VGND sg13g2_decap_4
XFILLER_5_163 VPWR VGND sg13g2_decap_8
XFILLER_9_56 VPWR VGND sg13g2_decap_8
X_061_ S2MID[3] net61 VPWR VGND sg13g2_buf_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_8
XFILLER_4_409 VPWR VGND sg13g2_decap_8
XFILLER_7_225 VPWR VGND sg13g2_decap_8
X_044_ FrameStrobe[11] net35 VPWR VGND sg13g2_buf_1
XFILLER_3_420 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_4
X_027_ FrameData[26] net19 VPWR VGND sg13g2_buf_1
XANTENNA_6 VPWR VGND FrameData[29] sg13g2_antennanp
XFILLER_6_35 VPWR VGND sg13g2_decap_8
Xoutput21 net21 FrameData_O[28] VPWR VGND sg13g2_buf_1
Xoutput43 net43 FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
Xoutput98 net98 NN4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput76 net76 N4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput87 net87 N4BEG[8] VPWR VGND sg13g2_buf_1
Xoutput65 net65 N2BEGb[0] VPWR VGND sg13g2_buf_1
Xoutput54 net54 N1BEG[1] VPWR VGND sg13g2_buf_1
Xoutput10 net10 FrameData_O[18] VPWR VGND sg13g2_buf_1
Xoutput8 net8 FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_0_231 VPWR VGND sg13g2_decap_8
Xoutput32 net32 FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_5_345 VPWR VGND sg13g2_fill_2
XFILLER_8_161 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_2_337 VPWR VGND sg13g2_decap_8
XFILLER_2_359 VPWR VGND sg13g2_decap_8
XFILLER_1_381 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_7_429 VPWR VGND sg13g2_decap_8
X_060_ S2MID[4] net60 VPWR VGND sg13g2_buf_1
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_189 VPWR VGND sg13g2_decap_4
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_7_204 VPWR VGND sg13g2_decap_8
X_043_ FrameStrobe[10] net34 VPWR VGND sg13g2_buf_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
X_026_ FrameData[25] net18 VPWR VGND sg13g2_buf_1
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XANTENNA_7 VPWR VGND FrameData[16] sg13g2_antennanp
XFILLER_3_295 VPWR VGND sg13g2_decap_8
Xoutput22 net22 FrameData_O[29] VPWR VGND sg13g2_buf_1
Xoutput44 net44 FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
Xoutput33 net33 FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
Xoutput99 net99 NN4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput77 net77 N4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput88 net88 N4BEG[9] VPWR VGND sg13g2_buf_1
Xoutput66 net66 N2BEGb[1] VPWR VGND sg13g2_buf_1
Xoutput55 net55 N1BEG[2] VPWR VGND sg13g2_buf_1
Xoutput11 net11 FrameData_O[19] VPWR VGND sg13g2_buf_1
Xoutput9 net9 FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_8_365 VPWR VGND sg13g2_fill_2
XFILLER_8_343 VPWR VGND sg13g2_fill_1
XFILLER_8_332 VPWR VGND sg13g2_decap_8
X_009_ FrameData[8] net31 VPWR VGND sg13g2_buf_1
XFILLER_8_140 VPWR VGND sg13g2_decap_8
XFILLER_5_335 VPWR VGND sg13g2_decap_4
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_5_121 VPWR VGND sg13g2_decap_4
XFILLER_1_360 VPWR VGND sg13g2_decap_8
XFILLER_4_80 VPWR VGND sg13g2_decap_8
XFILLER_7_408 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_9_14 VPWR VGND sg13g2_decap_8
X_042_ FrameStrobe[9] net52 VPWR VGND sg13g2_buf_1
XFILLER_6_293 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
X_025_ FrameData[24] net17 VPWR VGND sg13g2_buf_1
XANTENNA_8 VPWR VGND FrameData[21] sg13g2_antennanp
XFILLER_3_274 VPWR VGND sg13g2_decap_8
Xoutput34 net34 FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
Xoutput45 net45 FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
Xoutput89 net89 NN4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput78 net78 N4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput67 net67 N2BEGb[2] VPWR VGND sg13g2_buf_1
Xoutput56 net56 N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_0_266 VPWR VGND sg13g2_decap_8
Xoutput23 net23 FrameData_O[2] VPWR VGND sg13g2_buf_1
Xoutput12 net12 FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_8_311 VPWR VGND sg13g2_decap_8
X_008_ FrameData[7] net30 VPWR VGND sg13g2_buf_1
XFILLER_5_347 VPWR VGND sg13g2_fill_1
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_8_196 VPWR VGND sg13g2_decap_8
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_4
XFILLER_6_442 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_9_291 VPWR VGND sg13g2_decap_8
XFILLER_7_239 VPWR VGND sg13g2_decap_8
X_041_ FrameStrobe[8] net51 VPWR VGND sg13g2_buf_1
XFILLER_3_434 VPWR VGND sg13g2_decap_8
XFILLER_6_272 VPWR VGND sg13g2_decap_8
XFILLER_4_209 VPWR VGND sg13g2_decap_8
XFILLER_10_91 VPWR VGND sg13g2_decap_8
XANTENNA_9 VPWR VGND FrameData[24] sg13g2_antennanp
X_024_ FrameData[23] net16 VPWR VGND sg13g2_buf_1
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_3_231 VPWR VGND sg13g2_decap_4
XFILLER_3_253 VPWR VGND sg13g2_fill_2
Xoutput24 net24 FrameData_O[30] VPWR VGND sg13g2_buf_1
Xoutput35 net35 FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
Xoutput46 net46 FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
Xoutput57 net57 N2BEG[0] VPWR VGND sg13g2_buf_1
Xoutput13 net13 FrameData_O[20] VPWR VGND sg13g2_buf_1
Xoutput79 net79 N4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput68 net68 N2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_0_245 VPWR VGND sg13g2_decap_8
X_007_ FrameData[6] net29 VPWR VGND sg13g2_buf_1
XFILLER_7_92 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_4
XFILLER_5_359 VPWR VGND sg13g2_decap_8
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_8_175 VPWR VGND sg13g2_decap_8
XFILLER_4_381 VPWR VGND sg13g2_decap_8
XFILLER_2_307 VPWR VGND sg13g2_decap_8
XFILLER_2_318 VPWR VGND sg13g2_fill_1
XFILLER_5_156 VPWR VGND sg13g2_decap_8
XFILLER_1_395 VPWR VGND sg13g2_decap_8
XFILLER_9_49 VPWR VGND sg13g2_decap_8
XFILLER_6_421 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_7_218 VPWR VGND sg13g2_decap_8
X_040_ FrameStrobe[7] net50 VPWR VGND sg13g2_buf_1
XFILLER_3_413 VPWR VGND sg13g2_decap_8
XFILLER_6_251 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_0_438 VPWR VGND sg13g2_fill_1
X_023_ FrameData[22] net15 VPWR VGND sg13g2_buf_1
XFILLER_10_70 VPWR VGND sg13g2_decap_8
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_3_210 VPWR VGND sg13g2_decap_8
Xoutput25 net25 FrameData_O[31] VPWR VGND sg13g2_buf_1
Xoutput36 net36 FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
Xoutput47 net47 FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
Xoutput69 net69 N2BEGb[4] VPWR VGND sg13g2_buf_1
Xoutput58 net58 N2BEG[1] VPWR VGND sg13g2_buf_1
Xoutput14 net14 FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_0_224 VPWR VGND sg13g2_decap_8
X_006_ FrameData[5] net28 VPWR VGND sg13g2_buf_1
XFILLER_8_154 VPWR VGND sg13g2_decap_8
XFILLER_4_360 VPWR VGND sg13g2_decap_8
XFILLER_1_374 VPWR VGND sg13g2_decap_8
XFILLER_4_94 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_6_400 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_1_193 VPWR VGND sg13g2_decap_8
XFILLER_10_292 VPWR VGND sg13g2_decap_8
X_099_ SS4END[5] net90 VPWR VGND sg13g2_buf_1
XFILLER_6_230 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
X_022_ FrameData[21] net14 VPWR VGND sg13g2_buf_1
XFILLER_3_255 VPWR VGND sg13g2_fill_1
XFILLER_3_288 VPWR VGND sg13g2_decap_8
Xoutput15 net15 FrameData_O[22] VPWR VGND sg13g2_buf_1
Xoutput37 net37 FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
Xoutput48 net48 FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
Xoutput59 net59 N2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_8_325 VPWR VGND sg13g2_fill_2
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xoutput26 net26 FrameData_O[3] VPWR VGND sg13g2_buf_1
X_005_ FrameData[4] net27 VPWR VGND sg13g2_buf_1
XFILLER_7_380 VPWR VGND sg13g2_decap_8
XFILLER_5_339 VPWR VGND sg13g2_fill_2
XFILLER_5_317 VPWR VGND sg13g2_decap_4
XFILLER_8_133 VPWR VGND sg13g2_decap_8
XFILLER_5_114 VPWR VGND sg13g2_decap_8
XFILLER_1_353 VPWR VGND sg13g2_decap_8
XFILLER_9_442 VPWR VGND sg13g2_fill_1
XFILLER_9_431 VPWR VGND sg13g2_decap_8
XFILLER_9_261 VPWR VGND sg13g2_fill_2
XFILLER_1_172 VPWR VGND sg13g2_fill_2
XFILLER_10_271 VPWR VGND sg13g2_decap_8
X_098_ SS4END[6] net104 VPWR VGND sg13g2_buf_1
XFILLER_6_286 VPWR VGND sg13g2_decap_8
XFILLER_3_448 VPWR VGND sg13g2_fill_2
XFILLER_1_63 VPWR VGND sg13g2_decap_8
X_021_ FrameData[20] net13 VPWR VGND sg13g2_buf_1
XFILLER_3_267 VPWR VGND sg13g2_decap_8
Xoutput16 net16 FrameData_O[23] VPWR VGND sg13g2_buf_1
Xoutput38 net38 FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
Xoutput49 net49 FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_0_259 VPWR VGND sg13g2_decap_8
Xoutput27 net27 FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_8_304 VPWR VGND sg13g2_decap_8
X_004_ FrameData[3] net26 VPWR VGND sg13g2_buf_1
XFILLER_8_189 VPWR VGND sg13g2_decap_8
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_5_329 VPWR VGND sg13g2_fill_2
XFILLER_4_395 VPWR VGND sg13g2_decap_8
XFILLER_1_332 VPWR VGND sg13g2_decap_8
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_4_74 VPWR VGND sg13g2_fill_2
XFILLER_6_435 VPWR VGND sg13g2_decap_8
XFILLER_1_151 VPWR VGND sg13g2_decap_8
XFILLER_10_250 VPWR VGND sg13g2_decap_8
XFILLER_3_427 VPWR VGND sg13g2_decap_8
X_097_ SS4END[7] net103 VPWR VGND sg13g2_buf_1
XFILLER_6_265 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_020_ FrameData[19] net11 VPWR VGND sg13g2_buf_1
XFILLER_3_224 VPWR VGND sg13g2_decap_8
XFILLER_3_246 VPWR VGND sg13g2_decap_8
XFILLER_10_84 VPWR VGND sg13g2_decap_8
Xoutput17 net17 FrameData_O[24] VPWR VGND sg13g2_buf_1
Xoutput39 net39 FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
XFILLER_0_238 VPWR VGND sg13g2_decap_8
Xoutput28 net28 FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_8_327 VPWR VGND sg13g2_fill_1
X_003_ FrameData[2] net23 VPWR VGND sg13g2_buf_1
XFILLER_7_85 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_8_168 VPWR VGND sg13g2_decap_8
XFILLER_4_374 VPWR VGND sg13g2_decap_8
XFILLER_7_190 VPWR VGND sg13g2_decap_8
XFILLER_5_149 VPWR VGND sg13g2_decap_8
XFILLER_1_311 VPWR VGND sg13g2_decap_8
XFILLER_1_388 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_fill_1
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_6_414 VPWR VGND sg13g2_decap_8
XFILLER_1_174 VPWR VGND sg13g2_fill_1
XFILLER_1_130 VPWR VGND sg13g2_decap_8
XFILLER_9_241 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_3_406 VPWR VGND sg13g2_decap_8
X_096_ SS4END[8] net102 VPWR VGND sg13g2_buf_1
XFILLER_6_244 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_2_450 VPWR VGND sg13g2_fill_1
XFILLER_10_63 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_decap_8
Xoutput18 net18 FrameData_O[25] VPWR VGND sg13g2_buf_1
X_079_ S4END[9] net85 VPWR VGND sg13g2_buf_1
XFILLER_0_217 VPWR VGND sg13g2_decap_8
Xoutput29 net29 FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_8_339 VPWR VGND sg13g2_decap_4
X_002_ FrameData[1] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_394 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_decap_8
XFILLER_4_353 VPWR VGND sg13g2_decap_8
XFILLER_1_367 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_4_87 VPWR VGND sg13g2_fill_2
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_10_433 VPWR VGND sg13g2_fill_2
XFILLER_10_422 VPWR VGND sg13g2_decap_8
XFILLER_9_220 VPWR VGND sg13g2_decap_8
XFILLER_1_186 VPWR VGND sg13g2_decap_8
XFILLER_10_285 VPWR VGND sg13g2_decap_8
X_095_ SS4END[9] net101 VPWR VGND sg13g2_buf_1
XFILLER_6_223 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_10_42 VPWR VGND sg13g2_decap_8
X_078_ S4END[10] net84 VPWR VGND sg13g2_buf_1
XFILLER_2_270 VPWR VGND sg13g2_decap_4
Xoutput19 net19 FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_8_318 VPWR VGND sg13g2_decap_8
X_001_ FrameData[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_7_373 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_4_332 VPWR VGND sg13g2_decap_8
XFILLER_1_346 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_6_449 VPWR VGND sg13g2_fill_2
XFILLER_9_298 VPWR VGND sg13g2_decap_8
XFILLER_1_165 VPWR VGND sg13g2_decap_8
XFILLER_10_264 VPWR VGND sg13g2_decap_8
X_094_ SS4END[10] net100 VPWR VGND sg13g2_buf_1
XFILLER_6_279 VPWR VGND sg13g2_decap_8
XFILLER_6_202 VPWR VGND sg13g2_decap_8
XFILLER_5_290 VPWR VGND sg13g2_decap_4
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_10_98 VPWR VGND sg13g2_fill_1
XFILLER_10_21 VPWR VGND sg13g2_decap_8
X_077_ S4END[11] net83 VPWR VGND sg13g2_buf_1
XFILLER_2_293 VPWR VGND sg13g2_decap_8
XFILLER_7_352 VPWR VGND sg13g2_decap_8
XFILLER_7_99 VPWR VGND sg13g2_decap_8
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_4_388 VPWR VGND sg13g2_decap_8
XFILLER_1_325 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_4_89 VPWR VGND sg13g2_fill_1
XFILLER_9_255 VPWR VGND sg13g2_fill_2
XFILLER_6_428 VPWR VGND sg13g2_decap_8
XFILLER_1_144 VPWR VGND sg13g2_decap_8
XFILLER_5_450 VPWR VGND sg13g2_fill_1
XFILLER_10_243 VPWR VGND sg13g2_decap_8
X_093_ SS4END[11] net99 VPWR VGND sg13g2_buf_1
XFILLER_6_258 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_10_77 VPWR VGND sg13g2_decap_8
XFILLER_3_217 VPWR VGND sg13g2_decap_8
XFILLER_3_239 VPWR VGND sg13g2_decap_8
XFILLER_2_250 VPWR VGND sg13g2_decap_8
XFILLER_2_261 VPWR VGND sg13g2_decap_4
X_076_ S4END[12] net82 VPWR VGND sg13g2_buf_1
XFILLER_7_78 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
X_059_ S2MID[5] net59 VPWR VGND sg13g2_buf_1
XFILLER_4_312 VPWR VGND sg13g2_decap_4
XFILLER_7_183 VPWR VGND sg13g2_decap_8
XFILLER_4_367 VPWR VGND sg13g2_decap_8
XFILLER_1_304 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_fill_2
XFILLER_6_407 VPWR VGND sg13g2_decap_8
XFILLER_1_123 VPWR VGND sg13g2_decap_8
XFILLER_9_267 VPWR VGND sg13g2_decap_4
XFILLER_9_234 VPWR VGND sg13g2_decap_8
XFILLER_10_222 VPWR VGND sg13g2_decap_8
XFILLER_10_299 VPWR VGND sg13g2_decap_8
X_092_ SS4END[12] net98 VPWR VGND sg13g2_buf_1
XFILLER_6_237 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_2_443 VPWR VGND sg13g2_decap_8
XFILLER_10_56 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_fill_2
X_075_ S4END[13] net81 VPWR VGND sg13g2_buf_1
XANTENNA_40 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_7_387 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_058_ S2MID[6] net58 VPWR VGND sg13g2_buf_1
XFILLER_4_346 VPWR VGND sg13g2_decap_8
XFILLER_7_162 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_4
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_10_415 VPWR VGND sg13g2_decap_8
XFILLER_1_179 VPWR VGND sg13g2_decap_8
XFILLER_9_213 VPWR VGND sg13g2_decap_8
XFILLER_8_290 VPWR VGND sg13g2_decap_8
XFILLER_10_278 VPWR VGND sg13g2_decap_8
X_091_ SS4END[13] net97 VPWR VGND sg13g2_buf_1
XFILLER_6_216 VPWR VGND sg13g2_decap_8
XFILLER_2_422 VPWR VGND sg13g2_decap_8
XFILLER_10_35 VPWR VGND sg13g2_decap_8
X_074_ S4END[14] net80 VPWR VGND sg13g2_buf_1
XFILLER_2_274 VPWR VGND sg13g2_fill_1
XANTENNA_30 VPWR VGND FrameData[24] sg13g2_antennanp
XANTENNA_41 VPWR VGND FrameData[27] sg13g2_antennanp
XFILLER_2_91 VPWR VGND sg13g2_decap_8
XFILLER_7_366 VPWR VGND sg13g2_decap_8
XFILLER_7_333 VPWR VGND sg13g2_fill_1
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_057_ S2MID[7] net57 VPWR VGND sg13g2_buf_1
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_4_325 VPWR VGND sg13g2_decap_8
XFILLER_7_141 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_1_339 VPWR VGND sg13g2_decap_8
XFILLER_8_450 VPWR VGND sg13g2_fill_1
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_4_122 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_4_188 VPWR VGND sg13g2_fill_1
XFILLER_1_158 VPWR VGND sg13g2_decap_8
X_090_ SS4END[14] net96 VPWR VGND sg13g2_buf_1
XFILLER_10_257 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_2_401 VPWR VGND sg13g2_decap_8
XFILLER_5_283 VPWR VGND sg13g2_decap_8
XFILLER_10_14 VPWR VGND sg13g2_decap_8
X_073_ S4END[15] net73 VPWR VGND sg13g2_buf_1
XFILLER_2_286 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XANTENNA_31 VPWR VGND FrameData[25] sg13g2_antennanp
XANTENNA_42 VPWR VGND FrameData[24] sg13g2_antennanp
XANTENNA_20 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XFILLER_7_345 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_decap_8
X_056_ S1END[0] net56 VPWR VGND sg13g2_buf_1
XFILLER_7_197 VPWR VGND sg13g2_decap_8
XFILLER_7_120 VPWR VGND sg13g2_decap_8
XFILLER_3_392 VPWR VGND sg13g2_decap_8
X_039_ FrameStrobe[6] net49 VPWR VGND sg13g2_buf_1
XFILLER_8_91 VPWR VGND sg13g2_decap_8
XFILLER_1_318 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_4_101 VPWR VGND sg13g2_decap_8
XFILLER_9_248 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_5_443 VPWR VGND sg13g2_decap_8
XFILLER_1_137 VPWR VGND sg13g2_decap_8
XFILLER_5_81 VPWR VGND sg13g2_fill_1
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_10_236 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
X_072_ S2END[0] net72 VPWR VGND sg13g2_buf_1
XFILLER_2_265 VPWR VGND sg13g2_fill_1
XANTENNA_21 VPWR VGND FrameData[27] sg13g2_antennanp
XANTENNA_10 VPWR VGND FrameData[25] sg13g2_antennanp
XANTENNA_43 VPWR VGND FrameData[25] sg13g2_antennanp
XANTENNA_32 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_7_49 VPWR VGND sg13g2_decap_8
X_055_ S1END[1] net55 VPWR VGND sg13g2_buf_1
XFILLER_4_305 VPWR VGND sg13g2_decap_8
XFILLER_4_316 VPWR VGND sg13g2_fill_1
XFILLER_7_176 VPWR VGND sg13g2_decap_8
X_038_ FrameStrobe[5] net48 VPWR VGND sg13g2_buf_1
XFILLER_3_371 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_8_441 VPWR VGND sg13g2_decap_8
XFILLER_10_429 VPWR VGND sg13g2_decap_4
XFILLER_9_227 VPWR VGND sg13g2_decap_8
XFILLER_1_116 VPWR VGND sg13g2_decap_8
XFILLER_5_422 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_10_215 VPWR VGND sg13g2_decap_8
XFILLER_2_436 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_decap_8
XFILLER_10_49 VPWR VGND sg13g2_decap_8
X_071_ S2END[1] net71 VPWR VGND sg13g2_buf_1
XFILLER_2_222 VPWR VGND sg13g2_fill_1
XANTENNA_22 VPWR VGND FrameData[24] sg13g2_antennanp
XANTENNA_33 VPWR VGND FrameData[27] sg13g2_antennanp
XANTENNA_44 VPWR VGND FrameData[26] sg13g2_antennanp
XANTENNA_11 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_054_ S1END[2] net54 VPWR VGND sg13g2_buf_1
XFILLER_4_339 VPWR VGND sg13g2_decap_8
XFILLER_7_155 VPWR VGND sg13g2_decap_8
X_037_ FrameStrobe[4] net47 VPWR VGND sg13g2_buf_1
XFILLER_3_350 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_8_431 VPWR VGND sg13g2_decap_4
XFILLER_9_206 VPWR VGND sg13g2_decap_8
XFILLER_5_401 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_8_283 VPWR VGND sg13g2_decap_8
XFILLER_6_209 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_2_415 VPWR VGND sg13g2_decap_8
XFILLER_10_28 VPWR VGND sg13g2_decap_8
X_070_ S2END[2] net70 VPWR VGND sg13g2_buf_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
XANTENNA_12 VPWR VGND FrameData[27] sg13g2_antennanp
XANTENNA_23 VPWR VGND FrameData[25] sg13g2_antennanp
XANTENNA_34 VPWR VGND FrameData[24] sg13g2_antennanp
XANTENNA_45 VPWR VGND FrameData[27] sg13g2_antennanp
XFILLER_7_315 VPWR VGND sg13g2_decap_8
X_053_ S1END[3] net53 VPWR VGND sg13g2_buf_1
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_7_134 VPWR VGND sg13g2_decap_8
X_105_ UserCLK net105 VPWR VGND sg13g2_buf_1
X_036_ FrameStrobe[3] net46 VPWR VGND sg13g2_buf_1
XFILLER_4_115 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
X_019_ FrameData[18] net10 VPWR VGND sg13g2_buf_1
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_5_276 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_fill_2
XFILLER_2_279 VPWR VGND sg13g2_decap_8
XANTENNA_13 VPWR VGND FrameData[29] sg13g2_antennanp
XANTENNA_35 VPWR VGND FrameData[25] sg13g2_antennanp
XANTENNA_24 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_1_290 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
XFILLER_7_338 VPWR VGND sg13g2_decap_8
X_052_ FrameStrobe[19] net43 VPWR VGND sg13g2_buf_1
XFILLER_6_393 VPWR VGND sg13g2_decap_8
X_104_ SS4END[0] net95 VPWR VGND sg13g2_buf_1
XFILLER_7_113 VPWR VGND sg13g2_decap_8
XFILLER_3_330 VPWR VGND sg13g2_decap_8
XFILLER_3_385 VPWR VGND sg13g2_decap_8
X_035_ FrameStrobe[2] net45 VPWR VGND sg13g2_buf_1
XFILLER_8_84 VPWR VGND sg13g2_decap_8
X_018_ FrameData[17] net9 VPWR VGND sg13g2_buf_1
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_3_182 VPWR VGND sg13g2_decap_8
XFILLER_5_436 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
XFILLER_5_63 VPWR VGND sg13g2_decap_8
XFILLER_10_229 VPWR VGND sg13g2_decap_8
XANTENNA_25 VPWR VGND FrameData[27] sg13g2_antennanp
XANTENNA_14 VPWR VGND FrameData[24] sg13g2_antennanp
XANTENNA_36 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_2_42 VPWR VGND sg13g2_decap_8
X_051_ FrameStrobe[18] net42 VPWR VGND sg13g2_buf_1
XFILLER_6_372 VPWR VGND sg13g2_decap_8
XFILLER_6_350 VPWR VGND sg13g2_decap_8
X_103_ SS4END[1] net94 VPWR VGND sg13g2_buf_1
XFILLER_7_169 VPWR VGND sg13g2_decap_8
X_034_ FrameStrobe[1] net44 VPWR VGND sg13g2_buf_1
XFILLER_3_364 VPWR VGND sg13g2_decap_8
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_6_191 VPWR VGND sg13g2_fill_2
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_3_161 VPWR VGND sg13g2_decap_8
X_017_ FrameData[16] net8 VPWR VGND sg13g2_buf_1
XFILLER_5_415 VPWR VGND sg13g2_decap_8
XFILLER_1_109 VPWR VGND sg13g2_decap_8
XFILLER_8_297 VPWR VGND sg13g2_decap_8
XFILLER_8_231 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_2_429 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_2_204 VPWR VGND sg13g2_fill_2
XFILLER_2_237 VPWR VGND sg13g2_fill_1
XANTENNA_26 VPWR VGND FrameData[24] sg13g2_antennanp
XANTENNA_37 VPWR VGND FrameData[27] sg13g2_antennanp
XANTENNA_15 VPWR VGND FrameData[25] sg13g2_antennanp
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
Xoutput100 net100 NN4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_7_329 VPWR VGND sg13g2_decap_4
X_050_ FrameStrobe[17] net41 VPWR VGND sg13g2_buf_1
X_102_ SS4END[2] net93 VPWR VGND sg13g2_buf_1
XFILLER_7_148 VPWR VGND sg13g2_decap_8
X_033_ FrameStrobe[0] net33 VPWR VGND sg13g2_buf_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_4_129 VPWR VGND sg13g2_decap_4
XFILLER_8_435 VPWR VGND sg13g2_fill_2
XFILLER_8_424 VPWR VGND sg13g2_decap_8
X_016_ FrameData[15] net7 VPWR VGND sg13g2_buf_1
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_8_210 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_2_408 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_1_430 VPWR VGND sg13g2_decap_8
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XANTENNA_27 VPWR VGND FrameData[25] sg13g2_antennanp
XANTENNA_38 VPWR VGND FrameData[24] sg13g2_antennanp
Xoutput101 net101 NN4BEG[6] VPWR VGND sg13g2_buf_1
XANTENNA_16 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_7_308 VPWR VGND sg13g2_decap_8
X_101_ SS4END[3] net92 VPWR VGND sg13g2_buf_1
X_032_ FrameData[31] net25 VPWR VGND sg13g2_buf_1
XFILLER_7_127 VPWR VGND sg13g2_decap_8
XFILLER_3_344 VPWR VGND sg13g2_fill_2
XFILLER_8_98 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_6_193 VPWR VGND sg13g2_fill_1
XFILLER_3_399 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_4_108 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
X_015_ FrameData[14] net6 VPWR VGND sg13g2_buf_1
XFILLER_3_196 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_5_77 VPWR VGND sg13g2_decap_4
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_4_291 VPWR VGND sg13g2_decap_8
XFILLER_1_283 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XANTENNA_17 VPWR VGND FrameData[27] sg13g2_antennanp
XANTENNA_39 VPWR VGND FrameData[25] sg13g2_antennanp
Xoutput102 net102 NN4BEG[7] VPWR VGND sg13g2_buf_1
XANTENNA_28 VPWR VGND FrameData[26] sg13g2_antennanp
XFILLER_6_386 VPWR VGND sg13g2_decap_8
X_100_ SS4END[4] net91 VPWR VGND sg13g2_buf_1
X_031_ FrameData[30] net24 VPWR VGND sg13g2_buf_1
XFILLER_7_106 VPWR VGND sg13g2_decap_8
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_6_183 VPWR VGND sg13g2_decap_4
XFILLER_3_323 VPWR VGND sg13g2_decap_8
XFILLER_3_378 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_8_448 VPWR VGND sg13g2_fill_2
X_014_ FrameData[13] net5 VPWR VGND sg13g2_buf_1
XFILLER_3_175 VPWR VGND sg13g2_decap_8
XFILLER_5_429 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_8_278 VPWR VGND sg13g2_fill_1
XFILLER_8_245 VPWR VGND sg13g2_decap_4
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_2_218 VPWR VGND sg13g2_decap_4
XFILLER_4_270 VPWR VGND sg13g2_decap_8
XANTENNA_29 VPWR VGND FrameData[27] sg13g2_antennanp
Xoutput103 net103 NN4BEG[8] VPWR VGND sg13g2_buf_1
XANTENNA_18 VPWR VGND FrameData[24] sg13g2_antennanp
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XFILLER_6_365 VPWR VGND sg13g2_decap_8
XFILLER_6_343 VPWR VGND sg13g2_decap_8
XFILLER_6_321 VPWR VGND sg13g2_decap_8
X_030_ FrameData[29] net22 VPWR VGND sg13g2_buf_1
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_3_302 VPWR VGND sg13g2_decap_8
XFILLER_3_357 VPWR VGND sg13g2_decap_8
XFILLER_6_162 VPWR VGND sg13g2_decap_8
X_013_ FrameData[12] net4 VPWR VGND sg13g2_buf_1
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_5_408 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_8_224 VPWR VGND sg13g2_decap_8
XFILLER_4_430 VPWR VGND sg13g2_decap_8
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_1_444 VPWR VGND sg13g2_fill_2
XANTENNA_19 VPWR VGND FrameData[25] sg13g2_antennanp
XFILLER_9_374 VPWR VGND sg13g2_fill_1
Xoutput104 net104 NN4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_1_274 VPWR VGND sg13g2_decap_4
XFILLER_1_263 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_6_300 VPWR VGND sg13g2_decap_8
X_089_ SS4END[15] net89 VPWR VGND sg13g2_buf_1
XFILLER_8_35 VPWR VGND sg13g2_decap_8
XFILLER_6_141 VPWR VGND sg13g2_decap_8
XFILLER_2_380 VPWR VGND sg13g2_decap_8
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_7_450 VPWR VGND sg13g2_fill_1
X_012_ FrameData[11] net3 VPWR VGND sg13g2_buf_1
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_8_203 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_7_280 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_1_423 VPWR VGND sg13g2_decap_8
XFILLER_1_297 VPWR VGND sg13g2_decap_8
XFILLER_1_242 VPWR VGND sg13g2_decap_8
Xoutput105 net105 UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_3_91 VPWR VGND sg13g2_decap_8
XFILLER_3_337 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
X_088_ S4END[0] net79 VPWR VGND sg13g2_buf_1
XFILLER_0_329 VPWR VGND sg13g2_decap_8
X_011_ FrameData[10] net2 VPWR VGND sg13g2_buf_1
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_189 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
XFILLER_1_402 VPWR VGND sg13g2_decap_8
XFILLER_1_446 VPWR VGND sg13g2_fill_1
XFILLER_4_251 VPWR VGND sg13g2_decap_8
XFILLER_4_284 VPWR VGND sg13g2_decap_8
XFILLER_1_221 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_6_335 VPWR VGND sg13g2_decap_4
XFILLER_6_379 VPWR VGND sg13g2_decap_8
XFILLER_6_357 VPWR VGND sg13g2_fill_2
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_3_316 VPWR VGND sg13g2_decap_8
XFILLER_6_176 VPWR VGND sg13g2_decap_8
X_087_ S4END[1] net78 VPWR VGND sg13g2_buf_1
XFILLER_0_308 VPWR VGND sg13g2_decap_8
X_010_ FrameData[9] net32 VPWR VGND sg13g2_buf_1
XFILLER_3_168 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_fill_1
XFILLER_8_238 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_444 VPWR VGND sg13g2_decap_8
XFILLER_4_230 VPWR VGND sg13g2_decap_8
XFILLER_4_263 VPWR VGND sg13g2_decap_8
XFILLER_1_200 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_6_314 VPWR VGND sg13g2_decap_8
XFILLER_5_380 VPWR VGND sg13g2_decap_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_6_155 VPWR VGND sg13g2_decap_8
XFILLER_6_122 VPWR VGND sg13g2_decap_8
X_086_ S4END[2] net77 VPWR VGND sg13g2_buf_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_2_394 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
X_069_ S2END[3] net69 VPWR VGND sg13g2_buf_1
XFILLER_9_70 VPWR VGND sg13g2_decap_8
XFILLER_8_217 VPWR VGND sg13g2_decap_8
XFILLER_4_423 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_7_294 VPWR VGND sg13g2_decap_8
XFILLER_1_437 VPWR VGND sg13g2_decap_8
XFILLER_1_256 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_decap_8
Xoutput90 net90 NN4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_1_278 VPWR VGND sg13g2_fill_1
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_6_101 VPWR VGND sg13g2_decap_8
XFILLER_6_134 VPWR VGND sg13g2_decap_8
X_085_ S4END[3] net76 VPWR VGND sg13g2_buf_1
XFILLER_2_373 VPWR VGND sg13g2_decap_8
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_7_443 VPWR VGND sg13g2_decap_8
X_068_ S2END[4] net68 VPWR VGND sg13g2_buf_1
XS_term_single_106 VPWR VGND Co sg13g2_tielo
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_7_273 VPWR VGND sg13g2_decap_8
XFILLER_1_416 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_6_94 VPWR VGND sg13g2_decap_8
XFILLER_6_72 VPWR VGND sg13g2_fill_2
XFILLER_1_235 VPWR VGND sg13g2_decap_8
Xoutput1 net1 FrameData_O[0] VPWR VGND sg13g2_buf_1
Xoutput91 net91 NN4BEG[11] VPWR VGND sg13g2_buf_1
Xoutput80 net80 N4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_3_84 VPWR VGND sg13g2_decap_8
XFILLER_2_330 VPWR VGND sg13g2_decap_8
XFILLER_2_352 VPWR VGND sg13g2_decap_8
X_084_ S4END[4] net75 VPWR VGND sg13g2_buf_1
XFILLER_7_422 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
X_067_ S2END[5] net67 VPWR VGND sg13g2_buf_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_2_182 VPWR VGND sg13g2_fill_2
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_4_244 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_decap_8
XFILLER_1_214 VPWR VGND sg13g2_decap_8
Xoutput92 net92 NN4BEG[12] VPWR VGND sg13g2_buf_1
Xoutput81 net81 N4BEG[2] VPWR VGND sg13g2_buf_1
Xoutput70 net70 N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_0_280 VPWR VGND sg13g2_decap_8
Xoutput2 net2 FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_6_328 VPWR VGND sg13g2_decap_8
XFILLER_9_199 VPWR VGND sg13g2_decap_8
XFILLER_5_394 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
XFILLER_3_309 VPWR VGND sg13g2_decap_8
X_083_ S4END[5] net74 VPWR VGND sg13g2_buf_1
XFILLER_6_169 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_9_84 VPWR VGND sg13g2_decap_8
XFILLER_7_401 VPWR VGND sg13g2_decap_8
X_066_ S2END[6] net66 VPWR VGND sg13g2_buf_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_2_161 VPWR VGND sg13g2_decap_8
XFILLER_4_437 VPWR VGND sg13g2_decap_8
XFILLER_7_253 VPWR VGND sg13g2_fill_2
X_049_ FrameStrobe[16] net40 VPWR VGND sg13g2_buf_1
XFILLER_4_223 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_fill_1
XFILLER_6_63 VPWR VGND sg13g2_fill_1
XANTENNA_1 VPWR VGND FrameData[16] sg13g2_antennanp
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_9_359 VPWR VGND sg13g2_fill_1
Xoutput93 net93 NN4BEG[13] VPWR VGND sg13g2_buf_1
Xoutput82 net82 N4BEG[3] VPWR VGND sg13g2_buf_1
Xoutput71 net71 N2BEGb[6] VPWR VGND sg13g2_buf_1
Xoutput60 net60 N2BEG[3] VPWR VGND sg13g2_buf_1
Xoutput3 net3 FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_8_392 VPWR VGND sg13g2_decap_8
XFILLER_6_307 VPWR VGND sg13g2_decap_8
XFILLER_5_373 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_6_148 VPWR VGND sg13g2_decap_8
XFILLER_6_115 VPWR VGND sg13g2_decap_8
X_082_ S4END[6] net88 VPWR VGND sg13g2_buf_1
XFILLER_2_387 VPWR VGND sg13g2_decap_8
XFILLER_5_170 VPWR VGND sg13g2_decap_4
X_065_ S2END[7] net65 VPWR VGND sg13g2_buf_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_140 VPWR VGND sg13g2_decap_8
XFILLER_2_184 VPWR VGND sg13g2_fill_1
XFILLER_9_63 VPWR VGND sg13g2_decap_8
XFILLER_7_232 VPWR VGND sg13g2_decap_8
XFILLER_4_416 VPWR VGND sg13g2_decap_8
XFILLER_7_287 VPWR VGND sg13g2_decap_8
X_048_ FrameStrobe[15] net39 VPWR VGND sg13g2_buf_1
XFILLER_4_202 VPWR VGND sg13g2_decap_8
XANTENNA_2 VPWR VGND FrameData[21] sg13g2_antennanp
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XFILLER_1_249 VPWR VGND sg13g2_decap_8
Xoutput50 net50 FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_9_305 VPWR VGND sg13g2_decap_8
Xoutput94 net94 NN4BEG[14] VPWR VGND sg13g2_buf_1
Xoutput83 net83 N4BEG[4] VPWR VGND sg13g2_buf_1
Xoutput72 net72 N2BEGb[7] VPWR VGND sg13g2_buf_1
Xoutput61 net61 N2BEG[4] VPWR VGND sg13g2_buf_1
Xoutput4 net4 FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_9_102 VPWR VGND sg13g2_fill_1
XFILLER_5_352 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
XFILLER_2_300 VPWR VGND sg13g2_decap_8
X_081_ S4END[7] net87 VPWR VGND sg13g2_buf_1
XFILLER_2_344 VPWR VGND sg13g2_fill_2
XFILLER_2_366 VPWR VGND sg13g2_decap_8
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_7_436 VPWR VGND sg13g2_decap_8
X_064_ S2MID[0] net64 VPWR VGND sg13g2_buf_1
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_decap_8
XFILLER_7_211 VPWR VGND sg13g2_decap_8
XFILLER_3_450 VPWR VGND sg13g2_fill_1
X_047_ FrameStrobe[14] net38 VPWR VGND sg13g2_buf_1
XFILLER_1_409 VPWR VGND sg13g2_decap_8
XANTENNA_3 VPWR VGND FrameData[24] sg13g2_antennanp
XFILLER_6_87 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_4_258 VPWR VGND sg13g2_fill_1
XFILLER_1_228 VPWR VGND sg13g2_decap_8
Xoutput40 net40 FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
XFILLER_9_339 VPWR VGND sg13g2_fill_1
Xoutput51 net51 FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
Xoutput95 net95 NN4BEG[15] VPWR VGND sg13g2_buf_1
Xoutput84 net84 N4BEG[5] VPWR VGND sg13g2_buf_1
Xoutput73 net73 N4BEG[0] VPWR VGND sg13g2_buf_1
Xoutput62 net62 N2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_0_294 VPWR VGND sg13g2_decap_8
Xoutput5 net5 FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_3_77 VPWR VGND sg13g2_decap_8
X_080_ S4END[8] net86 VPWR VGND sg13g2_buf_1
XFILLER_2_323 VPWR VGND sg13g2_decap_8
XFILLER_7_415 VPWR VGND sg13g2_decap_8
X_063_ S2MID[1] net63 VPWR VGND sg13g2_buf_1
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_2_197 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_9_98 VPWR VGND sg13g2_decap_4
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
X_046_ FrameStrobe[13] net37 VPWR VGND sg13g2_buf_1
XFILLER_4_237 VPWR VGND sg13g2_decap_8
XANTENNA_4 VPWR VGND FrameData[25] sg13g2_antennanp
X_029_ FrameData[28] net21 VPWR VGND sg13g2_buf_1
XFILLER_3_281 VPWR VGND sg13g2_decap_8
Xoutput41 net41 FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
Xoutput52 net52 FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
Xoutput6 net6 FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_1_207 VPWR VGND sg13g2_decap_8
Xoutput30 net30 FrameData_O[7] VPWR VGND sg13g2_buf_1
Xoutput96 net96 NN4BEG[1] VPWR VGND sg13g2_buf_1
Xoutput74 net74 N4BEG[10] VPWR VGND sg13g2_buf_1
Xoutput85 net85 N4BEG[6] VPWR VGND sg13g2_buf_1
Xoutput63 net63 N2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_0_273 VPWR VGND sg13g2_decap_8
.ends

