module S_CPU_IF (Co,
    I_top0,
    I_top1,
    I_top10,
    I_top11,
    I_top12,
    I_top13,
    I_top14,
    I_top15,
    I_top2,
    I_top3,
    I_top4,
    I_top5,
    I_top6,
    I_top7,
    I_top8,
    I_top9,
    O_top0,
    O_top1,
    O_top10,
    O_top11,
    O_top12,
    O_top13,
    O_top14,
    O_top15,
    O_top2,
    O_top3,
    O_top4,
    O_top5,
    O_top6,
    O_top7,
    O_top8,
    O_top9,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output Co;
 output I_top0;
 output I_top1;
 output I_top10;
 output I_top11;
 output I_top12;
 output I_top13;
 output I_top14;
 output I_top15;
 output I_top2;
 output I_top3;
 output I_top4;
 output I_top5;
 output I_top6;
 output I_top7;
 output I_top8;
 output I_top9;
 input O_top0;
 input O_top1;
 input O_top10;
 input O_top11;
 input O_top12;
 input O_top13;
 input O_top14;
 input O_top15;
 input O_top2;
 input O_top3;
 input O_top4;
 input O_top5;
 input O_top6;
 input O_top7;
 input O_top8;
 input O_top9;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N1BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG4 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG5 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG6 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEG7 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb4 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb5 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb6 ;
 wire \Inst_S_CPU_IF_switch_matrix.N2BEGb7 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG10 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG11 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG12 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG13 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG14 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG15 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG4 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG5 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG6 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG7 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG8 ;
 wire \Inst_S_CPU_IF_switch_matrix.N4BEG9 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG0 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG1 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG10 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG11 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG12 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG13 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG14 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG15 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG2 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG3 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG4 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG5 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG6 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG7 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG8 ;
 wire \Inst_S_CPU_IF_switch_matrix.NN4BEG9 ;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net237;

 sg13g2_mux4_1 _000_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .A0(net67),
    .A1(net83),
    .A2(net90),
    .A3(net106),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .X(net175));
 sg13g2_mux4_1 _001_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .A0(net66),
    .A1(net82),
    .A2(net89),
    .A3(net105),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .X(net174));
 sg13g2_mux4_1 _002_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .A0(net65),
    .A1(net81),
    .A2(net88),
    .A3(net104),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .X(net173));
 sg13g2_mux4_1 _003_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .A0(net64),
    .A1(net80),
    .A2(net87),
    .A3(net103),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .X(net172));
 sg13g2_mux4_1 _004_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(net67),
    .A1(net75),
    .A2(net86),
    .A3(net102),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q ),
    .X(net171));
 sg13g2_mux4_1 _005_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(net66),
    .A1(net74),
    .A2(net85),
    .A3(net101),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q ),
    .X(net170));
 sg13g2_mux4_1 _006_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(net65),
    .A1(net73),
    .A2(net99),
    .A3(net115),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q ),
    .X(net183));
 sg13g2_mux4_1 _007_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(net64),
    .A1(net72),
    .A2(net98),
    .A3(net114),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q ),
    .X(net182));
 sg13g2_mux4_1 _008_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q ),
    .A0(net67),
    .A1(net71),
    .A2(net97),
    .A3(net113),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q ),
    .X(net181));
 sg13g2_mux4_1 _009_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(net66),
    .A1(net70),
    .A2(net96),
    .A3(net112),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q ),
    .X(net180));
 sg13g2_mux4_1 _010_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(net65),
    .A1(net69),
    .A2(net95),
    .A3(net111),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q ),
    .X(net179));
 sg13g2_mux4_1 _011_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(net64),
    .A1(net68),
    .A2(net94),
    .A3(net110),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q ),
    .X(net178));
 sg13g2_mux4_1 _012_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(net67),
    .A1(net79),
    .A2(net93),
    .A3(net109),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q ),
    .X(net177));
 sg13g2_mux4_1 _013_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(net66),
    .A1(net78),
    .A2(net92),
    .A3(net108),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q ),
    .X(net176));
 sg13g2_mux4_1 _014_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(net65),
    .A1(net77),
    .A2(net91),
    .A3(net107),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q ),
    .X(net169));
 sg13g2_mux4_1 _015_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(net64),
    .A1(net76),
    .A2(net84),
    .A3(net100),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q ),
    .X(net168));
 sg13g2_mux2_1 _016_ (.A0(net100),
    .A1(net33),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG15 ));
 sg13g2_mux2_1 _017_ (.A0(net107),
    .A1(net34),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG14 ));
 sg13g2_mux2_1 _018_ (.A0(net108),
    .A1(net41),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG13 ));
 sg13g2_mux2_1 _019_ (.A0(net109),
    .A1(net42),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG12 ));
 sg13g2_mux2_1 _020_ (.A0(net110),
    .A1(net43),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG11 ));
 sg13g2_mux2_1 _021_ (.A0(net111),
    .A1(net59),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG10 ));
 sg13g2_mux2_1 _022_ (.A0(net112),
    .A1(net60),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG9 ));
 sg13g2_mux2_1 _023_ (.A0(net113),
    .A1(net61),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG8 ));
 sg13g2_mux2_1 _024_ (.A0(net114),
    .A1(net62),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG7 ));
 sg13g2_mux2_1 _025_ (.A0(net115),
    .A1(net63),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG6 ));
 sg13g2_mux2_1 _026_ (.A0(net101),
    .A1(net35),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG5 ));
 sg13g2_mux2_1 _027_ (.A0(net102),
    .A1(net36),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG4 ));
 sg13g2_mux2_1 _028_ (.A0(net103),
    .A1(net37),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG3 ));
 sg13g2_mux2_1 _029_ (.A0(net104),
    .A1(net38),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG2 ));
 sg13g2_mux2_1 _030_ (.A0(net105),
    .A1(net39),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG1 ));
 sg13g2_mux2_1 _031_ (.A0(net106),
    .A1(net40),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.NN4BEG0 ));
 sg13g2_mux2_1 _032_ (.A0(net84),
    .A1(net33),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG15 ));
 sg13g2_mux2_1 _033_ (.A0(net91),
    .A1(net34),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG14 ));
 sg13g2_mux2_1 _034_ (.A0(net92),
    .A1(net41),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG13 ));
 sg13g2_mux2_1 _035_ (.A0(net93),
    .A1(net42),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG12 ));
 sg13g2_mux2_1 _036_ (.A0(net94),
    .A1(net43),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG11 ));
 sg13g2_mux2_1 _037_ (.A0(net95),
    .A1(net59),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG10 ));
 sg13g2_mux2_1 _038_ (.A0(net96),
    .A1(net60),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG9 ));
 sg13g2_mux2_1 _039_ (.A0(net97),
    .A1(net61),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG8 ));
 sg13g2_mux2_1 _040_ (.A0(net98),
    .A1(net62),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG7 ));
 sg13g2_mux2_1 _041_ (.A0(net99),
    .A1(net63),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG6 ));
 sg13g2_mux2_1 _042_ (.A0(net85),
    .A1(net35),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG5 ));
 sg13g2_mux2_1 _043_ (.A0(net86),
    .A1(net36),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG4 ));
 sg13g2_mux2_1 _044_ (.A0(net87),
    .A1(net37),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG3 ));
 sg13g2_mux2_1 _045_ (.A0(net88),
    .A1(net38),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG2 ));
 sg13g2_mux2_1 _046_ (.A0(net89),
    .A1(net39),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG1 ));
 sg13g2_mux2_1 _047_ (.A0(net90),
    .A1(net40),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N4BEG0 ));
 sg13g2_mux2_1 _048_ (.A0(net68),
    .A1(net62),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb7 ));
 sg13g2_mux2_1 _049_ (.A0(net69),
    .A1(net63),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb6 ));
 sg13g2_mux2_1 _050_ (.A0(net70),
    .A1(net35),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb5 ));
 sg13g2_mux2_1 _051_ (.A0(net71),
    .A1(net36),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb4 ));
 sg13g2_mux2_1 _052_ (.A0(net72),
    .A1(net37),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb3 ));
 sg13g2_mux2_1 _053_ (.A0(net73),
    .A1(net38),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb2 ));
 sg13g2_mux2_1 _054_ (.A0(net74),
    .A1(net39),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb1 ));
 sg13g2_mux2_1 _055_ (.A0(net75),
    .A1(net40),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEGb0 ));
 sg13g2_mux2_1 _056_ (.A0(net76),
    .A1(net33),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG7 ));
 sg13g2_mux2_1 _057_ (.A0(net77),
    .A1(net34),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG6 ));
 sg13g2_mux2_1 _058_ (.A0(net78),
    .A1(net41),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG5 ));
 sg13g2_mux2_1 _059_ (.A0(net79),
    .A1(net42),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG4 ));
 sg13g2_mux2_1 _060_ (.A0(net80),
    .A1(net43),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG3 ));
 sg13g2_mux2_1 _061_ (.A0(net81),
    .A1(net59),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG2 ));
 sg13g2_mux2_1 _062_ (.A0(net82),
    .A1(net60),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG1 ));
 sg13g2_mux2_1 _063_ (.A0(net83),
    .A1(net61),
    .S(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N2BEG0 ));
 sg13g2_mux4_1 _064_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(net64),
    .A1(net33),
    .A2(net43),
    .A3(net37),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _065_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net65),
    .A1(net34),
    .A2(net59),
    .A3(net38),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG2 ));
 sg13g2_mux4_1 _066_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(net66),
    .A1(net41),
    .A2(net60),
    .A3(net39),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG1 ));
 sg13g2_mux4_1 _067_ (.S0(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(net67),
    .A1(net42),
    .A2(net61),
    .A3(net40),
    .S1(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_S_CPU_IF_switch_matrix.N1BEG0 ));
 sg13g2_dlhq_1 _068_ (.D(net31),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _069_ (.D(net32),
    .GATE(net46),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _070_ (.D(net2),
    .GATE(net47),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _071_ (.D(net3),
    .GATE(net46),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _072_ (.D(net4),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _073_ (.D(net5),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _074_ (.D(net6),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _075_ (.D(net7),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _076_ (.D(net8),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _077_ (.D(net9),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _078_ (.D(net10),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _079_ (.D(net11),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _080_ (.D(net13),
    .GATE(net45),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _081_ (.D(net14),
    .GATE(net46),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _082_ (.D(net15),
    .GATE(net46),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _083_ (.D(net16),
    .GATE(net46),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _084_ (.D(net17),
    .GATE(net47),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _085_ (.D(net18),
    .GATE(net47),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _086_ (.D(net19),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _087_ (.D(net20),
    .GATE(net44),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _088_ (.D(net21),
    .GATE(net47),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _089_ (.D(net22),
    .GATE(net47),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _090_ (.D(net24),
    .GATE(net47),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _091_ (.D(net25),
    .GATE(net46),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _092_ (.D(net1),
    .GATE(net52),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _093_ (.D(net12),
    .GATE(net52),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _094_ (.D(net23),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _095_ (.D(net26),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _096_ (.D(net27),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _097_ (.D(net28),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _098_ (.D(net29),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _099_ (.D(net30),
    .GATE(net50),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _100_ (.D(net31),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _101_ (.D(net32),
    .GATE(net53),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _102_ (.D(net2),
    .GATE(net53),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _103_ (.D(net3),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _104_ (.D(net4),
    .GATE(net50),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _105_ (.D(net5),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _106_ (.D(net6),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _107_ (.D(net7),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _108_ (.D(net8),
    .GATE(net52),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _109_ (.D(net9),
    .GATE(net52),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _110_ (.D(net10),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _111_ (.D(net11),
    .GATE(net48),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _112_ (.D(net13),
    .GATE(net52),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _113_ (.D(net14),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _114_ (.D(net15),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _115_ (.D(net16),
    .GATE(net50),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _116_ (.D(net17),
    .GATE(net51),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _117_ (.D(net18),
    .GATE(net50),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _118_ (.D(net19),
    .GATE(net50),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _119_ (.D(net20),
    .GATE(net49),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _120_ (.D(net21),
    .GATE(net50),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _121_ (.D(net22),
    .GATE(net49),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _122_ (.D(net24),
    .GATE(net49),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _123_ (.D(net25),
    .GATE(net49),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _124_ (.D(net1),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _125_ (.D(net12),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _126_ (.D(net23),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _127_ (.D(net26),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _128_ (.D(net27),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _129_ (.D(net28),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _130_ (.D(net29),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _131_ (.D(net30),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _132_ (.D(net31),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _133_ (.D(net32),
    .GATE(net55),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _134_ (.D(net2),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _135_ (.D(net3),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _136_ (.D(net4),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _137_ (.D(net5),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _138_ (.D(net6),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _139_ (.D(net7),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _140_ (.D(net8),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _141_ (.D(net9),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _142_ (.D(net10),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _143_ (.D(net11),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _144_ (.D(net13),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _145_ (.D(net14),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _146_ (.D(net15),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _147_ (.D(net16),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _148_ (.D(net17),
    .GATE(net54),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _149_ (.D(net18),
    .GATE(net58),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _150_ (.D(net19),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _151_ (.D(net20),
    .GATE(net57),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _152_ (.D(net21),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _153_ (.D(net22),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _154_ (.D(net24),
    .GATE(net58),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _155_ (.D(net25),
    .GATE(net56),
    .Q(\Inst_S_CPU_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_antennanp ANTENNA_1 (.A(net121));
 sg13g2_buf_1 _157_ (.A(net1),
    .X(net116));
 sg13g2_buf_1 _158_ (.A(net12),
    .X(net127));
 sg13g2_buf_1 _159_ (.A(net23),
    .X(net138));
 sg13g2_buf_1 _160_ (.A(net26),
    .X(net141));
 sg13g2_buf_1 _161_ (.A(net27),
    .X(net142));
 sg13g2_buf_1 _162_ (.A(net28),
    .X(net143));
 sg13g2_buf_1 _163_ (.A(net29),
    .X(net144));
 sg13g2_buf_1 _164_ (.A(net30),
    .X(net145));
 sg13g2_buf_1 _165_ (.A(net31),
    .X(net146));
 sg13g2_buf_1 _166_ (.A(net32),
    .X(net147));
 sg13g2_buf_1 _167_ (.A(net2),
    .X(net117));
 sg13g2_buf_1 _168_ (.A(net3),
    .X(net118));
 sg13g2_buf_1 _169_ (.A(net4),
    .X(net119));
 sg13g2_buf_1 _170_ (.A(net5),
    .X(net120));
 sg13g2_buf_1 _171_ (.A(net6),
    .X(net121));
 sg13g2_buf_1 _172_ (.A(net7),
    .X(net122));
 sg13g2_buf_1 _173_ (.A(net8),
    .X(net123));
 sg13g2_buf_1 _174_ (.A(net9),
    .X(net124));
 sg13g2_buf_1 _175_ (.A(net10),
    .X(net125));
 sg13g2_buf_1 _176_ (.A(net11),
    .X(net126));
 sg13g2_buf_1 _177_ (.A(net13),
    .X(net128));
 sg13g2_buf_1 _178_ (.A(net14),
    .X(net129));
 sg13g2_buf_1 _179_ (.A(net15),
    .X(net130));
 sg13g2_buf_1 _180_ (.A(net16),
    .X(net131));
 sg13g2_buf_1 _181_ (.A(net17),
    .X(net132));
 sg13g2_buf_1 _182_ (.A(net18),
    .X(net133));
 sg13g2_buf_1 _183_ (.A(net19),
    .X(net134));
 sg13g2_buf_1 _184_ (.A(net20),
    .X(net135));
 sg13g2_buf_1 _185_ (.A(net21),
    .X(net136));
 sg13g2_buf_1 _186_ (.A(net22),
    .X(net137));
 sg13g2_buf_1 _187_ (.A(net24),
    .X(net139));
 sg13g2_buf_1 _188_ (.A(net25),
    .X(net140));
 sg13g2_buf_1 _189_ (.A(net56),
    .X(net148));
 sg13g2_buf_1 _190_ (.A(net51),
    .X(net159));
 sg13g2_buf_1 _191_ (.A(net47),
    .X(net160));
 sg13g2_buf_1 _192_ (.A(FrameStrobe[3]),
    .X(net161));
 sg13g2_buf_1 _193_ (.A(FrameStrobe[4]),
    .X(net162));
 sg13g2_buf_1 _194_ (.A(FrameStrobe[5]),
    .X(net163));
 sg13g2_buf_1 _195_ (.A(FrameStrobe[6]),
    .X(net164));
 sg13g2_buf_1 _196_ (.A(FrameStrobe[7]),
    .X(net165));
 sg13g2_buf_1 _197_ (.A(FrameStrobe[8]),
    .X(net166));
 sg13g2_buf_1 _198_ (.A(FrameStrobe[9]),
    .X(net167));
 sg13g2_buf_1 _199_ (.A(FrameStrobe[10]),
    .X(net149));
 sg13g2_buf_1 _200_ (.A(FrameStrobe[11]),
    .X(net150));
 sg13g2_buf_1 _201_ (.A(FrameStrobe[12]),
    .X(net151));
 sg13g2_buf_1 _202_ (.A(FrameStrobe[13]),
    .X(net152));
 sg13g2_buf_1 _203_ (.A(FrameStrobe[14]),
    .X(net153));
 sg13g2_buf_1 _204_ (.A(FrameStrobe[15]),
    .X(net154));
 sg13g2_buf_1 _205_ (.A(FrameStrobe[16]),
    .X(net155));
 sg13g2_buf_1 _206_ (.A(FrameStrobe[17]),
    .X(net156));
 sg13g2_buf_1 _207_ (.A(FrameStrobe[18]),
    .X(net157));
 sg13g2_buf_1 _208_ (.A(FrameStrobe[19]),
    .X(net158));
 sg13g2_buf_1 _209_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG0 ),
    .X(net184));
 sg13g2_buf_1 _210_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG1 ),
    .X(net185));
 sg13g2_buf_1 _211_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG2 ),
    .X(net186));
 sg13g2_buf_1 _212_ (.A(\Inst_S_CPU_IF_switch_matrix.N1BEG3 ),
    .X(net187));
 sg13g2_buf_1 _213_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG0 ),
    .X(net188));
 sg13g2_buf_1 _214_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG1 ),
    .X(net189));
 sg13g2_buf_1 _215_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG2 ),
    .X(net190));
 sg13g2_buf_1 _216_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG3 ),
    .X(net191));
 sg13g2_buf_1 _217_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG4 ),
    .X(net192));
 sg13g2_buf_1 _218_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG5 ),
    .X(net193));
 sg13g2_buf_1 _219_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG6 ),
    .X(net194));
 sg13g2_buf_1 _220_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEG7 ),
    .X(net195));
 sg13g2_buf_1 _221_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb0 ),
    .X(net196));
 sg13g2_buf_1 _222_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb1 ),
    .X(net197));
 sg13g2_buf_1 _223_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb2 ),
    .X(net198));
 sg13g2_buf_1 _224_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb3 ),
    .X(net199));
 sg13g2_buf_1 _225_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb4 ),
    .X(net200));
 sg13g2_buf_1 _226_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb5 ),
    .X(net201));
 sg13g2_buf_1 _227_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb6 ),
    .X(net202));
 sg13g2_buf_1 _228_ (.A(\Inst_S_CPU_IF_switch_matrix.N2BEGb7 ),
    .X(net203));
 sg13g2_buf_1 _229_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG0 ),
    .X(net204));
 sg13g2_buf_1 _230_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG1 ),
    .X(net211));
 sg13g2_buf_1 _231_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG2 ),
    .X(net212));
 sg13g2_buf_1 _232_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG3 ),
    .X(net213));
 sg13g2_buf_1 _233_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG4 ),
    .X(net214));
 sg13g2_buf_1 _234_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG5 ),
    .X(net215));
 sg13g2_buf_1 _235_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG6 ),
    .X(net216));
 sg13g2_buf_1 _236_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG7 ),
    .X(net217));
 sg13g2_buf_1 _237_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG8 ),
    .X(net218));
 sg13g2_buf_1 _238_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG9 ),
    .X(net219));
 sg13g2_buf_1 _239_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG10 ),
    .X(net205));
 sg13g2_buf_1 _240_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG11 ),
    .X(net206));
 sg13g2_buf_1 _241_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG12 ),
    .X(net207));
 sg13g2_buf_1 _242_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG13 ),
    .X(net208));
 sg13g2_buf_1 _243_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG14 ),
    .X(net209));
 sg13g2_buf_1 _244_ (.A(\Inst_S_CPU_IF_switch_matrix.N4BEG15 ),
    .X(net210));
 sg13g2_buf_1 _245_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG0 ),
    .X(net220));
 sg13g2_buf_1 _246_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG1 ),
    .X(net227));
 sg13g2_buf_1 _247_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG2 ),
    .X(net228));
 sg13g2_buf_1 _248_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG3 ),
    .X(net229));
 sg13g2_buf_1 _249_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG4 ),
    .X(net230));
 sg13g2_buf_1 _250_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG5 ),
    .X(net231));
 sg13g2_buf_1 _251_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG6 ),
    .X(net232));
 sg13g2_buf_1 _252_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG7 ),
    .X(net233));
 sg13g2_buf_1 _253_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG8 ),
    .X(net234));
 sg13g2_buf_1 _254_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG9 ),
    .X(net235));
 sg13g2_buf_1 _255_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG10 ),
    .X(net221));
 sg13g2_buf_1 _256_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG11 ),
    .X(net222));
 sg13g2_buf_1 _257_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG12 ),
    .X(net223));
 sg13g2_buf_1 _258_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG13 ),
    .X(net224));
 sg13g2_buf_1 _259_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG14 ),
    .X(net225));
 sg13g2_buf_1 _260_ (.A(\Inst_S_CPU_IF_switch_matrix.NN4BEG15 ),
    .X(net226));
 sg13g2_buf_1 _261_ (.A(UserCLK),
    .X(net236));
 sg13g2_buf_1 fanout44 (.A(net46),
    .X(net44));
 sg13g2_buf_1 fanout45 (.A(net46),
    .X(net45));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_1 fanout47 (.A(FrameStrobe[2]),
    .X(net47));
 sg13g2_buf_1 fanout48 (.A(net50),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_1 fanout50 (.A(net53),
    .X(net50));
 sg13g2_buf_1 fanout51 (.A(net53),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(net53),
    .X(net52));
 sg13g2_buf_1 fanout53 (.A(FrameStrobe[1]),
    .X(net53));
 sg13g2_buf_1 fanout54 (.A(net58),
    .X(net54));
 sg13g2_buf_1 fanout55 (.A(net58),
    .X(net55));
 sg13g2_buf_1 fanout56 (.A(net57),
    .X(net56));
 sg13g2_buf_1 fanout57 (.A(net58),
    .X(net57));
 sg13g2_buf_1 fanout58 (.A(FrameStrobe[0]),
    .X(net58));
 sg13g2_buf_1 input1 (.A(FrameData[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(FrameData[10]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(FrameData[11]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(FrameData[12]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(FrameData[13]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(FrameData[14]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(FrameData[15]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(FrameData[16]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(FrameData[17]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(FrameData[18]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(FrameData[19]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(FrameData[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(FrameData[20]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(FrameData[21]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(FrameData[22]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(FrameData[23]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(FrameData[24]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(FrameData[25]),
    .X(net18));
 sg13g2_buf_1 input19 (.A(FrameData[26]),
    .X(net19));
 sg13g2_buf_1 input20 (.A(FrameData[27]),
    .X(net20));
 sg13g2_buf_1 input21 (.A(FrameData[28]),
    .X(net21));
 sg13g2_buf_1 input22 (.A(FrameData[29]),
    .X(net22));
 sg13g2_buf_1 input23 (.A(FrameData[2]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(FrameData[30]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(FrameData[31]),
    .X(net25));
 sg13g2_buf_1 input26 (.A(FrameData[3]),
    .X(net26));
 sg13g2_buf_1 input27 (.A(FrameData[4]),
    .X(net27));
 sg13g2_buf_1 input28 (.A(FrameData[5]),
    .X(net28));
 sg13g2_buf_1 input29 (.A(FrameData[6]),
    .X(net29));
 sg13g2_buf_1 input30 (.A(FrameData[7]),
    .X(net30));
 sg13g2_buf_1 input31 (.A(FrameData[8]),
    .X(net31));
 sg13g2_buf_1 input32 (.A(FrameData[9]),
    .X(net32));
 sg13g2_buf_1 input33 (.A(O_top0),
    .X(net33));
 sg13g2_buf_1 input34 (.A(O_top1),
    .X(net34));
 sg13g2_buf_1 input35 (.A(O_top10),
    .X(net35));
 sg13g2_buf_1 input36 (.A(O_top11),
    .X(net36));
 sg13g2_buf_1 input37 (.A(O_top12),
    .X(net37));
 sg13g2_buf_1 input38 (.A(O_top13),
    .X(net38));
 sg13g2_buf_1 input39 (.A(O_top14),
    .X(net39));
 sg13g2_buf_1 input40 (.A(O_top15),
    .X(net40));
 sg13g2_buf_1 input41 (.A(O_top2),
    .X(net41));
 sg13g2_buf_1 input42 (.A(O_top3),
    .X(net42));
 sg13g2_buf_1 input43 (.A(O_top4),
    .X(net43));
 sg13g2_buf_1 input44 (.A(O_top5),
    .X(net59));
 sg13g2_buf_1 input45 (.A(O_top6),
    .X(net60));
 sg13g2_buf_1 input46 (.A(O_top7),
    .X(net61));
 sg13g2_buf_1 input47 (.A(O_top8),
    .X(net62));
 sg13g2_buf_1 input48 (.A(O_top9),
    .X(net63));
 sg13g2_buf_1 input49 (.A(S1END[0]),
    .X(net64));
 sg13g2_buf_1 input50 (.A(S1END[1]),
    .X(net65));
 sg13g2_buf_1 input51 (.A(S1END[2]),
    .X(net66));
 sg13g2_buf_1 input52 (.A(S1END[3]),
    .X(net67));
 sg13g2_buf_1 input53 (.A(S2END[0]),
    .X(net68));
 sg13g2_buf_1 input54 (.A(S2END[1]),
    .X(net69));
 sg13g2_buf_1 input55 (.A(S2END[2]),
    .X(net70));
 sg13g2_buf_1 input56 (.A(S2END[3]),
    .X(net71));
 sg13g2_buf_1 input57 (.A(S2END[4]),
    .X(net72));
 sg13g2_buf_1 input58 (.A(S2END[5]),
    .X(net73));
 sg13g2_buf_1 input59 (.A(S2END[6]),
    .X(net74));
 sg13g2_buf_1 input60 (.A(S2END[7]),
    .X(net75));
 sg13g2_buf_1 input61 (.A(S2MID[0]),
    .X(net76));
 sg13g2_buf_1 input62 (.A(S2MID[1]),
    .X(net77));
 sg13g2_buf_1 input63 (.A(S2MID[2]),
    .X(net78));
 sg13g2_buf_1 input64 (.A(S2MID[3]),
    .X(net79));
 sg13g2_buf_1 input65 (.A(S2MID[4]),
    .X(net80));
 sg13g2_buf_1 input66 (.A(S2MID[5]),
    .X(net81));
 sg13g2_buf_1 input67 (.A(S2MID[6]),
    .X(net82));
 sg13g2_buf_1 input68 (.A(S2MID[7]),
    .X(net83));
 sg13g2_buf_1 input69 (.A(S4END[0]),
    .X(net84));
 sg13g2_buf_1 input70 (.A(S4END[10]),
    .X(net85));
 sg13g2_buf_1 input71 (.A(S4END[11]),
    .X(net86));
 sg13g2_buf_1 input72 (.A(S4END[12]),
    .X(net87));
 sg13g2_buf_1 input73 (.A(S4END[13]),
    .X(net88));
 sg13g2_buf_1 input74 (.A(S4END[14]),
    .X(net89));
 sg13g2_buf_1 input75 (.A(S4END[15]),
    .X(net90));
 sg13g2_buf_1 input76 (.A(S4END[1]),
    .X(net91));
 sg13g2_buf_1 input77 (.A(S4END[2]),
    .X(net92));
 sg13g2_buf_1 input78 (.A(S4END[3]),
    .X(net93));
 sg13g2_buf_1 input79 (.A(S4END[4]),
    .X(net94));
 sg13g2_buf_1 input80 (.A(S4END[5]),
    .X(net95));
 sg13g2_buf_1 input81 (.A(S4END[6]),
    .X(net96));
 sg13g2_buf_1 input82 (.A(S4END[7]),
    .X(net97));
 sg13g2_buf_1 input83 (.A(S4END[8]),
    .X(net98));
 sg13g2_buf_1 input84 (.A(S4END[9]),
    .X(net99));
 sg13g2_buf_1 input85 (.A(SS4END[0]),
    .X(net100));
 sg13g2_buf_1 input86 (.A(SS4END[10]),
    .X(net101));
 sg13g2_buf_1 input87 (.A(SS4END[11]),
    .X(net102));
 sg13g2_buf_1 input88 (.A(SS4END[12]),
    .X(net103));
 sg13g2_buf_1 input89 (.A(SS4END[13]),
    .X(net104));
 sg13g2_buf_1 input90 (.A(SS4END[14]),
    .X(net105));
 sg13g2_buf_1 input91 (.A(SS4END[15]),
    .X(net106));
 sg13g2_buf_1 input92 (.A(SS4END[1]),
    .X(net107));
 sg13g2_buf_1 input93 (.A(SS4END[2]),
    .X(net108));
 sg13g2_buf_1 input94 (.A(SS4END[3]),
    .X(net109));
 sg13g2_buf_1 input95 (.A(SS4END[4]),
    .X(net110));
 sg13g2_buf_1 input96 (.A(SS4END[5]),
    .X(net111));
 sg13g2_buf_1 input97 (.A(SS4END[6]),
    .X(net112));
 sg13g2_buf_1 input98 (.A(SS4END[7]),
    .X(net113));
 sg13g2_buf_1 input99 (.A(SS4END[8]),
    .X(net114));
 sg13g2_buf_1 input100 (.A(SS4END[9]),
    .X(net115));
 sg13g2_buf_1 output101 (.A(net116),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output102 (.A(net117),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output103 (.A(net118),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output104 (.A(net119),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output105 (.A(net120),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output106 (.A(net121),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output107 (.A(net122),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output108 (.A(net123),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output109 (.A(net124),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output110 (.A(net125),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output111 (.A(net126),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output112 (.A(net127),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output113 (.A(net128),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output114 (.A(net129),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output115 (.A(net130),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output116 (.A(net131),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output117 (.A(net132),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output118 (.A(net133),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output119 (.A(net134),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output120 (.A(net135),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output121 (.A(net136),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output122 (.A(net137),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output123 (.A(net138),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output124 (.A(net139),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output125 (.A(net140),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output126 (.A(net141),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output127 (.A(net142),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output128 (.A(net143),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output129 (.A(net144),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output130 (.A(net145),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output131 (.A(net146),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output132 (.A(net147),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output133 (.A(net148),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output134 (.A(net149),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output135 (.A(net150),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output136 (.A(net151),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output137 (.A(net152),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output138 (.A(net153),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output139 (.A(net154),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output140 (.A(net155),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output141 (.A(net156),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output142 (.A(net157),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output143 (.A(net158),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output144 (.A(net159),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output145 (.A(net160),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output146 (.A(net161),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output147 (.A(net162),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output148 (.A(net163),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output149 (.A(net164),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output150 (.A(net165),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output151 (.A(net166),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output152 (.A(net167),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output153 (.A(net168),
    .X(I_top0));
 sg13g2_buf_1 output154 (.A(net169),
    .X(I_top1));
 sg13g2_buf_1 output155 (.A(net170),
    .X(I_top10));
 sg13g2_buf_1 output156 (.A(net171),
    .X(I_top11));
 sg13g2_buf_1 output157 (.A(net172),
    .X(I_top12));
 sg13g2_buf_1 output158 (.A(net173),
    .X(I_top13));
 sg13g2_buf_1 output159 (.A(net174),
    .X(I_top14));
 sg13g2_buf_1 output160 (.A(net175),
    .X(I_top15));
 sg13g2_buf_1 output161 (.A(net176),
    .X(I_top2));
 sg13g2_buf_1 output162 (.A(net177),
    .X(I_top3));
 sg13g2_buf_1 output163 (.A(net178),
    .X(I_top4));
 sg13g2_buf_1 output164 (.A(net179),
    .X(I_top5));
 sg13g2_buf_1 output165 (.A(net180),
    .X(I_top6));
 sg13g2_buf_1 output166 (.A(net181),
    .X(I_top7));
 sg13g2_buf_1 output167 (.A(net182),
    .X(I_top8));
 sg13g2_buf_1 output168 (.A(net183),
    .X(I_top9));
 sg13g2_buf_1 output169 (.A(net184),
    .X(N1BEG[0]));
 sg13g2_buf_1 output170 (.A(net185),
    .X(N1BEG[1]));
 sg13g2_buf_1 output171 (.A(net186),
    .X(N1BEG[2]));
 sg13g2_buf_1 output172 (.A(net187),
    .X(N1BEG[3]));
 sg13g2_buf_1 output173 (.A(net188),
    .X(N2BEG[0]));
 sg13g2_buf_1 output174 (.A(net189),
    .X(N2BEG[1]));
 sg13g2_buf_1 output175 (.A(net190),
    .X(N2BEG[2]));
 sg13g2_buf_1 output176 (.A(net191),
    .X(N2BEG[3]));
 sg13g2_buf_1 output177 (.A(net192),
    .X(N2BEG[4]));
 sg13g2_buf_1 output178 (.A(net193),
    .X(N2BEG[5]));
 sg13g2_buf_1 output179 (.A(net194),
    .X(N2BEG[6]));
 sg13g2_buf_1 output180 (.A(net195),
    .X(N2BEG[7]));
 sg13g2_buf_1 output181 (.A(net196),
    .X(N2BEGb[0]));
 sg13g2_buf_1 output182 (.A(net197),
    .X(N2BEGb[1]));
 sg13g2_buf_1 output183 (.A(net198),
    .X(N2BEGb[2]));
 sg13g2_buf_1 output184 (.A(net199),
    .X(N2BEGb[3]));
 sg13g2_buf_1 output185 (.A(net200),
    .X(N2BEGb[4]));
 sg13g2_buf_1 output186 (.A(net201),
    .X(N2BEGb[5]));
 sg13g2_buf_1 output187 (.A(net202),
    .X(N2BEGb[6]));
 sg13g2_buf_1 output188 (.A(net203),
    .X(N2BEGb[7]));
 sg13g2_buf_1 output189 (.A(net204),
    .X(N4BEG[0]));
 sg13g2_buf_1 output190 (.A(net205),
    .X(N4BEG[10]));
 sg13g2_buf_1 output191 (.A(net206),
    .X(N4BEG[11]));
 sg13g2_buf_1 output192 (.A(net207),
    .X(N4BEG[12]));
 sg13g2_buf_1 output193 (.A(net208),
    .X(N4BEG[13]));
 sg13g2_buf_1 output194 (.A(net209),
    .X(N4BEG[14]));
 sg13g2_buf_1 output195 (.A(net210),
    .X(N4BEG[15]));
 sg13g2_buf_1 output196 (.A(net211),
    .X(N4BEG[1]));
 sg13g2_buf_1 output197 (.A(net212),
    .X(N4BEG[2]));
 sg13g2_buf_1 output198 (.A(net213),
    .X(N4BEG[3]));
 sg13g2_buf_1 output199 (.A(net214),
    .X(N4BEG[4]));
 sg13g2_buf_1 output200 (.A(net215),
    .X(N4BEG[5]));
 sg13g2_buf_1 output201 (.A(net216),
    .X(N4BEG[6]));
 sg13g2_buf_1 output202 (.A(net217),
    .X(N4BEG[7]));
 sg13g2_buf_1 output203 (.A(net218),
    .X(N4BEG[8]));
 sg13g2_buf_1 output204 (.A(net219),
    .X(N4BEG[9]));
 sg13g2_buf_1 output205 (.A(net220),
    .X(NN4BEG[0]));
 sg13g2_buf_1 output206 (.A(net221),
    .X(NN4BEG[10]));
 sg13g2_buf_1 output207 (.A(net222),
    .X(NN4BEG[11]));
 sg13g2_buf_1 output208 (.A(net223),
    .X(NN4BEG[12]));
 sg13g2_buf_1 output209 (.A(net224),
    .X(NN4BEG[13]));
 sg13g2_buf_1 output210 (.A(net225),
    .X(NN4BEG[14]));
 sg13g2_buf_1 output211 (.A(net226),
    .X(NN4BEG[15]));
 sg13g2_buf_1 output212 (.A(net227),
    .X(NN4BEG[1]));
 sg13g2_buf_1 output213 (.A(net228),
    .X(NN4BEG[2]));
 sg13g2_buf_1 output214 (.A(net229),
    .X(NN4BEG[3]));
 sg13g2_buf_1 output215 (.A(net230),
    .X(NN4BEG[4]));
 sg13g2_buf_1 output216 (.A(net231),
    .X(NN4BEG[5]));
 sg13g2_buf_1 output217 (.A(net232),
    .X(NN4BEG[6]));
 sg13g2_buf_1 output218 (.A(net233),
    .X(NN4BEG[7]));
 sg13g2_buf_1 output219 (.A(net234),
    .X(NN4BEG[8]));
 sg13g2_buf_1 output220 (.A(net235),
    .X(NN4BEG[9]));
 sg13g2_buf_1 output221 (.A(net236),
    .X(UserCLKo));
 sg13g2_tielo S_CPU_IF_222 (.L_LO(net237));
 sg13g2_antennanp ANTENNA_2 (.A(net125));
 sg13g2_antennanp ANTENNA_3 (.A(net130));
 sg13g2_antennanp ANTENNA_4 (.A(net134));
 sg13g2_antennanp ANTENNA_5 (.A(net135));
 sg13g2_antennanp ANTENNA_6 (.A(net138));
 sg13g2_antennanp ANTENNA_7 (.A(net144));
 sg13g2_antennanp ANTENNA_8 (.A(net121));
 sg13g2_antennanp ANTENNA_9 (.A(net125));
 sg13g2_antennanp ANTENNA_10 (.A(net130));
 sg13g2_antennanp ANTENNA_11 (.A(net134));
 sg13g2_antennanp ANTENNA_12 (.A(net135));
 sg13g2_antennanp ANTENNA_13 (.A(net138));
 sg13g2_antennanp ANTENNA_14 (.A(net144));
 sg13g2_antennanp ANTENNA_15 (.A(net121));
 sg13g2_antennanp ANTENNA_16 (.A(net125));
 sg13g2_antennanp ANTENNA_17 (.A(net130));
 sg13g2_antennanp ANTENNA_18 (.A(net134));
 sg13g2_antennanp ANTENNA_19 (.A(net135));
 sg13g2_antennanp ANTENNA_20 (.A(net138));
 sg13g2_antennanp ANTENNA_21 (.A(net144));
 sg13g2_antennanp ANTENNA_22 (.A(net121));
 sg13g2_antennanp ANTENNA_23 (.A(net125));
 sg13g2_antennanp ANTENNA_24 (.A(net130));
 sg13g2_antennanp ANTENNA_25 (.A(net134));
 sg13g2_antennanp ANTENNA_26 (.A(net135));
 sg13g2_antennanp ANTENNA_27 (.A(net138));
 sg13g2_antennanp ANTENNA_28 (.A(net144));
 sg13g2_antennanp ANTENNA_29 (.A(net121));
 sg13g2_antennanp ANTENNA_30 (.A(net125));
 sg13g2_antennanp ANTENNA_31 (.A(net130));
 sg13g2_antennanp ANTENNA_32 (.A(net134));
 sg13g2_antennanp ANTENNA_33 (.A(net135));
 sg13g2_antennanp ANTENNA_34 (.A(net138));
 sg13g2_antennanp ANTENNA_35 (.A(net144));
 sg13g2_antennanp ANTENNA_36 (.A(net121));
 sg13g2_antennanp ANTENNA_37 (.A(net125));
 sg13g2_antennanp ANTENNA_38 (.A(net130));
 sg13g2_antennanp ANTENNA_39 (.A(net134));
 sg13g2_antennanp ANTENNA_40 (.A(net135));
 sg13g2_antennanp ANTENNA_41 (.A(net138));
 sg13g2_antennanp ANTENNA_42 (.A(net144));
 sg13g2_antennanp ANTENNA_43 (.A(net121));
 sg13g2_antennanp ANTENNA_44 (.A(net125));
 sg13g2_antennanp ANTENNA_45 (.A(net130));
 sg13g2_antennanp ANTENNA_46 (.A(net134));
 sg13g2_antennanp ANTENNA_47 (.A(net135));
 sg13g2_antennanp ANTENNA_48 (.A(net138));
 sg13g2_antennanp ANTENNA_49 (.A(net144));
 sg13g2_antennanp ANTENNA_50 (.A(net121));
 sg13g2_antennanp ANTENNA_51 (.A(net125));
 sg13g2_antennanp ANTENNA_52 (.A(net130));
 sg13g2_antennanp ANTENNA_53 (.A(net134));
 sg13g2_antennanp ANTENNA_54 (.A(net135));
 sg13g2_antennanp ANTENNA_55 (.A(net138));
 sg13g2_antennanp ANTENNA_56 (.A(net144));
 sg13g2_antennanp ANTENNA_57 (.A(net121));
 sg13g2_antennanp ANTENNA_58 (.A(net125));
 sg13g2_antennanp ANTENNA_59 (.A(net130));
 sg13g2_antennanp ANTENNA_60 (.A(net134));
 sg13g2_antennanp ANTENNA_61 (.A(net135));
 sg13g2_antennanp ANTENNA_62 (.A(net138));
 sg13g2_antennanp ANTENNA_63 (.A(net144));
 sg13g2_antennanp ANTENNA_64 (.A(net121));
 sg13g2_antennanp ANTENNA_65 (.A(net125));
 sg13g2_antennanp ANTENNA_66 (.A(net130));
 sg13g2_antennanp ANTENNA_67 (.A(net134));
 sg13g2_antennanp ANTENNA_68 (.A(net135));
 sg13g2_antennanp ANTENNA_69 (.A(net138));
 sg13g2_antennanp ANTENNA_70 (.A(net144));
 sg13g2_decap_4 FILLER_0_16 ();
 sg13g2_fill_1 FILLER_0_20 ();
 sg13g2_decap_4 FILLER_0_25 ();
 sg13g2_fill_2 FILLER_0_33 ();
 sg13g2_fill_2 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_145 ();
 sg13g2_fill_1 FILLER_0_147 ();
 sg13g2_fill_1 FILLER_0_193 ();
 sg13g2_fill_2 FILLER_0_219 ();
 sg13g2_fill_2 FILLER_0_225 ();
 sg13g2_fill_1 FILLER_0_227 ();
 sg13g2_fill_2 FILLER_0_275 ();
 sg13g2_fill_1 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_4 FILLER_0_309 ();
 sg13g2_fill_1 FILLER_0_313 ();
 sg13g2_fill_1 FILLER_0_318 ();
 sg13g2_decap_4 FILLER_0_323 ();
 sg13g2_fill_2 FILLER_0_327 ();
 sg13g2_decap_4 FILLER_0_346 ();
 sg13g2_fill_1 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_fill_1 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_4 FILLER_0_388 ();
 sg13g2_fill_2 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_fill_1 FILLER_0_405 ();
 sg13g2_fill_2 FILLER_0_413 ();
 sg13g2_fill_1 FILLER_0_451 ();
 sg13g2_decap_8 FILLER_1_12 ();
 sg13g2_decap_8 FILLER_1_19 ();
 sg13g2_decap_8 FILLER_1_26 ();
 sg13g2_decap_8 FILLER_1_33 ();
 sg13g2_fill_2 FILLER_1_40 ();
 sg13g2_fill_1 FILLER_1_42 ();
 sg13g2_fill_2 FILLER_1_64 ();
 sg13g2_fill_2 FILLER_1_83 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_207 ();
 sg13g2_fill_2 FILLER_1_225 ();
 sg13g2_fill_1 FILLER_1_258 ();
 sg13g2_fill_1 FILLER_1_280 ();
 sg13g2_decap_4 FILLER_1_344 ();
 sg13g2_fill_2 FILLER_1_348 ();
 sg13g2_fill_1 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_decap_4 FILLER_1_407 ();
 sg13g2_fill_1 FILLER_1_411 ();
 sg13g2_fill_2 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_2_8 ();
 sg13g2_decap_8 FILLER_2_15 ();
 sg13g2_decap_4 FILLER_2_22 ();
 sg13g2_fill_2 FILLER_2_26 ();
 sg13g2_decap_8 FILLER_2_45 ();
 sg13g2_decap_8 FILLER_2_52 ();
 sg13g2_decap_4 FILLER_2_59 ();
 sg13g2_fill_1 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_82 ();
 sg13g2_decap_8 FILLER_2_89 ();
 sg13g2_decap_8 FILLER_2_96 ();
 sg13g2_fill_2 FILLER_2_103 ();
 sg13g2_fill_1 FILLER_2_105 ();
 sg13g2_fill_2 FILLER_2_137 ();
 sg13g2_fill_1 FILLER_2_139 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_4 FILLER_2_231 ();
 sg13g2_fill_1 FILLER_2_235 ();
 sg13g2_fill_2 FILLER_2_250 ();
 sg13g2_fill_1 FILLER_2_252 ();
 sg13g2_decap_4 FILLER_2_257 ();
 sg13g2_fill_1 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_286 ();
 sg13g2_fill_1 FILLER_2_297 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_304 ();
 sg13g2_decap_4 FILLER_2_322 ();
 sg13g2_fill_2 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_fill_1 FILLER_2_363 ();
 sg13g2_fill_2 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_404 ();
 sg13g2_decap_8 FILLER_2_411 ();
 sg13g2_fill_1 FILLER_2_442 ();
 sg13g2_fill_1 FILLER_2_454 ();
 sg13g2_decap_8 FILLER_3_8 ();
 sg13g2_decap_8 FILLER_3_15 ();
 sg13g2_decap_8 FILLER_3_22 ();
 sg13g2_fill_1 FILLER_3_29 ();
 sg13g2_fill_2 FILLER_3_34 ();
 sg13g2_fill_1 FILLER_3_36 ();
 sg13g2_fill_2 FILLER_3_58 ();
 sg13g2_fill_2 FILLER_3_99 ();
 sg13g2_fill_1 FILLER_3_101 ();
 sg13g2_decap_8 FILLER_3_106 ();
 sg13g2_fill_2 FILLER_3_113 ();
 sg13g2_fill_1 FILLER_3_132 ();
 sg13g2_decap_4 FILLER_3_137 ();
 sg13g2_fill_2 FILLER_3_141 ();
 sg13g2_decap_8 FILLER_3_153 ();
 sg13g2_fill_2 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_222 ();
 sg13g2_decap_4 FILLER_3_229 ();
 sg13g2_fill_2 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_273 ();
 sg13g2_fill_1 FILLER_3_296 ();
 sg13g2_decap_8 FILLER_3_314 ();
 sg13g2_decap_4 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_fill_2 FILLER_3_373 ();
 sg13g2_fill_1 FILLER_3_439 ();
 sg13g2_fill_2 FILLER_3_446 ();
 sg13g2_decap_8 FILLER_4_8 ();
 sg13g2_decap_8 FILLER_4_15 ();
 sg13g2_decap_8 FILLER_4_22 ();
 sg13g2_decap_8 FILLER_4_29 ();
 sg13g2_decap_8 FILLER_4_36 ();
 sg13g2_fill_2 FILLER_4_63 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_fill_2 FILLER_4_104 ();
 sg13g2_fill_1 FILLER_4_106 ();
 sg13g2_fill_1 FILLER_4_115 ();
 sg13g2_fill_2 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_decap_4 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_4 FILLER_4_189 ();
 sg13g2_decap_4 FILLER_4_201 ();
 sg13g2_fill_2 FILLER_4_205 ();
 sg13g2_fill_2 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_243 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_fill_1 FILLER_4_257 ();
 sg13g2_decap_8 FILLER_4_262 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_8 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_fill_1 FILLER_4_290 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_fill_1 FILLER_4_330 ();
 sg13g2_decap_4 FILLER_4_345 ();
 sg13g2_fill_2 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_fill_1 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_fill_2 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_421 ();
 sg13g2_decap_8 FILLER_4_428 ();
 sg13g2_fill_2 FILLER_4_441 ();
 sg13g2_fill_1 FILLER_4_446 ();
 sg13g2_decap_8 FILLER_5_12 ();
 sg13g2_decap_4 FILLER_5_19 ();
 sg13g2_fill_1 FILLER_5_23 ();
 sg13g2_decap_4 FILLER_5_41 ();
 sg13g2_decap_8 FILLER_5_59 ();
 sg13g2_decap_8 FILLER_5_66 ();
 sg13g2_fill_2 FILLER_5_73 ();
 sg13g2_fill_1 FILLER_5_75 ();
 sg13g2_decap_8 FILLER_5_86 ();
 sg13g2_fill_1 FILLER_5_93 ();
 sg13g2_fill_1 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_4 FILLER_5_192 ();
 sg13g2_decap_4 FILLER_5_213 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_fill_1 FILLER_5_250 ();
 sg13g2_fill_2 FILLER_5_272 ();
 sg13g2_fill_1 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_296 ();
 sg13g2_fill_2 FILLER_5_302 ();
 sg13g2_fill_1 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_fill_1 FILLER_5_374 ();
 sg13g2_decap_4 FILLER_5_379 ();
 sg13g2_fill_2 FILLER_5_387 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_426 ();
 sg13g2_fill_1 FILLER_5_442 ();
 sg13g2_fill_2 FILLER_5_446 ();
 sg13g2_decap_8 FILLER_6_8 ();
 sg13g2_decap_8 FILLER_6_15 ();
 sg13g2_decap_4 FILLER_6_22 ();
 sg13g2_fill_2 FILLER_6_43 ();
 sg13g2_fill_1 FILLER_6_45 ();
 sg13g2_fill_2 FILLER_6_84 ();
 sg13g2_fill_2 FILLER_6_144 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_fill_1 FILLER_6_151 ();
 sg13g2_fill_1 FILLER_6_202 ();
 sg13g2_fill_2 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_decap_4 FILLER_6_265 ();
 sg13g2_fill_1 FILLER_6_269 ();
 sg13g2_decap_4 FILLER_6_274 ();
 sg13g2_fill_1 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_fill_2 FILLER_6_301 ();
 sg13g2_fill_2 FILLER_6_357 ();
 sg13g2_fill_1 FILLER_6_359 ();
 sg13g2_decap_4 FILLER_6_387 ();
 sg13g2_fill_2 FILLER_6_391 ();
 sg13g2_fill_1 FILLER_6_414 ();
 sg13g2_fill_1 FILLER_6_439 ();
 sg13g2_fill_1 FILLER_6_450 ();
 sg13g2_decap_8 FILLER_7_8 ();
 sg13g2_decap_8 FILLER_7_15 ();
 sg13g2_fill_2 FILLER_7_22 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_4 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_57 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_fill_1 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_94 ();
 sg13g2_fill_1 FILLER_7_96 ();
 sg13g2_fill_2 FILLER_7_107 ();
 sg13g2_fill_2 FILLER_7_182 ();
 sg13g2_fill_1 FILLER_7_236 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_fill_1 FILLER_7_248 ();
 sg13g2_fill_2 FILLER_7_253 ();
 sg13g2_decap_4 FILLER_7_263 ();
 sg13g2_fill_2 FILLER_7_267 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_fill_2 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_415 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_8 ();
 sg13g2_decap_8 FILLER_8_15 ();
 sg13g2_decap_8 FILLER_8_22 ();
 sg13g2_fill_1 FILLER_8_29 ();
 sg13g2_decap_8 FILLER_8_51 ();
 sg13g2_decap_8 FILLER_8_58 ();
 sg13g2_fill_1 FILLER_8_65 ();
 sg13g2_fill_2 FILLER_8_83 ();
 sg13g2_fill_1 FILLER_8_85 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_fill_1 FILLER_8_135 ();
 sg13g2_fill_2 FILLER_8_153 ();
 sg13g2_fill_1 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_185 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_fill_2 FILLER_8_259 ();
 sg13g2_fill_2 FILLER_8_311 ();
 sg13g2_fill_1 FILLER_8_313 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_fill_2 FILLER_8_376 ();
 sg13g2_fill_2 FILLER_8_395 ();
 sg13g2_fill_1 FILLER_8_397 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_4 FILLER_8_409 ();
 sg13g2_fill_1 FILLER_8_413 ();
 sg13g2_fill_2 FILLER_8_421 ();
 sg13g2_decap_8 FILLER_9_16 ();
 sg13g2_decap_8 FILLER_9_23 ();
 sg13g2_fill_2 FILLER_9_30 ();
 sg13g2_fill_1 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_50 ();
 sg13g2_fill_1 FILLER_9_57 ();
 sg13g2_fill_1 FILLER_9_75 ();
 sg13g2_fill_2 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_103 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_fill_2 FILLER_9_151 ();
 sg13g2_fill_1 FILLER_9_174 ();
 sg13g2_fill_2 FILLER_9_263 ();
 sg13g2_fill_1 FILLER_9_265 ();
 sg13g2_fill_2 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_332 ();
 sg13g2_fill_2 FILLER_9_343 ();
 sg13g2_fill_2 FILLER_9_359 ();
 sg13g2_fill_1 FILLER_9_361 ();
 sg13g2_fill_1 FILLER_9_407 ();
 sg13g2_fill_1 FILLER_9_451 ();
 sg13g2_decap_8 FILLER_10_24 ();
 sg13g2_decap_8 FILLER_10_31 ();
 sg13g2_decap_8 FILLER_10_38 ();
 sg13g2_decap_8 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_52 ();
 sg13g2_fill_2 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_134 ();
 sg13g2_fill_2 FILLER_10_199 ();
 sg13g2_fill_1 FILLER_10_201 ();
 sg13g2_fill_2 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_349 ();
 sg13g2_fill_2 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_439 ();
 assign Co = net237;
endmodule
