magic
tech sky130A
magscale 1 2
timestamp 1740383619
<< viali >>
rect 2789 8585 2823 8619
rect 4169 8585 4203 8619
rect 4905 8585 4939 8619
rect 5549 8585 5583 8619
rect 5825 8585 5859 8619
rect 6101 8585 6135 8619
rect 6561 8585 6595 8619
rect 7297 8585 7331 8619
rect 7665 8585 7699 8619
rect 8033 8585 8067 8619
rect 8677 8585 8711 8619
rect 9413 8585 9447 8619
rect 9689 8585 9723 8619
rect 10057 8585 10091 8619
rect 10425 8585 10459 8619
rect 10793 8585 10827 8619
rect 11253 8585 11287 8619
rect 11989 8585 12023 8619
rect 12265 8585 12299 8619
rect 12633 8585 12667 8619
rect 13001 8585 13035 8619
rect 13461 8585 13495 8619
rect 14473 8585 14507 8619
rect 14841 8585 14875 8619
rect 15209 8585 15243 8619
rect 15577 8585 15611 8619
rect 16037 8585 16071 8619
rect 16405 8585 16439 8619
rect 16957 8585 16991 8619
rect 17509 8585 17543 8619
rect 17969 8585 18003 8619
rect 18521 8585 18555 8619
rect 19073 8585 19107 8619
rect 20177 8585 20211 8619
rect 20453 8585 20487 8619
rect 26249 8585 26283 8619
rect 31585 8585 31619 8619
rect 32137 8585 32171 8619
rect 32781 8585 32815 8619
rect 33149 8585 33183 8619
rect 33517 8585 33551 8619
rect 34253 8585 34287 8619
rect 34805 8585 34839 8619
rect 35633 8585 35667 8619
rect 36645 8585 36679 8619
rect 37749 8585 37783 8619
rect 38577 8585 38611 8619
rect 39037 8585 39071 8619
rect 29101 8517 29135 8551
rect 29285 8517 29319 8551
rect 31677 8517 31711 8551
rect 1409 8449 1443 8483
rect 2513 8449 2547 8483
rect 2605 8449 2639 8483
rect 3249 8449 3283 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 5365 8449 5399 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 6745 8449 6779 8483
rect 7113 8449 7147 8483
rect 7481 8449 7515 8483
rect 7849 8449 7883 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 8493 8449 8527 8483
rect 9137 8449 9171 8483
rect 9229 8449 9263 8483
rect 9873 8449 9907 8483
rect 9965 8449 9999 8483
rect 10609 8449 10643 8483
rect 10977 8449 11011 8483
rect 11069 8449 11103 8483
rect 11805 8449 11839 8483
rect 12449 8449 12483 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 13277 8449 13311 8483
rect 13921 8449 13955 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 15853 8449 15887 8483
rect 16221 8449 16255 8483
rect 17141 8449 17175 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 18337 8449 18371 8483
rect 18613 8449 18647 8483
rect 18889 8449 18923 8483
rect 19533 8449 19567 8483
rect 19625 8449 19659 8483
rect 20085 8449 20119 8483
rect 20361 8449 20395 8483
rect 20637 8449 20671 8483
rect 20729 8449 20763 8483
rect 21189 8449 21223 8483
rect 21281 8449 21315 8483
rect 22017 8449 22051 8483
rect 22109 8449 22143 8483
rect 22569 8449 22603 8483
rect 22661 8449 22695 8483
rect 23121 8449 23155 8483
rect 23213 8449 23247 8483
rect 23673 8449 23707 8483
rect 23765 8449 23799 8483
rect 24225 8449 24259 8483
rect 24409 8449 24443 8483
rect 25329 8449 25363 8483
rect 26433 8449 26467 8483
rect 27905 8449 27939 8483
rect 28181 8449 28215 8483
rect 28457 8449 28491 8483
rect 29561 8449 29595 8483
rect 30481 8449 30515 8483
rect 32321 8449 32355 8483
rect 32597 8449 32631 8483
rect 32965 8449 32999 8483
rect 33333 8449 33367 8483
rect 33701 8449 33735 8483
rect 34069 8449 34103 8483
rect 34989 8449 35023 8483
rect 35357 8449 35391 8483
rect 35449 8449 35483 8483
rect 35817 8449 35851 8483
rect 36461 8449 36495 8483
rect 36829 8449 36863 8483
rect 37289 8449 37323 8483
rect 37933 8449 37967 8483
rect 38301 8449 38335 8483
rect 38393 8449 38427 8483
rect 38853 8449 38887 8483
rect 39221 8449 39255 8483
rect 1685 8381 1719 8415
rect 24685 8381 24719 8415
rect 25605 8381 25639 8415
rect 29837 8381 29871 8415
rect 30757 8381 30791 8415
rect 3065 8313 3099 8347
rect 6929 8313 6963 8347
rect 13737 8313 13771 8347
rect 20913 8313 20947 8347
rect 21005 8313 21039 8347
rect 21465 8313 21499 8347
rect 21833 8313 21867 8347
rect 23489 8313 23523 8347
rect 23949 8313 23983 8347
rect 28089 8313 28123 8347
rect 33885 8313 33919 8347
rect 35173 8313 35207 8347
rect 36001 8313 36035 8347
rect 36277 8313 36311 8347
rect 38117 8313 38151 8347
rect 39405 8313 39439 8347
rect 3433 8245 3467 8279
rect 4537 8245 4571 8279
rect 18797 8245 18831 8279
rect 19349 8245 19383 8279
rect 19809 8245 19843 8279
rect 19901 8245 19935 8279
rect 22293 8245 22327 8279
rect 22385 8245 22419 8279
rect 22845 8245 22879 8279
rect 22937 8245 22971 8279
rect 23397 8245 23431 8279
rect 24041 8245 24075 8279
rect 37473 8245 37507 8279
rect 3433 8041 3467 8075
rect 4261 8041 4295 8075
rect 5089 8041 5123 8075
rect 6193 8041 6227 8075
rect 6745 8041 6779 8075
rect 7389 8041 7423 8075
rect 8401 8041 8435 8075
rect 9045 8041 9079 8075
rect 9597 8041 9631 8075
rect 10057 8041 10091 8075
rect 10609 8041 10643 8075
rect 11437 8041 11471 8075
rect 11989 8041 12023 8075
rect 12909 8041 12943 8075
rect 13645 8041 13679 8075
rect 14565 8041 14599 8075
rect 15117 8041 15151 8075
rect 15485 8041 15519 8075
rect 16221 8041 16255 8075
rect 17693 8041 17727 8075
rect 20177 8041 20211 8075
rect 29009 8041 29043 8075
rect 32137 8041 32171 8075
rect 32413 8041 32447 8075
rect 34805 8041 34839 8075
rect 35725 8041 35759 8075
rect 36369 8041 36403 8075
rect 36921 8041 36955 8075
rect 38025 8041 38059 8075
rect 38209 8041 38243 8075
rect 38669 8041 38703 8075
rect 2973 7973 3007 8007
rect 14105 7973 14139 8007
rect 24685 7973 24719 8007
rect 30113 7973 30147 8007
rect 37565 7973 37599 8007
rect 9321 7905 9355 7939
rect 25605 7905 25639 7939
rect 30941 7905 30975 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 2789 7837 2823 7871
rect 3065 7837 3099 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 4445 7837 4479 7871
rect 5273 7837 5307 7871
rect 6377 7837 6411 7871
rect 6929 7837 6963 7871
rect 7205 7837 7239 7871
rect 8585 7837 8619 7871
rect 9229 7837 9263 7871
rect 9781 7837 9815 7871
rect 10241 7837 10275 7871
rect 10793 7837 10827 7871
rect 11621 7837 11655 7871
rect 12173 7837 12207 7871
rect 12725 7837 12759 7871
rect 13829 7837 13863 7871
rect 14265 7837 14299 7871
rect 14381 7837 14415 7871
rect 14933 7837 14967 7871
rect 15301 7837 15335 7871
rect 16037 7837 16071 7871
rect 18153 7837 18187 7871
rect 18429 7837 18463 7871
rect 19625 7837 19659 7871
rect 20361 7837 20395 7871
rect 20913 7837 20947 7871
rect 24593 7837 24627 7871
rect 24869 7837 24903 7871
rect 25145 7837 25179 7871
rect 25881 7837 25915 7871
rect 28641 7837 28675 7871
rect 29193 7837 29227 7871
rect 29561 7837 29595 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 30849 7837 30883 7871
rect 31217 7837 31251 7871
rect 32045 7837 32079 7871
rect 32321 7837 32355 7871
rect 32597 7837 32631 7871
rect 34989 7837 35023 7871
rect 35909 7837 35943 7871
rect 36185 7837 36219 7871
rect 36737 7837 36771 7871
rect 37749 7837 37783 7871
rect 37841 7837 37875 7871
rect 38393 7837 38427 7871
rect 38485 7837 38519 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 2421 7769 2455 7803
rect 2513 7701 2547 7735
rect 3249 7701 3283 7735
rect 3985 7701 4019 7735
rect 17969 7701 18003 7735
rect 18245 7701 18279 7735
rect 19441 7701 19475 7735
rect 20729 7701 20763 7735
rect 24409 7701 24443 7735
rect 25329 7701 25363 7735
rect 26617 7701 26651 7735
rect 28457 7701 28491 7735
rect 29745 7701 29779 7735
rect 29837 7701 29871 7735
rect 30665 7701 30699 7735
rect 31861 7701 31895 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 7941 7497 7975 7531
rect 11897 7497 11931 7531
rect 13553 7497 13587 7531
rect 15577 7497 15611 7531
rect 15853 7497 15887 7531
rect 19533 7497 19567 7531
rect 24961 7497 24995 7531
rect 26433 7497 26467 7531
rect 30849 7497 30883 7531
rect 34345 7497 34379 7531
rect 36829 7497 36863 7531
rect 38301 7497 38335 7531
rect 38669 7497 38703 7531
rect 39037 7497 39071 7531
rect 2329 7361 2363 7395
rect 2697 7361 2731 7395
rect 2973 7361 3007 7395
rect 7757 7361 7791 7395
rect 8033 7361 8067 7395
rect 8309 7361 8343 7395
rect 9229 7361 9263 7395
rect 11069 7361 11103 7395
rect 11713 7361 11747 7395
rect 12633 7361 12667 7395
rect 15393 7361 15427 7395
rect 15761 7361 15795 7395
rect 16037 7361 16071 7395
rect 16313 7361 16347 7395
rect 18613 7361 18647 7395
rect 19717 7361 19751 7395
rect 20453 7361 20487 7395
rect 20729 7361 20763 7395
rect 21649 7361 21683 7395
rect 24777 7361 24811 7395
rect 25329 7361 25363 7395
rect 26157 7361 26191 7395
rect 26617 7361 26651 7395
rect 27721 7361 27755 7395
rect 30389 7361 30423 7395
rect 30665 7361 30699 7395
rect 34161 7361 34195 7395
rect 36369 7361 36403 7395
rect 36645 7361 36679 7395
rect 37657 7361 37691 7395
rect 37749 7361 37783 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 38853 7361 38887 7395
rect 39221 7361 39255 7395
rect 1409 7293 1443 7327
rect 1685 7293 1719 7327
rect 8493 7293 8527 7327
rect 9346 7293 9380 7327
rect 9505 7293 9539 7327
rect 11345 7293 11379 7327
rect 12357 7293 12391 7327
rect 14197 7293 14231 7327
rect 14356 7293 14390 7327
rect 14473 7293 14507 7327
rect 15209 7293 15243 7327
rect 18337 7293 18371 7327
rect 20591 7293 20625 7327
rect 21465 7293 21499 7327
rect 25053 7293 25087 7327
rect 27997 7293 28031 7327
rect 2881 7225 2915 7259
rect 8217 7225 8251 7259
rect 8953 7225 8987 7259
rect 10333 7225 10367 7259
rect 13369 7225 13403 7259
rect 14749 7225 14783 7259
rect 16129 7225 16163 7259
rect 21005 7225 21039 7259
rect 26065 7225 26099 7259
rect 26985 7225 27019 7259
rect 30573 7225 30607 7259
rect 36553 7225 36587 7259
rect 37933 7225 37967 7259
rect 2513 7157 2547 7191
rect 3157 7157 3191 7191
rect 10149 7157 10183 7191
rect 19349 7157 19383 7191
rect 19809 7157 19843 7191
rect 26341 7157 26375 7191
rect 37473 7157 37507 7191
rect 39405 7157 39439 7191
rect 8769 6953 8803 6987
rect 24501 6953 24535 6987
rect 11437 6885 11471 6919
rect 13921 6885 13955 6919
rect 21373 6885 21407 6919
rect 27997 6885 28031 6919
rect 36737 6885 36771 6919
rect 37013 6885 37047 6919
rect 5641 6817 5675 6851
rect 7757 6817 7791 6851
rect 10032 6817 10066 6851
rect 10149 6817 10183 6851
rect 10425 6817 10459 6851
rect 10885 6817 10919 6851
rect 11805 6817 11839 6851
rect 15301 6817 15335 6851
rect 15945 6817 15979 6851
rect 20223 6817 20257 6851
rect 20361 6817 20395 6851
rect 20637 6817 20671 6851
rect 21097 6817 21131 6851
rect 23121 6817 23155 6851
rect 25789 6817 25823 6851
rect 26433 6817 26467 6851
rect 26847 6817 26881 6851
rect 37289 6817 37323 6851
rect 38025 6817 38059 6851
rect 38393 6817 38427 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 1961 6749 1995 6783
rect 2237 6749 2271 6783
rect 5825 6749 5859 6783
rect 6101 6749 6135 6783
rect 6377 6749 6411 6783
rect 7481 6749 7515 6783
rect 8033 6749 8067 6783
rect 9137 6749 9171 6783
rect 9873 6749 9907 6783
rect 11069 6749 11103 6783
rect 11529 6749 11563 6783
rect 12081 6749 12115 6783
rect 12912 6749 12946 6783
rect 13185 6749 13219 6783
rect 14749 6749 14783 6783
rect 14887 6749 14921 6783
rect 15025 6749 15059 6783
rect 15761 6749 15795 6783
rect 16221 6749 16255 6783
rect 18061 6749 18095 6783
rect 18337 6749 18371 6783
rect 20085 6749 20119 6783
rect 21281 6749 21315 6783
rect 22109 6749 22143 6783
rect 22385 6749 22419 6783
rect 22477 6749 22511 6783
rect 23397 6749 23431 6783
rect 25237 6749 25271 6783
rect 25513 6749 25547 6783
rect 25973 6749 26007 6783
rect 26709 6749 26743 6783
rect 26985 6749 27019 6783
rect 27721 6749 27755 6783
rect 28181 6749 28215 6783
rect 28457 6749 28491 6783
rect 28733 6749 28767 6783
rect 29009 6749 29043 6783
rect 36921 6749 36955 6783
rect 37197 6749 37231 6783
rect 37841 6749 37875 6783
rect 38209 6749 38243 6783
rect 38945 6749 38979 6783
rect 5457 6681 5491 6715
rect 6009 6681 6043 6715
rect 9229 6681 9263 6715
rect 11253 6681 11287 6715
rect 17785 6681 17819 6715
rect 17969 6681 18003 6715
rect 27629 6681 27663 6715
rect 37473 6681 37507 6715
rect 38577 6681 38611 6715
rect 1593 6613 1627 6647
rect 1869 6613 1903 6647
rect 2145 6613 2179 6647
rect 2421 6613 2455 6647
rect 7113 6613 7147 6647
rect 7665 6613 7699 6647
rect 8953 6613 8987 6647
rect 11713 6613 11747 6647
rect 12817 6613 12851 6647
rect 14105 6613 14139 6647
rect 16037 6613 16071 6647
rect 19073 6613 19107 6647
rect 19441 6613 19475 6647
rect 22661 6613 22695 6647
rect 24133 6613 24167 6647
rect 27905 6613 27939 6647
rect 28273 6613 28307 6647
rect 28549 6613 28583 6647
rect 28825 6613 28859 6647
rect 38761 6613 38795 6647
rect 39129 6613 39163 6647
rect 10333 6409 10367 6443
rect 12817 6409 12851 6443
rect 13921 6409 13955 6443
rect 21833 6409 21867 6443
rect 26617 6409 26651 6443
rect 28825 6409 28859 6443
rect 29101 6409 29135 6443
rect 38117 6409 38151 6443
rect 39037 6409 39071 6443
rect 39405 6409 39439 6443
rect 20269 6341 20303 6375
rect 25513 6341 25547 6375
rect 26249 6341 26283 6375
rect 37657 6341 37691 6375
rect 38209 6341 38243 6375
rect 1685 6273 1719 6307
rect 6653 6273 6687 6307
rect 8376 6273 8410 6307
rect 9413 6273 9447 6307
rect 9781 6273 9815 6307
rect 9965 6273 9999 6307
rect 11069 6273 11103 6307
rect 12081 6273 12115 6307
rect 13185 6273 13219 6307
rect 14816 6273 14850 6307
rect 15669 6273 15703 6307
rect 18153 6273 18187 6307
rect 18429 6273 18463 6307
rect 19367 6273 19401 6307
rect 19487 6273 19521 6307
rect 20545 6273 20579 6307
rect 20637 6273 20671 6307
rect 20913 6273 20947 6307
rect 22017 6273 22051 6307
rect 24961 6273 24995 6307
rect 25881 6273 25915 6307
rect 26341 6273 26375 6307
rect 26985 6273 27019 6307
rect 27905 6273 27939 6307
rect 28917 6273 28951 6307
rect 37841 6273 37875 6307
rect 38485 6273 38519 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 1409 6205 1443 6239
rect 6377 6205 6411 6239
rect 8217 6205 8251 6239
rect 8493 6205 8527 6239
rect 8769 6205 8803 6239
rect 9229 6205 9263 6239
rect 10149 6205 10183 6239
rect 11345 6205 11379 6239
rect 11805 6205 11839 6239
rect 12909 6205 12943 6239
rect 14657 6205 14691 6239
rect 14933 6205 14967 6239
rect 15209 6205 15243 6239
rect 15853 6205 15887 6239
rect 18613 6205 18647 6239
rect 19073 6205 19107 6239
rect 19625 6205 19659 6239
rect 27169 6205 27203 6239
rect 27629 6205 27663 6239
rect 28022 6205 28056 6239
rect 28181 6205 28215 6239
rect 7389 6137 7423 6171
rect 18337 6137 18371 6171
rect 20361 6137 20395 6171
rect 21649 6137 21683 6171
rect 7573 6069 7607 6103
rect 9597 6069 9631 6103
rect 14013 6069 14047 6103
rect 25145 6069 25179 6103
rect 25329 6069 25363 6103
rect 38669 6069 38703 6103
rect 1869 5865 1903 5899
rect 2145 5865 2179 5899
rect 9965 5865 9999 5899
rect 12173 5865 12207 5899
rect 20269 5865 20303 5899
rect 37933 5865 37967 5899
rect 38209 5865 38243 5899
rect 39405 5865 39439 5899
rect 1593 5797 1627 5831
rect 27077 5797 27111 5831
rect 39037 5797 39071 5831
rect 8953 5729 8987 5763
rect 24961 5729 24995 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 9229 5661 9263 5695
rect 11161 5661 11195 5695
rect 11437 5661 11471 5695
rect 13093 5661 13127 5695
rect 14105 5661 14139 5695
rect 19257 5661 19291 5695
rect 19533 5661 19567 5695
rect 20361 5661 20395 5695
rect 25237 5661 25271 5695
rect 26065 5661 26099 5695
rect 26341 5661 26375 5695
rect 38117 5661 38151 5695
rect 38393 5661 38427 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 13645 5593 13679 5627
rect 13829 5593 13863 5627
rect 13185 5525 13219 5559
rect 14289 5525 14323 5559
rect 20545 5525 20579 5559
rect 25973 5525 26007 5559
rect 5733 5321 5767 5355
rect 20821 5321 20855 5355
rect 39405 5321 39439 5355
rect 20913 5253 20947 5287
rect 21281 5253 21315 5287
rect 1409 5185 1443 5219
rect 1685 5185 1719 5219
rect 5181 5185 5215 5219
rect 5273 5185 5307 5219
rect 5549 5185 5583 5219
rect 20729 5185 20763 5219
rect 28549 5185 28583 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 28273 5117 28307 5151
rect 1593 5049 1627 5083
rect 5457 5049 5491 5083
rect 1869 4981 1903 5015
rect 5181 4981 5215 5015
rect 21373 4981 21407 5015
rect 29285 4981 29319 5015
rect 39037 4981 39071 5015
rect 4905 4777 4939 4811
rect 39405 4777 39439 4811
rect 6193 4709 6227 4743
rect 29745 4709 29779 4743
rect 39037 4709 39071 4743
rect 5641 4641 5675 4675
rect 5800 4641 5834 4675
rect 6653 4641 6687 4675
rect 6929 4641 6963 4675
rect 11115 4641 11149 4675
rect 11253 4641 11287 4675
rect 11529 4641 11563 4675
rect 11989 4641 12023 4675
rect 12173 4641 12207 4675
rect 18521 4641 18555 4675
rect 21649 4641 21683 4675
rect 21833 4641 21867 4675
rect 22293 4641 22327 4675
rect 22845 4641 22879 4675
rect 1409 4573 1443 4607
rect 1685 4573 1719 4607
rect 5917 4573 5951 4607
rect 6837 4573 6871 4607
rect 7192 4563 7226 4597
rect 10977 4573 11011 4607
rect 16681 4573 16715 4607
rect 18245 4573 18279 4607
rect 18613 4573 18647 4607
rect 22569 4573 22603 4607
rect 22707 4573 22741 4607
rect 29009 4573 29043 4607
rect 29285 4573 29319 4607
rect 29929 4573 29963 4607
rect 38853 4573 38887 4607
rect 39221 4573 39255 4607
rect 4169 4505 4203 4539
rect 16865 4505 16899 4539
rect 1593 4437 1627 4471
rect 1869 4437 1903 4471
rect 4261 4437 4295 4471
rect 4997 4437 5031 4471
rect 7941 4437 7975 4471
rect 10333 4437 10367 4471
rect 18797 4437 18831 4471
rect 23489 4437 23523 4471
rect 28273 4437 28307 4471
rect 5089 4233 5123 4267
rect 8309 4233 8343 4267
rect 11529 4233 11563 4267
rect 19165 4233 19199 4267
rect 30665 4233 30699 4267
rect 3801 4165 3835 4199
rect 5549 4165 5583 4199
rect 11069 4165 11103 4199
rect 11253 4165 11287 4199
rect 15117 4165 15151 4199
rect 19073 4165 19107 4199
rect 29561 4165 29595 4199
rect 29929 4165 29963 4199
rect 30297 4165 30331 4199
rect 1409 4097 1443 4131
rect 1685 4097 1719 4131
rect 4077 4097 4111 4131
rect 4353 4097 4387 4131
rect 5181 4097 5215 4131
rect 6193 4097 6227 4131
rect 6377 4097 6411 4131
rect 7021 4097 7055 4131
rect 7159 4097 7193 4131
rect 7297 4097 7331 4131
rect 8217 4097 8251 4131
rect 9781 4097 9815 4131
rect 12265 4097 12299 4131
rect 12541 4097 12575 4131
rect 16221 4097 16255 4131
rect 17049 4097 17083 4131
rect 18153 4097 18187 4131
rect 21833 4097 21867 4131
rect 22109 4097 22143 4131
rect 23121 4097 23155 4131
rect 23397 4097 23431 4131
rect 23673 4097 23707 4131
rect 23765 4097 23799 4131
rect 24225 4097 24259 4131
rect 28641 4097 28675 4131
rect 29837 4097 29871 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 8033 4029 8067 4063
rect 8401 4029 8435 4063
rect 16497 4029 16531 4063
rect 16773 4029 16807 4063
rect 17877 4029 17911 4063
rect 27445 4029 27479 4063
rect 27629 4029 27663 4063
rect 28089 4029 28123 4063
rect 28365 4029 28399 4063
rect 28482 4029 28516 4063
rect 1869 3961 1903 3995
rect 5365 3961 5399 3995
rect 6009 3961 6043 3995
rect 7573 3961 7607 3995
rect 9965 3961 9999 3995
rect 15301 3961 15335 3995
rect 15485 3961 15519 3995
rect 22937 3961 22971 3995
rect 23213 3961 23247 3995
rect 23489 3961 23523 3995
rect 23949 3961 23983 3995
rect 39405 3961 39439 3995
rect 1593 3893 1627 3927
rect 3893 3893 3927 3927
rect 5641 3893 5675 3927
rect 17785 3893 17819 3927
rect 18889 3893 18923 3927
rect 22845 3893 22879 3927
rect 24041 3893 24075 3927
rect 29285 3893 29319 3927
rect 30849 3893 30883 3927
rect 39037 3893 39071 3927
rect 2145 3689 2179 3723
rect 4997 3689 5031 3723
rect 9597 3689 9631 3723
rect 9689 3689 9723 3723
rect 19073 3689 19107 3723
rect 24133 3689 24167 3723
rect 24409 3689 24443 3723
rect 27261 3689 27295 3723
rect 29377 3689 29411 3723
rect 30021 3689 30055 3723
rect 30297 3689 30331 3723
rect 32965 3689 32999 3723
rect 33241 3689 33275 3723
rect 33793 3689 33827 3723
rect 34345 3689 34379 3723
rect 37473 3689 37507 3723
rect 38117 3689 38151 3723
rect 39405 3689 39439 3723
rect 1593 3621 1627 3655
rect 5549 3621 5583 3655
rect 6653 3621 6687 3655
rect 7941 3621 7975 3655
rect 14105 3621 14139 3655
rect 15485 3621 15519 3655
rect 17969 3621 18003 3655
rect 28181 3621 28215 3655
rect 33425 3621 33459 3655
rect 38669 3621 38703 3655
rect 39037 3621 39071 3655
rect 3985 3553 4019 3587
rect 5641 3553 5675 3587
rect 7548 3553 7582 3587
rect 10241 3553 10275 3587
rect 10425 3553 10459 3587
rect 10885 3553 10919 3587
rect 15117 3553 15151 3587
rect 16681 3553 16715 3587
rect 21189 3553 21223 3587
rect 22293 3553 22327 3587
rect 22477 3553 22511 3587
rect 22937 3553 22971 3587
rect 23330 3553 23364 3587
rect 23489 3553 23523 3587
rect 27721 3553 27755 3587
rect 28457 3553 28491 3587
rect 28574 3553 28608 3587
rect 28733 3553 28767 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 1961 3485 1995 3519
rect 4261 3485 4295 3519
rect 5365 3485 5399 3519
rect 5917 3485 5951 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 9413 3485 9447 3519
rect 9873 3485 9907 3519
rect 9965 3485 9999 3519
rect 11161 3485 11195 3519
rect 11299 3485 11333 3519
rect 11437 3485 11471 3519
rect 12081 3485 12115 3519
rect 12357 3485 12391 3519
rect 14841 3485 14875 3519
rect 16405 3485 16439 3519
rect 16957 3485 16991 3519
rect 17233 3485 17267 3519
rect 18061 3485 18095 3519
rect 18337 3485 18371 3519
rect 21465 3485 21499 3519
rect 23213 3485 23247 3519
rect 24593 3485 24627 3519
rect 27445 3485 27479 3519
rect 27537 3485 27571 3519
rect 29745 3485 29779 3519
rect 30481 3485 30515 3519
rect 30573 3485 30607 3519
rect 32597 3485 32631 3519
rect 32781 3485 32815 3519
rect 33057 3485 33091 3519
rect 33517 3485 33551 3519
rect 33609 3485 33643 3519
rect 33885 3485 33919 3519
rect 34161 3485 34195 3519
rect 37197 3485 37231 3519
rect 37381 3485 37415 3519
rect 37657 3485 37691 3519
rect 38025 3485 38059 3519
rect 38301 3485 38335 3519
rect 38577 3485 38611 3519
rect 38669 3485 38703 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 15301 3417 15335 3451
rect 30113 3417 30147 3451
rect 1869 3349 1903 3383
rect 6745 3349 6779 3383
rect 10149 3349 10183 3383
rect 12173 3349 12207 3383
rect 15669 3349 15703 3383
rect 22201 3349 22235 3383
rect 29653 3349 29687 3383
rect 30757 3349 30791 3383
rect 34069 3349 34103 3383
rect 37013 3349 37047 3383
rect 37289 3349 37323 3383
rect 37933 3349 37967 3383
rect 38393 3349 38427 3383
rect 2513 3145 2547 3179
rect 6193 3145 6227 3179
rect 6561 3145 6595 3179
rect 7757 3145 7791 3179
rect 7941 3145 7975 3179
rect 8401 3145 8435 3179
rect 11529 3145 11563 3179
rect 16681 3145 16715 3179
rect 21649 3145 21683 3179
rect 28273 3145 28307 3179
rect 37933 3145 37967 3179
rect 39405 3145 39439 3179
rect 15301 3077 15335 3111
rect 22477 3077 22511 3111
rect 22845 3077 22879 3111
rect 23213 3077 23247 3111
rect 23581 3077 23615 3111
rect 2329 3009 2363 3043
rect 2605 3009 2639 3043
rect 5181 3009 5215 3043
rect 5457 3009 5491 3043
rect 6377 3009 6411 3043
rect 7021 3009 7055 3043
rect 8125 3009 8159 3043
rect 9321 3009 9355 3043
rect 10057 3009 10091 3043
rect 12265 3009 12299 3043
rect 15669 3009 15703 3043
rect 17417 3009 17451 3043
rect 17693 3009 17727 3043
rect 17785 3009 17819 3043
rect 18061 3009 18095 3043
rect 18337 3009 18371 3043
rect 21465 3009 21499 3043
rect 21925 3009 21959 3043
rect 23305 3009 23339 3043
rect 23857 3009 23891 3043
rect 27537 3009 27571 3043
rect 28641 3009 28675 3043
rect 29469 3009 29503 3043
rect 37749 3009 37783 3043
rect 38301 3009 38335 3043
rect 38761 3009 38795 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 6745 2941 6779 2975
rect 9045 2941 9079 2975
rect 9204 2941 9238 2975
rect 9597 2941 9631 2975
rect 10241 2941 10275 2975
rect 12541 2941 12575 2975
rect 15853 2941 15887 2975
rect 27261 2941 27295 2975
rect 28365 2941 28399 2975
rect 2789 2873 2823 2907
rect 19073 2873 19107 2907
rect 22109 2873 22143 2907
rect 24041 2873 24075 2907
rect 29377 2873 29411 2907
rect 15393 2805 15427 2839
rect 17969 2805 18003 2839
rect 22293 2805 22327 2839
rect 29653 2805 29687 2839
rect 38485 2805 38519 2839
rect 39037 2805 39071 2839
rect 2513 2601 2547 2635
rect 39405 2601 39439 2635
rect 3065 2533 3099 2567
rect 23029 2533 23063 2567
rect 22017 2465 22051 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 2329 2397 2363 2431
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 4261 2397 4295 2431
rect 5641 2397 5675 2431
rect 7021 2397 7055 2431
rect 8125 2397 8159 2431
rect 9413 2397 9447 2431
rect 9781 2397 9815 2431
rect 11161 2397 11195 2431
rect 22293 2397 22327 2431
rect 28549 2397 28583 2431
rect 37749 2397 37783 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 2697 2261 2731 2295
rect 4077 2261 4111 2295
rect 5457 2261 5491 2295
rect 6837 2261 6871 2295
rect 8309 2261 8343 2295
rect 9597 2261 9631 2295
rect 10977 2261 11011 2295
rect 28365 2261 28399 2295
rect 37933 2261 37967 2295
rect 38301 2261 38335 2295
rect 38669 2261 38703 2295
rect 39037 2261 39071 2295
<< metal1 >>
rect 26970 11160 26976 11212
rect 27028 11200 27034 11212
rect 37366 11200 37372 11212
rect 27028 11172 37372 11200
rect 27028 11160 27034 11172
rect 37366 11160 37372 11172
rect 37424 11160 37430 11212
rect 27246 11092 27252 11144
rect 27304 11132 27310 11144
rect 37550 11132 37556 11144
rect 27304 11104 37556 11132
rect 27304 11092 27310 11104
rect 37550 11092 37556 11104
rect 37608 11092 37614 11144
rect 26694 11024 26700 11076
rect 26752 11064 26758 11076
rect 35986 11064 35992 11076
rect 26752 11036 35992 11064
rect 26752 11024 26758 11036
rect 35986 11024 35992 11036
rect 36044 11024 36050 11076
rect 25866 10956 25872 11008
rect 25924 10996 25930 11008
rect 34606 10996 34612 11008
rect 25924 10968 34612 10996
rect 25924 10956 25930 10968
rect 34606 10956 34612 10968
rect 34664 10956 34670 11008
rect 19426 10344 19432 10396
rect 19484 10384 19490 10396
rect 24118 10384 24124 10396
rect 19484 10356 24124 10384
rect 19484 10344 19490 10356
rect 24118 10344 24124 10356
rect 24176 10344 24182 10396
rect 9950 10276 9956 10328
rect 10008 10316 10014 10328
rect 10008 10288 31754 10316
rect 10008 10276 10014 10288
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 24394 10248 24400 10260
rect 5592 10220 24400 10248
rect 5592 10208 5598 10220
rect 24394 10208 24400 10220
rect 24452 10208 24458 10260
rect 31726 10248 31754 10288
rect 36538 10248 36544 10260
rect 31726 10220 36544 10248
rect 36538 10208 36544 10220
rect 36596 10208 36602 10260
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 26878 10180 26884 10192
rect 10836 10152 26884 10180
rect 10836 10140 10842 10152
rect 26878 10140 26884 10152
rect 26936 10140 26942 10192
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 23566 10112 23572 10124
rect 7892 10084 23572 10112
rect 7892 10072 7898 10084
rect 23566 10072 23572 10084
rect 23624 10072 23630 10124
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 28718 10044 28724 10056
rect 8168 10016 28724 10044
rect 8168 10004 8174 10016
rect 28718 10004 28724 10016
rect 28776 10004 28782 10056
rect 6730 9936 6736 9988
rect 6788 9976 6794 9988
rect 19426 9976 19432 9988
rect 6788 9948 19432 9976
rect 6788 9936 6794 9948
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 24118 9936 24124 9988
rect 24176 9976 24182 9988
rect 29638 9976 29644 9988
rect 24176 9948 29644 9976
rect 24176 9936 24182 9948
rect 29638 9936 29644 9948
rect 29696 9936 29702 9988
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 19334 9908 19340 9920
rect 9548 9880 19340 9908
rect 9548 9868 9554 9880
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 34330 9908 34336 9920
rect 19944 9880 34336 9908
rect 19944 9868 19950 9880
rect 34330 9868 34336 9880
rect 34388 9868 34394 9920
rect 10042 9800 10048 9852
rect 10100 9840 10106 9852
rect 35618 9840 35624 9852
rect 10100 9812 19564 9840
rect 10100 9800 10106 9812
rect 9674 9732 9680 9784
rect 9732 9772 9738 9784
rect 18874 9772 18880 9784
rect 9732 9744 18880 9772
rect 9732 9732 9738 9744
rect 18874 9732 18880 9744
rect 18932 9732 18938 9784
rect 19536 9772 19564 9812
rect 28966 9812 35624 9840
rect 28966 9772 28994 9812
rect 35618 9800 35624 9812
rect 35676 9800 35682 9852
rect 19536 9744 28994 9772
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 37090 9704 37096 9716
rect 8444 9676 37096 9704
rect 8444 9664 8450 9676
rect 37090 9664 37096 9676
rect 37148 9664 37154 9716
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 17218 9636 17224 9648
rect 7524 9608 17224 9636
rect 7524 9596 7530 9608
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 37458 9596 37464 9648
rect 37516 9636 37522 9648
rect 38378 9636 38384 9648
rect 37516 9608 38384 9636
rect 37516 9596 37522 9608
rect 38378 9596 38384 9608
rect 38436 9596 38442 9648
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 10928 9472 12664 9500
rect 10928 9460 10934 9472
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 12636 9432 12664 9472
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 23474 9500 23480 9512
rect 12768 9472 23480 9500
rect 12768 9460 12774 9472
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 19886 9432 19892 9444
rect 4764 9404 12572 9432
rect 12636 9404 19892 9432
rect 4764 9392 4770 9404
rect 12544 9364 12572 9404
rect 19886 9392 19892 9404
rect 19944 9392 19950 9444
rect 15746 9364 15752 9376
rect 12544 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 21634 9364 21640 9376
rect 15856 9336 21640 9364
rect 12526 9256 12532 9308
rect 12584 9296 12590 9308
rect 15856 9296 15884 9336
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 12584 9268 15884 9296
rect 12584 9256 12590 9268
rect 16298 9256 16304 9308
rect 16356 9296 16362 9308
rect 32122 9296 32128 9308
rect 16356 9268 32128 9296
rect 16356 9256 16362 9268
rect 32122 9256 32128 9268
rect 32180 9256 32186 9308
rect 7282 9188 7288 9240
rect 7340 9228 7346 9240
rect 7340 9200 9674 9228
rect 7340 9188 7346 9200
rect 9646 9160 9674 9200
rect 17034 9188 17040 9240
rect 17092 9228 17098 9240
rect 17862 9228 17868 9240
rect 17092 9200 17868 9228
rect 17092 9188 17098 9200
rect 17862 9188 17868 9200
rect 17920 9188 17926 9240
rect 18782 9188 18788 9240
rect 18840 9228 18846 9240
rect 28810 9228 28816 9240
rect 18840 9200 28816 9228
rect 18840 9188 18846 9200
rect 28810 9188 28816 9200
rect 28868 9188 28874 9240
rect 15562 9160 15568 9172
rect 9646 9132 15568 9160
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 29086 9160 29092 9172
rect 17276 9132 29092 9160
rect 17276 9120 17282 9132
rect 29086 9120 29092 9132
rect 29144 9120 29150 9172
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 9766 9092 9772 9104
rect 8352 9064 9772 9092
rect 8352 9052 8358 9064
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 10376 9064 11560 9092
rect 10376 9052 10382 9064
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 11422 9024 11428 9036
rect 4580 8996 11428 9024
rect 4580 8984 4586 8996
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11532 9024 11560 9064
rect 14642 9052 14648 9104
rect 14700 9092 14706 9104
rect 23198 9092 23204 9104
rect 14700 9064 23204 9092
rect 14700 9052 14706 9064
rect 23198 9052 23204 9064
rect 23256 9052 23262 9104
rect 24118 9052 24124 9104
rect 24176 9092 24182 9104
rect 29546 9092 29552 9104
rect 24176 9064 29552 9092
rect 24176 9052 24182 9064
rect 29546 9052 29552 9064
rect 29604 9052 29610 9104
rect 35250 9052 35256 9104
rect 35308 9092 35314 9104
rect 36262 9092 36268 9104
rect 35308 9064 36268 9092
rect 35308 9052 35314 9064
rect 36262 9052 36268 9064
rect 36320 9052 36326 9104
rect 17770 9024 17776 9036
rect 11532 8996 17776 9024
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 18598 8984 18604 9036
rect 18656 9024 18662 9036
rect 27246 9024 27252 9036
rect 18656 8996 27252 9024
rect 18656 8984 18662 8996
rect 27246 8984 27252 8996
rect 27304 8984 27310 9036
rect 27522 8984 27528 9036
rect 27580 9024 27586 9036
rect 36446 9024 36452 9036
rect 27580 8996 36452 9024
rect 27580 8984 27586 8996
rect 36446 8984 36452 8996
rect 36504 8984 36510 9036
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 11054 8956 11060 8968
rect 5960 8928 11060 8956
rect 5960 8916 5966 8928
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 24118 8956 24124 8968
rect 18564 8928 24124 8956
rect 18564 8916 18570 8928
rect 24118 8916 24124 8928
rect 24176 8916 24182 8968
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 29822 8956 29828 8968
rect 27488 8928 29828 8956
rect 27488 8916 27494 8928
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 31570 8916 31576 8968
rect 31628 8956 31634 8968
rect 38838 8956 38844 8968
rect 31628 8928 38844 8956
rect 31628 8916 31634 8928
rect 38838 8916 38844 8928
rect 38896 8916 38902 8968
rect 3602 8848 3608 8900
rect 3660 8888 3666 8900
rect 20806 8888 20812 8900
rect 3660 8860 20812 8888
rect 3660 8848 3666 8860
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 38562 8888 38568 8900
rect 21468 8860 38568 8888
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 8570 8820 8576 8832
rect 5132 8792 8576 8820
rect 5132 8780 5138 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 16390 8820 16396 8832
rect 13320 8792 16396 8820
rect 13320 8780 13326 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 21468 8820 21496 8860
rect 38562 8848 38568 8860
rect 38620 8848 38626 8900
rect 16632 8792 21496 8820
rect 16632 8780 16638 8792
rect 33042 8780 33048 8832
rect 33100 8820 33106 8832
rect 33502 8820 33508 8832
rect 33100 8792 33508 8820
rect 33100 8780 33106 8792
rect 33502 8780 33508 8792
rect 33560 8780 33566 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 37274 8820 37280 8832
rect 34572 8792 37280 8820
rect 34572 8780 34578 8792
rect 37274 8780 37280 8792
rect 37332 8780 37338 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 3510 8616 3516 8628
rect 2823 8588 3516 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 4614 8616 4620 8628
rect 4203 8588 4620 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5442 8616 5448 8628
rect 4939 8588 5448 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5537 8619 5595 8625
rect 5537 8585 5549 8619
rect 5583 8616 5595 8619
rect 5718 8616 5724 8628
rect 5583 8588 5724 8616
rect 5583 8585 5595 8588
rect 5537 8579 5595 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5810 8576 5816 8628
rect 5868 8576 5874 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6270 8616 6276 8628
rect 6135 8588 6276 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6549 8619 6607 8625
rect 6549 8585 6561 8619
rect 6595 8616 6607 8619
rect 6822 8616 6828 8628
rect 6595 8588 6828 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7285 8619 7343 8625
rect 7285 8585 7297 8619
rect 7331 8616 7343 8619
rect 7558 8616 7564 8628
rect 7331 8588 7564 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7653 8619 7711 8625
rect 7653 8585 7665 8619
rect 7699 8616 7711 8619
rect 7926 8616 7932 8628
rect 7699 8588 7932 8616
rect 7699 8585 7711 8588
rect 7653 8579 7711 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8478 8616 8484 8628
rect 8067 8588 8484 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8846 8616 8852 8628
rect 8711 8588 8852 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 9582 8616 9588 8628
rect 9447 8588 9588 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9858 8616 9864 8628
rect 9723 8588 9864 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10042 8576 10048 8628
rect 10100 8576 10106 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11514 8616 11520 8628
rect 11287 8588 11520 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11977 8619 12035 8625
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12066 8616 12072 8628
rect 12023 8588 12072 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 12894 8616 12900 8628
rect 12667 8588 12900 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13170 8616 13176 8628
rect 13035 8588 13176 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13449 8619 13507 8625
rect 13449 8585 13461 8619
rect 13495 8616 13507 8619
rect 13722 8616 13728 8628
rect 13495 8588 13728 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14550 8616 14556 8628
rect 14507 8588 14556 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15654 8616 15660 8628
rect 15611 8588 15660 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16206 8616 16212 8628
rect 16071 8588 16212 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16482 8616 16488 8628
rect 16439 8588 16488 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 16945 8619 17003 8625
rect 16945 8616 16957 8619
rect 16816 8588 16957 8616
rect 16816 8576 16822 8588
rect 16945 8585 16957 8588
rect 16991 8585 17003 8619
rect 16945 8579 17003 8585
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17368 8588 17509 8616
rect 17368 8576 17374 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 17920 8588 17969 8616
rect 17920 8576 17926 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 18506 8576 18512 8628
rect 18564 8576 18570 8628
rect 19061 8619 19119 8625
rect 19061 8585 19073 8619
rect 19107 8616 19119 8619
rect 19150 8616 19156 8628
rect 19107 8588 19156 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 19392 8588 20177 8616
rect 19392 8576 19398 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 20441 8619 20499 8625
rect 20441 8616 20453 8619
rect 20312 8588 20453 8616
rect 20312 8576 20318 8588
rect 20441 8585 20453 8588
rect 20487 8585 20499 8619
rect 20441 8579 20499 8585
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 21818 8616 21824 8628
rect 20680 8588 20760 8616
rect 20680 8576 20686 8588
rect 8294 8548 8300 8560
rect 2746 8520 8300 8548
rect 750 8440 756 8492
rect 808 8480 814 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 808 8452 1409 8480
rect 808 8440 814 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 2590 8480 2596 8492
rect 2547 8452 2596 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2746 8412 2774 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 10318 8548 10324 8560
rect 9646 8520 10324 8548
rect 9646 8492 9674 8520
rect 10318 8508 10324 8520
rect 10376 8508 10382 8560
rect 12526 8548 12532 8560
rect 10612 8520 12532 8548
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3510 8480 3516 8492
rect 3283 8452 3516 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4522 8480 4528 8492
rect 4387 8452 4528 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 1719 8384 2774 8412
rect 3620 8412 3648 8443
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 5307 8452 5365 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5353 8449 5365 8452
rect 5399 8480 5411 8483
rect 5534 8480 5540 8492
rect 5399 8452 5540 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5859 8452 5917 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 7282 8480 7288 8492
rect 7147 8452 7288 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7742 8480 7748 8492
rect 7515 8452 7748 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7834 8440 7840 8492
rect 7892 8440 7898 8492
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8168 8452 8217 8480
rect 8168 8440 8174 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8444 8452 8493 8480
rect 8444 8440 8450 8452
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9171 8452 9229 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9217 8449 9229 8452
rect 9263 8480 9275 8483
rect 9490 8480 9496 8492
rect 9263 8452 9496 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9582 8440 9588 8492
rect 9640 8452 9674 8492
rect 10612 8489 10640 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 14734 8548 14740 8560
rect 12820 8520 14740 8548
rect 9861 8483 9919 8489
rect 9640 8440 9646 8452
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9907 8452 9965 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8480 12495 8483
rect 12710 8480 12716 8492
rect 12483 8452 12716 8480
rect 12483 8449 12495 8452
rect 12437 8443 12495 8449
rect 9674 8412 9680 8424
rect 3620 8384 4476 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3786 8344 3792 8356
rect 3099 8316 3792 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 4338 8344 4344 8356
rect 3896 8316 4344 8344
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 3896 8276 3924 8316
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4448 8344 4476 8384
rect 6656 8384 9680 8412
rect 6656 8344 6684 8384
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 11808 8412 11836 8443
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12820 8489 12848 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 18782 8548 18788 8560
rect 15764 8520 18788 8548
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 9784 8384 11836 8412
rect 4448 8316 6684 8344
rect 6917 8347 6975 8353
rect 6917 8313 6929 8347
rect 6963 8344 6975 8347
rect 7374 8344 7380 8356
rect 6963 8316 7380 8344
rect 6963 8313 6975 8316
rect 6917 8307 6975 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 9784 8344 9812 8384
rect 13078 8372 13084 8424
rect 13136 8412 13142 8424
rect 13280 8412 13308 8443
rect 13136 8384 13308 8412
rect 13924 8412 13952 8443
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 15764 8489 15792 8520
rect 18782 8508 18788 8520
rect 18840 8508 18846 8560
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 14918 8412 14924 8424
rect 13924 8384 14924 8412
rect 13136 8372 13142 8384
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 7892 8316 9812 8344
rect 13725 8347 13783 8353
rect 7892 8304 7898 8316
rect 13725 8313 13737 8347
rect 13771 8344 13783 8347
rect 13998 8344 14004 8356
rect 13771 8316 14004 8344
rect 13771 8313 13783 8316
rect 13725 8307 13783 8313
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 15028 8344 15056 8443
rect 14700 8316 15056 8344
rect 15396 8344 15424 8443
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 16172 8452 16221 8480
rect 16172 8440 16178 8452
rect 16209 8449 16221 8452
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17696 8412 17724 8443
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 18325 8483 18383 8489
rect 18325 8449 18337 8483
rect 18371 8480 18383 8483
rect 18414 8480 18420 8492
rect 18371 8452 18420 8480
rect 18371 8449 18383 8452
rect 18325 8443 18383 8449
rect 18414 8440 18420 8452
rect 18472 8440 18478 8492
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 18690 8480 18696 8492
rect 18647 8452 18696 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18966 8480 18972 8492
rect 18923 8452 18972 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19242 8464 19248 8516
rect 19300 8504 19306 8516
rect 19300 8480 19334 8504
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 19300 8464 19533 8480
rect 19306 8452 19533 8464
rect 19521 8449 19533 8452
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 19852 8452 20085 8480
rect 19852 8440 19858 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20349 8483 20407 8489
rect 20349 8480 20361 8483
rect 20220 8452 20361 8480
rect 20220 8440 20226 8452
rect 20349 8449 20361 8452
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 20438 8440 20444 8492
rect 20496 8480 20502 8492
rect 20732 8489 20760 8588
rect 21652 8588 21824 8616
rect 20806 8508 20812 8560
rect 20864 8548 20870 8560
rect 21652 8548 21680 8588
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22060 8588 22232 8616
rect 22060 8576 22066 8588
rect 20864 8520 21680 8548
rect 20864 8508 20870 8520
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 21784 8520 22140 8548
rect 21784 8508 21790 8520
rect 20625 8483 20683 8489
rect 20625 8480 20637 8483
rect 20496 8452 20637 8480
rect 20496 8440 20502 8452
rect 20625 8449 20637 8452
rect 20671 8449 20683 8483
rect 20625 8443 20683 8449
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 20898 8440 20904 8492
rect 20956 8480 20962 8492
rect 21177 8483 21235 8489
rect 21177 8480 21189 8483
rect 20956 8452 21189 8480
rect 20956 8440 20962 8452
rect 21177 8449 21189 8452
rect 21223 8449 21235 8483
rect 21177 8443 21235 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21358 8480 21364 8492
rect 21315 8452 21364 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 21450 8440 21456 8492
rect 21508 8480 21514 8492
rect 22112 8489 22140 8520
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21508 8452 22017 8480
rect 21508 8440 21514 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22204 8480 22232 8588
rect 22554 8576 22560 8628
rect 22612 8616 22618 8628
rect 22612 8588 22784 8616
rect 22612 8576 22618 8588
rect 22278 8508 22284 8560
rect 22336 8548 22342 8560
rect 22336 8520 22692 8548
rect 22336 8508 22342 8520
rect 22664 8489 22692 8520
rect 22557 8483 22615 8489
rect 22557 8480 22569 8483
rect 22204 8452 22569 8480
rect 22097 8443 22155 8449
rect 22557 8449 22569 8452
rect 22603 8449 22615 8483
rect 22557 8443 22615 8449
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22756 8480 22784 8588
rect 23106 8576 23112 8628
rect 23164 8616 23170 8628
rect 23164 8588 23336 8616
rect 23164 8576 23170 8588
rect 22830 8508 22836 8560
rect 22888 8548 22894 8560
rect 22888 8520 23244 8548
rect 22888 8508 22894 8520
rect 23216 8489 23244 8520
rect 23109 8483 23167 8489
rect 23109 8480 23121 8483
rect 22756 8452 23121 8480
rect 22649 8443 22707 8449
rect 23109 8449 23121 8452
rect 23155 8449 23167 8483
rect 23109 8443 23167 8449
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23308 8480 23336 8588
rect 23658 8576 23664 8628
rect 23716 8616 23722 8628
rect 23716 8588 24440 8616
rect 23716 8576 23722 8588
rect 23382 8508 23388 8560
rect 23440 8548 23446 8560
rect 23440 8520 23796 8548
rect 23440 8508 23446 8520
rect 23768 8489 23796 8520
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23308 8452 23673 8480
rect 23201 8443 23259 8449
rect 23661 8449 23673 8452
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 23753 8483 23811 8489
rect 23753 8449 23765 8483
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24412 8489 24440 8588
rect 24578 8576 24584 8628
rect 24636 8616 24642 8628
rect 26237 8619 26295 8625
rect 26237 8616 26249 8619
rect 24636 8588 26249 8616
rect 24636 8576 24642 8588
rect 26237 8585 26249 8588
rect 26283 8585 26295 8619
rect 26237 8579 26295 8585
rect 30374 8576 30380 8628
rect 30432 8616 30438 8628
rect 31573 8619 31631 8625
rect 31573 8616 31585 8619
rect 30432 8588 31585 8616
rect 30432 8576 30438 8588
rect 31573 8585 31585 8588
rect 31619 8585 31631 8619
rect 31573 8579 31631 8585
rect 32122 8576 32128 8628
rect 32180 8576 32186 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32548 8588 32781 8616
rect 32548 8576 32554 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 32858 8576 32864 8628
rect 32916 8616 32922 8628
rect 33137 8619 33195 8625
rect 33137 8616 33149 8619
rect 32916 8588 33149 8616
rect 32916 8576 32922 8588
rect 33137 8585 33149 8588
rect 33183 8585 33195 8619
rect 33137 8579 33195 8585
rect 33502 8576 33508 8628
rect 33560 8576 33566 8628
rect 33594 8576 33600 8628
rect 33652 8616 33658 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 33652 8588 34253 8616
rect 33652 8576 33658 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 34793 8619 34851 8625
rect 34793 8585 34805 8619
rect 34839 8585 34851 8619
rect 34793 8579 34851 8585
rect 25498 8508 25504 8560
rect 25556 8548 25562 8560
rect 25556 8520 28488 8548
rect 25556 8508 25562 8520
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 23992 8452 24225 8480
rect 23992 8440 23998 8452
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8449 24455 8483
rect 24397 8443 24455 8449
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 25317 8483 25375 8489
rect 25317 8480 25329 8483
rect 24820 8452 25329 8480
rect 24820 8440 24826 8452
rect 25317 8449 25329 8452
rect 25363 8449 25375 8483
rect 25317 8443 25375 8449
rect 25406 8440 25412 8492
rect 25464 8480 25470 8492
rect 26421 8483 26479 8489
rect 26421 8480 26433 8483
rect 25464 8452 26433 8480
rect 25464 8440 25470 8452
rect 26421 8449 26433 8452
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 27856 8452 27905 8480
rect 27856 8440 27862 8452
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 28074 8440 28080 8492
rect 28132 8480 28138 8492
rect 28460 8489 28488 8520
rect 29086 8508 29092 8560
rect 29144 8508 29150 8560
rect 29178 8508 29184 8560
rect 29236 8548 29242 8560
rect 29273 8551 29331 8557
rect 29273 8548 29285 8551
rect 29236 8520 29285 8548
rect 29236 8508 29242 8520
rect 29273 8517 29285 8520
rect 29319 8517 29331 8551
rect 29273 8511 29331 8517
rect 31386 8508 31392 8560
rect 31444 8548 31450 8560
rect 31665 8551 31723 8557
rect 31665 8548 31677 8551
rect 31444 8520 31677 8548
rect 31444 8508 31450 8520
rect 31665 8517 31677 8520
rect 31711 8517 31723 8551
rect 31665 8511 31723 8517
rect 33870 8508 33876 8560
rect 33928 8548 33934 8560
rect 34808 8548 34836 8579
rect 34882 8576 34888 8628
rect 34940 8616 34946 8628
rect 35621 8619 35679 8625
rect 35621 8616 35633 8619
rect 34940 8588 35633 8616
rect 34940 8576 34946 8588
rect 35621 8585 35633 8588
rect 35667 8585 35679 8619
rect 35621 8579 35679 8585
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36633 8619 36691 8625
rect 36633 8616 36645 8619
rect 35860 8588 36645 8616
rect 35860 8576 35866 8588
rect 36633 8585 36645 8588
rect 36679 8585 36691 8619
rect 36633 8579 36691 8585
rect 36906 8576 36912 8628
rect 36964 8616 36970 8628
rect 37737 8619 37795 8625
rect 37737 8616 37749 8619
rect 36964 8588 37749 8616
rect 36964 8576 36970 8588
rect 37737 8585 37749 8588
rect 37783 8585 37795 8619
rect 37737 8579 37795 8585
rect 38378 8576 38384 8628
rect 38436 8616 38442 8628
rect 38565 8619 38623 8625
rect 38565 8616 38577 8619
rect 38436 8588 38577 8616
rect 38436 8576 38442 8588
rect 38565 8585 38577 8588
rect 38611 8585 38623 8619
rect 38565 8579 38623 8585
rect 39025 8619 39083 8625
rect 39025 8585 39037 8619
rect 39071 8616 39083 8619
rect 39574 8616 39580 8628
rect 39071 8588 39580 8616
rect 39071 8585 39083 8588
rect 39025 8579 39083 8585
rect 39574 8576 39580 8588
rect 39632 8576 39638 8628
rect 33928 8520 34836 8548
rect 33928 8508 33934 8520
rect 28169 8483 28227 8489
rect 28169 8480 28181 8483
rect 28132 8452 28181 8480
rect 28132 8440 28138 8452
rect 28169 8449 28181 8452
rect 28215 8449 28227 8483
rect 28169 8443 28227 8449
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8449 28503 8483
rect 28445 8443 28503 8449
rect 28626 8440 28632 8492
rect 28684 8480 28690 8492
rect 29549 8483 29607 8489
rect 29549 8480 29561 8483
rect 28684 8452 29561 8480
rect 28684 8440 28690 8452
rect 29549 8449 29561 8452
rect 29595 8449 29607 8483
rect 29549 8443 29607 8449
rect 30282 8440 30288 8492
rect 30340 8480 30346 8492
rect 30469 8483 30527 8489
rect 30469 8480 30481 8483
rect 30340 8452 30481 8480
rect 30340 8440 30346 8452
rect 30469 8449 30481 8452
rect 30515 8449 30527 8483
rect 30469 8443 30527 8449
rect 31110 8440 31116 8492
rect 31168 8480 31174 8492
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 31168 8452 32321 8480
rect 31168 8440 31174 8452
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 32585 8483 32643 8489
rect 32585 8449 32597 8483
rect 32631 8449 32643 8483
rect 32585 8443 32643 8449
rect 17696 8384 19196 8412
rect 18690 8344 18696 8356
rect 15396 8316 18696 8344
rect 14700 8304 14706 8316
rect 18690 8304 18696 8316
rect 18748 8304 18754 8356
rect 19168 8344 19196 8384
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 19300 8384 20668 8412
rect 19300 8372 19306 8384
rect 20346 8344 20352 8356
rect 19168 8316 20352 8344
rect 20346 8304 20352 8316
rect 20404 8304 20410 8356
rect 3467 8248 3924 8276
rect 4525 8279 4583 8285
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 4525 8245 4537 8279
rect 4571 8276 4583 8279
rect 5166 8276 5172 8288
rect 4571 8248 5172 8276
rect 4571 8245 4583 8248
rect 4525 8239 4583 8245
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 10042 8276 10048 8288
rect 8444 8248 10048 8276
rect 8444 8236 8450 8248
rect 10042 8236 10048 8248
rect 10100 8276 10106 8288
rect 17218 8276 17224 8288
rect 10100 8248 17224 8276
rect 10100 8236 10106 8248
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 18782 8236 18788 8288
rect 18840 8236 18846 8288
rect 19337 8279 19395 8285
rect 19337 8245 19349 8279
rect 19383 8276 19395 8279
rect 19426 8276 19432 8288
rect 19383 8248 19432 8276
rect 19383 8245 19395 8248
rect 19337 8239 19395 8245
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 19794 8236 19800 8288
rect 19852 8236 19858 8288
rect 19886 8236 19892 8288
rect 19944 8236 19950 8288
rect 20640 8276 20668 8384
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 21600 8384 22094 8412
rect 21600 8372 21606 8384
rect 20806 8304 20812 8356
rect 20864 8344 20870 8356
rect 20901 8347 20959 8353
rect 20901 8344 20913 8347
rect 20864 8316 20913 8344
rect 20864 8304 20870 8316
rect 20901 8313 20913 8316
rect 20947 8313 20959 8347
rect 20901 8307 20959 8313
rect 20990 8304 20996 8356
rect 21048 8304 21054 8356
rect 21450 8304 21456 8356
rect 21508 8304 21514 8356
rect 21726 8304 21732 8356
rect 21784 8344 21790 8356
rect 21821 8347 21879 8353
rect 21821 8344 21833 8347
rect 21784 8316 21833 8344
rect 21784 8304 21790 8316
rect 21821 8313 21833 8316
rect 21867 8313 21879 8347
rect 22066 8344 22094 8384
rect 24670 8372 24676 8424
rect 24728 8372 24734 8424
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 25593 8415 25651 8421
rect 25593 8412 25605 8415
rect 24912 8384 25605 8412
rect 24912 8372 24918 8384
rect 25593 8381 25605 8384
rect 25639 8381 25651 8415
rect 25593 8375 25651 8381
rect 26510 8372 26516 8424
rect 26568 8412 26574 8424
rect 26568 8384 28212 8412
rect 26568 8372 26574 8384
rect 23477 8347 23535 8353
rect 23477 8344 23489 8347
rect 22066 8316 23489 8344
rect 21821 8307 21879 8313
rect 23477 8313 23489 8316
rect 23523 8313 23535 8347
rect 23477 8307 23535 8313
rect 23937 8347 23995 8353
rect 23937 8313 23949 8347
rect 23983 8344 23995 8347
rect 25682 8344 25688 8356
rect 23983 8316 25688 8344
rect 23983 8313 23995 8316
rect 23937 8307 23995 8313
rect 25682 8304 25688 8316
rect 25740 8304 25746 8356
rect 27522 8304 27528 8356
rect 27580 8344 27586 8356
rect 28077 8347 28135 8353
rect 28077 8344 28089 8347
rect 27580 8316 28089 8344
rect 27580 8304 27586 8316
rect 28077 8313 28089 8316
rect 28123 8313 28135 8347
rect 28184 8344 28212 8384
rect 28534 8372 28540 8424
rect 28592 8412 28598 8424
rect 29825 8415 29883 8421
rect 29825 8412 29837 8415
rect 28592 8384 29837 8412
rect 28592 8372 28598 8384
rect 29825 8381 29837 8384
rect 29871 8381 29883 8415
rect 29825 8375 29883 8381
rect 30745 8415 30803 8421
rect 30745 8381 30757 8415
rect 30791 8381 30803 8415
rect 30745 8375 30803 8381
rect 28184 8316 29224 8344
rect 28077 8307 28135 8313
rect 21358 8276 21364 8288
rect 20640 8248 21364 8276
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 22278 8236 22284 8288
rect 22336 8236 22342 8288
rect 22370 8236 22376 8288
rect 22428 8236 22434 8288
rect 22830 8236 22836 8288
rect 22888 8236 22894 8288
rect 22922 8236 22928 8288
rect 22980 8236 22986 8288
rect 23014 8236 23020 8288
rect 23072 8276 23078 8288
rect 23385 8279 23443 8285
rect 23385 8276 23397 8279
rect 23072 8248 23397 8276
rect 23072 8236 23078 8248
rect 23385 8245 23397 8248
rect 23431 8245 23443 8279
rect 23385 8239 23443 8245
rect 23842 8236 23848 8288
rect 23900 8276 23906 8288
rect 24029 8279 24087 8285
rect 24029 8276 24041 8279
rect 23900 8248 24041 8276
rect 23900 8236 23906 8248
rect 24029 8245 24041 8248
rect 24075 8245 24087 8279
rect 24029 8239 24087 8245
rect 24118 8236 24124 8288
rect 24176 8276 24182 8288
rect 29086 8276 29092 8288
rect 24176 8248 29092 8276
rect 24176 8236 24182 8248
rect 29086 8236 29092 8248
rect 29144 8236 29150 8288
rect 29196 8276 29224 8316
rect 29362 8304 29368 8356
rect 29420 8344 29426 8356
rect 30760 8344 30788 8375
rect 30926 8372 30932 8424
rect 30984 8412 30990 8424
rect 32600 8412 32628 8443
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 32953 8483 33011 8489
rect 32953 8480 32965 8483
rect 32732 8452 32965 8480
rect 32732 8440 32738 8452
rect 32953 8449 32965 8452
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 33321 8483 33379 8489
rect 33321 8449 33333 8483
rect 33367 8449 33379 8483
rect 33321 8443 33379 8449
rect 30984 8384 32628 8412
rect 30984 8372 30990 8384
rect 32858 8372 32864 8424
rect 32916 8412 32922 8424
rect 33336 8412 33364 8443
rect 33686 8440 33692 8492
rect 33744 8440 33750 8492
rect 34054 8440 34060 8492
rect 34112 8440 34118 8492
rect 34977 8483 35035 8489
rect 34977 8449 34989 8483
rect 35023 8480 35035 8483
rect 35158 8480 35164 8492
rect 35023 8452 35164 8480
rect 35023 8449 35035 8452
rect 34977 8443 35035 8449
rect 35158 8440 35164 8452
rect 35216 8440 35222 8492
rect 35342 8440 35348 8492
rect 35400 8440 35406 8492
rect 35434 8440 35440 8492
rect 35492 8440 35498 8492
rect 35802 8440 35808 8492
rect 35860 8440 35866 8492
rect 36449 8483 36507 8489
rect 36449 8449 36461 8483
rect 36495 8449 36507 8483
rect 36449 8443 36507 8449
rect 36817 8483 36875 8489
rect 36817 8449 36829 8483
rect 36863 8480 36875 8483
rect 36998 8480 37004 8492
rect 36863 8452 37004 8480
rect 36863 8449 36875 8452
rect 36817 8443 36875 8449
rect 32916 8384 33364 8412
rect 32916 8372 32922 8384
rect 35066 8372 35072 8424
rect 35124 8412 35130 8424
rect 36464 8412 36492 8443
rect 36998 8440 37004 8452
rect 37056 8440 37062 8492
rect 37274 8440 37280 8492
rect 37332 8440 37338 8492
rect 37826 8440 37832 8492
rect 37884 8480 37890 8492
rect 37921 8483 37979 8489
rect 37921 8480 37933 8483
rect 37884 8452 37933 8480
rect 37884 8440 37890 8452
rect 37921 8449 37933 8452
rect 37967 8449 37979 8483
rect 37921 8443 37979 8449
rect 38286 8440 38292 8492
rect 38344 8440 38350 8492
rect 38378 8440 38384 8492
rect 38436 8440 38442 8492
rect 38838 8440 38844 8492
rect 38896 8440 38902 8492
rect 39206 8440 39212 8492
rect 39264 8440 39270 8492
rect 37642 8412 37648 8424
rect 35124 8384 36032 8412
rect 36464 8384 37648 8412
rect 35124 8372 35130 8384
rect 29420 8316 30788 8344
rect 31496 8316 31708 8344
rect 29420 8304 29426 8316
rect 31496 8276 31524 8316
rect 29196 8248 31524 8276
rect 31680 8276 31708 8316
rect 33410 8304 33416 8356
rect 33468 8344 33474 8356
rect 33873 8347 33931 8353
rect 33873 8344 33885 8347
rect 33468 8316 33885 8344
rect 33468 8304 33474 8316
rect 33873 8313 33885 8316
rect 33919 8313 33931 8347
rect 33873 8307 33931 8313
rect 34146 8304 34152 8356
rect 34204 8344 34210 8356
rect 36004 8353 36032 8384
rect 37642 8372 37648 8384
rect 37700 8372 37706 8424
rect 35161 8347 35219 8353
rect 35161 8344 35173 8347
rect 34204 8316 35173 8344
rect 34204 8304 34210 8316
rect 35161 8313 35173 8316
rect 35207 8313 35219 8347
rect 35161 8307 35219 8313
rect 35989 8347 36047 8353
rect 35989 8313 36001 8347
rect 36035 8313 36047 8347
rect 35989 8307 36047 8313
rect 36262 8304 36268 8356
rect 36320 8304 36326 8356
rect 36354 8304 36360 8356
rect 36412 8344 36418 8356
rect 36412 8316 37136 8344
rect 36412 8304 36418 8316
rect 34698 8276 34704 8288
rect 31680 8248 34704 8276
rect 34698 8236 34704 8248
rect 34756 8236 34762 8288
rect 37108 8276 37136 8316
rect 37182 8304 37188 8356
rect 37240 8344 37246 8356
rect 38105 8347 38163 8353
rect 38105 8344 38117 8347
rect 37240 8316 38117 8344
rect 37240 8304 37246 8316
rect 38105 8313 38117 8316
rect 38151 8313 38163 8347
rect 38105 8307 38163 8313
rect 39390 8304 39396 8356
rect 39448 8304 39454 8356
rect 37461 8279 37519 8285
rect 37461 8276 37473 8279
rect 37108 8248 37473 8276
rect 37461 8245 37473 8248
rect 37507 8245 37519 8279
rect 37461 8239 37519 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 3418 8032 3424 8084
rect 3476 8032 3482 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4120 8044 4261 8072
rect 4120 8032 4126 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4890 8032 4896 8084
rect 4948 8072 4954 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4948 8044 5089 8072
rect 4948 8032 4954 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5077 8035 5135 8041
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 6052 8044 6193 8072
rect 6052 8032 6058 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6604 8044 6745 8072
rect 6604 8032 6610 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7377 8075 7435 8081
rect 7377 8072 7389 8075
rect 7156 8044 7389 8072
rect 7156 8032 7162 8044
rect 7377 8041 7389 8044
rect 7423 8041 7435 8075
rect 7377 8035 7435 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8389 8075 8447 8081
rect 8389 8072 8401 8075
rect 8352 8044 8401 8072
rect 8352 8032 8358 8044
rect 8389 8041 8401 8044
rect 8435 8041 8447 8075
rect 8389 8035 8447 8041
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8812 8044 9045 8072
rect 8812 8032 8818 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 9456 8044 9597 8072
rect 9456 8032 9462 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10134 8072 10140 8084
rect 10091 8044 10140 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10468 8044 10609 8072
rect 10468 8032 10474 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11425 8075 11483 8081
rect 11425 8072 11437 8075
rect 11296 8044 11437 8072
rect 11296 8032 11302 8044
rect 11425 8041 11437 8044
rect 11471 8041 11483 8075
rect 11425 8035 11483 8041
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11848 8044 11989 8072
rect 11848 8032 11854 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12676 8044 12909 8072
rect 12676 8032 12682 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13504 8044 13645 8072
rect 13504 8032 13510 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14182 8072 14188 8084
rect 13780 8044 14188 8072
rect 13780 8032 13786 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14553 8075 14611 8081
rect 14553 8072 14565 8075
rect 14332 8044 14565 8072
rect 14332 8032 14338 8044
rect 14553 8041 14565 8044
rect 14599 8041 14611 8075
rect 14553 8035 14611 8041
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14884 8044 15117 8072
rect 14884 8032 14890 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 15473 8075 15531 8081
rect 15473 8041 15485 8075
rect 15519 8072 15531 8075
rect 15838 8072 15844 8084
rect 15519 8044 15844 8072
rect 15519 8041 15531 8044
rect 15473 8035 15531 8041
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 15988 8044 16221 8072
rect 15988 8032 15994 8044
rect 16209 8041 16221 8044
rect 16255 8041 16267 8075
rect 16209 8035 16267 8041
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 17644 8044 17693 8072
rect 17644 8032 17650 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 20165 8075 20223 8081
rect 20165 8072 20177 8075
rect 18748 8044 20177 8072
rect 18748 8032 18754 8044
rect 20165 8041 20177 8044
rect 20211 8041 20223 8075
rect 20165 8035 20223 8041
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 23106 8072 23112 8084
rect 20312 8044 23112 8072
rect 20312 8032 20318 8044
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 28997 8075 29055 8081
rect 28997 8072 29009 8075
rect 24412 8044 29009 8072
rect 2961 8007 3019 8013
rect 2961 7973 2973 8007
rect 3007 8004 3019 8007
rect 6362 8004 6368 8016
rect 3007 7976 6368 8004
rect 3007 7973 3019 7976
rect 2961 7967 3019 7973
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 7984 7976 12572 8004
rect 7984 7964 7990 7976
rect 566 7896 572 7948
rect 624 7936 630 7948
rect 6178 7936 6184 7948
rect 624 7908 3832 7936
rect 624 7896 630 7908
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 1670 7828 1676 7880
rect 1728 7828 1734 7880
rect 2774 7828 2780 7880
rect 2832 7828 2838 7880
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2924 7840 3065 7868
rect 2924 7828 2930 7840
rect 3053 7837 3065 7840
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 3804 7877 3832 7908
rect 3896 7908 6184 7936
rect 3789 7871 3847 7877
rect 3789 7837 3801 7871
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 2409 7803 2467 7809
rect 2409 7800 2421 7803
rect 992 7772 2421 7800
rect 992 7760 998 7772
rect 2409 7769 2421 7772
rect 2455 7769 2467 7803
rect 3896 7800 3924 7908
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 7374 7936 7380 7948
rect 6380 7908 7380 7936
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5994 7868 6000 7880
rect 5307 7840 6000 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 2409 7763 2467 7769
rect 2746 7772 3924 7800
rect 4448 7800 4476 7831
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6380 7877 6408 7908
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 8720 7908 9321 7936
rect 8720 7896 8726 7908
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 9232 7877 9260 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10870 7936 10876 7948
rect 9732 7908 10876 7936
rect 9732 7896 9738 7908
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 12544 7936 12572 7976
rect 14090 7964 14096 8016
rect 14148 7964 14154 8016
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 14516 7976 16068 8004
rect 14516 7964 14522 7976
rect 10980 7908 12434 7936
rect 12544 7908 14412 7936
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9769 7871 9827 7877
rect 9263 7840 9297 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 9950 7868 9956 7880
rect 9815 7840 9956 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 8202 7800 8208 7812
rect 4448 7772 8208 7800
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 2746 7732 2774 7772
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 8588 7800 8616 7831
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 8588 7772 9812 7800
rect 9784 7744 9812 7772
rect 2547 7704 2774 7732
rect 3237 7735 3295 7741
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3878 7732 3884 7744
rect 3283 7704 3884 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 3973 7735 4031 7741
rect 3973 7701 3985 7735
rect 4019 7732 4031 7735
rect 8846 7732 8852 7744
rect 4019 7704 8852 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 9766 7692 9772 7744
rect 9824 7692 9830 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 10980 7732 11008 7908
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12406 7868 12434 7908
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 12406 7840 12725 7868
rect 12161 7831 12219 7837
rect 12713 7837 12725 7840
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 10284 7704 11008 7732
rect 11624 7732 11652 7831
rect 12176 7800 12204 7831
rect 13814 7828 13820 7880
rect 13872 7828 13878 7880
rect 14090 7868 14096 7880
rect 13924 7840 14096 7868
rect 13924 7800 13952 7840
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14274 7877 14280 7880
rect 14253 7871 14280 7877
rect 14253 7837 14265 7871
rect 14253 7831 14280 7837
rect 14274 7828 14280 7831
rect 14332 7828 14338 7880
rect 14384 7877 14412 7908
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 14792 7908 15424 7936
rect 14792 7896 14798 7908
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14921 7871 14979 7877
rect 14921 7837 14933 7871
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 12176 7772 13952 7800
rect 13538 7732 13544 7744
rect 11624 7704 13544 7732
rect 10284 7692 10290 7704
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 14936 7732 14964 7831
rect 13688 7704 14964 7732
rect 15304 7732 15332 7831
rect 15396 7800 15424 7908
rect 16040 7877 16068 7976
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 21910 8004 21916 8016
rect 17276 7976 21916 8004
rect 17276 7964 17282 7976
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16264 7908 19564 7936
rect 16264 7896 16270 7908
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 17954 7828 17960 7880
rect 18012 7868 18018 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 18012 7840 18153 7868
rect 18012 7828 18018 7840
rect 18141 7837 18153 7840
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 18417 7871 18475 7877
rect 18417 7868 18429 7871
rect 18288 7840 18429 7868
rect 18288 7828 18294 7840
rect 18417 7837 18429 7840
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 19536 7800 19564 7908
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 20036 7908 21036 7936
rect 20036 7896 20042 7908
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 20254 7800 20260 7812
rect 15396 7772 19472 7800
rect 19536 7772 20260 7800
rect 15378 7732 15384 7744
rect 15304 7704 15384 7732
rect 13688 7692 13694 7704
rect 15378 7692 15384 7704
rect 15436 7732 15442 7744
rect 16206 7732 16212 7744
rect 15436 7704 16212 7732
rect 15436 7692 15442 7704
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 19444 7741 19472 7772
rect 20254 7760 20260 7772
rect 20312 7760 20318 7812
rect 20916 7800 20944 7831
rect 20364 7772 20944 7800
rect 21008 7800 21036 7908
rect 23106 7896 23112 7948
rect 23164 7936 23170 7948
rect 24412 7936 24440 8044
rect 28997 8041 29009 8044
rect 29043 8041 29055 8075
rect 28997 8035 29055 8041
rect 29086 8032 29092 8084
rect 29144 8072 29150 8084
rect 32125 8075 32183 8081
rect 32125 8072 32137 8075
rect 29144 8044 32137 8072
rect 29144 8032 29150 8044
rect 32125 8041 32137 8044
rect 32171 8041 32183 8075
rect 32125 8035 32183 8041
rect 32306 8032 32312 8084
rect 32364 8072 32370 8084
rect 32401 8075 32459 8081
rect 32401 8072 32413 8075
rect 32364 8044 32413 8072
rect 32364 8032 32370 8044
rect 32401 8041 32413 8044
rect 32447 8041 32459 8075
rect 32401 8035 32459 8041
rect 34422 8032 34428 8084
rect 34480 8072 34486 8084
rect 34793 8075 34851 8081
rect 34793 8072 34805 8075
rect 34480 8044 34805 8072
rect 34480 8032 34486 8044
rect 34793 8041 34805 8044
rect 34839 8041 34851 8075
rect 34793 8035 34851 8041
rect 35526 8032 35532 8084
rect 35584 8072 35590 8084
rect 35713 8075 35771 8081
rect 35713 8072 35725 8075
rect 35584 8044 35725 8072
rect 35584 8032 35590 8044
rect 35713 8041 35725 8044
rect 35759 8041 35771 8075
rect 35713 8035 35771 8041
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36357 8075 36415 8081
rect 36357 8072 36369 8075
rect 36136 8044 36369 8072
rect 36136 8032 36142 8044
rect 36357 8041 36369 8044
rect 36403 8041 36415 8075
rect 36357 8035 36415 8041
rect 36630 8032 36636 8084
rect 36688 8072 36694 8084
rect 36909 8075 36967 8081
rect 36909 8072 36921 8075
rect 36688 8044 36921 8072
rect 36688 8032 36694 8044
rect 36909 8041 36921 8044
rect 36955 8041 36967 8075
rect 36909 8035 36967 8041
rect 37734 8032 37740 8084
rect 37792 8072 37798 8084
rect 38013 8075 38071 8081
rect 38013 8072 38025 8075
rect 37792 8044 38025 8072
rect 37792 8032 37798 8044
rect 38013 8041 38025 8044
rect 38059 8041 38071 8075
rect 38013 8035 38071 8041
rect 38197 8075 38255 8081
rect 38197 8041 38209 8075
rect 38243 8072 38255 8075
rect 38286 8072 38292 8084
rect 38243 8044 38292 8072
rect 38243 8041 38255 8044
rect 38197 8035 38255 8041
rect 38286 8032 38292 8044
rect 38344 8032 38350 8084
rect 38654 8032 38660 8084
rect 38712 8032 38718 8084
rect 24673 8007 24731 8013
rect 24673 7973 24685 8007
rect 24719 7973 24731 8007
rect 24673 7967 24731 7973
rect 23164 7908 24440 7936
rect 23164 7896 23170 7908
rect 24210 7828 24216 7880
rect 24268 7868 24274 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24268 7840 24593 7868
rect 24268 7828 24274 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24688 7800 24716 7967
rect 28166 7964 28172 8016
rect 28224 8004 28230 8016
rect 30101 8007 30159 8013
rect 30101 8004 30113 8007
rect 28224 7976 30113 8004
rect 28224 7964 28230 7976
rect 30101 7973 30113 7976
rect 30147 7973 30159 8007
rect 30101 7967 30159 7973
rect 30834 7964 30840 8016
rect 30892 7964 30898 8016
rect 36814 8004 36820 8016
rect 34992 7976 36820 8004
rect 25590 7896 25596 7948
rect 25648 7896 25654 7948
rect 27706 7896 27712 7948
rect 27764 7936 27770 7948
rect 30852 7936 30880 7964
rect 30929 7939 30987 7945
rect 30929 7936 30941 7939
rect 27764 7908 30420 7936
rect 30852 7908 30941 7936
rect 27764 7896 27770 7908
rect 24857 7871 24915 7877
rect 24857 7837 24869 7871
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 21008 7772 24716 7800
rect 18233 7735 18291 7741
rect 18233 7732 18245 7735
rect 18104 7704 18245 7732
rect 18104 7692 18110 7704
rect 18233 7701 18245 7704
rect 18279 7701 18291 7735
rect 18233 7695 18291 7701
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 19702 7692 19708 7744
rect 19760 7732 19766 7744
rect 20364 7732 20392 7772
rect 19760 7704 20392 7732
rect 19760 7692 19766 7704
rect 20714 7692 20720 7744
rect 20772 7692 20778 7744
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 21968 7704 24409 7732
rect 21968 7692 21974 7704
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 24486 7692 24492 7744
rect 24544 7732 24550 7744
rect 24872 7732 24900 7831
rect 25038 7828 25044 7880
rect 25096 7868 25102 7880
rect 25133 7871 25191 7877
rect 25133 7868 25145 7871
rect 25096 7840 25145 7868
rect 25096 7828 25102 7840
rect 25133 7837 25145 7840
rect 25179 7837 25191 7871
rect 25133 7831 25191 7837
rect 25222 7828 25228 7880
rect 25280 7868 25286 7880
rect 25869 7871 25927 7877
rect 25869 7868 25881 7871
rect 25280 7840 25881 7868
rect 25280 7828 25286 7840
rect 25869 7837 25881 7840
rect 25915 7837 25927 7871
rect 25869 7831 25927 7837
rect 25958 7828 25964 7880
rect 26016 7868 26022 7880
rect 28258 7868 28264 7880
rect 26016 7840 28264 7868
rect 26016 7828 26022 7840
rect 28258 7828 28264 7840
rect 28316 7828 28322 7880
rect 28350 7828 28356 7880
rect 28408 7868 28414 7880
rect 28629 7871 28687 7877
rect 28629 7868 28641 7871
rect 28408 7840 28641 7868
rect 28408 7828 28414 7840
rect 28629 7837 28641 7840
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 28902 7828 28908 7880
rect 28960 7868 28966 7880
rect 29181 7871 29239 7877
rect 29181 7868 29193 7871
rect 28960 7840 29193 7868
rect 28960 7828 28966 7840
rect 29181 7837 29193 7840
rect 29227 7837 29239 7871
rect 29181 7831 29239 7837
rect 29454 7828 29460 7880
rect 29512 7868 29518 7880
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 29512 7840 29561 7868
rect 29512 7828 29518 7840
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 29730 7828 29736 7880
rect 29788 7868 29794 7880
rect 30009 7871 30067 7877
rect 30009 7868 30021 7871
rect 29788 7840 30021 7868
rect 29788 7828 29794 7840
rect 30009 7837 30021 7840
rect 30055 7837 30067 7871
rect 30009 7831 30067 7837
rect 30098 7828 30104 7880
rect 30156 7868 30162 7880
rect 30285 7871 30343 7877
rect 30285 7868 30297 7871
rect 30156 7840 30297 7868
rect 30156 7828 30162 7840
rect 30285 7837 30297 7840
rect 30331 7837 30343 7871
rect 30285 7831 30343 7837
rect 24946 7760 24952 7812
rect 25004 7800 25010 7812
rect 30392 7800 30420 7908
rect 30929 7905 30941 7908
rect 30975 7905 30987 7939
rect 30929 7899 30987 7905
rect 31846 7896 31852 7948
rect 31904 7936 31910 7948
rect 31904 7908 32352 7936
rect 31904 7896 31910 7908
rect 30558 7828 30564 7880
rect 30616 7868 30622 7880
rect 30837 7871 30895 7877
rect 30837 7868 30849 7871
rect 30616 7840 30849 7868
rect 30616 7828 30622 7840
rect 30837 7837 30849 7840
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 31205 7871 31263 7877
rect 31205 7837 31217 7871
rect 31251 7837 31263 7871
rect 31205 7831 31263 7837
rect 31220 7800 31248 7831
rect 31662 7828 31668 7880
rect 31720 7868 31726 7880
rect 32324 7877 32352 7908
rect 34992 7877 35020 7976
rect 36814 7964 36820 7976
rect 36872 7964 36878 8016
rect 37553 8007 37611 8013
rect 37553 7973 37565 8007
rect 37599 7973 37611 8007
rect 37553 7967 37611 7973
rect 37568 7936 37596 7967
rect 35912 7908 37596 7936
rect 35912 7877 35940 7908
rect 38286 7896 38292 7948
rect 38344 7936 38350 7948
rect 38344 7908 38516 7936
rect 38344 7896 38350 7908
rect 32033 7871 32091 7877
rect 32033 7868 32045 7871
rect 31720 7840 32045 7868
rect 31720 7828 31726 7840
rect 32033 7837 32045 7840
rect 32079 7837 32091 7871
rect 32033 7831 32091 7837
rect 32309 7871 32367 7877
rect 32309 7837 32321 7871
rect 32355 7837 32367 7871
rect 32309 7831 32367 7837
rect 32585 7871 32643 7877
rect 32585 7837 32597 7871
rect 32631 7837 32643 7871
rect 32585 7831 32643 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7837 35035 7871
rect 34977 7831 35035 7837
rect 35897 7871 35955 7877
rect 35897 7837 35909 7871
rect 35943 7837 35955 7871
rect 35897 7831 35955 7837
rect 25004 7772 29868 7800
rect 30392 7772 31248 7800
rect 32600 7800 32628 7831
rect 36170 7828 36176 7880
rect 36228 7828 36234 7880
rect 36722 7828 36728 7880
rect 36780 7828 36786 7880
rect 38488 7877 38516 7908
rect 37737 7871 37795 7877
rect 37737 7868 37749 7871
rect 36832 7840 37749 7868
rect 36262 7800 36268 7812
rect 32600 7772 36268 7800
rect 25004 7760 25010 7772
rect 24544 7704 24900 7732
rect 25317 7735 25375 7741
rect 24544 7692 24550 7704
rect 25317 7701 25329 7735
rect 25363 7732 25375 7735
rect 26418 7732 26424 7744
rect 25363 7704 26424 7732
rect 25363 7701 25375 7704
rect 25317 7695 25375 7701
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 26605 7735 26663 7741
rect 26605 7701 26617 7735
rect 26651 7732 26663 7735
rect 27614 7732 27620 7744
rect 26651 7704 27620 7732
rect 26651 7701 26663 7704
rect 26605 7695 26663 7701
rect 27614 7692 27620 7704
rect 27672 7692 27678 7744
rect 28442 7692 28448 7744
rect 28500 7692 28506 7744
rect 29730 7692 29736 7744
rect 29788 7692 29794 7744
rect 29840 7741 29868 7772
rect 36262 7760 36268 7772
rect 36320 7760 36326 7812
rect 29825 7735 29883 7741
rect 29825 7701 29837 7735
rect 29871 7701 29883 7735
rect 29825 7695 29883 7701
rect 30006 7692 30012 7744
rect 30064 7732 30070 7744
rect 30653 7735 30711 7741
rect 30653 7732 30665 7735
rect 30064 7704 30665 7732
rect 30064 7692 30070 7704
rect 30653 7701 30665 7704
rect 30699 7701 30711 7735
rect 30653 7695 30711 7701
rect 30742 7692 30748 7744
rect 30800 7732 30806 7744
rect 31849 7735 31907 7741
rect 31849 7732 31861 7735
rect 30800 7704 31861 7732
rect 30800 7692 30806 7704
rect 31849 7701 31861 7704
rect 31895 7701 31907 7735
rect 31849 7695 31907 7701
rect 34790 7692 34796 7744
rect 34848 7732 34854 7744
rect 36832 7732 36860 7840
rect 37737 7837 37749 7840
rect 37783 7837 37795 7871
rect 37737 7831 37795 7837
rect 37829 7871 37887 7877
rect 37829 7837 37841 7871
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 38381 7871 38439 7877
rect 38381 7837 38393 7871
rect 38427 7837 38439 7871
rect 38381 7831 38439 7837
rect 38473 7871 38531 7877
rect 38473 7837 38485 7871
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 37274 7760 37280 7812
rect 37332 7800 37338 7812
rect 37844 7800 37872 7831
rect 37332 7772 37872 7800
rect 37332 7760 37338 7772
rect 34848 7704 36860 7732
rect 34848 7692 34854 7704
rect 36906 7692 36912 7744
rect 36964 7732 36970 7744
rect 38396 7732 38424 7831
rect 38838 7828 38844 7880
rect 38896 7828 38902 7880
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 38654 7760 38660 7812
rect 38712 7800 38718 7812
rect 39224 7800 39252 7831
rect 38712 7772 39252 7800
rect 38712 7760 38718 7772
rect 36964 7704 38424 7732
rect 36964 7692 36970 7704
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 1210 7488 1216 7540
rect 1268 7528 1274 7540
rect 1268 7500 3004 7528
rect 1268 7488 1274 7500
rect 1302 7420 1308 7472
rect 1360 7460 1366 7472
rect 1360 7432 2728 7460
rect 1360 7420 1366 7432
rect 1118 7352 1124 7404
rect 1176 7392 1182 7404
rect 2700 7401 2728 7432
rect 2976 7401 3004 7500
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 8404 7500 11100 7528
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 1176 7364 2329 7392
rect 1176 7352 1182 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 7926 7392 7932 7404
rect 7791 7364 7932 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 8294 7392 8300 7404
rect 8067 7364 8300 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 290 7284 296 7336
rect 348 7324 354 7336
rect 1397 7327 1455 7333
rect 1397 7324 1409 7327
rect 348 7296 1409 7324
rect 348 7284 354 7296
rect 1397 7293 1409 7296
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 7006 7324 7012 7336
rect 1719 7296 7012 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 8404 7324 8432 7500
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 11072 7401 11100 7500
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 13541 7531 13599 7537
rect 13541 7497 13553 7531
rect 13587 7528 13599 7531
rect 13587 7500 15516 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 15488 7460 15516 7500
rect 15562 7488 15568 7540
rect 15620 7488 15626 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15804 7500 15853 7528
rect 15804 7488 15810 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 19521 7531 19579 7537
rect 19521 7528 19533 7531
rect 16448 7500 19533 7528
rect 16448 7488 16454 7500
rect 19521 7497 19533 7500
rect 19567 7497 19579 7531
rect 20346 7528 20352 7540
rect 19521 7491 19579 7497
rect 19720 7500 20352 7528
rect 19334 7460 19340 7472
rect 11532 7432 12434 7460
rect 15488 7432 16068 7460
rect 11532 7404 11560 7432
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7392 11115 7395
rect 11514 7392 11520 7404
rect 11103 7364 11520 7392
rect 11103 7361 11115 7364
rect 11057 7355 11115 7361
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 12406 7392 12434 7432
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 12406 7364 12633 7392
rect 11701 7355 11759 7361
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 16040 7401 16068 7432
rect 16224 7432 19340 7460
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 15528 7364 15761 7392
rect 15528 7352 15534 7364
rect 15749 7361 15761 7364
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 7116 7296 8432 7324
rect 8481 7327 8539 7333
rect 2869 7259 2927 7265
rect 2869 7225 2881 7259
rect 2915 7256 2927 7259
rect 7116 7256 7144 7296
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8527 7296 9076 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 2915 7228 7144 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 8205 7259 8263 7265
rect 8205 7256 8217 7259
rect 7892 7228 8217 7256
rect 7892 7216 7898 7228
rect 8205 7225 8217 7228
rect 8251 7225 8263 7259
rect 8205 7219 8263 7225
rect 8938 7216 8944 7268
rect 8996 7216 9002 7268
rect 2498 7148 2504 7200
rect 2556 7148 2562 7200
rect 3145 7191 3203 7197
rect 3145 7157 3157 7191
rect 3191 7188 3203 7191
rect 7282 7188 7288 7200
rect 3191 7160 7288 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 9048 7188 9076 7296
rect 9306 7284 9312 7336
rect 9364 7333 9370 7336
rect 9364 7327 9392 7333
rect 9380 7293 9392 7327
rect 9364 7287 9392 7293
rect 9493 7327 9551 7333
rect 9493 7293 9505 7327
rect 9539 7324 9551 7327
rect 9674 7324 9680 7336
rect 9539 7296 9680 7324
rect 9539 7293 9551 7296
rect 9493 7287 9551 7293
rect 9364 7284 9370 7287
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 11333 7327 11391 7333
rect 11333 7293 11345 7327
rect 11379 7324 11391 7327
rect 11790 7324 11796 7336
rect 11379 7296 11796 7324
rect 11379 7293 11391 7296
rect 11333 7287 11391 7293
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 12308 7296 12357 7324
rect 12308 7284 12314 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 14366 7333 14372 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 13044 7296 14197 7324
rect 13044 7284 13050 7296
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14344 7327 14372 7333
rect 14344 7293 14356 7327
rect 14344 7287 14372 7293
rect 14366 7284 14372 7287
rect 14424 7284 14430 7336
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 15010 7324 15016 7336
rect 14507 7296 15016 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7324 15255 7327
rect 16224 7324 16252 7432
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 16298 7352 16304 7404
rect 16356 7352 16362 7404
rect 17770 7352 17776 7404
rect 17828 7392 17834 7404
rect 19720 7401 19748 7500
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 24210 7528 24216 7540
rect 20588 7500 24216 7528
rect 20588 7488 20594 7500
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 24949 7531 25007 7537
rect 24949 7497 24961 7531
rect 24995 7497 25007 7531
rect 24949 7491 25007 7497
rect 24578 7460 24584 7472
rect 21468 7432 24584 7460
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17828 7364 18613 7392
rect 17828 7352 17834 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 18601 7355 18659 7361
rect 19352 7364 19717 7392
rect 19352 7336 19380 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 20438 7352 20444 7404
rect 20496 7352 20502 7404
rect 20714 7352 20720 7404
rect 20772 7352 20778 7404
rect 21468 7392 21496 7432
rect 24578 7420 24584 7432
rect 24636 7420 24642 7472
rect 24964 7460 24992 7491
rect 25774 7488 25780 7540
rect 25832 7528 25838 7540
rect 26421 7531 26479 7537
rect 26421 7528 26433 7531
rect 25832 7500 26433 7528
rect 25832 7488 25838 7500
rect 26421 7497 26433 7500
rect 26467 7497 26479 7531
rect 26421 7491 26479 7497
rect 28258 7488 28264 7540
rect 28316 7528 28322 7540
rect 30374 7528 30380 7540
rect 28316 7500 30380 7528
rect 28316 7488 28322 7500
rect 30374 7488 30380 7500
rect 30432 7488 30438 7540
rect 30837 7531 30895 7537
rect 30837 7497 30849 7531
rect 30883 7528 30895 7531
rect 34333 7531 34391 7537
rect 30883 7500 31754 7528
rect 30883 7497 30895 7500
rect 30837 7491 30895 7497
rect 27890 7460 27896 7472
rect 24964 7432 27896 7460
rect 27890 7420 27896 7432
rect 27948 7420 27954 7472
rect 28350 7420 28356 7472
rect 28408 7460 28414 7472
rect 31570 7460 31576 7472
rect 28408 7432 31576 7460
rect 28408 7420 28414 7432
rect 31570 7420 31576 7432
rect 31628 7420 31634 7472
rect 31726 7460 31754 7500
rect 34333 7497 34345 7531
rect 34379 7528 34391 7531
rect 36722 7528 36728 7540
rect 34379 7500 36728 7528
rect 34379 7497 34391 7500
rect 34333 7491 34391 7497
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 36817 7531 36875 7537
rect 36817 7497 36829 7531
rect 36863 7528 36875 7531
rect 37274 7528 37280 7540
rect 36863 7500 37280 7528
rect 36863 7497 36875 7500
rect 36817 7491 36875 7497
rect 37274 7488 37280 7500
rect 37332 7488 37338 7540
rect 38289 7531 38347 7537
rect 38289 7497 38301 7531
rect 38335 7528 38347 7531
rect 38470 7528 38476 7540
rect 38335 7500 38476 7528
rect 38335 7497 38347 7500
rect 38289 7491 38347 7497
rect 38470 7488 38476 7500
rect 38528 7488 38534 7540
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7497 38715 7531
rect 38657 7491 38715 7497
rect 39025 7531 39083 7537
rect 39025 7497 39037 7531
rect 39071 7528 39083 7531
rect 39482 7528 39488 7540
rect 39071 7500 39488 7528
rect 39071 7497 39083 7500
rect 39025 7491 39083 7497
rect 36170 7460 36176 7472
rect 31726 7432 36176 7460
rect 36170 7420 36176 7432
rect 36228 7420 36234 7472
rect 38672 7460 38700 7491
rect 39482 7488 39488 7500
rect 39540 7488 39546 7540
rect 39850 7460 39856 7472
rect 36280 7432 37688 7460
rect 38672 7432 39856 7460
rect 21284 7364 21496 7392
rect 21637 7395 21695 7401
rect 15243 7296 16252 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 18322 7284 18328 7336
rect 18380 7284 18386 7336
rect 19334 7284 19340 7336
rect 19392 7284 19398 7336
rect 19610 7284 19616 7336
rect 19668 7324 19674 7336
rect 20579 7327 20637 7333
rect 20579 7324 20591 7327
rect 19668 7296 20591 7324
rect 19668 7284 19674 7296
rect 20579 7293 20591 7296
rect 20625 7324 20637 7327
rect 21082 7324 21088 7336
rect 20625 7296 21088 7324
rect 20625 7293 20637 7296
rect 20579 7287 20637 7293
rect 21082 7284 21088 7296
rect 21140 7324 21146 7336
rect 21284 7324 21312 7364
rect 21637 7361 21649 7395
rect 21683 7392 21695 7395
rect 21910 7392 21916 7404
rect 21683 7364 21916 7392
rect 21683 7361 21695 7364
rect 21637 7355 21695 7361
rect 21910 7352 21916 7364
rect 21968 7392 21974 7404
rect 22370 7392 22376 7404
rect 21968 7364 22376 7392
rect 21968 7352 21974 7364
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 24765 7395 24823 7401
rect 24765 7361 24777 7395
rect 24811 7392 24823 7395
rect 25222 7392 25228 7404
rect 24811 7364 25228 7392
rect 24811 7361 24823 7364
rect 24765 7355 24823 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 25314 7352 25320 7404
rect 25372 7392 25378 7404
rect 26145 7395 26203 7401
rect 26145 7392 26157 7395
rect 25372 7364 26157 7392
rect 25372 7352 25378 7364
rect 26145 7361 26157 7364
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 26326 7352 26332 7404
rect 26384 7392 26390 7404
rect 26605 7395 26663 7401
rect 26605 7392 26617 7395
rect 26384 7364 26617 7392
rect 26384 7352 26390 7364
rect 26605 7361 26617 7364
rect 26651 7392 26663 7395
rect 27430 7392 27436 7404
rect 26651 7364 27436 7392
rect 26651 7361 26663 7364
rect 26605 7355 26663 7361
rect 27430 7352 27436 7364
rect 27488 7352 27494 7404
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7392 27767 7395
rect 27798 7392 27804 7404
rect 27755 7364 27804 7392
rect 27755 7361 27767 7364
rect 27709 7355 27767 7361
rect 27798 7352 27804 7364
rect 27856 7352 27862 7404
rect 30377 7395 30435 7401
rect 30377 7361 30389 7395
rect 30423 7361 30435 7395
rect 30377 7355 30435 7361
rect 30653 7395 30711 7401
rect 30653 7361 30665 7395
rect 30699 7392 30711 7395
rect 31478 7392 31484 7404
rect 30699 7364 31484 7392
rect 30699 7361 30711 7364
rect 30653 7355 30711 7361
rect 21140 7296 21312 7324
rect 21140 7284 21146 7296
rect 21358 7284 21364 7336
rect 21416 7324 21422 7336
rect 21453 7327 21511 7333
rect 21453 7324 21465 7327
rect 21416 7296 21465 7324
rect 21416 7284 21422 7296
rect 21453 7293 21465 7296
rect 21499 7293 21511 7327
rect 21453 7287 21511 7293
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 24946 7324 24952 7336
rect 22060 7296 24952 7324
rect 22060 7284 22066 7296
rect 24946 7284 24952 7296
rect 25004 7284 25010 7336
rect 25038 7284 25044 7336
rect 25096 7284 25102 7336
rect 27985 7327 28043 7333
rect 25700 7296 27016 7324
rect 10321 7259 10379 7265
rect 10321 7256 10333 7259
rect 9876 7228 10333 7256
rect 9876 7200 9904 7228
rect 10321 7225 10333 7228
rect 10367 7225 10379 7259
rect 10321 7219 10379 7225
rect 13357 7259 13415 7265
rect 13357 7225 13369 7259
rect 13403 7256 13415 7259
rect 14737 7259 14795 7265
rect 13403 7228 13860 7256
rect 13403 7225 13415 7228
rect 13357 7219 13415 7225
rect 9582 7188 9588 7200
rect 9048 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 10134 7148 10140 7200
rect 10192 7148 10198 7200
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 13630 7188 13636 7200
rect 10652 7160 13636 7188
rect 10652 7148 10658 7160
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13832 7188 13860 7228
rect 14737 7225 14749 7259
rect 14783 7225 14795 7259
rect 14737 7219 14795 7225
rect 14752 7188 14780 7219
rect 14918 7216 14924 7268
rect 14976 7256 14982 7268
rect 16117 7259 16175 7265
rect 16117 7256 16129 7259
rect 14976 7228 16129 7256
rect 14976 7216 14982 7228
rect 16117 7225 16129 7228
rect 16163 7225 16175 7259
rect 19978 7256 19984 7268
rect 16117 7219 16175 7225
rect 18984 7228 19984 7256
rect 13832 7160 14780 7188
rect 14826 7148 14832 7200
rect 14884 7188 14890 7200
rect 18984 7188 19012 7228
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 20993 7259 21051 7265
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 24486 7256 24492 7268
rect 21039 7228 24492 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 24486 7216 24492 7228
rect 24544 7216 24550 7268
rect 14884 7160 19012 7188
rect 14884 7148 14890 7160
rect 19058 7148 19064 7200
rect 19116 7188 19122 7200
rect 19337 7191 19395 7197
rect 19337 7188 19349 7191
rect 19116 7160 19349 7188
rect 19116 7148 19122 7160
rect 19337 7157 19349 7160
rect 19383 7157 19395 7191
rect 19337 7151 19395 7157
rect 19610 7148 19616 7200
rect 19668 7188 19674 7200
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 19668 7160 19809 7188
rect 19668 7148 19674 7160
rect 19797 7157 19809 7160
rect 19843 7157 19855 7191
rect 19797 7151 19855 7157
rect 20346 7148 20352 7200
rect 20404 7188 20410 7200
rect 24118 7188 24124 7200
rect 20404 7160 24124 7188
rect 20404 7148 20410 7160
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24210 7148 24216 7200
rect 24268 7188 24274 7200
rect 25700 7188 25728 7296
rect 26053 7259 26111 7265
rect 26053 7225 26065 7259
rect 26099 7256 26111 7259
rect 26510 7256 26516 7268
rect 26099 7228 26516 7256
rect 26099 7225 26111 7228
rect 26053 7219 26111 7225
rect 26510 7216 26516 7228
rect 26568 7216 26574 7268
rect 26988 7265 27016 7296
rect 27985 7293 27997 7327
rect 28031 7324 28043 7327
rect 28902 7324 28908 7336
rect 28031 7296 28908 7324
rect 28031 7293 28043 7296
rect 27985 7287 28043 7293
rect 28902 7284 28908 7296
rect 28960 7284 28966 7336
rect 30392 7324 30420 7355
rect 31478 7352 31484 7364
rect 31536 7352 31542 7404
rect 34149 7395 34207 7401
rect 34149 7361 34161 7395
rect 34195 7392 34207 7395
rect 34238 7392 34244 7404
rect 34195 7364 34244 7392
rect 34195 7361 34207 7364
rect 34149 7355 34207 7361
rect 34238 7352 34244 7364
rect 34296 7352 34302 7404
rect 34698 7352 34704 7404
rect 34756 7392 34762 7404
rect 36280 7392 36308 7432
rect 34756 7364 36308 7392
rect 34756 7352 34762 7364
rect 36354 7352 36360 7404
rect 36412 7352 36418 7404
rect 36630 7352 36636 7404
rect 36688 7352 36694 7404
rect 37660 7401 37688 7432
rect 39850 7420 39856 7432
rect 39908 7420 39914 7472
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7361 37703 7395
rect 37645 7355 37703 7361
rect 37734 7352 37740 7404
rect 37792 7352 37798 7404
rect 38102 7352 38108 7404
rect 38160 7352 38166 7404
rect 38473 7395 38531 7401
rect 38473 7361 38485 7395
rect 38519 7392 38531 7395
rect 38562 7392 38568 7404
rect 38519 7364 38568 7392
rect 38519 7361 38531 7364
rect 38473 7355 38531 7361
rect 38562 7352 38568 7364
rect 38620 7352 38626 7404
rect 38838 7352 38844 7404
rect 38896 7352 38902 7404
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7392 39267 7395
rect 39574 7392 39580 7404
rect 39255 7364 39580 7392
rect 39255 7361 39267 7364
rect 39209 7355 39267 7361
rect 39574 7352 39580 7364
rect 39632 7352 39638 7404
rect 38378 7324 38384 7336
rect 30392 7296 31524 7324
rect 26973 7259 27031 7265
rect 26973 7225 26985 7259
rect 27019 7225 27031 7259
rect 26973 7219 27031 7225
rect 30561 7259 30619 7265
rect 30561 7225 30573 7259
rect 30607 7256 30619 7259
rect 31496 7256 31524 7296
rect 36556 7296 38384 7324
rect 32766 7256 32772 7268
rect 30607 7228 31156 7256
rect 31496 7228 32772 7256
rect 30607 7225 30619 7228
rect 30561 7219 30619 7225
rect 24268 7160 25728 7188
rect 26329 7191 26387 7197
rect 24268 7148 24274 7160
rect 26329 7157 26341 7191
rect 26375 7188 26387 7191
rect 27246 7188 27252 7200
rect 26375 7160 27252 7188
rect 26375 7157 26387 7160
rect 26329 7151 26387 7157
rect 27246 7148 27252 7160
rect 27304 7148 27310 7200
rect 31128 7188 31156 7228
rect 32766 7216 32772 7228
rect 32824 7216 32830 7268
rect 36556 7265 36584 7296
rect 38378 7284 38384 7296
rect 38436 7284 38442 7336
rect 36541 7259 36599 7265
rect 36541 7225 36553 7259
rect 36587 7225 36599 7259
rect 36541 7219 36599 7225
rect 37921 7259 37979 7265
rect 37921 7225 37933 7259
rect 37967 7256 37979 7259
rect 39482 7256 39488 7268
rect 37967 7228 39488 7256
rect 37967 7225 37979 7228
rect 37921 7219 37979 7225
rect 39482 7216 39488 7228
rect 39540 7216 39546 7268
rect 34514 7188 34520 7200
rect 31128 7160 34520 7188
rect 34514 7148 34520 7160
rect 34572 7148 34578 7200
rect 35618 7148 35624 7200
rect 35676 7188 35682 7200
rect 37461 7191 37519 7197
rect 37461 7188 37473 7191
rect 35676 7160 37473 7188
rect 35676 7148 35682 7160
rect 37461 7157 37473 7160
rect 37507 7157 37519 7191
rect 37461 7151 37519 7157
rect 39390 7148 39396 7200
rect 39448 7148 39454 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8757 6987 8815 6993
rect 7800 6956 8432 6984
rect 7800 6944 7806 6956
rect 1210 6876 1216 6928
rect 1268 6916 1274 6928
rect 1268 6888 1808 6916
rect 1268 6876 1274 6888
rect 842 6808 848 6860
rect 900 6848 906 6860
rect 1780 6848 1808 6888
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 7616 6888 7788 6916
rect 7616 6876 7622 6888
rect 900 6820 1716 6848
rect 1780 6820 2268 6848
rect 900 6808 906 6820
rect 750 6740 756 6792
rect 808 6780 814 6792
rect 1688 6789 1716 6820
rect 2240 6789 2268 6820
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 7760 6857 7788 6888
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6817 7803 6851
rect 8404 6848 8432 6956
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 8938 6984 8944 6996
rect 8803 6956 8944 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9306 6944 9312 6996
rect 9364 6984 9370 6996
rect 22554 6984 22560 6996
rect 9364 6956 22560 6984
rect 9364 6944 9370 6956
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 9324 6916 9352 6944
rect 8536 6888 9352 6916
rect 8536 6876 8542 6888
rect 8404 6820 9352 6848
rect 7745 6811 7803 6817
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 808 6752 1409 6780
rect 808 6740 814 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2332 6752 2774 6780
rect 1026 6672 1032 6724
rect 1084 6712 1090 6724
rect 1964 6712 1992 6743
rect 1084 6684 1992 6712
rect 1084 6672 1090 6684
rect 1578 6604 1584 6656
rect 1636 6604 1642 6656
rect 1762 6604 1768 6656
rect 1820 6644 1826 6656
rect 1857 6647 1915 6653
rect 1857 6644 1869 6647
rect 1820 6616 1869 6644
rect 1820 6604 1826 6616
rect 1857 6613 1869 6616
rect 1903 6613 1915 6647
rect 1857 6607 1915 6613
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 2332 6644 2360 6752
rect 2746 6712 2774 6752
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5592 6752 5825 6780
rect 5592 6740 5598 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6270 6780 6276 6792
rect 6135 6752 6276 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 2746 6684 3648 6712
rect 2179 6616 2360 6644
rect 2409 6647 2467 6653
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 3510 6644 3516 6656
rect 2455 6616 3516 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3620 6644 3648 6684
rect 3694 6672 3700 6724
rect 3752 6712 3758 6724
rect 5442 6712 5448 6724
rect 3752 6684 5448 6712
rect 3752 6672 3758 6684
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 5718 6644 5724 6656
rect 3620 6616 5724 6644
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 5828 6644 5856 6743
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 7469 6783 7527 6789
rect 6411 6752 6592 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 5997 6715 6055 6721
rect 5997 6681 6009 6715
rect 6043 6712 6055 6715
rect 6454 6712 6460 6724
rect 6043 6684 6460 6712
rect 6043 6681 6055 6684
rect 5997 6675 6055 6681
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 6564 6644 6592 6752
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 7650 6780 7656 6792
rect 7515 6752 7656 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8168 6752 9137 6780
rect 8168 6740 8174 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 7282 6672 7288 6724
rect 7340 6712 7346 6724
rect 8036 6712 8064 6740
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 7340 6684 8064 6712
rect 8864 6684 9229 6712
rect 7340 6672 7346 6684
rect 5828 6616 6592 6644
rect 7098 6604 7104 6656
rect 7156 6604 7162 6656
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8864 6644 8892 6684
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 9217 6675 9275 6681
rect 8352 6616 8892 6644
rect 8941 6647 8999 6653
rect 8352 6604 8358 6616
rect 8941 6613 8953 6647
rect 8987 6644 8999 6647
rect 9324 6644 9352 6820
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 10042 6857 10048 6860
rect 10020 6851 10048 6857
rect 10020 6848 10032 6851
rect 9548 6820 10032 6848
rect 9548 6808 9554 6820
rect 10020 6817 10032 6820
rect 10020 6811 10048 6817
rect 10042 6808 10048 6811
rect 10100 6808 10106 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10336 6848 10364 6956
rect 22554 6944 22560 6956
rect 22612 6944 22618 6996
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 22704 6956 23796 6984
rect 22704 6944 22710 6956
rect 11422 6876 11428 6928
rect 11480 6876 11486 6928
rect 13909 6919 13967 6925
rect 13909 6885 13921 6919
rect 13955 6885 13967 6919
rect 13909 6879 13967 6885
rect 10183 6820 10364 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10410 6808 10416 6860
rect 10468 6808 10474 6860
rect 10870 6808 10876 6860
rect 10928 6808 10934 6860
rect 11790 6808 11796 6860
rect 11848 6808 11854 6860
rect 13924 6848 13952 6879
rect 15194 6876 15200 6928
rect 15252 6916 15258 6928
rect 16298 6916 16304 6928
rect 15252 6888 16304 6916
rect 15252 6876 15258 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 18874 6876 18880 6928
rect 18932 6916 18938 6928
rect 19610 6916 19616 6928
rect 18932 6888 19616 6916
rect 18932 6876 18938 6888
rect 19610 6876 19616 6888
rect 19668 6876 19674 6928
rect 21361 6919 21419 6925
rect 21361 6916 21373 6919
rect 20824 6888 21373 6916
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 13924 6820 15301 6848
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15933 6851 15991 6857
rect 15933 6848 15945 6851
rect 15436 6820 15945 6848
rect 15436 6808 15442 6820
rect 15933 6817 15945 6820
rect 15979 6817 15991 6851
rect 15933 6811 15991 6817
rect 17954 6808 17960 6860
rect 18012 6808 18018 6860
rect 19518 6808 19524 6860
rect 19576 6848 19582 6860
rect 20254 6857 20260 6860
rect 20211 6851 20260 6857
rect 20211 6848 20223 6851
rect 19576 6820 20223 6848
rect 19576 6808 19582 6820
rect 20211 6817 20223 6820
rect 20257 6817 20260 6851
rect 20211 6811 20260 6817
rect 20254 6808 20260 6811
rect 20312 6808 20318 6860
rect 20346 6808 20352 6860
rect 20404 6808 20410 6860
rect 20625 6851 20683 6857
rect 20625 6817 20637 6851
rect 20671 6848 20683 6851
rect 20824 6848 20852 6888
rect 21361 6885 21373 6888
rect 21407 6885 21419 6919
rect 23768 6916 23796 6956
rect 24486 6944 24492 6996
rect 24544 6944 24550 6996
rect 25866 6984 25872 6996
rect 24596 6956 25872 6984
rect 24596 6916 24624 6956
rect 25866 6944 25872 6956
rect 25924 6944 25930 6996
rect 26878 6944 26884 6996
rect 26936 6984 26942 6996
rect 26936 6956 28396 6984
rect 26936 6944 26942 6956
rect 23768 6888 24624 6916
rect 21361 6879 21419 6885
rect 27430 6876 27436 6928
rect 27488 6916 27494 6928
rect 27985 6919 28043 6925
rect 27985 6916 27997 6919
rect 27488 6888 27997 6916
rect 27488 6876 27494 6888
rect 27985 6885 27997 6888
rect 28031 6885 28043 6919
rect 27985 6879 28043 6885
rect 20671 6820 20852 6848
rect 20671 6817 20683 6820
rect 20625 6811 20683 6817
rect 20898 6808 20904 6860
rect 20956 6848 20962 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 20956 6820 21097 6848
rect 20956 6808 20962 6820
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 21085 6811 21143 6817
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21542 6848 21548 6860
rect 21232 6820 21548 6848
rect 21232 6808 21238 6820
rect 21542 6808 21548 6820
rect 21600 6808 21606 6860
rect 23106 6808 23112 6860
rect 23164 6808 23170 6860
rect 25682 6808 25688 6860
rect 25740 6848 25746 6860
rect 25777 6851 25835 6857
rect 25777 6848 25789 6851
rect 25740 6820 25789 6848
rect 25740 6808 25746 6820
rect 25777 6817 25789 6820
rect 25823 6817 25835 6851
rect 25777 6811 25835 6817
rect 26421 6851 26479 6857
rect 26421 6817 26433 6851
rect 26467 6848 26479 6851
rect 26510 6848 26516 6860
rect 26467 6820 26516 6848
rect 26467 6817 26479 6820
rect 26421 6811 26479 6817
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 26835 6851 26893 6857
rect 26835 6817 26847 6851
rect 26881 6848 26893 6851
rect 27522 6848 27528 6860
rect 26881 6820 27528 6848
rect 26881 6817 26893 6820
rect 26835 6811 26893 6817
rect 27522 6808 27528 6820
rect 27580 6808 27586 6860
rect 28258 6848 28264 6860
rect 27816 6820 28264 6848
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 11054 6740 11060 6792
rect 11112 6740 11118 6792
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 11624 6752 12081 6780
rect 11241 6715 11299 6721
rect 11241 6681 11253 6715
rect 11287 6712 11299 6715
rect 11624 6712 11652 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12894 6780 12900 6792
rect 12069 6743 12127 6749
rect 12176 6752 12900 6780
rect 11287 6684 11652 6712
rect 11287 6681 11299 6684
rect 11241 6675 11299 6681
rect 8987 6616 9352 6644
rect 8987 6613 8999 6616
rect 8941 6607 8999 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 11256 6644 11284 6675
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 12176 6712 12204 6752
rect 12894 6740 12900 6752
rect 12952 6780 12958 6792
rect 13173 6783 13231 6789
rect 12952 6752 13124 6780
rect 12952 6740 12958 6752
rect 11848 6684 12204 6712
rect 13096 6712 13124 6752
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13262 6780 13268 6792
rect 13219 6752 13268 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 14734 6740 14740 6792
rect 14792 6740 14798 6792
rect 14826 6740 14832 6792
rect 14884 6789 14890 6792
rect 14884 6783 14933 6789
rect 14884 6749 14887 6783
rect 14921 6749 14933 6783
rect 14884 6743 14933 6749
rect 14884 6740 14890 6743
rect 15010 6740 15016 6792
rect 15068 6740 15074 6792
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 17972 6780 18000 6808
rect 27816 6792 27844 6820
rect 28258 6808 28264 6820
rect 28316 6808 28322 6860
rect 28368 6848 28396 6956
rect 36630 6944 36636 6996
rect 36688 6984 36694 6996
rect 39850 6984 39856 6996
rect 36688 6956 39856 6984
rect 36688 6944 36694 6956
rect 39850 6944 39856 6956
rect 39908 6944 39914 6996
rect 36725 6919 36783 6925
rect 36725 6885 36737 6919
rect 36771 6885 36783 6919
rect 36725 6879 36783 6885
rect 36740 6848 36768 6879
rect 36998 6876 37004 6928
rect 37056 6876 37062 6928
rect 28368 6820 36768 6848
rect 37090 6808 37096 6860
rect 37148 6848 37154 6860
rect 37277 6851 37335 6857
rect 37277 6848 37289 6851
rect 37148 6820 37289 6848
rect 37148 6808 37154 6820
rect 37277 6817 37289 6820
rect 37323 6817 37335 6851
rect 37277 6811 37335 6817
rect 37458 6808 37464 6860
rect 37516 6848 37522 6860
rect 37918 6848 37924 6860
rect 37516 6820 37924 6848
rect 37516 6808 37522 6820
rect 37918 6808 37924 6820
rect 37976 6808 37982 6860
rect 38010 6808 38016 6860
rect 38068 6808 38074 6860
rect 38378 6808 38384 6860
rect 38436 6808 38442 6860
rect 16264 6752 18000 6780
rect 18049 6783 18107 6789
rect 16264 6740 16270 6752
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 14182 6712 14188 6724
rect 13096 6684 14188 6712
rect 11848 6672 11854 6684
rect 14182 6672 14188 6684
rect 14240 6672 14246 6724
rect 17770 6672 17776 6724
rect 17828 6672 17834 6724
rect 17954 6672 17960 6724
rect 18012 6672 18018 6724
rect 18064 6712 18092 6743
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 18288 6752 18337 6780
rect 18288 6740 18294 6752
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 20070 6740 20076 6792
rect 20128 6740 20134 6792
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 22002 6780 22008 6792
rect 21324 6752 22008 6780
rect 21324 6740 21330 6752
rect 22002 6740 22008 6752
rect 22060 6740 22066 6792
rect 22094 6740 22100 6792
rect 22152 6740 22158 6792
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 22465 6783 22523 6789
rect 22465 6749 22477 6783
rect 22511 6780 22523 6783
rect 23385 6783 23443 6789
rect 23385 6780 23397 6783
rect 22511 6752 23397 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 23385 6749 23397 6752
rect 23431 6749 23443 6783
rect 23385 6743 23443 6749
rect 18064 6684 18368 6712
rect 18340 6656 18368 6684
rect 9456 6616 11284 6644
rect 9456 6604 9462 6616
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6644 14151 6647
rect 15470 6644 15476 6656
rect 14139 6616 15476 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 16022 6604 16028 6656
rect 16080 6604 16086 6656
rect 18322 6604 18328 6656
rect 18380 6604 18386 6656
rect 19061 6647 19119 6653
rect 19061 6613 19073 6647
rect 19107 6644 19119 6647
rect 19242 6644 19248 6656
rect 19107 6616 19248 6644
rect 19107 6613 19119 6616
rect 19061 6607 19119 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 20438 6644 20444 6656
rect 19475 6616 20444 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 21284 6644 21312 6740
rect 21542 6672 21548 6724
rect 21600 6712 21606 6724
rect 22388 6712 22416 6743
rect 21600 6684 22416 6712
rect 21600 6672 21606 6684
rect 20680 6616 21312 6644
rect 20680 6604 20686 6616
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22480 6644 22508 6743
rect 25222 6740 25228 6792
rect 25280 6740 25286 6792
rect 25314 6740 25320 6792
rect 25372 6780 25378 6792
rect 25501 6783 25559 6789
rect 25501 6780 25513 6783
rect 25372 6752 25513 6780
rect 25372 6740 25378 6752
rect 25501 6749 25513 6752
rect 25547 6749 25559 6783
rect 25501 6743 25559 6749
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6749 26019 6783
rect 25961 6743 26019 6749
rect 23750 6672 23756 6724
rect 23808 6712 23814 6724
rect 25976 6712 26004 6743
rect 26694 6740 26700 6792
rect 26752 6740 26758 6792
rect 26970 6740 26976 6792
rect 27028 6740 27034 6792
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6780 27767 6783
rect 27798 6780 27804 6792
rect 27755 6752 27804 6780
rect 27755 6749 27767 6752
rect 27709 6743 27767 6749
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 28166 6740 28172 6792
rect 28224 6740 28230 6792
rect 28350 6740 28356 6792
rect 28408 6780 28414 6792
rect 28445 6783 28503 6789
rect 28445 6780 28457 6783
rect 28408 6752 28457 6780
rect 28408 6740 28414 6752
rect 28445 6749 28457 6752
rect 28491 6749 28503 6783
rect 28445 6743 28503 6749
rect 28721 6783 28779 6789
rect 28721 6749 28733 6783
rect 28767 6749 28779 6783
rect 28721 6743 28779 6749
rect 23808 6684 26004 6712
rect 27617 6715 27675 6721
rect 23808 6672 23814 6684
rect 27617 6681 27629 6715
rect 27663 6712 27675 6715
rect 28736 6712 28764 6743
rect 28810 6740 28816 6792
rect 28868 6780 28874 6792
rect 28997 6783 29055 6789
rect 28997 6780 29009 6783
rect 28868 6752 29009 6780
rect 28868 6740 28874 6752
rect 28997 6749 29009 6752
rect 29043 6749 29055 6783
rect 28997 6743 29055 6749
rect 34606 6740 34612 6792
rect 34664 6780 34670 6792
rect 36909 6783 36967 6789
rect 36909 6780 36921 6783
rect 34664 6752 36921 6780
rect 34664 6740 34670 6752
rect 36909 6749 36921 6752
rect 36955 6749 36967 6783
rect 36909 6743 36967 6749
rect 37185 6783 37243 6789
rect 37185 6749 37197 6783
rect 37231 6749 37243 6783
rect 37829 6783 37887 6789
rect 37829 6780 37841 6783
rect 37185 6743 37243 6749
rect 37292 6752 37841 6780
rect 27663 6684 28764 6712
rect 27663 6681 27675 6684
rect 27617 6675 27675 6681
rect 30098 6672 30104 6724
rect 30156 6712 30162 6724
rect 37200 6712 37228 6743
rect 30156 6684 37228 6712
rect 30156 6672 30162 6684
rect 22152 6616 22508 6644
rect 22649 6647 22707 6653
rect 22152 6604 22158 6616
rect 22649 6613 22661 6647
rect 22695 6644 22707 6647
rect 24026 6644 24032 6656
rect 22695 6616 24032 6644
rect 22695 6613 22707 6616
rect 22649 6607 22707 6613
rect 24026 6604 24032 6616
rect 24084 6604 24090 6656
rect 24118 6604 24124 6656
rect 24176 6604 24182 6656
rect 25682 6604 25688 6656
rect 25740 6644 25746 6656
rect 26602 6644 26608 6656
rect 25740 6616 26608 6644
rect 25740 6604 25746 6616
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 26694 6604 26700 6656
rect 26752 6644 26758 6656
rect 27798 6644 27804 6656
rect 26752 6616 27804 6644
rect 26752 6604 26758 6616
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 27890 6604 27896 6656
rect 27948 6604 27954 6656
rect 27982 6604 27988 6656
rect 28040 6644 28046 6656
rect 28261 6647 28319 6653
rect 28261 6644 28273 6647
rect 28040 6616 28273 6644
rect 28040 6604 28046 6616
rect 28261 6613 28273 6616
rect 28307 6613 28319 6647
rect 28261 6607 28319 6613
rect 28537 6647 28595 6653
rect 28537 6613 28549 6647
rect 28583 6644 28595 6647
rect 28626 6644 28632 6656
rect 28583 6616 28632 6644
rect 28583 6613 28595 6616
rect 28537 6607 28595 6613
rect 28626 6604 28632 6616
rect 28684 6604 28690 6656
rect 28718 6604 28724 6656
rect 28776 6644 28782 6656
rect 28813 6647 28871 6653
rect 28813 6644 28825 6647
rect 28776 6616 28825 6644
rect 28776 6604 28782 6616
rect 28813 6613 28825 6616
rect 28859 6613 28871 6647
rect 28813 6607 28871 6613
rect 28994 6604 29000 6656
rect 29052 6644 29058 6656
rect 37292 6644 37320 6752
rect 37829 6749 37841 6752
rect 37875 6780 37887 6783
rect 38197 6783 38255 6789
rect 38197 6780 38209 6783
rect 37875 6752 38209 6780
rect 37875 6749 37887 6752
rect 37829 6743 37887 6749
rect 38197 6749 38209 6752
rect 38243 6749 38255 6783
rect 38197 6743 38255 6749
rect 38746 6740 38752 6792
rect 38804 6780 38810 6792
rect 38933 6783 38991 6789
rect 38933 6780 38945 6783
rect 38804 6752 38945 6780
rect 38804 6740 38810 6752
rect 38933 6749 38945 6752
rect 38979 6749 38991 6783
rect 38933 6743 38991 6749
rect 37461 6715 37519 6721
rect 37461 6681 37473 6715
rect 37507 6712 37519 6715
rect 37550 6712 37556 6724
rect 37507 6684 37556 6712
rect 37507 6681 37519 6684
rect 37461 6675 37519 6681
rect 37550 6672 37556 6684
rect 37608 6672 37614 6724
rect 38565 6715 38623 6721
rect 38565 6681 38577 6715
rect 38611 6712 38623 6715
rect 38611 6684 38645 6712
rect 38611 6681 38623 6684
rect 38565 6675 38623 6681
rect 29052 6616 37320 6644
rect 29052 6604 29058 6616
rect 38470 6604 38476 6656
rect 38528 6644 38534 6656
rect 38580 6644 38608 6675
rect 38749 6647 38807 6653
rect 38749 6644 38761 6647
rect 38528 6616 38761 6644
rect 38528 6604 38534 6616
rect 38749 6613 38761 6616
rect 38795 6613 38807 6647
rect 38749 6607 38807 6613
rect 39117 6647 39175 6653
rect 39117 6613 39129 6647
rect 39163 6644 39175 6647
rect 39666 6644 39672 6656
rect 39163 6616 39672 6644
rect 39163 6613 39175 6616
rect 39117 6607 39175 6613
rect 39666 6604 39672 6616
rect 39724 6604 39730 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 3510 6400 3516 6452
rect 3568 6440 3574 6452
rect 6638 6440 6644 6452
rect 3568 6412 6644 6440
rect 3568 6400 3574 6412
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 10321 6443 10379 6449
rect 7708 6412 10272 6440
rect 7708 6400 7714 6412
rect 10134 6372 10140 6384
rect 9784 6344 10140 6372
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 8386 6313 8392 6316
rect 6641 6307 6699 6313
rect 6641 6304 6653 6307
rect 5500 6276 6653 6304
rect 5500 6264 5506 6276
rect 6641 6273 6653 6276
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 8364 6307 8392 6313
rect 8364 6273 8376 6307
rect 8364 6267 8392 6273
rect 8386 6264 8392 6267
rect 8444 6264 8450 6316
rect 9401 6307 9459 6313
rect 9140 6276 9352 6304
rect 566 6196 572 6248
rect 624 6236 630 6248
rect 1397 6239 1455 6245
rect 1397 6236 1409 6239
rect 624 6208 1409 6236
rect 624 6196 630 6208
rect 1397 6205 1409 6208
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6365 6239 6423 6245
rect 6365 6236 6377 6239
rect 6328 6208 6377 6236
rect 6328 6196 6334 6208
rect 6365 6205 6377 6208
rect 6411 6205 6423 6239
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 6365 6199 6423 6205
rect 7392 6208 8217 6236
rect 7392 6177 7420 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8662 6236 8668 6248
rect 8527 6208 8668 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 8754 6196 8760 6248
rect 8812 6196 8818 6248
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 9140 6236 9168 6276
rect 8904 6208 9168 6236
rect 9217 6239 9275 6245
rect 8904 6196 8910 6208
rect 9217 6205 9229 6239
rect 9263 6205 9275 6239
rect 9324 6236 9352 6276
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9490 6304 9496 6316
rect 9447 6276 9496 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9784 6313 9812 6344
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 10244 6372 10272 6412
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10410 6440 10416 6452
rect 10367 6412 10416 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11882 6440 11888 6452
rect 11112 6412 11888 6440
rect 11112 6400 11118 6412
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 12986 6440 12992 6452
rect 12851 6412 12992 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14734 6440 14740 6452
rect 13955 6412 14740 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 18966 6440 18972 6452
rect 18340 6412 18972 6440
rect 10244 6344 14136 6372
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 9968 6236 9996 6267
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 10468 6276 11069 6304
rect 10468 6264 10474 6276
rect 11057 6273 11069 6276
rect 11103 6304 11115 6307
rect 11606 6304 11612 6316
rect 11103 6276 11612 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 11606 6264 11612 6276
rect 11664 6304 11670 6316
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 11664 6276 12081 6304
rect 11664 6264 11670 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 13170 6304 13176 6316
rect 12492 6276 13176 6304
rect 12492 6264 12498 6276
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 9324 6208 9996 6236
rect 10137 6239 10195 6245
rect 9217 6199 9275 6205
rect 10137 6205 10149 6239
rect 10183 6236 10195 6239
rect 10502 6236 10508 6248
rect 10183 6208 10508 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 7377 6171 7435 6177
rect 7377 6137 7389 6171
rect 7423 6137 7435 6171
rect 9232 6168 9260 6199
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 11698 6236 11704 6248
rect 11379 6208 11704 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 9232 6140 10732 6168
rect 7377 6131 7435 6137
rect 10704 6112 10732 6140
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 8110 6100 8116 6112
rect 7607 6072 8116 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 9585 6103 9643 6109
rect 9585 6100 9597 6103
rect 8720 6072 9597 6100
rect 8720 6060 8726 6072
rect 9585 6069 9597 6072
rect 9631 6069 9643 6103
rect 9585 6063 9643 6069
rect 10686 6060 10692 6112
rect 10744 6060 10750 6112
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11808 6100 11836 6199
rect 12894 6196 12900 6248
rect 12952 6196 12958 6248
rect 14108 6236 14136 6344
rect 14826 6313 14832 6316
rect 14804 6307 14832 6313
rect 14804 6273 14816 6307
rect 14804 6267 14832 6273
rect 14826 6264 14832 6267
rect 14884 6264 14890 6316
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 16206 6304 16212 6316
rect 15703 6276 16212 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6304 18199 6307
rect 18230 6304 18236 6316
rect 18187 6276 18236 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 14458 6236 14464 6248
rect 14108 6208 14464 6236
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 14642 6196 14648 6248
rect 14700 6196 14706 6248
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6236 14979 6239
rect 14967 6208 15148 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15120 6168 15148 6208
rect 15194 6196 15200 6248
rect 15252 6196 15258 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 18340 6236 18368 6412
rect 18966 6400 18972 6412
rect 19024 6400 19030 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 19208 6412 20208 6440
rect 19208 6400 19214 6412
rect 18417 6307 18475 6313
rect 18417 6273 18429 6307
rect 18463 6304 18475 6307
rect 18463 6276 18828 6304
rect 18463 6273 18475 6276
rect 18417 6267 18475 6273
rect 15887 6208 18368 6236
rect 18601 6239 18659 6245
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 18601 6205 18613 6239
rect 18647 6236 18659 6239
rect 18690 6236 18696 6248
rect 18647 6208 18696 6236
rect 18647 6205 18659 6208
rect 18601 6199 18659 6205
rect 15378 6168 15384 6180
rect 15120 6140 15384 6168
rect 15378 6128 15384 6140
rect 15436 6128 15442 6180
rect 18325 6171 18383 6177
rect 18325 6137 18337 6171
rect 18371 6168 18383 6171
rect 18506 6168 18512 6180
rect 18371 6140 18512 6168
rect 18371 6137 18383 6140
rect 18325 6131 18383 6137
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 12250 6100 12256 6112
rect 11112 6072 12256 6100
rect 11112 6060 11118 6072
rect 12250 6060 12256 6072
rect 12308 6100 12314 6112
rect 13630 6100 13636 6112
rect 12308 6072 13636 6100
rect 12308 6060 12314 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 14001 6103 14059 6109
rect 14001 6069 14013 6103
rect 14047 6100 14059 6103
rect 14458 6100 14464 6112
rect 14047 6072 14464 6100
rect 14047 6069 14059 6072
rect 14001 6063 14059 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 16114 6100 16120 6112
rect 14608 6072 16120 6100
rect 14608 6060 14614 6072
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 18616 6100 18644 6199
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 16724 6072 18644 6100
rect 18800 6100 18828 6276
rect 19334 6264 19340 6316
rect 19392 6313 19398 6316
rect 19518 6313 19524 6316
rect 19392 6307 19413 6313
rect 19401 6273 19413 6307
rect 19392 6267 19413 6273
rect 19475 6307 19524 6313
rect 19475 6273 19487 6307
rect 19521 6273 19524 6307
rect 19475 6267 19524 6273
rect 19392 6264 19398 6267
rect 19518 6264 19524 6267
rect 19576 6264 19582 6316
rect 20180 6304 20208 6412
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 21450 6440 21456 6452
rect 20864 6412 21456 6440
rect 20864 6400 20870 6412
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 21818 6400 21824 6452
rect 21876 6400 21882 6452
rect 26160 6412 26464 6440
rect 20254 6332 20260 6384
rect 20312 6332 20318 6384
rect 25501 6375 25559 6381
rect 25501 6372 25513 6375
rect 21284 6344 25513 6372
rect 20180 6276 20484 6304
rect 19058 6196 19064 6248
rect 19116 6196 19122 6248
rect 19608 6196 19614 6248
rect 19666 6236 19672 6248
rect 19666 6208 19711 6236
rect 19666 6196 19672 6208
rect 19794 6196 19800 6248
rect 19852 6236 19858 6248
rect 19852 6208 20392 6236
rect 19852 6196 19858 6208
rect 20364 6177 20392 6208
rect 20349 6171 20407 6177
rect 20349 6137 20361 6171
rect 20395 6137 20407 6171
rect 20456 6168 20484 6276
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6304 20683 6307
rect 20806 6304 20812 6316
rect 20671 6276 20812 6304
rect 20671 6273 20683 6276
rect 20625 6267 20683 6273
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 20898 6264 20904 6316
rect 20956 6264 20962 6316
rect 20456 6140 20760 6168
rect 20349 6131 20407 6137
rect 20622 6100 20628 6112
rect 18800 6072 20628 6100
rect 16724 6060 16730 6072
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 20732 6100 20760 6140
rect 21284 6100 21312 6344
rect 25501 6341 25513 6344
rect 25547 6372 25559 6375
rect 26160 6372 26188 6412
rect 25547 6344 26188 6372
rect 25547 6341 25559 6344
rect 25501 6335 25559 6341
rect 26234 6332 26240 6384
rect 26292 6332 26298 6384
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21416 6276 22017 6304
rect 21416 6264 21422 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22830 6264 22836 6316
rect 22888 6304 22894 6316
rect 23382 6304 23388 6316
rect 22888 6276 23388 6304
rect 22888 6264 22894 6276
rect 23382 6264 23388 6276
rect 23440 6304 23446 6316
rect 23440 6276 23888 6304
rect 23440 6264 23446 6276
rect 21450 6196 21456 6248
rect 21508 6236 21514 6248
rect 23750 6236 23756 6248
rect 21508 6208 23756 6236
rect 21508 6196 21514 6208
rect 23750 6196 23756 6208
rect 23808 6196 23814 6248
rect 23860 6236 23888 6276
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 24949 6307 25007 6313
rect 24949 6304 24961 6307
rect 24912 6276 24961 6304
rect 24912 6264 24918 6276
rect 24949 6273 24961 6276
rect 24995 6273 25007 6307
rect 25869 6307 25927 6313
rect 25869 6304 25881 6307
rect 24949 6267 25007 6273
rect 25056 6276 25881 6304
rect 25056 6236 25084 6276
rect 25869 6273 25881 6276
rect 25915 6273 25927 6307
rect 25869 6267 25927 6273
rect 26326 6264 26332 6316
rect 26384 6264 26390 6316
rect 26436 6304 26464 6412
rect 26602 6400 26608 6452
rect 26660 6400 26666 6452
rect 27890 6400 27896 6452
rect 27948 6440 27954 6452
rect 27948 6412 28764 6440
rect 27948 6400 27954 6412
rect 26620 6372 26648 6400
rect 26620 6344 27016 6372
rect 26988 6313 27016 6344
rect 26973 6307 27031 6313
rect 26436 6276 26924 6304
rect 26896 6236 26924 6276
rect 26973 6273 26985 6307
rect 27019 6304 27031 6307
rect 27019 6276 27384 6304
rect 27019 6273 27031 6276
rect 26973 6267 27031 6273
rect 27157 6239 27215 6245
rect 27157 6236 27169 6239
rect 23860 6208 25084 6236
rect 25148 6208 25622 6236
rect 26896 6208 27169 6236
rect 21637 6171 21695 6177
rect 21637 6137 21649 6171
rect 21683 6168 21695 6171
rect 25148 6168 25176 6208
rect 27157 6205 27169 6208
rect 27203 6205 27215 6239
rect 27157 6199 27215 6205
rect 21683 6140 25176 6168
rect 21683 6137 21695 6140
rect 21637 6131 21695 6137
rect 20732 6072 21312 6100
rect 25133 6103 25191 6109
rect 25133 6069 25145 6103
rect 25179 6100 25191 6103
rect 25222 6100 25228 6112
rect 25179 6072 25228 6100
rect 25179 6069 25191 6072
rect 25133 6063 25191 6069
rect 25222 6060 25228 6072
rect 25280 6060 25286 6112
rect 25314 6060 25320 6112
rect 25372 6060 25378 6112
rect 27356 6100 27384 6276
rect 27890 6264 27896 6316
rect 27948 6264 27954 6316
rect 27614 6196 27620 6248
rect 27672 6196 27678 6248
rect 28010 6239 28068 6245
rect 28010 6236 28022 6239
rect 27724 6208 28022 6236
rect 27522 6128 27528 6180
rect 27580 6168 27586 6180
rect 27724 6168 27752 6208
rect 28010 6205 28022 6208
rect 28056 6205 28068 6239
rect 28010 6199 28068 6205
rect 28166 6196 28172 6248
rect 28224 6196 28230 6248
rect 27580 6140 27752 6168
rect 28736 6168 28764 6412
rect 28810 6400 28816 6452
rect 28868 6400 28874 6452
rect 29089 6443 29147 6449
rect 29089 6409 29101 6443
rect 29135 6440 29147 6443
rect 30926 6440 30932 6452
rect 29135 6412 30932 6440
rect 29135 6409 29147 6412
rect 29089 6403 29147 6409
rect 30926 6400 30932 6412
rect 30984 6400 30990 6452
rect 36538 6400 36544 6452
rect 36596 6440 36602 6452
rect 38105 6443 38163 6449
rect 38105 6440 38117 6443
rect 36596 6412 38117 6440
rect 36596 6400 36602 6412
rect 38105 6409 38117 6412
rect 38151 6409 38163 6443
rect 38105 6403 38163 6409
rect 39022 6400 39028 6452
rect 39080 6400 39086 6452
rect 39393 6443 39451 6449
rect 39393 6409 39405 6443
rect 39439 6440 39451 6443
rect 39758 6440 39764 6452
rect 39439 6412 39764 6440
rect 39439 6409 39451 6412
rect 39393 6403 39451 6409
rect 39758 6400 39764 6412
rect 39816 6400 39822 6452
rect 34330 6332 34336 6384
rect 34388 6372 34394 6384
rect 37645 6375 37703 6381
rect 37645 6372 37657 6375
rect 34388 6344 37657 6372
rect 34388 6332 34394 6344
rect 37645 6341 37657 6344
rect 37691 6341 37703 6375
rect 37645 6335 37703 6341
rect 37918 6332 37924 6384
rect 37976 6372 37982 6384
rect 38197 6375 38255 6381
rect 38197 6372 38209 6375
rect 37976 6344 38209 6372
rect 37976 6332 37982 6344
rect 38197 6341 38209 6344
rect 38243 6341 38255 6375
rect 39666 6372 39672 6384
rect 38197 6335 38255 6341
rect 38856 6344 39672 6372
rect 28902 6264 28908 6316
rect 28960 6264 28966 6316
rect 35986 6264 35992 6316
rect 36044 6304 36050 6316
rect 38856 6313 38884 6344
rect 39666 6332 39672 6344
rect 39724 6332 39730 6384
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 36044 6276 37841 6304
rect 36044 6264 36050 6276
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 38473 6307 38531 6313
rect 38473 6273 38485 6307
rect 38519 6273 38531 6307
rect 38473 6267 38531 6273
rect 38841 6307 38899 6313
rect 38841 6273 38853 6307
rect 38887 6273 38899 6307
rect 38841 6267 38899 6273
rect 39209 6307 39267 6313
rect 39209 6273 39221 6307
rect 39255 6273 39267 6307
rect 39209 6267 39267 6273
rect 34422 6196 34428 6248
rect 34480 6236 34486 6248
rect 38488 6236 38516 6267
rect 34480 6208 38516 6236
rect 34480 6196 34486 6208
rect 38562 6196 38568 6248
rect 38620 6236 38626 6248
rect 39224 6236 39252 6267
rect 38620 6208 39252 6236
rect 38620 6196 38626 6208
rect 38286 6168 38292 6180
rect 28736 6140 38292 6168
rect 27580 6128 27586 6140
rect 38286 6128 38292 6140
rect 38344 6128 38350 6180
rect 28350 6100 28356 6112
rect 27356 6072 28356 6100
rect 28350 6060 28356 6072
rect 28408 6060 28414 6112
rect 36446 6060 36452 6112
rect 36504 6100 36510 6112
rect 38470 6100 38476 6112
rect 36504 6072 38476 6100
rect 36504 6060 36510 6072
rect 38470 6060 38476 6072
rect 38528 6060 38534 6112
rect 38654 6060 38660 6112
rect 38712 6060 38718 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 2133 5899 2191 5905
rect 2133 5865 2145 5899
rect 2179 5896 2191 5899
rect 2314 5896 2320 5908
rect 2179 5868 2320 5896
rect 2179 5865 2191 5868
rect 2133 5859 2191 5865
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 8956 5868 9628 5896
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 6822 5828 6828 5840
rect 1627 5800 6828 5828
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 8386 5828 8392 5840
rect 7064 5800 8392 5828
rect 7064 5788 7070 5800
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 842 5720 848 5772
rect 900 5760 906 5772
rect 900 5732 1992 5760
rect 900 5720 906 5732
rect 198 5652 204 5704
rect 256 5692 262 5704
rect 1964 5701 1992 5732
rect 2498 5720 2504 5772
rect 2556 5760 2562 5772
rect 6914 5760 6920 5772
rect 2556 5732 6920 5760
rect 2556 5720 2562 5732
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 8956 5769 8984 5868
rect 9600 5828 9628 5868
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 9953 5899 10011 5905
rect 9953 5896 9965 5899
rect 9732 5868 9965 5896
rect 9732 5856 9738 5868
rect 9953 5865 9965 5868
rect 9999 5865 10011 5899
rect 9953 5859 10011 5865
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 12161 5899 12219 5905
rect 10744 5868 11836 5896
rect 10744 5856 10750 5868
rect 11054 5828 11060 5840
rect 9600 5800 11060 5828
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11146 5788 11152 5840
rect 11204 5788 11210 5840
rect 11808 5828 11836 5868
rect 12161 5865 12173 5899
rect 12207 5896 12219 5899
rect 14642 5896 14648 5908
rect 12207 5868 14648 5896
rect 12207 5865 12219 5868
rect 12161 5859 12219 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 20257 5899 20315 5905
rect 17236 5868 20208 5896
rect 17236 5828 17264 5868
rect 11808 5800 17264 5828
rect 17954 5788 17960 5840
rect 18012 5828 18018 5840
rect 18690 5828 18696 5840
rect 18012 5800 18696 5828
rect 18012 5788 18018 5800
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 20180 5828 20208 5868
rect 20257 5865 20269 5899
rect 20303 5896 20315 5899
rect 20346 5896 20352 5908
rect 20303 5868 20352 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 25222 5856 25228 5908
rect 25280 5896 25286 5908
rect 25280 5868 31754 5896
rect 25280 5856 25286 5868
rect 21910 5828 21916 5840
rect 20180 5800 21916 5828
rect 21910 5788 21916 5800
rect 21968 5788 21974 5840
rect 27065 5831 27123 5837
rect 27065 5797 27077 5831
rect 27111 5828 27123 5831
rect 28166 5828 28172 5840
rect 27111 5800 28172 5828
rect 27111 5797 27123 5800
rect 27065 5791 27123 5797
rect 28166 5788 28172 5800
rect 28224 5788 28230 5840
rect 31726 5828 31754 5868
rect 37826 5856 37832 5908
rect 37884 5896 37890 5908
rect 37921 5899 37979 5905
rect 37921 5896 37933 5899
rect 37884 5868 37933 5896
rect 37884 5856 37890 5868
rect 37921 5865 37933 5868
rect 37967 5865 37979 5899
rect 37921 5859 37979 5865
rect 38194 5856 38200 5908
rect 38252 5856 38258 5908
rect 39393 5899 39451 5905
rect 39393 5865 39405 5899
rect 39439 5896 39451 5899
rect 39574 5896 39580 5908
rect 39439 5868 39580 5896
rect 39439 5865 39451 5868
rect 39393 5859 39451 5865
rect 39574 5856 39580 5868
rect 39632 5856 39638 5908
rect 39025 5831 39083 5837
rect 31726 5800 38884 5828
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 7616 5732 8953 5760
rect 7616 5720 7622 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 10778 5760 10784 5772
rect 9732 5732 10784 5760
rect 9732 5720 9738 5732
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11164 5760 11192 5788
rect 10888 5732 11192 5760
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 256 5664 1409 5692
rect 256 5652 262 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 658 5584 664 5636
rect 716 5624 722 5636
rect 1688 5624 1716 5655
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 7742 5692 7748 5704
rect 3660 5664 7748 5692
rect 3660 5652 3666 5664
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8904 5664 9229 5692
rect 8904 5652 8910 5664
rect 9217 5661 9229 5664
rect 9263 5692 9275 5695
rect 10888 5692 10916 5732
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 12434 5760 12440 5772
rect 11940 5732 12440 5760
rect 11940 5720 11946 5732
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 16758 5760 16764 5772
rect 13096 5732 16764 5760
rect 9263 5664 10916 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 11256 5664 11437 5692
rect 11256 5636 11284 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 13096 5701 13124 5732
rect 16758 5720 16764 5732
rect 16816 5720 16822 5772
rect 19150 5760 19156 5772
rect 18524 5732 19156 5760
rect 13081 5695 13139 5701
rect 13081 5692 13093 5695
rect 11756 5664 13093 5692
rect 11756 5652 11762 5664
rect 13081 5661 13093 5664
rect 13127 5661 13139 5695
rect 13081 5655 13139 5661
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13228 5664 14105 5692
rect 13228 5652 13234 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 18524 5692 18552 5732
rect 19150 5720 19156 5732
rect 19208 5720 19214 5772
rect 20898 5760 20904 5772
rect 20364 5732 20904 5760
rect 14792 5664 18552 5692
rect 14792 5652 14798 5664
rect 18598 5652 18604 5704
rect 18656 5692 18662 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 18656 5664 19257 5692
rect 18656 5652 18662 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 20364 5701 20392 5732
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 24946 5720 24952 5772
rect 25004 5720 25010 5772
rect 29270 5720 29276 5772
rect 29328 5760 29334 5772
rect 29328 5732 38424 5760
rect 29328 5720 29334 5732
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 19576 5664 20361 5692
rect 19576 5652 19582 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 23382 5692 23388 5704
rect 20349 5655 20407 5661
rect 20456 5664 23388 5692
rect 716 5596 1716 5624
rect 716 5584 722 5596
rect 1762 5584 1768 5636
rect 1820 5624 1826 5636
rect 10778 5624 10784 5636
rect 1820 5596 10784 5624
rect 1820 5584 1826 5596
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 11238 5584 11244 5636
rect 11296 5584 11302 5636
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 13262 5624 13268 5636
rect 11388 5596 13268 5624
rect 11388 5584 11394 5596
rect 13262 5584 13268 5596
rect 13320 5624 13326 5636
rect 13633 5627 13691 5633
rect 13633 5624 13645 5627
rect 13320 5596 13645 5624
rect 13320 5584 13326 5596
rect 13633 5593 13645 5596
rect 13679 5593 13691 5627
rect 13633 5587 13691 5593
rect 13814 5584 13820 5636
rect 13872 5584 13878 5636
rect 15654 5624 15660 5636
rect 13924 5596 15660 5624
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 10410 5556 10416 5568
rect 1636 5528 10416 5556
rect 1636 5516 1642 5528
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11698 5556 11704 5568
rect 11204 5528 11704 5556
rect 11204 5516 11210 5528
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 13173 5559 13231 5565
rect 13173 5556 13185 5559
rect 12952 5528 13185 5556
rect 12952 5516 12958 5528
rect 13173 5525 13185 5528
rect 13219 5525 13231 5559
rect 13173 5519 13231 5525
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 13924 5556 13952 5596
rect 15654 5584 15660 5596
rect 15712 5584 15718 5636
rect 15746 5584 15752 5636
rect 15804 5624 15810 5636
rect 20456 5624 20484 5664
rect 23382 5652 23388 5664
rect 23440 5652 23446 5704
rect 25222 5652 25228 5704
rect 25280 5652 25286 5704
rect 26050 5652 26056 5704
rect 26108 5652 26114 5704
rect 26329 5695 26387 5701
rect 26329 5661 26341 5695
rect 26375 5692 26387 5695
rect 28258 5692 28264 5704
rect 26375 5664 28264 5692
rect 26375 5661 26387 5664
rect 26329 5655 26387 5661
rect 28258 5652 28264 5664
rect 28316 5652 28322 5704
rect 35618 5652 35624 5704
rect 35676 5692 35682 5704
rect 38396 5701 38424 5732
rect 38856 5701 38884 5800
rect 39025 5797 39037 5831
rect 39071 5828 39083 5831
rect 39942 5828 39948 5840
rect 39071 5800 39948 5828
rect 39071 5797 39083 5800
rect 39025 5791 39083 5797
rect 39942 5788 39948 5800
rect 40000 5788 40006 5840
rect 38105 5695 38163 5701
rect 38105 5692 38117 5695
rect 35676 5664 38117 5692
rect 35676 5652 35682 5664
rect 38105 5661 38117 5664
rect 38151 5661 38163 5695
rect 38105 5655 38163 5661
rect 38381 5695 38439 5701
rect 38381 5661 38393 5695
rect 38427 5661 38439 5695
rect 38381 5655 38439 5661
rect 38841 5695 38899 5701
rect 38841 5661 38853 5695
rect 38887 5661 38899 5695
rect 38841 5655 38899 5661
rect 39209 5695 39267 5701
rect 39209 5661 39221 5695
rect 39255 5661 39267 5695
rect 39209 5655 39267 5661
rect 15804 5596 20484 5624
rect 15804 5584 15810 5596
rect 21450 5584 21456 5636
rect 21508 5624 21514 5636
rect 24670 5624 24676 5636
rect 21508 5596 24676 5624
rect 21508 5584 21514 5596
rect 24670 5584 24676 5596
rect 24728 5584 24734 5636
rect 38654 5584 38660 5636
rect 38712 5624 38718 5636
rect 39224 5624 39252 5655
rect 38712 5596 39252 5624
rect 38712 5584 38718 5596
rect 13596 5528 13952 5556
rect 14277 5559 14335 5565
rect 13596 5516 13602 5528
rect 14277 5525 14289 5559
rect 14323 5556 14335 5559
rect 14642 5556 14648 5568
rect 14323 5528 14648 5556
rect 14323 5525 14335 5528
rect 14277 5519 14335 5525
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 16666 5556 16672 5568
rect 14792 5528 16672 5556
rect 14792 5516 14798 5528
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 20438 5556 20444 5568
rect 16816 5528 20444 5556
rect 16816 5516 16822 5528
rect 20438 5516 20444 5528
rect 20496 5516 20502 5568
rect 20530 5516 20536 5568
rect 20588 5516 20594 5568
rect 25961 5559 26019 5565
rect 25961 5525 25973 5559
rect 26007 5556 26019 5559
rect 26878 5556 26884 5568
rect 26007 5528 26884 5556
rect 26007 5525 26019 5528
rect 25961 5519 26019 5525
rect 26878 5516 26884 5528
rect 26936 5516 26942 5568
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5902 5352 5908 5364
rect 5767 5324 5908 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 13722 5352 13728 5364
rect 6880 5324 13728 5352
rect 6880 5312 6886 5324
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 20714 5352 20720 5364
rect 20496 5324 20720 5352
rect 20496 5312 20502 5324
rect 20714 5312 20720 5324
rect 20772 5352 20778 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20772 5324 20821 5352
rect 20772 5312 20778 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 20809 5315 20867 5321
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 28442 5352 28448 5364
rect 23164 5324 28448 5352
rect 23164 5312 23170 5324
rect 28442 5312 28448 5324
rect 28500 5312 28506 5364
rect 28718 5312 28724 5364
rect 28776 5352 28782 5364
rect 34790 5352 34796 5364
rect 28776 5324 34796 5352
rect 28776 5312 28782 5324
rect 34790 5312 34796 5324
rect 34848 5312 34854 5364
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 6638 5244 6644 5296
rect 6696 5284 6702 5296
rect 6696 5256 9674 5284
rect 6696 5244 6702 5256
rect 382 5176 388 5228
rect 440 5216 446 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 440 5188 1409 5216
rect 440 5176 446 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 5215 5188 5273 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 5810 5216 5816 5228
rect 5583 5188 5816 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 842 5108 848 5160
rect 900 5148 906 5160
rect 1688 5148 1716 5179
rect 5810 5176 5816 5188
rect 5868 5216 5874 5228
rect 7098 5216 7104 5228
rect 5868 5188 7104 5216
rect 5868 5176 5874 5188
rect 7098 5176 7104 5188
rect 7156 5216 7162 5228
rect 7558 5216 7564 5228
rect 7156 5188 7564 5216
rect 7156 5176 7162 5188
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 9646 5216 9674 5256
rect 11974 5244 11980 5296
rect 12032 5284 12038 5296
rect 19334 5284 19340 5296
rect 12032 5256 19340 5284
rect 12032 5244 12038 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 20901 5287 20959 5293
rect 20901 5253 20913 5287
rect 20947 5284 20959 5287
rect 21269 5287 21327 5293
rect 21269 5284 21281 5287
rect 20947 5256 21281 5284
rect 20947 5253 20959 5256
rect 20901 5247 20959 5253
rect 21269 5253 21281 5256
rect 21315 5253 21327 5287
rect 21269 5247 21327 5253
rect 21542 5244 21548 5296
rect 21600 5284 21606 5296
rect 25590 5284 25596 5296
rect 21600 5256 25596 5284
rect 21600 5244 21606 5256
rect 25590 5244 25596 5256
rect 25648 5284 25654 5296
rect 26050 5284 26056 5296
rect 25648 5256 26056 5284
rect 25648 5244 25654 5256
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 27338 5244 27344 5296
rect 27396 5284 27402 5296
rect 38930 5284 38936 5296
rect 27396 5256 38936 5284
rect 27396 5244 27402 5256
rect 38930 5244 38936 5256
rect 38988 5244 38994 5296
rect 12250 5216 12256 5228
rect 9646 5188 12256 5216
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 13538 5176 13544 5228
rect 13596 5216 13602 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 13596 5188 20729 5216
rect 13596 5176 13602 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 27430 5216 27436 5228
rect 20864 5188 27436 5216
rect 20864 5176 20870 5188
rect 27430 5176 27436 5188
rect 27488 5176 27494 5228
rect 28166 5176 28172 5228
rect 28224 5216 28230 5228
rect 28537 5219 28595 5225
rect 28537 5216 28549 5219
rect 28224 5188 28549 5216
rect 28224 5176 28230 5188
rect 28537 5185 28549 5188
rect 28583 5185 28595 5219
rect 28537 5179 28595 5185
rect 38838 5176 38844 5228
rect 38896 5176 38902 5228
rect 39209 5219 39267 5225
rect 39209 5185 39221 5219
rect 39255 5185 39267 5219
rect 39209 5179 39267 5185
rect 900 5120 1716 5148
rect 900 5108 906 5120
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 12342 5148 12348 5160
rect 5776 5120 12348 5148
rect 5776 5108 5782 5120
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 18046 5148 18052 5160
rect 12492 5120 18052 5148
rect 12492 5108 12498 5120
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 28074 5148 28080 5160
rect 18932 5120 28080 5148
rect 18932 5108 18938 5120
rect 28074 5108 28080 5120
rect 28132 5108 28138 5160
rect 28261 5151 28319 5157
rect 28261 5117 28273 5151
rect 28307 5117 28319 5151
rect 28261 5111 28319 5117
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5080 1639 5083
rect 5350 5080 5356 5092
rect 1627 5052 5356 5080
rect 1627 5049 1639 5052
rect 1581 5043 1639 5049
rect 5350 5040 5356 5052
rect 5408 5040 5414 5092
rect 5445 5083 5503 5089
rect 5445 5049 5457 5083
rect 5491 5080 5503 5083
rect 13078 5080 13084 5092
rect 5491 5052 13084 5080
rect 5491 5049 5503 5052
rect 5445 5043 5503 5049
rect 13078 5040 13084 5052
rect 13136 5040 13142 5092
rect 13170 5040 13176 5092
rect 13228 5080 13234 5092
rect 25498 5080 25504 5092
rect 13228 5052 25504 5080
rect 13228 5040 13234 5052
rect 25498 5040 25504 5052
rect 25556 5040 25562 5092
rect 27890 5040 27896 5092
rect 27948 5080 27954 5092
rect 28276 5080 28304 5111
rect 37274 5108 37280 5160
rect 37332 5148 37338 5160
rect 39224 5148 39252 5179
rect 37332 5120 39252 5148
rect 37332 5108 37338 5120
rect 27948 5052 28304 5080
rect 27948 5040 27954 5052
rect 1857 5015 1915 5021
rect 1857 4981 1869 5015
rect 1903 5012 1915 5015
rect 4798 5012 4804 5024
rect 1903 4984 4804 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5169 5015 5227 5021
rect 5169 5012 5181 5015
rect 4948 4984 5181 5012
rect 4948 4972 4954 4984
rect 5169 4981 5181 4984
rect 5215 5012 5227 5015
rect 5902 5012 5908 5024
rect 5215 4984 5908 5012
rect 5215 4981 5227 4984
rect 5169 4975 5227 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 15378 5012 15384 5024
rect 7064 4984 15384 5012
rect 7064 4972 7070 4984
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 21358 4972 21364 5024
rect 21416 4972 21422 5024
rect 28276 5012 28304 5052
rect 28902 5012 28908 5024
rect 28276 4984 28908 5012
rect 28902 4972 28908 4984
rect 28960 4972 28966 5024
rect 29270 4972 29276 5024
rect 29328 4972 29334 5024
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 4890 4768 4896 4820
rect 4948 4768 4954 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5132 4780 6224 4808
rect 5132 4768 5138 4780
rect 6196 4749 6224 4780
rect 6270 4768 6276 4820
rect 6328 4808 6334 4820
rect 10502 4808 10508 4820
rect 6328 4780 10508 4808
rect 6328 4768 6334 4780
rect 6181 4743 6239 4749
rect 6181 4709 6193 4743
rect 6227 4709 6239 4743
rect 6181 4703 6239 4709
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5810 4681 5816 4684
rect 5629 4675 5687 4681
rect 5629 4672 5641 4675
rect 5040 4644 5641 4672
rect 5040 4632 5046 4644
rect 5629 4641 5641 4644
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5788 4675 5816 4681
rect 5788 4641 5800 4675
rect 5788 4635 5816 4641
rect 5810 4632 5816 4635
rect 5868 4632 5874 4684
rect 6638 4632 6644 4684
rect 6696 4632 6702 4684
rect 6932 4681 6960 4780
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10612 4780 11468 4808
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4641 6975 4675
rect 6917 4635 6975 4641
rect 750 4564 756 4616
rect 808 4604 814 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 808 4576 1409 4604
rect 808 4564 814 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 2746 4576 4476 4604
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 1688 4536 1716 4567
rect 900 4508 1716 4536
rect 900 4496 906 4508
rect 1578 4428 1584 4480
rect 1636 4428 1642 4480
rect 1857 4471 1915 4477
rect 1857 4437 1869 4471
rect 1903 4468 1915 4471
rect 2746 4468 2774 4576
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 4338 4536 4344 4548
rect 4203 4508 4344 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 4448 4536 4476 4576
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6788 4576 6837 4604
rect 6788 4564 6794 4576
rect 6825 4573 6837 4576
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 4448 4508 5212 4536
rect 1903 4440 2774 4468
rect 1903 4437 1915 4440
rect 1857 4431 1915 4437
rect 4246 4428 4252 4480
rect 4304 4428 4310 4480
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 4985 4471 5043 4477
rect 4985 4468 4997 4471
rect 4948 4440 4997 4468
rect 4948 4428 4954 4440
rect 4985 4437 4997 4440
rect 5031 4437 5043 4471
rect 5184 4468 5212 4508
rect 6638 4496 6644 4548
rect 6696 4536 6702 4548
rect 6932 4536 6960 4635
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 10612 4672 10640 4780
rect 11440 4740 11468 4780
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 13170 4808 13176 4820
rect 11572 4780 13176 4808
rect 11572 4768 11578 4780
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 22278 4808 22284 4820
rect 21928 4780 22284 4808
rect 21450 4740 21456 4752
rect 11440 4712 21456 4740
rect 21450 4700 21456 4712
rect 21508 4700 21514 4752
rect 21928 4740 21956 4780
rect 22278 4768 22284 4780
rect 22336 4808 22342 4820
rect 23842 4808 23848 4820
rect 22336 4780 23848 4808
rect 22336 4768 22342 4780
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 30282 4808 30288 4820
rect 23952 4780 30288 4808
rect 21744 4712 21956 4740
rect 11103 4675 11161 4681
rect 11103 4672 11115 4675
rect 10284 4644 11115 4672
rect 10284 4632 10290 4644
rect 11103 4641 11115 4644
rect 11149 4641 11161 4675
rect 11103 4635 11161 4641
rect 11241 4675 11299 4681
rect 11241 4641 11253 4675
rect 11287 4672 11299 4675
rect 11422 4672 11428 4684
rect 11287 4644 11428 4672
rect 11287 4641 11299 4644
rect 11241 4635 11299 4641
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 11514 4632 11520 4684
rect 11572 4632 11578 4684
rect 11974 4632 11980 4684
rect 12032 4632 12038 4684
rect 12158 4632 12164 4684
rect 12216 4632 12222 4684
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 18509 4675 18567 4681
rect 18509 4672 18521 4675
rect 14792 4644 18521 4672
rect 14792 4632 14798 4644
rect 18509 4641 18521 4644
rect 18555 4672 18567 4675
rect 19058 4672 19064 4684
rect 18555 4644 19064 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 21637 4675 21695 4681
rect 21637 4641 21649 4675
rect 21683 4672 21695 4675
rect 21744 4672 21772 4712
rect 23290 4700 23296 4752
rect 23348 4740 23354 4752
rect 23952 4740 23980 4780
rect 30282 4768 30288 4780
rect 30340 4768 30346 4820
rect 39390 4768 39396 4820
rect 39448 4768 39454 4820
rect 23348 4712 23980 4740
rect 23348 4700 23354 4712
rect 29638 4700 29644 4752
rect 29696 4740 29702 4752
rect 29733 4743 29791 4749
rect 29733 4740 29745 4743
rect 29696 4712 29745 4740
rect 29696 4700 29702 4712
rect 29733 4709 29745 4712
rect 29779 4709 29791 4743
rect 29733 4703 29791 4709
rect 39025 4743 39083 4749
rect 39025 4709 39037 4743
rect 39071 4740 39083 4743
rect 39942 4740 39948 4752
rect 39071 4712 39948 4740
rect 39071 4709 39083 4712
rect 39025 4703 39083 4709
rect 39942 4700 39948 4712
rect 40000 4700 40006 4752
rect 21683 4644 21772 4672
rect 21683 4641 21695 4644
rect 21637 4635 21695 4641
rect 21818 4632 21824 4684
rect 21876 4632 21882 4684
rect 22186 4632 22192 4684
rect 22244 4672 22250 4684
rect 22281 4675 22339 4681
rect 22281 4672 22293 4675
rect 22244 4644 22293 4672
rect 22244 4632 22250 4644
rect 22281 4641 22293 4644
rect 22327 4641 22339 4675
rect 22281 4635 22339 4641
rect 22830 4632 22836 4684
rect 22888 4632 22894 4684
rect 7180 4597 7238 4603
rect 7180 4594 7192 4597
rect 7162 4563 7192 4594
rect 7226 4563 7238 4597
rect 10962 4564 10968 4616
rect 11020 4564 11026 4616
rect 14826 4564 14832 4616
rect 14884 4604 14890 4616
rect 16206 4604 16212 4616
rect 14884 4576 16212 4604
rect 14884 4564 14890 4576
rect 16206 4564 16212 4576
rect 16264 4604 16270 4616
rect 16669 4607 16727 4613
rect 16669 4604 16681 4607
rect 16264 4576 16681 4604
rect 16264 4564 16270 4576
rect 16669 4573 16681 4576
rect 16715 4573 16727 4607
rect 16669 4567 16727 4573
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 7162 4557 7238 4563
rect 6696 4508 6960 4536
rect 6696 4496 6702 4508
rect 7006 4496 7012 4548
rect 7064 4536 7070 4548
rect 7162 4536 7190 4557
rect 7064 4508 7190 4536
rect 7064 4496 7070 4508
rect 7466 4496 7472 4548
rect 7524 4536 7530 4548
rect 8202 4536 8208 4548
rect 7524 4508 8208 4536
rect 7524 4496 7530 4508
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 16850 4496 16856 4548
rect 16908 4496 16914 4548
rect 17862 4496 17868 4548
rect 17920 4536 17926 4548
rect 18248 4536 18276 4567
rect 18598 4564 18604 4616
rect 18656 4564 18662 4616
rect 22554 4564 22560 4616
rect 22612 4564 22618 4616
rect 22738 4613 22744 4616
rect 22695 4607 22744 4613
rect 22695 4573 22707 4607
rect 22741 4573 22744 4607
rect 22695 4567 22744 4573
rect 22738 4564 22744 4567
rect 22796 4564 22802 4616
rect 28994 4564 29000 4616
rect 29052 4564 29058 4616
rect 29086 4564 29092 4616
rect 29144 4604 29150 4616
rect 29273 4607 29331 4613
rect 29273 4604 29285 4607
rect 29144 4576 29285 4604
rect 29144 4564 29150 4576
rect 29273 4573 29285 4576
rect 29319 4573 29331 4607
rect 29273 4567 29331 4573
rect 29914 4564 29920 4616
rect 29972 4564 29978 4616
rect 37458 4564 37464 4616
rect 37516 4604 37522 4616
rect 38841 4607 38899 4613
rect 38841 4604 38853 4607
rect 37516 4576 38853 4604
rect 37516 4564 37522 4576
rect 38841 4573 38853 4576
rect 38887 4573 38899 4607
rect 38841 4567 38899 4573
rect 38930 4564 38936 4616
rect 38988 4604 38994 4616
rect 39209 4607 39267 4613
rect 39209 4604 39221 4607
rect 38988 4576 39221 4604
rect 38988 4564 38994 4576
rect 39209 4573 39221 4576
rect 39255 4573 39267 4607
rect 39209 4567 39267 4573
rect 21542 4536 21548 4548
rect 17920 4508 21548 4536
rect 17920 4496 17926 4508
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 23382 4496 23388 4548
rect 23440 4536 23446 4548
rect 30006 4536 30012 4548
rect 23440 4508 30012 4536
rect 23440 4496 23446 4508
rect 30006 4496 30012 4508
rect 30064 4496 30070 4548
rect 5718 4468 5724 4480
rect 5184 4440 5724 4468
rect 4985 4431 5043 4437
rect 5718 4428 5724 4440
rect 5776 4428 5782 4480
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 7484 4468 7512 4496
rect 6788 4440 7512 4468
rect 6788 4428 6794 4440
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 7892 4440 7941 4468
rect 7892 4428 7898 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 10318 4428 10324 4480
rect 10376 4428 10382 4480
rect 10410 4428 10416 4480
rect 10468 4468 10474 4480
rect 11974 4468 11980 4480
rect 10468 4440 11980 4468
rect 10468 4428 10474 4440
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 15378 4428 15384 4480
rect 15436 4468 15442 4480
rect 18322 4468 18328 4480
rect 15436 4440 18328 4468
rect 15436 4428 15442 4440
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 18782 4428 18788 4480
rect 18840 4428 18846 4480
rect 21818 4428 21824 4480
rect 21876 4468 21882 4480
rect 22462 4468 22468 4480
rect 21876 4440 22468 4468
rect 21876 4428 21882 4440
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 22554 4428 22560 4480
rect 22612 4468 22618 4480
rect 23400 4468 23428 4496
rect 22612 4440 23428 4468
rect 23477 4471 23535 4477
rect 22612 4428 22618 4440
rect 23477 4437 23489 4471
rect 23523 4468 23535 4471
rect 24578 4468 24584 4480
rect 23523 4440 24584 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 24578 4428 24584 4440
rect 24636 4428 24642 4480
rect 28258 4428 28264 4480
rect 28316 4428 28322 4480
rect 29546 4428 29552 4480
rect 29604 4468 29610 4480
rect 30650 4468 30656 4480
rect 29604 4440 30656 4468
rect 29604 4428 29610 4440
rect 30650 4428 30656 4440
rect 30708 4428 30714 4480
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 5074 4224 5080 4276
rect 5132 4224 5138 4276
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 7282 4264 7288 4276
rect 5960 4236 7288 4264
rect 5960 4224 5966 4236
rect 7282 4224 7288 4236
rect 7340 4264 7346 4276
rect 8297 4267 8355 4273
rect 8297 4264 8309 4267
rect 7340 4236 8309 4264
rect 7340 4224 7346 4236
rect 8297 4233 8309 4236
rect 8343 4233 8355 4267
rect 8297 4227 8355 4233
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 11020 4236 11529 4264
rect 11020 4224 11026 4236
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 12526 4264 12532 4276
rect 11517 4227 11575 4233
rect 11992 4236 12532 4264
rect 3786 4156 3792 4208
rect 3844 4156 3850 4208
rect 5184 4196 5212 4224
rect 4080 4168 5212 4196
rect 382 4088 388 4140
rect 440 4128 446 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 440 4100 1409 4128
rect 440 4088 446 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 842 4020 848 4072
rect 900 4060 906 4072
rect 1688 4060 1716 4091
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4080 4137 4108 4168
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 5537 4199 5595 4205
rect 5537 4196 5549 4199
rect 5408 4168 5549 4196
rect 5408 4156 5414 4168
rect 5537 4165 5549 4168
rect 5583 4165 5595 4199
rect 5537 4159 5595 4165
rect 10502 4156 10508 4208
rect 10560 4196 10566 4208
rect 11057 4199 11115 4205
rect 11057 4196 11069 4199
rect 10560 4168 11069 4196
rect 10560 4156 10566 4168
rect 11057 4165 11069 4168
rect 11103 4165 11115 4199
rect 11057 4159 11115 4165
rect 11241 4199 11299 4205
rect 11241 4165 11253 4199
rect 11287 4196 11299 4199
rect 11698 4196 11704 4208
rect 11287 4168 11704 4196
rect 11287 4165 11299 4168
rect 11241 4159 11299 4165
rect 4065 4131 4123 4137
rect 4065 4128 4077 4131
rect 4028 4100 4077 4128
rect 4028 4088 4034 4100
rect 4065 4097 4077 4100
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 4338 4088 4344 4140
rect 4396 4088 4402 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4948 4100 5181 4128
rect 4948 4088 4954 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 6227 4100 6377 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 7006 4088 7012 4140
rect 7064 4088 7070 4140
rect 7098 4088 7104 4140
rect 7156 4137 7162 4140
rect 7156 4131 7205 4137
rect 7156 4097 7159 4131
rect 7193 4097 7205 4131
rect 7156 4091 7205 4097
rect 7156 4088 7162 4091
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 8202 4088 8208 4140
rect 8260 4088 8266 4140
rect 9398 4088 9404 4140
rect 9456 4128 9462 4140
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9456 4100 9781 4128
rect 9456 4088 9462 4100
rect 9769 4097 9781 4100
rect 9815 4128 9827 4131
rect 11072 4128 11100 4159
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 11992 4128 12020 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 17678 4224 17684 4276
rect 17736 4264 17742 4276
rect 18598 4264 18604 4276
rect 17736 4236 18604 4264
rect 17736 4224 17742 4236
rect 18598 4224 18604 4236
rect 18656 4264 18662 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 18656 4236 19165 4264
rect 18656 4224 18662 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19153 4227 19211 4233
rect 21376 4236 23520 4264
rect 15105 4199 15163 4205
rect 15105 4196 15117 4199
rect 12360 4168 15117 4196
rect 12360 4140 12388 4168
rect 15105 4165 15117 4168
rect 15151 4196 15163 4199
rect 15151 4168 18276 4196
rect 15151 4165 15163 4168
rect 15105 4159 15163 4165
rect 12342 4138 12348 4140
rect 12268 4137 12348 4138
rect 9815 4100 10732 4128
rect 11072 4100 12020 4128
rect 12253 4131 12348 4137
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 900 4032 1716 4060
rect 900 4020 906 4032
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8021 4063 8079 4069
rect 8021 4060 8033 4063
rect 7708 4032 8033 4060
rect 7708 4020 7714 4032
rect 8021 4029 8033 4032
rect 8067 4029 8079 4063
rect 8021 4023 8079 4029
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 10502 4060 10508 4072
rect 8435 4032 10508 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 5353 3995 5411 4001
rect 1903 3964 4200 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 3694 3924 3700 3936
rect 1627 3896 3700 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4062 3924 4068 3936
rect 3927 3896 4068 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4172 3924 4200 3964
rect 5353 3961 5365 3995
rect 5399 3992 5411 3995
rect 5399 3964 5948 3992
rect 5399 3961 5411 3964
rect 5353 3955 5411 3961
rect 5534 3924 5540 3936
rect 4172 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5626 3884 5632 3936
rect 5684 3884 5690 3936
rect 5920 3924 5948 3964
rect 5994 3952 6000 4004
rect 6052 3952 6058 4004
rect 7561 3995 7619 4001
rect 7561 3961 7573 3995
rect 7607 3992 7619 3995
rect 9582 3992 9588 4004
rect 7607 3964 9588 3992
rect 7607 3961 7619 3964
rect 7561 3955 7619 3961
rect 9582 3952 9588 3964
rect 9640 3952 9646 4004
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10594 3992 10600 4004
rect 9999 3964 10600 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10704 3992 10732 4100
rect 12253 4097 12265 4131
rect 12299 4110 12348 4131
rect 12299 4097 12311 4110
rect 12253 4091 12311 4097
rect 12342 4088 12348 4110
rect 12400 4088 12406 4140
rect 12526 4088 12532 4140
rect 12584 4088 12590 4140
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 17037 4131 17095 4137
rect 17037 4128 17049 4131
rect 16264 4100 17049 4128
rect 16264 4088 16270 4100
rect 17037 4097 17049 4100
rect 17083 4097 17095 4131
rect 17037 4091 17095 4097
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 18248 4128 18276 4168
rect 19058 4156 19064 4208
rect 19116 4156 19122 4208
rect 18187 4100 18276 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18414 4088 18420 4140
rect 18472 4128 18478 4140
rect 21376 4128 21404 4236
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 21508 4168 22232 4196
rect 21508 4156 21514 4168
rect 18472 4100 21404 4128
rect 21821 4131 21879 4137
rect 18472 4088 18478 4100
rect 21821 4097 21833 4131
rect 21867 4128 21879 4131
rect 22002 4128 22008 4140
rect 21867 4100 22008 4128
rect 21867 4097 21879 4100
rect 21821 4091 21879 4097
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11422 4060 11428 4072
rect 10836 4032 11428 4060
rect 10836 4020 10842 4032
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 16485 4063 16543 4069
rect 16485 4029 16497 4063
rect 16531 4060 16543 4063
rect 16574 4060 16580 4072
rect 16531 4032 16580 4060
rect 16531 4029 16543 4032
rect 16485 4023 16543 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16758 4020 16764 4072
rect 16816 4020 16822 4072
rect 17862 4020 17868 4072
rect 17920 4020 17926 4072
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 20346 4060 20352 4072
rect 19852 4032 20352 4060
rect 19852 4020 19858 4032
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 21174 4020 21180 4072
rect 21232 4060 21238 4072
rect 21358 4060 21364 4072
rect 21232 4032 21364 4060
rect 21232 4020 21238 4032
rect 21358 4020 21364 4032
rect 21416 4060 21422 4072
rect 21836 4060 21864 4091
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22097 4132 22155 4137
rect 22204 4132 22232 4168
rect 22370 4156 22376 4208
rect 22428 4196 22434 4208
rect 22554 4196 22560 4208
rect 22428 4168 22560 4196
rect 22428 4156 22434 4168
rect 22554 4156 22560 4168
rect 22612 4196 22618 4208
rect 23290 4196 23296 4208
rect 22612 4168 23296 4196
rect 22612 4156 22618 4168
rect 23290 4156 23296 4168
rect 23348 4156 23354 4208
rect 22097 4131 22232 4132
rect 22097 4097 22109 4131
rect 22143 4104 22232 4131
rect 22143 4097 22155 4104
rect 22097 4091 22155 4097
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 23106 4128 23112 4140
rect 22796 4100 23112 4128
rect 22796 4088 22802 4100
rect 23106 4088 23112 4100
rect 23164 4088 23170 4140
rect 23382 4088 23388 4140
rect 23440 4088 23446 4140
rect 21416 4032 21864 4060
rect 23492 4060 23520 4236
rect 28350 4224 28356 4276
rect 28408 4264 28414 4276
rect 28408 4236 29960 4264
rect 28408 4224 28414 4236
rect 23842 4196 23848 4208
rect 23676 4168 23848 4196
rect 23566 4088 23572 4140
rect 23624 4128 23630 4140
rect 23676 4137 23704 4168
rect 23842 4156 23848 4168
rect 23900 4156 23906 4208
rect 27614 4196 27620 4208
rect 23952 4168 27620 4196
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23624 4100 23673 4128
rect 23624 4088 23630 4100
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 23661 4091 23719 4097
rect 23750 4088 23756 4140
rect 23808 4128 23814 4140
rect 23952 4128 23980 4168
rect 27614 4156 27620 4168
rect 27672 4156 27678 4208
rect 29932 4205 29960 4236
rect 30006 4224 30012 4276
rect 30064 4264 30070 4276
rect 30650 4264 30656 4276
rect 30064 4236 30656 4264
rect 30064 4224 30070 4236
rect 30650 4224 30656 4236
rect 30708 4224 30714 4276
rect 29549 4199 29607 4205
rect 29549 4196 29561 4199
rect 29196 4168 29561 4196
rect 23808 4100 23980 4128
rect 23808 4088 23814 4100
rect 24118 4088 24124 4140
rect 24176 4128 24182 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 24176 4100 24225 4128
rect 24176 4088 24182 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 27798 4128 27804 4140
rect 24213 4091 24271 4097
rect 24320 4100 27804 4128
rect 24320 4060 24348 4100
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 28626 4088 28632 4140
rect 28684 4088 28690 4140
rect 23492 4032 24348 4060
rect 21416 4020 21422 4032
rect 25130 4020 25136 4072
rect 25188 4060 25194 4072
rect 27433 4063 27491 4069
rect 25188 4032 27384 4060
rect 25188 4020 25194 4032
rect 10704 3964 11192 3992
rect 11164 3936 11192 3964
rect 15286 3952 15292 4004
rect 15344 3952 15350 4004
rect 15470 3952 15476 4004
rect 15528 3952 15534 4004
rect 18800 3964 19334 3992
rect 7190 3924 7196 3936
rect 5920 3896 7196 3924
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 11054 3924 11060 3936
rect 7340 3896 11060 3924
rect 7340 3884 7346 3896
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 15654 3924 15660 3936
rect 11204 3896 15660 3924
rect 11204 3884 11210 3896
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 17773 3927 17831 3933
rect 17773 3893 17785 3927
rect 17819 3924 17831 3927
rect 18800 3924 18828 3964
rect 17819 3896 18828 3924
rect 17819 3893 17831 3896
rect 17773 3887 17831 3893
rect 18874 3884 18880 3936
rect 18932 3884 18938 3936
rect 19306 3924 19334 3964
rect 20714 3952 20720 4004
rect 20772 3992 20778 4004
rect 21634 3992 21640 4004
rect 20772 3964 21640 3992
rect 20772 3952 20778 3964
rect 21634 3952 21640 3964
rect 21692 3952 21698 4004
rect 22925 3995 22983 4001
rect 22925 3992 22937 3995
rect 22480 3964 22937 3992
rect 21726 3924 21732 3936
rect 19306 3896 21732 3924
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22480 3924 22508 3964
rect 22925 3961 22937 3964
rect 22971 3961 22983 3995
rect 22925 3955 22983 3961
rect 23198 3952 23204 4004
rect 23256 3952 23262 4004
rect 23474 3952 23480 4004
rect 23532 3952 23538 4004
rect 23937 3995 23995 4001
rect 23937 3961 23949 3995
rect 23983 3992 23995 3995
rect 26234 3992 26240 4004
rect 23983 3964 26240 3992
rect 23983 3961 23995 3964
rect 23937 3955 23995 3961
rect 26234 3952 26240 3964
rect 26292 3952 26298 4004
rect 27356 3992 27384 4032
rect 27433 4029 27445 4063
rect 27479 4060 27491 4063
rect 27522 4060 27528 4072
rect 27479 4032 27528 4060
rect 27479 4029 27491 4032
rect 27433 4023 27491 4029
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 27617 4063 27675 4069
rect 27617 4029 27629 4063
rect 27663 4029 27675 4063
rect 27617 4023 27675 4029
rect 27632 3992 27660 4023
rect 28074 4020 28080 4072
rect 28132 4020 28138 4072
rect 28353 4063 28411 4069
rect 28353 4060 28365 4063
rect 28184 4032 28365 4060
rect 27356 3964 27660 3992
rect 27982 3952 27988 4004
rect 28040 3992 28046 4004
rect 28184 3992 28212 4032
rect 28353 4029 28365 4032
rect 28399 4029 28411 4063
rect 28353 4023 28411 4029
rect 28442 4020 28448 4072
rect 28500 4069 28506 4072
rect 28500 4063 28528 4069
rect 28516 4060 28528 4063
rect 29196 4060 29224 4168
rect 29549 4165 29561 4168
rect 29595 4165 29607 4199
rect 29549 4159 29607 4165
rect 29917 4199 29975 4205
rect 29917 4165 29929 4199
rect 29963 4165 29975 4199
rect 29917 4159 29975 4165
rect 30282 4156 30288 4208
rect 30340 4156 30346 4208
rect 29454 4088 29460 4140
rect 29512 4128 29518 4140
rect 29730 4128 29736 4140
rect 29512 4100 29736 4128
rect 29512 4088 29518 4100
rect 29730 4088 29736 4100
rect 29788 4128 29794 4140
rect 29825 4131 29883 4137
rect 29825 4128 29837 4131
rect 29788 4100 29837 4128
rect 29788 4088 29794 4100
rect 29825 4097 29837 4100
rect 29871 4097 29883 4131
rect 29825 4091 29883 4097
rect 38841 4131 38899 4137
rect 38841 4097 38853 4131
rect 38887 4128 38899 4131
rect 38887 4100 39160 4128
rect 38887 4097 38899 4100
rect 38841 4091 38899 4097
rect 28516 4032 29224 4060
rect 29368 4072 29420 4078
rect 28516 4029 28528 4032
rect 28500 4023 28528 4029
rect 28500 4020 28506 4023
rect 39132 4060 39160 4100
rect 39206 4088 39212 4140
rect 39264 4088 39270 4140
rect 40034 4060 40040 4072
rect 39132 4032 40040 4060
rect 40034 4020 40040 4032
rect 40092 4020 40098 4072
rect 29368 4014 29420 4020
rect 28040 3964 28212 3992
rect 39393 3995 39451 4001
rect 28040 3952 28046 3964
rect 39393 3961 39405 3995
rect 39439 3992 39451 3995
rect 39482 3992 39488 4004
rect 39439 3964 39488 3992
rect 39439 3961 39451 3964
rect 39393 3955 39451 3961
rect 39482 3952 39488 3964
rect 39540 3952 39546 4004
rect 22244 3896 22508 3924
rect 22244 3884 22250 3896
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 22833 3927 22891 3933
rect 22833 3924 22845 3927
rect 22796 3896 22845 3924
rect 22796 3884 22802 3896
rect 22833 3893 22845 3896
rect 22879 3893 22891 3927
rect 22833 3887 22891 3893
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 24029 3927 24087 3933
rect 24029 3924 24041 3927
rect 23716 3896 24041 3924
rect 23716 3884 23722 3896
rect 24029 3893 24041 3896
rect 24075 3893 24087 3927
rect 24029 3887 24087 3893
rect 26326 3884 26332 3936
rect 26384 3924 26390 3936
rect 28626 3924 28632 3936
rect 26384 3896 28632 3924
rect 26384 3884 26390 3896
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 29273 3927 29331 3933
rect 29273 3893 29285 3927
rect 29319 3924 29331 3927
rect 29546 3924 29552 3936
rect 29319 3896 29552 3924
rect 29319 3893 29331 3896
rect 29273 3887 29331 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 30834 3884 30840 3936
rect 30892 3884 30898 3936
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 3786 3720 3792 3732
rect 2179 3692 3792 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 4982 3680 4988 3732
rect 5040 3680 5046 3732
rect 6730 3720 6736 3732
rect 5644 3692 6736 3720
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 2406 3652 2412 3664
rect 1627 3624 2412 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 5534 3612 5540 3664
rect 5592 3612 5598 3664
rect 1026 3544 1032 3596
rect 1084 3584 1090 3596
rect 1084 3556 1992 3584
rect 1084 3544 1090 3556
rect 198 3476 204 3528
rect 256 3516 262 3528
rect 1964 3525 1992 3556
rect 3970 3544 3976 3596
rect 4028 3544 4034 3596
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5644 3593 5672 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 9490 3720 9496 3732
rect 7064 3692 9496 3720
rect 7064 3680 7070 3692
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9582 3680 9588 3732
rect 9640 3680 9646 3732
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9766 3720 9772 3732
rect 9723 3692 9772 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 12434 3720 12440 3732
rect 9876 3692 12440 3720
rect 6641 3655 6699 3661
rect 6641 3621 6653 3655
rect 6687 3652 6699 3655
rect 6914 3652 6920 3664
rect 6687 3624 6920 3652
rect 6687 3621 6699 3624
rect 6641 3615 6699 3621
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 7834 3612 7840 3664
rect 7892 3652 7898 3664
rect 7929 3655 7987 3661
rect 7929 3652 7941 3655
rect 7892 3624 7941 3652
rect 7892 3612 7898 3624
rect 7929 3621 7941 3624
rect 7975 3621 7987 3655
rect 9876 3652 9904 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 16574 3720 16580 3732
rect 13688 3692 16580 3720
rect 13688 3680 13694 3692
rect 10778 3652 10784 3664
rect 7929 3615 7987 3621
rect 9646 3624 9904 3652
rect 9968 3624 10784 3652
rect 7558 3593 7564 3596
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 5224 3556 5641 3584
rect 5224 3544 5230 3556
rect 5629 3553 5641 3556
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 7536 3587 7564 3593
rect 7536 3553 7548 3587
rect 7536 3547 7564 3553
rect 7558 3544 7564 3547
rect 7616 3544 7622 3596
rect 9646 3584 9674 3624
rect 9968 3584 9996 3624
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 12544 3624 14105 3652
rect 8496 3556 9674 3584
rect 9784 3556 9996 3584
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 256 3488 1409 3516
rect 256 3476 262 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 842 3408 848 3460
rect 900 3448 906 3460
rect 1688 3448 1716 3479
rect 3786 3476 3792 3528
rect 3844 3516 3850 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 3844 3488 4261 3516
rect 3844 3476 3850 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 4856 3488 5365 3516
rect 4856 3476 4862 3488
rect 5353 3485 5365 3488
rect 5399 3516 5411 3519
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5399 3512 5580 3516
rect 5736 3512 5917 3516
rect 5399 3488 5917 3512
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5552 3484 5764 3488
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 8496 3516 8524 3556
rect 9784 3528 9812 3556
rect 10226 3544 10232 3596
rect 10284 3544 10290 3596
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 12544 3584 12572 3624
rect 14093 3621 14105 3624
rect 14139 3621 14151 3655
rect 14093 3615 14151 3621
rect 15120 3593 15148 3692
rect 16574 3680 16580 3692
rect 16632 3720 16638 3732
rect 17678 3720 17684 3732
rect 16632 3692 17684 3720
rect 16632 3680 16638 3692
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 15562 3652 15568 3664
rect 15519 3624 15568 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 15562 3612 15568 3624
rect 15620 3612 15626 3664
rect 10919 3556 12572 3584
rect 15105 3587 15163 3593
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 15105 3553 15117 3587
rect 15151 3553 15163 3587
rect 16022 3584 16028 3596
rect 15105 3547 15163 3553
rect 15212 3556 16028 3584
rect 8444 3488 8524 3516
rect 8573 3519 8631 3525
rect 8444 3476 8450 3488
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9766 3516 9772 3528
rect 9447 3488 9772 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 900 3420 1716 3448
rect 8588 3448 8616 3479
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10244 3516 10272 3544
rect 9999 3488 10272 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 11330 3525 11336 3528
rect 11287 3519 11336 3525
rect 11287 3485 11299 3519
rect 11333 3485 11336 3519
rect 11287 3479 11336 3485
rect 11330 3476 11336 3479
rect 11388 3476 11394 3528
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3516 12127 3519
rect 12345 3519 12403 3525
rect 12345 3516 12357 3519
rect 12115 3488 12357 3516
rect 12115 3485 12127 3488
rect 12069 3479 12127 3485
rect 12345 3485 12357 3488
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 15212 3516 15240 3556
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 16684 3593 16712 3692
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 19061 3723 19119 3729
rect 17788 3692 18736 3720
rect 16669 3587 16727 3593
rect 16669 3553 16681 3587
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 17586 3544 17592 3596
rect 17644 3584 17650 3596
rect 17788 3584 17816 3692
rect 17957 3655 18015 3661
rect 17957 3621 17969 3655
rect 18003 3652 18015 3655
rect 18046 3652 18052 3664
rect 18003 3624 18052 3652
rect 18003 3621 18015 3624
rect 17957 3615 18015 3621
rect 18046 3612 18052 3624
rect 18104 3612 18110 3664
rect 18708 3652 18736 3692
rect 19061 3689 19073 3723
rect 19107 3720 19119 3723
rect 19107 3692 22094 3720
rect 19107 3689 19119 3692
rect 19061 3683 19119 3689
rect 20714 3652 20720 3664
rect 18708 3624 20720 3652
rect 20714 3612 20720 3624
rect 20772 3612 20778 3664
rect 22066 3596 22094 3692
rect 22848 3692 23888 3720
rect 17644 3556 17816 3584
rect 17644 3544 17650 3556
rect 21174 3544 21180 3596
rect 21232 3544 21238 3596
rect 22066 3556 22100 3596
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 22278 3544 22284 3596
rect 22336 3544 22342 3596
rect 22465 3587 22523 3593
rect 22465 3553 22477 3587
rect 22511 3584 22523 3587
rect 22554 3584 22560 3596
rect 22511 3556 22560 3584
rect 22511 3553 22523 3556
rect 22465 3547 22523 3553
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 22848 3584 22876 3692
rect 22664 3556 22876 3584
rect 22925 3587 22983 3593
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 14936 3488 15240 3516
rect 15580 3488 16405 3516
rect 10042 3448 10048 3460
rect 8588 3420 10048 3448
rect 900 3408 906 3420
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 14936 3448 14964 3488
rect 12032 3420 14964 3448
rect 12032 3408 12038 3420
rect 15286 3408 15292 3460
rect 15344 3408 15350 3460
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 6638 3380 6644 3392
rect 1903 3352 6644 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 7466 3380 7472 3392
rect 6779 3352 7472 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9582 3380 9588 3392
rect 8904 3352 9588 3380
rect 8904 3340 8910 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 10134 3340 10140 3392
rect 10192 3340 10198 3392
rect 12158 3340 12164 3392
rect 12216 3340 12222 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 15580 3380 15608 3488
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 13780 3352 15608 3380
rect 13780 3340 13786 3352
rect 15654 3340 15660 3392
rect 15712 3340 15718 3392
rect 16408 3380 16436 3479
rect 16942 3476 16948 3528
rect 17000 3476 17006 3528
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 17184 3488 17233 3516
rect 17184 3476 17190 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18049 3519 18107 3525
rect 17920 3512 18000 3516
rect 18049 3512 18061 3519
rect 17920 3488 18061 3512
rect 17920 3476 17926 3488
rect 17972 3485 18061 3488
rect 18095 3485 18107 3519
rect 17972 3484 18107 3485
rect 18049 3479 18107 3484
rect 18322 3476 18328 3528
rect 18380 3476 18386 3528
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 21910 3516 21916 3528
rect 21499 3488 21916 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22664 3516 22692 3556
rect 22925 3553 22937 3587
rect 22971 3584 22983 3587
rect 23014 3584 23020 3596
rect 22971 3556 23020 3584
rect 22971 3553 22983 3556
rect 22925 3547 22983 3553
rect 23014 3544 23020 3556
rect 23072 3544 23078 3596
rect 23290 3544 23296 3596
rect 23348 3593 23354 3596
rect 23348 3587 23376 3593
rect 23364 3553 23376 3587
rect 23348 3547 23376 3553
rect 23477 3587 23535 3593
rect 23477 3553 23489 3587
rect 23523 3584 23535 3587
rect 23860 3584 23888 3692
rect 24118 3680 24124 3732
rect 24176 3680 24182 3732
rect 24394 3680 24400 3732
rect 24452 3680 24458 3732
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 27249 3723 27307 3729
rect 27249 3720 27261 3723
rect 25924 3692 27261 3720
rect 25924 3680 25930 3692
rect 27249 3689 27261 3692
rect 27295 3689 27307 3723
rect 29365 3723 29423 3729
rect 27249 3683 27307 3689
rect 27816 3692 29132 3720
rect 25774 3612 25780 3664
rect 25832 3652 25838 3664
rect 25832 3624 27752 3652
rect 25832 3612 25838 3624
rect 27724 3593 27752 3624
rect 23523 3556 23888 3584
rect 27709 3587 27767 3593
rect 23523 3553 23535 3556
rect 23477 3547 23535 3553
rect 27709 3553 27721 3587
rect 27755 3553 27767 3587
rect 27709 3547 27767 3553
rect 23348 3544 23354 3547
rect 22204 3488 22692 3516
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 21542 3448 21548 3460
rect 18196 3420 21548 3448
rect 18196 3408 18202 3420
rect 21542 3408 21548 3420
rect 21600 3408 21606 3460
rect 17770 3380 17776 3392
rect 16408 3352 17776 3380
rect 17770 3340 17776 3352
rect 17828 3380 17834 3392
rect 21450 3380 21456 3392
rect 17828 3352 21456 3380
rect 17828 3340 17834 3352
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 21634 3340 21640 3392
rect 21692 3380 21698 3392
rect 22094 3380 22100 3392
rect 21692 3352 22100 3380
rect 21692 3340 21698 3352
rect 22094 3340 22100 3352
rect 22152 3340 22158 3392
rect 22204 3389 22232 3488
rect 23198 3476 23204 3528
rect 23256 3476 23262 3528
rect 24578 3476 24584 3528
rect 24636 3476 24642 3528
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 27430 3516 27436 3528
rect 26476 3488 27436 3516
rect 26476 3476 26482 3488
rect 27430 3476 27436 3488
rect 27488 3476 27494 3528
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27816 3516 27844 3692
rect 27982 3612 27988 3664
rect 28040 3612 28046 3664
rect 28169 3655 28227 3661
rect 28169 3621 28181 3655
rect 28215 3652 28227 3655
rect 28258 3652 28264 3664
rect 28215 3624 28264 3652
rect 28215 3621 28227 3624
rect 28169 3615 28227 3621
rect 28258 3612 28264 3624
rect 28316 3612 28322 3664
rect 29104 3652 29132 3692
rect 29365 3689 29377 3723
rect 29411 3720 29423 3723
rect 29914 3720 29920 3732
rect 29411 3692 29920 3720
rect 29411 3689 29423 3692
rect 29365 3683 29423 3689
rect 29914 3680 29920 3692
rect 29972 3680 29978 3732
rect 30009 3723 30067 3729
rect 30009 3689 30021 3723
rect 30055 3720 30067 3723
rect 30190 3720 30196 3732
rect 30055 3692 30196 3720
rect 30055 3689 30067 3692
rect 30009 3683 30067 3689
rect 30190 3680 30196 3692
rect 30248 3680 30254 3732
rect 30282 3680 30288 3732
rect 30340 3680 30346 3732
rect 32858 3680 32864 3732
rect 32916 3720 32922 3732
rect 32953 3723 33011 3729
rect 32953 3720 32965 3723
rect 32916 3692 32965 3720
rect 32916 3680 32922 3692
rect 32953 3689 32965 3692
rect 32999 3689 33011 3723
rect 32953 3683 33011 3689
rect 33229 3723 33287 3729
rect 33229 3689 33241 3723
rect 33275 3720 33287 3723
rect 33686 3720 33692 3732
rect 33275 3692 33692 3720
rect 33275 3689 33287 3692
rect 33229 3683 33287 3689
rect 33686 3680 33692 3692
rect 33744 3680 33750 3732
rect 33781 3723 33839 3729
rect 33781 3689 33793 3723
rect 33827 3720 33839 3723
rect 34054 3720 34060 3732
rect 33827 3692 34060 3720
rect 33827 3689 33839 3692
rect 33781 3683 33839 3689
rect 34054 3680 34060 3692
rect 34112 3680 34118 3732
rect 34333 3723 34391 3729
rect 34333 3689 34345 3723
rect 34379 3720 34391 3723
rect 35802 3720 35808 3732
rect 34379 3692 35808 3720
rect 34379 3689 34391 3692
rect 34333 3683 34391 3689
rect 35802 3680 35808 3692
rect 35860 3680 35866 3732
rect 37461 3723 37519 3729
rect 37461 3720 37473 3723
rect 36464 3692 37473 3720
rect 29454 3652 29460 3664
rect 29104 3624 29460 3652
rect 29454 3612 29460 3624
rect 29512 3612 29518 3664
rect 29638 3612 29644 3664
rect 29696 3652 29702 3664
rect 30834 3652 30840 3664
rect 29696 3624 30840 3652
rect 29696 3612 29702 3624
rect 30834 3612 30840 3624
rect 30892 3612 30898 3664
rect 31662 3612 31668 3664
rect 31720 3652 31726 3664
rect 33413 3655 33471 3661
rect 33413 3652 33425 3655
rect 31720 3624 33425 3652
rect 31720 3612 31726 3624
rect 33413 3621 33425 3624
rect 33459 3621 33471 3655
rect 33413 3615 33471 3621
rect 35342 3612 35348 3664
rect 35400 3652 35406 3664
rect 36464 3652 36492 3692
rect 37461 3689 37473 3692
rect 37507 3689 37519 3723
rect 37461 3683 37519 3689
rect 37642 3680 37648 3732
rect 37700 3720 37706 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 37700 3692 38117 3720
rect 37700 3680 37706 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 39390 3680 39396 3732
rect 39448 3680 39454 3732
rect 35400 3624 36492 3652
rect 35400 3612 35406 3624
rect 36998 3612 37004 3664
rect 37056 3652 37062 3664
rect 38657 3655 38715 3661
rect 38657 3652 38669 3655
rect 37056 3624 38669 3652
rect 37056 3612 37062 3624
rect 38657 3621 38669 3624
rect 38703 3621 38715 3655
rect 38657 3615 38715 3621
rect 39025 3655 39083 3661
rect 39025 3621 39037 3655
rect 39071 3652 39083 3655
rect 39942 3652 39948 3664
rect 39071 3624 39948 3652
rect 39071 3621 39083 3624
rect 39025 3615 39083 3621
rect 39942 3612 39948 3624
rect 40000 3612 40006 3664
rect 28000 3584 28028 3612
rect 28442 3584 28448 3596
rect 28000 3556 28448 3584
rect 28442 3544 28448 3556
rect 28500 3544 28506 3596
rect 28534 3544 28540 3596
rect 28592 3593 28598 3596
rect 28592 3587 28620 3593
rect 28608 3553 28620 3587
rect 28592 3547 28620 3553
rect 28721 3587 28779 3593
rect 28721 3553 28733 3587
rect 28767 3584 28779 3587
rect 29270 3584 29276 3596
rect 28767 3556 29276 3584
rect 28767 3553 28779 3556
rect 28721 3547 28779 3553
rect 28592 3544 28598 3547
rect 29270 3544 29276 3556
rect 29328 3544 29334 3596
rect 29380 3556 39252 3584
rect 27580 3488 27844 3516
rect 27580 3476 27586 3488
rect 22189 3383 22247 3389
rect 22189 3349 22201 3383
rect 22235 3349 22247 3383
rect 22189 3343 22247 3349
rect 22278 3340 22284 3392
rect 22336 3380 22342 3392
rect 29380 3380 29408 3556
rect 29546 3476 29552 3528
rect 29604 3516 29610 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29604 3488 29745 3516
rect 29604 3476 29610 3488
rect 29733 3485 29745 3488
rect 29779 3485 29791 3519
rect 29733 3479 29791 3485
rect 29822 3476 29828 3528
rect 29880 3516 29886 3528
rect 30469 3519 30527 3525
rect 30469 3516 30481 3519
rect 29880 3488 30481 3516
rect 29880 3476 29886 3488
rect 30469 3485 30481 3488
rect 30515 3485 30527 3519
rect 30469 3479 30527 3485
rect 30558 3476 30564 3528
rect 30616 3476 30622 3528
rect 31570 3476 31576 3528
rect 31628 3516 31634 3528
rect 32585 3519 32643 3525
rect 32585 3516 32597 3519
rect 31628 3488 32597 3516
rect 31628 3476 31634 3488
rect 32585 3485 32597 3488
rect 32631 3516 32643 3519
rect 32769 3519 32827 3525
rect 32769 3516 32781 3519
rect 32631 3488 32781 3516
rect 32631 3485 32643 3488
rect 32585 3479 32643 3485
rect 32769 3485 32781 3488
rect 32815 3485 32827 3519
rect 32769 3479 32827 3485
rect 32858 3476 32864 3528
rect 32916 3516 32922 3528
rect 33045 3519 33103 3525
rect 33045 3516 33057 3519
rect 32916 3488 33057 3516
rect 32916 3476 32922 3488
rect 33045 3485 33057 3488
rect 33091 3485 33103 3519
rect 33045 3479 33103 3485
rect 33505 3519 33563 3525
rect 33505 3485 33517 3519
rect 33551 3516 33563 3519
rect 33597 3519 33655 3525
rect 33597 3516 33609 3519
rect 33551 3488 33609 3516
rect 33551 3485 33563 3488
rect 33505 3479 33563 3485
rect 33597 3485 33609 3488
rect 33643 3485 33655 3519
rect 33597 3479 33655 3485
rect 33870 3476 33876 3528
rect 33928 3476 33934 3528
rect 34146 3476 34152 3528
rect 34204 3476 34210 3528
rect 35158 3476 35164 3528
rect 35216 3516 35222 3528
rect 35526 3516 35532 3528
rect 35216 3488 35532 3516
rect 35216 3476 35222 3488
rect 35526 3476 35532 3488
rect 35584 3476 35590 3528
rect 35710 3476 35716 3528
rect 35768 3516 35774 3528
rect 37185 3519 37243 3525
rect 37185 3516 37197 3519
rect 35768 3488 37197 3516
rect 35768 3476 35774 3488
rect 37185 3485 37197 3488
rect 37231 3485 37243 3519
rect 37185 3479 37243 3485
rect 37369 3519 37427 3525
rect 37369 3485 37381 3519
rect 37415 3516 37427 3519
rect 37645 3519 37703 3525
rect 37645 3516 37657 3519
rect 37415 3488 37657 3516
rect 37415 3485 37427 3488
rect 37369 3479 37427 3485
rect 37645 3485 37657 3488
rect 37691 3485 37703 3519
rect 37645 3479 37703 3485
rect 38013 3519 38071 3525
rect 38013 3485 38025 3519
rect 38059 3516 38071 3519
rect 38289 3519 38347 3525
rect 38289 3516 38301 3519
rect 38059 3488 38301 3516
rect 38059 3485 38071 3488
rect 38013 3479 38071 3485
rect 38289 3485 38301 3488
rect 38335 3485 38347 3519
rect 38289 3479 38347 3485
rect 38565 3519 38623 3525
rect 38565 3485 38577 3519
rect 38611 3516 38623 3519
rect 38657 3519 38715 3525
rect 38657 3516 38669 3519
rect 38611 3488 38669 3516
rect 38611 3485 38623 3488
rect 38565 3479 38623 3485
rect 38657 3485 38669 3488
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 38838 3476 38844 3528
rect 38896 3476 38902 3528
rect 39224 3525 39252 3556
rect 39209 3519 39267 3525
rect 39209 3485 39221 3519
rect 39255 3485 39267 3519
rect 39209 3479 39267 3485
rect 30006 3408 30012 3460
rect 30064 3448 30070 3460
rect 30101 3451 30159 3457
rect 30101 3448 30113 3451
rect 30064 3420 30113 3448
rect 30064 3408 30070 3420
rect 30101 3417 30113 3420
rect 30147 3417 30159 3451
rect 36538 3448 36544 3460
rect 30101 3411 30159 3417
rect 31726 3420 36544 3448
rect 22336 3352 29408 3380
rect 29641 3383 29699 3389
rect 22336 3340 22342 3352
rect 29641 3349 29653 3383
rect 29687 3380 29699 3383
rect 29914 3380 29920 3392
rect 29687 3352 29920 3380
rect 29687 3349 29699 3352
rect 29641 3343 29699 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 30745 3383 30803 3389
rect 30745 3349 30757 3383
rect 30791 3380 30803 3383
rect 31726 3380 31754 3420
rect 36538 3408 36544 3420
rect 36596 3408 36602 3460
rect 36814 3408 36820 3460
rect 36872 3448 36878 3460
rect 36872 3420 38424 3448
rect 36872 3408 36878 3420
rect 30791 3352 31754 3380
rect 34057 3383 34115 3389
rect 30791 3349 30803 3352
rect 30745 3343 30803 3349
rect 34057 3349 34069 3383
rect 34103 3380 34115 3383
rect 35434 3380 35440 3392
rect 34103 3352 35440 3380
rect 34103 3349 34115 3352
rect 34057 3343 34115 3349
rect 35434 3340 35440 3352
rect 35492 3340 35498 3392
rect 35526 3340 35532 3392
rect 35584 3380 35590 3392
rect 37001 3383 37059 3389
rect 37001 3380 37013 3383
rect 35584 3352 37013 3380
rect 35584 3340 35590 3352
rect 37001 3349 37013 3352
rect 37047 3349 37059 3383
rect 37001 3343 37059 3349
rect 37090 3340 37096 3392
rect 37148 3380 37154 3392
rect 37277 3383 37335 3389
rect 37277 3380 37289 3383
rect 37148 3352 37289 3380
rect 37148 3340 37154 3352
rect 37277 3349 37289 3352
rect 37323 3349 37335 3383
rect 37277 3343 37335 3349
rect 37642 3340 37648 3392
rect 37700 3380 37706 3392
rect 38396 3389 38424 3420
rect 37921 3383 37979 3389
rect 37921 3380 37933 3383
rect 37700 3352 37933 3380
rect 37700 3340 37706 3352
rect 37921 3349 37933 3352
rect 37967 3349 37979 3383
rect 37921 3343 37979 3349
rect 38381 3383 38439 3389
rect 38381 3349 38393 3383
rect 38427 3349 38439 3383
rect 38381 3343 38439 3349
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 4338 3176 4344 3188
rect 2547 3148 4344 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 6178 3136 6184 3188
rect 6236 3136 6242 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6595 3148 6684 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 3878 3068 3884 3120
rect 3936 3108 3942 3120
rect 6656 3108 6684 3148
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7432 3148 7757 3176
rect 7432 3136 7438 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 7929 3179 7987 3185
rect 7929 3176 7941 3179
rect 7892 3148 7941 3176
rect 7892 3136 7898 3148
rect 7929 3145 7941 3148
rect 7975 3145 7987 3179
rect 7929 3139 7987 3145
rect 8389 3179 8447 3185
rect 8389 3145 8401 3179
rect 8435 3176 8447 3179
rect 9858 3176 9864 3188
rect 8435 3148 9864 3176
rect 8435 3145 8447 3148
rect 8389 3139 8447 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11514 3136 11520 3188
rect 11572 3136 11578 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 11900 3148 16681 3176
rect 6822 3108 6828 3120
rect 3936 3080 6316 3108
rect 6656 3080 6828 3108
rect 3936 3068 3942 3080
rect 1210 3000 1216 3052
rect 1268 3040 1274 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 1268 3012 2329 3040
rect 1268 3000 1274 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 750 2932 756 2984
rect 808 2972 814 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 808 2944 1409 2972
rect 808 2932 814 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2498 2972 2504 2984
rect 1719 2944 2504 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2498 2932 2504 2944
rect 2556 2932 2562 2984
rect 382 2864 388 2916
rect 440 2904 446 2916
rect 2608 2904 2636 3003
rect 5166 3000 5172 3052
rect 5224 3000 5230 3052
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5408 3012 5457 3040
rect 5408 3000 5414 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 6288 2972 6316 3080
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 8478 3108 8484 3120
rect 7024 3080 8484 3108
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 7024 3049 7052 3080
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 11900 3108 11928 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 17402 3136 17408 3188
rect 17460 3176 17466 3188
rect 17460 3148 19334 3176
rect 17460 3136 17466 3148
rect 11480 3080 11928 3108
rect 11480 3068 11486 3080
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 15289 3111 15347 3117
rect 15289 3108 15301 3111
rect 12216 3080 15301 3108
rect 12216 3068 12222 3080
rect 15289 3077 15301 3080
rect 15335 3108 15347 3111
rect 19306 3108 19334 3148
rect 21634 3136 21640 3188
rect 21692 3136 21698 3188
rect 28261 3179 28319 3185
rect 22388 3148 23520 3176
rect 22388 3108 22416 3148
rect 15335 3080 18368 3108
rect 19306 3080 22416 3108
rect 15335 3077 15347 3080
rect 15289 3071 15347 3077
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6656 3012 7021 3040
rect 6656 2972 6684 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8386 3040 8392 3052
rect 8159 3012 8392 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 11974 3040 11980 3052
rect 10100 3012 11980 3040
rect 10100 3000 10106 3012
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12250 3000 12256 3052
rect 12308 3040 12314 3052
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 12308 3012 15669 3040
rect 12308 3000 12314 3012
rect 15657 3009 15669 3012
rect 15703 3040 15715 3043
rect 15703 3012 15976 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 6288 2944 6684 2972
rect 6730 2932 6736 2984
rect 6788 2932 6794 2984
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8260 2944 9045 2972
rect 8260 2932 8266 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9192 2975 9250 2981
rect 9192 2941 9204 2975
rect 9238 2972 9250 2975
rect 9238 2944 9536 2972
rect 9238 2941 9250 2944
rect 9192 2935 9250 2941
rect 440 2876 2636 2904
rect 440 2864 446 2876
rect 2774 2864 2780 2916
rect 2832 2864 2838 2916
rect 9508 2904 9536 2944
rect 9582 2932 9588 2984
rect 9640 2932 9646 2984
rect 10226 2932 10232 2984
rect 10284 2932 10290 2984
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 10560 2944 11468 2972
rect 10560 2932 10566 2944
rect 9766 2904 9772 2916
rect 9508 2876 9772 2904
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 6638 2796 6644 2848
rect 6696 2836 6702 2848
rect 9306 2836 9312 2848
rect 6696 2808 9312 2836
rect 6696 2796 6702 2808
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 11440 2836 11468 2944
rect 12526 2932 12532 2984
rect 12584 2932 12590 2984
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 15746 2972 15752 2984
rect 13780 2944 15752 2972
rect 13780 2932 13786 2944
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 15838 2932 15844 2984
rect 15896 2932 15902 2984
rect 15948 2972 15976 3012
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 17310 3040 17316 3052
rect 16080 3012 17316 3040
rect 16080 3000 16086 3012
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17402 3000 17408 3052
rect 17460 3000 17466 3052
rect 17678 3000 17684 3052
rect 17736 3000 17742 3052
rect 17770 3000 17776 3052
rect 17828 3000 17834 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18340 3049 18368 3080
rect 22462 3068 22468 3120
rect 22520 3068 22526 3120
rect 22830 3068 22836 3120
rect 22888 3068 22894 3120
rect 22922 3068 22928 3120
rect 22980 3108 22986 3120
rect 23201 3111 23259 3117
rect 23201 3108 23213 3111
rect 22980 3080 23213 3108
rect 22980 3068 22986 3080
rect 23201 3077 23213 3080
rect 23247 3077 23259 3111
rect 23201 3071 23259 3077
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17920 3012 18061 3040
rect 17920 3000 17926 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 21910 3000 21916 3052
rect 21968 3000 21974 3052
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 23293 3043 23351 3049
rect 23293 3040 23305 3043
rect 23164 3012 23305 3040
rect 23164 3000 23170 3012
rect 23293 3009 23305 3012
rect 23339 3009 23351 3043
rect 23492 3040 23520 3148
rect 28261 3145 28273 3179
rect 28307 3176 28319 3179
rect 28350 3176 28356 3188
rect 28307 3148 28356 3176
rect 28307 3145 28319 3148
rect 28261 3139 28319 3145
rect 28350 3136 28356 3148
rect 28408 3136 28414 3188
rect 28442 3136 28448 3188
rect 28500 3176 28506 3188
rect 30742 3176 30748 3188
rect 28500 3148 30748 3176
rect 28500 3136 28506 3148
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 36262 3136 36268 3188
rect 36320 3176 36326 3188
rect 37921 3179 37979 3185
rect 37921 3176 37933 3179
rect 36320 3148 37933 3176
rect 36320 3136 36326 3148
rect 37921 3145 37933 3148
rect 37967 3145 37979 3179
rect 37921 3139 37979 3145
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 23566 3068 23572 3120
rect 23624 3068 23630 3120
rect 27706 3068 27712 3120
rect 27764 3108 27770 3120
rect 37458 3108 37464 3120
rect 27764 3080 37464 3108
rect 27764 3068 27770 3080
rect 37458 3068 37464 3080
rect 37516 3068 37522 3120
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23492 3012 23857 3040
rect 23293 3003 23351 3009
rect 23845 3009 23857 3012
rect 23891 3040 23903 3043
rect 27525 3043 27583 3049
rect 27525 3040 27537 3043
rect 23891 3012 27537 3040
rect 23891 3009 23903 3012
rect 23845 3003 23903 3009
rect 27525 3009 27537 3012
rect 27571 3009 27583 3043
rect 27525 3003 27583 3009
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 28629 3043 28687 3049
rect 28629 3040 28641 3043
rect 27672 3012 28641 3040
rect 27672 3000 27678 3012
rect 28629 3009 28641 3012
rect 28675 3009 28687 3043
rect 28629 3003 28687 3009
rect 28994 3000 29000 3052
rect 29052 3040 29058 3052
rect 29454 3040 29460 3052
rect 29052 3012 29460 3040
rect 29052 3000 29058 3012
rect 29454 3000 29460 3012
rect 29512 3000 29518 3052
rect 29546 3000 29552 3052
rect 29604 3040 29610 3052
rect 32858 3040 32864 3052
rect 29604 3012 32864 3040
rect 29604 3000 29610 3012
rect 32858 3000 32864 3012
rect 32916 3000 32922 3052
rect 37734 3000 37740 3052
rect 37792 3000 37798 3052
rect 37826 3000 37832 3052
rect 37884 3040 37890 3052
rect 38289 3043 38347 3049
rect 38289 3040 38301 3043
rect 37884 3012 38301 3040
rect 37884 3000 37890 3012
rect 38289 3009 38301 3012
rect 38335 3009 38347 3043
rect 38289 3003 38347 3009
rect 38746 3000 38752 3052
rect 38804 3040 38810 3052
rect 38841 3043 38899 3049
rect 38841 3040 38853 3043
rect 38804 3012 38853 3040
rect 38804 3000 38810 3012
rect 38841 3009 38853 3012
rect 38887 3009 38899 3043
rect 38841 3003 38899 3009
rect 38930 3000 38936 3052
rect 38988 3040 38994 3052
rect 39209 3043 39267 3049
rect 39209 3040 39221 3043
rect 38988 3012 39221 3040
rect 38988 3000 38994 3012
rect 39209 3009 39221 3012
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 17034 2972 17040 2984
rect 15948 2944 17040 2972
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 22370 2972 22376 2984
rect 18708 2944 22376 2972
rect 15304 2876 15516 2904
rect 15304 2836 15332 2876
rect 11440 2808 15332 2836
rect 15378 2796 15384 2848
rect 15436 2796 15442 2848
rect 15488 2836 15516 2876
rect 15562 2864 15568 2916
rect 15620 2904 15626 2916
rect 16482 2904 16488 2916
rect 15620 2876 16488 2904
rect 15620 2864 15626 2876
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 17604 2876 18092 2904
rect 17604 2836 17632 2876
rect 15488 2808 17632 2836
rect 17954 2796 17960 2848
rect 18012 2796 18018 2848
rect 18064 2836 18092 2876
rect 18708 2836 18736 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 22738 2932 22744 2984
rect 22796 2932 22802 2984
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 27249 2975 27307 2981
rect 27249 2972 27261 2975
rect 25648 2944 27261 2972
rect 25648 2932 25654 2944
rect 27249 2941 27261 2944
rect 27295 2941 27307 2975
rect 27249 2935 27307 2941
rect 19061 2907 19119 2913
rect 19061 2873 19073 2907
rect 19107 2904 19119 2907
rect 20898 2904 20904 2916
rect 19107 2876 20904 2904
rect 19107 2873 19119 2876
rect 19061 2867 19119 2873
rect 20898 2864 20904 2876
rect 20956 2864 20962 2916
rect 22097 2907 22155 2913
rect 22097 2873 22109 2907
rect 22143 2904 22155 2907
rect 24029 2907 24087 2913
rect 22143 2876 22416 2904
rect 22143 2873 22155 2876
rect 22097 2867 22155 2873
rect 22388 2848 22416 2876
rect 24029 2873 24041 2907
rect 24075 2904 24087 2907
rect 26510 2904 26516 2916
rect 24075 2876 26516 2904
rect 24075 2873 24087 2876
rect 24029 2867 24087 2873
rect 26510 2864 26516 2876
rect 26568 2864 26574 2916
rect 18064 2808 18736 2836
rect 22186 2796 22192 2848
rect 22244 2836 22250 2848
rect 22281 2839 22339 2845
rect 22281 2836 22293 2839
rect 22244 2808 22293 2836
rect 22244 2796 22250 2808
rect 22281 2805 22293 2808
rect 22327 2805 22339 2839
rect 22281 2799 22339 2805
rect 22370 2796 22376 2848
rect 22428 2796 22434 2848
rect 27264 2836 27292 2935
rect 27890 2932 27896 2984
rect 27948 2972 27954 2984
rect 28353 2975 28411 2981
rect 28353 2972 28365 2975
rect 27948 2944 28365 2972
rect 27948 2932 27954 2944
rect 28353 2941 28365 2944
rect 28399 2941 28411 2975
rect 28353 2935 28411 2941
rect 27908 2836 27936 2932
rect 29362 2864 29368 2916
rect 29420 2864 29426 2916
rect 30558 2904 30564 2916
rect 29564 2876 30564 2904
rect 27264 2808 27936 2836
rect 28166 2796 28172 2848
rect 28224 2836 28230 2848
rect 29564 2836 29592 2876
rect 30558 2864 30564 2876
rect 30616 2864 30622 2916
rect 28224 2808 29592 2836
rect 29641 2839 29699 2845
rect 28224 2796 28230 2808
rect 29641 2805 29653 2839
rect 29687 2836 29699 2839
rect 33134 2836 33140 2848
rect 29687 2808 33140 2836
rect 29687 2805 29699 2808
rect 29641 2799 29699 2805
rect 33134 2796 33140 2808
rect 33192 2796 33198 2848
rect 38470 2796 38476 2848
rect 38528 2796 38534 2848
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2632 2559 2635
rect 2547 2604 6914 2632
rect 2547 2601 2559 2604
rect 2501 2595 2559 2601
rect 1118 2524 1124 2576
rect 1176 2564 1182 2576
rect 3053 2567 3111 2573
rect 3053 2564 3065 2567
rect 1176 2536 3065 2564
rect 1176 2524 1182 2536
rect 3053 2533 3065 2536
rect 3099 2533 3111 2567
rect 6886 2564 6914 2604
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 14182 2632 14188 2644
rect 7064 2604 14188 2632
rect 7064 2592 7070 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 14550 2632 14556 2644
rect 14332 2604 14556 2632
rect 14332 2592 14338 2604
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 14700 2604 39252 2632
rect 14700 2592 14706 2604
rect 6886 2536 16574 2564
rect 3053 2527 3111 2533
rect 16546 2496 16574 2536
rect 23014 2524 23020 2576
rect 23072 2524 23078 2576
rect 18230 2496 18236 2508
rect 4264 2468 11100 2496
rect 16546 2468 18236 2496
rect 198 2388 204 2440
rect 256 2428 262 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 256 2400 1409 2428
rect 256 2388 262 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2332 2360 2360 2391
rect 2866 2388 2872 2440
rect 2924 2388 2930 2440
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 4264 2437 4292 2468
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2397 4307 2431
rect 4249 2391 4307 2397
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5675 2400 6914 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 1268 2332 2360 2360
rect 6886 2360 6914 2400
rect 7006 2388 7012 2440
rect 7064 2388 7070 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7524 2400 8125 2428
rect 7524 2388 7530 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 9766 2428 9772 2440
rect 9447 2400 9772 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 8312 2360 8340 2388
rect 6886 2332 8340 2360
rect 11072 2360 11100 2468
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 22002 2456 22008 2508
rect 22060 2456 22066 2508
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 33192 2468 38884 2496
rect 33192 2456 33198 2468
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 19518 2428 19524 2440
rect 11195 2400 19524 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 22281 2431 22339 2437
rect 22281 2397 22293 2431
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 22186 2360 22192 2372
rect 11072 2332 22192 2360
rect 1268 2320 1274 2332
rect 22186 2320 22192 2332
rect 22244 2320 22250 2372
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 2685 2295 2743 2301
rect 2685 2292 2697 2295
rect 2648 2264 2697 2292
rect 2648 2252 2654 2264
rect 2685 2261 2697 2264
rect 2731 2261 2743 2295
rect 2685 2255 2743 2261
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5316 2264 5457 2292
rect 5316 2252 5322 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6825 2295 6883 2301
rect 6825 2292 6837 2295
rect 6696 2264 6837 2292
rect 6696 2252 6702 2264
rect 6825 2261 6837 2264
rect 6871 2261 6883 2295
rect 6825 2255 6883 2261
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 8076 2264 8309 2292
rect 8076 2252 8082 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 9585 2295 9643 2301
rect 9585 2292 9597 2295
rect 9456 2264 9597 2292
rect 9456 2252 9462 2264
rect 9585 2261 9597 2264
rect 9631 2261 9643 2295
rect 9585 2255 9643 2261
rect 10778 2252 10784 2304
rect 10836 2292 10842 2304
rect 10965 2295 11023 2301
rect 10965 2292 10977 2295
rect 10836 2264 10977 2292
rect 10836 2252 10842 2264
rect 10965 2261 10977 2264
rect 11011 2261 11023 2295
rect 10965 2255 11023 2261
rect 21450 2252 21456 2304
rect 21508 2292 21514 2304
rect 22296 2292 22324 2391
rect 22370 2388 22376 2440
rect 22428 2428 22434 2440
rect 27706 2428 27712 2440
rect 22428 2400 27712 2428
rect 22428 2388 22434 2400
rect 27706 2388 27712 2400
rect 27764 2388 27770 2440
rect 28442 2388 28448 2440
rect 28500 2428 28506 2440
rect 28537 2431 28595 2437
rect 28537 2428 28549 2431
rect 28500 2400 28549 2428
rect 28500 2388 28506 2400
rect 28537 2397 28549 2400
rect 28583 2397 28595 2431
rect 28537 2391 28595 2397
rect 36538 2388 36544 2440
rect 36596 2428 36602 2440
rect 37737 2431 37795 2437
rect 37737 2428 37749 2431
rect 36596 2400 37749 2428
rect 36596 2388 36602 2400
rect 37737 2397 37749 2400
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 38102 2388 38108 2440
rect 38160 2388 38166 2440
rect 38470 2388 38476 2440
rect 38528 2388 38534 2440
rect 38856 2437 38884 2468
rect 39224 2437 39252 2604
rect 39390 2592 39396 2644
rect 39448 2592 39454 2644
rect 38841 2431 38899 2437
rect 38841 2397 38853 2431
rect 38887 2397 38899 2431
rect 38841 2391 38899 2397
rect 39209 2431 39267 2437
rect 39209 2397 39221 2431
rect 39255 2397 39267 2431
rect 39209 2391 39267 2397
rect 25958 2320 25964 2372
rect 26016 2360 26022 2372
rect 34146 2360 34152 2372
rect 26016 2332 34152 2360
rect 26016 2320 26022 2332
rect 34146 2320 34152 2332
rect 34204 2320 34210 2372
rect 21508 2264 22324 2292
rect 21508 2252 21514 2264
rect 28350 2252 28356 2304
rect 28408 2252 28414 2304
rect 37918 2252 37924 2304
rect 37976 2252 37982 2304
rect 38286 2252 38292 2304
rect 38344 2252 38350 2304
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39025 2295 39083 2301
rect 39025 2261 39037 2295
rect 39071 2292 39083 2295
rect 39942 2292 39948 2304
rect 39071 2264 39948 2292
rect 39071 2261 39083 2264
rect 39025 2255 39083 2261
rect 39942 2252 39948 2264
rect 40000 2252 40006 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 10318 2088 10324 2100
rect 2924 2060 10324 2088
rect 2924 2048 2930 2060
rect 10318 2048 10324 2060
rect 10376 2048 10382 2100
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 28350 2088 28356 2100
rect 14608 2060 28356 2088
rect 14608 2048 14614 2060
rect 28350 2048 28356 2060
rect 28408 2048 28414 2100
rect 19058 1980 19064 2032
rect 19116 2020 19122 2032
rect 31662 2020 31668 2032
rect 19116 1992 31668 2020
rect 19116 1980 19122 1992
rect 31662 1980 31668 1992
rect 31720 1980 31726 2032
rect 1670 1912 1676 1964
rect 1728 1952 1734 1964
rect 29454 1952 29460 1964
rect 1728 1924 29460 1952
rect 1728 1912 1734 1924
rect 29454 1912 29460 1924
rect 29512 1912 29518 1964
rect 38470 1952 38476 1964
rect 33704 1924 38476 1952
rect 18506 1844 18512 1896
rect 18564 1884 18570 1896
rect 33704 1884 33732 1924
rect 38470 1912 38476 1924
rect 38528 1912 38534 1964
rect 18564 1856 33732 1884
rect 18564 1844 18570 1856
rect 18690 1776 18696 1828
rect 18748 1816 18754 1828
rect 38102 1816 38108 1828
rect 18748 1788 38108 1816
rect 18748 1776 18754 1788
rect 38102 1776 38108 1788
rect 38160 1776 38166 1828
rect 9766 1708 9772 1760
rect 9824 1748 9830 1760
rect 29638 1748 29644 1760
rect 9824 1720 29644 1748
rect 9824 1708 9830 1720
rect 29638 1708 29644 1720
rect 29696 1708 29702 1760
rect 5718 1640 5724 1692
rect 5776 1680 5782 1692
rect 21450 1680 21456 1692
rect 5776 1652 21456 1680
rect 5776 1640 5782 1652
rect 21450 1640 21456 1652
rect 21508 1640 21514 1692
rect 4246 1300 4252 1352
rect 4304 1340 4310 1352
rect 38746 1340 38752 1352
rect 4304 1312 38752 1340
rect 4304 1300 4310 1312
rect 38746 1300 38752 1312
rect 38804 1300 38810 1352
rect 2498 1232 2504 1284
rect 2556 1272 2562 1284
rect 28166 1272 28172 1284
rect 2556 1244 28172 1272
rect 2556 1232 2562 1244
rect 28166 1232 28172 1244
rect 28224 1232 28230 1284
rect 13814 1164 13820 1216
rect 13872 1204 13878 1216
rect 38838 1204 38844 1216
rect 13872 1176 38844 1204
rect 13872 1164 13878 1176
rect 38838 1164 38844 1176
rect 38896 1164 38902 1216
rect 1578 1096 1584 1148
rect 1636 1136 1642 1148
rect 21818 1136 21824 1148
rect 1636 1108 21824 1136
rect 1636 1096 1642 1108
rect 21818 1096 21824 1108
rect 21876 1096 21882 1148
rect 12250 8 12256 60
rect 12308 48 12314 60
rect 37734 48 37740 60
rect 12308 20 37740 48
rect 12308 8 12314 20
rect 37734 8 37740 20
rect 37792 8 37798 60
<< via1 >>
rect 26976 11160 27028 11212
rect 37372 11160 37424 11212
rect 27252 11092 27304 11144
rect 37556 11092 37608 11144
rect 26700 11024 26752 11076
rect 35992 11024 36044 11076
rect 25872 10956 25924 11008
rect 34612 10956 34664 11008
rect 19432 10344 19484 10396
rect 24124 10344 24176 10396
rect 9956 10276 10008 10328
rect 5540 10208 5592 10260
rect 24400 10208 24452 10260
rect 36544 10208 36596 10260
rect 10784 10140 10836 10192
rect 26884 10140 26936 10192
rect 7840 10072 7892 10124
rect 23572 10072 23624 10124
rect 8116 10004 8168 10056
rect 28724 10004 28776 10056
rect 6736 9936 6788 9988
rect 19432 9936 19484 9988
rect 24124 9936 24176 9988
rect 29644 9936 29696 9988
rect 9496 9868 9548 9920
rect 19340 9868 19392 9920
rect 19892 9868 19944 9920
rect 34336 9868 34388 9920
rect 10048 9800 10100 9852
rect 9680 9732 9732 9784
rect 18880 9732 18932 9784
rect 35624 9800 35676 9852
rect 8392 9664 8444 9716
rect 37096 9664 37148 9716
rect 7472 9596 7524 9648
rect 17224 9596 17276 9648
rect 37464 9596 37516 9648
rect 38384 9596 38436 9648
rect 10876 9460 10928 9512
rect 4712 9392 4764 9444
rect 12716 9460 12768 9512
rect 23480 9460 23532 9512
rect 19892 9392 19944 9444
rect 15752 9324 15804 9376
rect 12532 9256 12584 9308
rect 21640 9324 21692 9376
rect 16304 9256 16356 9308
rect 32128 9256 32180 9308
rect 7288 9188 7340 9240
rect 17040 9188 17092 9240
rect 17868 9188 17920 9240
rect 18788 9188 18840 9240
rect 28816 9188 28868 9240
rect 15568 9120 15620 9172
rect 17224 9120 17276 9172
rect 29092 9120 29144 9172
rect 8300 9052 8352 9104
rect 9772 9052 9824 9104
rect 10324 9052 10376 9104
rect 4528 8984 4580 9036
rect 11428 8984 11480 9036
rect 14648 9052 14700 9104
rect 23204 9052 23256 9104
rect 24124 9052 24176 9104
rect 29552 9052 29604 9104
rect 35256 9052 35308 9104
rect 36268 9052 36320 9104
rect 17776 8984 17828 9036
rect 18604 8984 18656 9036
rect 27252 8984 27304 9036
rect 27528 8984 27580 9036
rect 36452 8984 36504 9036
rect 5908 8916 5960 8968
rect 11060 8916 11112 8968
rect 18512 8916 18564 8968
rect 24124 8916 24176 8968
rect 27436 8916 27488 8968
rect 29828 8916 29880 8968
rect 31576 8916 31628 8968
rect 38844 8916 38896 8968
rect 3608 8848 3660 8900
rect 20812 8848 20864 8900
rect 5080 8780 5132 8832
rect 8576 8780 8628 8832
rect 13268 8780 13320 8832
rect 16396 8780 16448 8832
rect 16580 8780 16632 8832
rect 38568 8848 38620 8900
rect 33048 8780 33100 8832
rect 33508 8780 33560 8832
rect 34520 8780 34572 8832
rect 37280 8780 37332 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 3516 8576 3568 8628
rect 4620 8576 4672 8628
rect 5448 8576 5500 8628
rect 5724 8576 5776 8628
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7564 8576 7616 8628
rect 7932 8576 7984 8628
rect 8484 8576 8536 8628
rect 8852 8576 8904 8628
rect 9588 8576 9640 8628
rect 9864 8576 9916 8628
rect 10048 8619 10100 8628
rect 10048 8585 10057 8619
rect 10057 8585 10091 8619
rect 10091 8585 10100 8619
rect 10048 8576 10100 8585
rect 10692 8576 10744 8628
rect 10968 8576 11020 8628
rect 11520 8576 11572 8628
rect 12072 8576 12124 8628
rect 12348 8576 12400 8628
rect 12900 8576 12952 8628
rect 13176 8576 13228 8628
rect 13728 8576 13780 8628
rect 14556 8576 14608 8628
rect 14924 8576 14976 8628
rect 15384 8576 15436 8628
rect 15660 8576 15712 8628
rect 16212 8576 16264 8628
rect 16488 8576 16540 8628
rect 16764 8576 16816 8628
rect 17316 8576 17368 8628
rect 17868 8576 17920 8628
rect 18512 8619 18564 8628
rect 18512 8585 18521 8619
rect 18521 8585 18555 8619
rect 18555 8585 18564 8619
rect 18512 8576 18564 8585
rect 19156 8576 19208 8628
rect 19340 8576 19392 8628
rect 20260 8576 20312 8628
rect 20628 8576 20680 8628
rect 756 8440 808 8492
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 8300 8508 8352 8560
rect 10324 8508 10376 8560
rect 3516 8440 3568 8492
rect 4528 8440 4580 8492
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 5540 8440 5592 8492
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7288 8440 7340 8492
rect 7748 8440 7800 8492
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 8116 8440 8168 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 9496 8440 9548 8492
rect 9588 8440 9640 8492
rect 12532 8508 12584 8560
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 3792 8304 3844 8356
rect 4344 8304 4396 8356
rect 9680 8372 9732 8424
rect 12716 8440 12768 8492
rect 14740 8508 14792 8560
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 7380 8304 7432 8356
rect 7840 8304 7892 8356
rect 13084 8372 13136 8424
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 18788 8508 18840 8560
rect 14924 8372 14976 8424
rect 14004 8304 14056 8356
rect 14648 8304 14700 8356
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16120 8440 16172 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18420 8440 18472 8492
rect 18696 8440 18748 8492
rect 18972 8440 19024 8492
rect 19248 8464 19300 8516
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 19800 8440 19852 8492
rect 20168 8440 20220 8492
rect 20444 8440 20496 8492
rect 20812 8508 20864 8560
rect 21824 8576 21876 8628
rect 22008 8576 22060 8628
rect 21732 8508 21784 8560
rect 20904 8440 20956 8492
rect 21364 8440 21416 8492
rect 21456 8440 21508 8492
rect 22560 8576 22612 8628
rect 22284 8508 22336 8560
rect 23112 8576 23164 8628
rect 22836 8508 22888 8560
rect 23664 8576 23716 8628
rect 23388 8508 23440 8560
rect 23940 8440 23992 8492
rect 24584 8576 24636 8628
rect 30380 8576 30432 8628
rect 32128 8619 32180 8628
rect 32128 8585 32137 8619
rect 32137 8585 32171 8619
rect 32171 8585 32180 8619
rect 32128 8576 32180 8585
rect 32496 8576 32548 8628
rect 32864 8576 32916 8628
rect 33508 8619 33560 8628
rect 33508 8585 33517 8619
rect 33517 8585 33551 8619
rect 33551 8585 33560 8619
rect 33508 8576 33560 8585
rect 33600 8576 33652 8628
rect 25504 8508 25556 8560
rect 24768 8440 24820 8492
rect 25412 8440 25464 8492
rect 27804 8440 27856 8492
rect 28080 8440 28132 8492
rect 29092 8551 29144 8560
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 29184 8508 29236 8560
rect 31392 8508 31444 8560
rect 33876 8508 33928 8560
rect 34888 8576 34940 8628
rect 35808 8576 35860 8628
rect 36912 8576 36964 8628
rect 38384 8576 38436 8628
rect 39580 8576 39632 8628
rect 28632 8440 28684 8492
rect 30288 8440 30340 8492
rect 31116 8440 31168 8492
rect 18696 8304 18748 8356
rect 19248 8372 19300 8424
rect 20352 8304 20404 8356
rect 5172 8236 5224 8288
rect 8392 8236 8444 8288
rect 10048 8236 10100 8288
rect 17224 8236 17276 8288
rect 18788 8279 18840 8288
rect 18788 8245 18797 8279
rect 18797 8245 18831 8279
rect 18831 8245 18840 8279
rect 18788 8236 18840 8245
rect 19432 8236 19484 8288
rect 19800 8279 19852 8288
rect 19800 8245 19809 8279
rect 19809 8245 19843 8279
rect 19843 8245 19852 8279
rect 19800 8236 19852 8245
rect 19892 8279 19944 8288
rect 19892 8245 19901 8279
rect 19901 8245 19935 8279
rect 19935 8245 19944 8279
rect 19892 8236 19944 8245
rect 21548 8372 21600 8424
rect 20812 8304 20864 8356
rect 20996 8347 21048 8356
rect 20996 8313 21005 8347
rect 21005 8313 21039 8347
rect 21039 8313 21048 8347
rect 20996 8304 21048 8313
rect 21456 8347 21508 8356
rect 21456 8313 21465 8347
rect 21465 8313 21499 8347
rect 21499 8313 21508 8347
rect 21456 8304 21508 8313
rect 21732 8304 21784 8356
rect 24676 8415 24728 8424
rect 24676 8381 24685 8415
rect 24685 8381 24719 8415
rect 24719 8381 24728 8415
rect 24676 8372 24728 8381
rect 24860 8372 24912 8424
rect 26516 8372 26568 8424
rect 25688 8304 25740 8356
rect 27528 8304 27580 8356
rect 28540 8372 28592 8424
rect 21364 8236 21416 8288
rect 22284 8279 22336 8288
rect 22284 8245 22293 8279
rect 22293 8245 22327 8279
rect 22327 8245 22336 8279
rect 22284 8236 22336 8245
rect 22376 8279 22428 8288
rect 22376 8245 22385 8279
rect 22385 8245 22419 8279
rect 22419 8245 22428 8279
rect 22376 8236 22428 8245
rect 22836 8279 22888 8288
rect 22836 8245 22845 8279
rect 22845 8245 22879 8279
rect 22879 8245 22888 8279
rect 22836 8236 22888 8245
rect 22928 8279 22980 8288
rect 22928 8245 22937 8279
rect 22937 8245 22971 8279
rect 22971 8245 22980 8279
rect 22928 8236 22980 8245
rect 23020 8236 23072 8288
rect 23848 8236 23900 8288
rect 24124 8236 24176 8288
rect 29092 8236 29144 8288
rect 29368 8304 29420 8356
rect 30932 8372 30984 8424
rect 32680 8440 32732 8492
rect 32864 8372 32916 8424
rect 33692 8483 33744 8492
rect 33692 8449 33701 8483
rect 33701 8449 33735 8483
rect 33735 8449 33744 8483
rect 33692 8440 33744 8449
rect 34060 8483 34112 8492
rect 34060 8449 34069 8483
rect 34069 8449 34103 8483
rect 34103 8449 34112 8483
rect 34060 8440 34112 8449
rect 35164 8440 35216 8492
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 35072 8372 35124 8424
rect 37004 8440 37056 8492
rect 37280 8483 37332 8492
rect 37280 8449 37289 8483
rect 37289 8449 37323 8483
rect 37323 8449 37332 8483
rect 37280 8440 37332 8449
rect 37832 8440 37884 8492
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 38384 8483 38436 8492
rect 38384 8449 38393 8483
rect 38393 8449 38427 8483
rect 38427 8449 38436 8483
rect 38384 8440 38436 8449
rect 38844 8483 38896 8492
rect 38844 8449 38853 8483
rect 38853 8449 38887 8483
rect 38887 8449 38896 8483
rect 38844 8440 38896 8449
rect 39212 8483 39264 8492
rect 39212 8449 39221 8483
rect 39221 8449 39255 8483
rect 39255 8449 39264 8483
rect 39212 8440 39264 8449
rect 33416 8304 33468 8356
rect 34152 8304 34204 8356
rect 37648 8372 37700 8424
rect 36268 8347 36320 8356
rect 36268 8313 36277 8347
rect 36277 8313 36311 8347
rect 36311 8313 36320 8347
rect 36268 8304 36320 8313
rect 36360 8304 36412 8356
rect 34704 8236 34756 8288
rect 37188 8304 37240 8356
rect 39396 8347 39448 8356
rect 39396 8313 39405 8347
rect 39405 8313 39439 8347
rect 39439 8313 39448 8347
rect 39396 8304 39448 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 4068 8032 4120 8084
rect 4896 8032 4948 8084
rect 6000 8032 6052 8084
rect 6552 8032 6604 8084
rect 7104 8032 7156 8084
rect 8300 8032 8352 8084
rect 8760 8032 8812 8084
rect 9404 8032 9456 8084
rect 10140 8032 10192 8084
rect 10416 8032 10468 8084
rect 11244 8032 11296 8084
rect 11796 8032 11848 8084
rect 12624 8032 12676 8084
rect 13452 8032 13504 8084
rect 13728 8032 13780 8084
rect 14188 8032 14240 8084
rect 14280 8032 14332 8084
rect 14832 8032 14884 8084
rect 15844 8032 15896 8084
rect 15936 8032 15988 8084
rect 17592 8032 17644 8084
rect 18696 8032 18748 8084
rect 20260 8032 20312 8084
rect 23112 8032 23164 8084
rect 6368 7964 6420 8016
rect 7932 7964 7984 8016
rect 572 7896 624 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1676 7871 1728 7880
rect 1676 7837 1685 7871
rect 1685 7837 1719 7871
rect 1719 7837 1728 7871
rect 1676 7828 1728 7837
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 2872 7828 2924 7880
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 940 7760 992 7812
rect 6184 7896 6236 7948
rect 6000 7828 6052 7880
rect 7380 7896 7432 7948
rect 8668 7896 8720 7948
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 9680 7896 9732 7948
rect 10876 7896 10928 7948
rect 14096 8007 14148 8016
rect 14096 7973 14105 8007
rect 14105 7973 14139 8007
rect 14139 7973 14148 8007
rect 14096 7964 14148 7973
rect 14464 7964 14516 8016
rect 8208 7760 8260 7812
rect 9956 7828 10008 7880
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 3884 7692 3936 7744
rect 8852 7692 8904 7744
rect 9772 7692 9824 7744
rect 10232 7692 10284 7744
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 14096 7828 14148 7880
rect 14280 7871 14332 7880
rect 14280 7837 14299 7871
rect 14299 7837 14332 7871
rect 14280 7828 14332 7837
rect 14740 7896 14792 7948
rect 13544 7692 13596 7744
rect 13636 7692 13688 7744
rect 17224 7964 17276 8016
rect 21916 7964 21968 8016
rect 16212 7896 16264 7948
rect 17960 7828 18012 7880
rect 18236 7828 18288 7880
rect 19984 7896 20036 7948
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 15384 7692 15436 7744
rect 16212 7692 16264 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18052 7692 18104 7744
rect 20260 7760 20312 7812
rect 23112 7896 23164 7948
rect 29092 8032 29144 8084
rect 32312 8032 32364 8084
rect 34428 8032 34480 8084
rect 35532 8032 35584 8084
rect 36084 8032 36136 8084
rect 36636 8032 36688 8084
rect 37740 8032 37792 8084
rect 38292 8032 38344 8084
rect 38660 8075 38712 8084
rect 38660 8041 38669 8075
rect 38669 8041 38703 8075
rect 38703 8041 38712 8075
rect 38660 8032 38712 8041
rect 24216 7828 24268 7880
rect 28172 7964 28224 8016
rect 30840 7964 30892 8016
rect 25596 7939 25648 7948
rect 25596 7905 25605 7939
rect 25605 7905 25639 7939
rect 25639 7905 25648 7939
rect 25596 7896 25648 7905
rect 27712 7896 27764 7948
rect 19708 7692 19760 7744
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 21916 7692 21968 7744
rect 24492 7692 24544 7744
rect 25044 7828 25096 7880
rect 25228 7828 25280 7880
rect 25964 7828 26016 7880
rect 28264 7828 28316 7880
rect 28356 7828 28408 7880
rect 28908 7828 28960 7880
rect 29460 7828 29512 7880
rect 29736 7828 29788 7880
rect 30104 7828 30156 7880
rect 24952 7760 25004 7812
rect 31852 7896 31904 7948
rect 30564 7828 30616 7880
rect 31668 7828 31720 7880
rect 36820 7964 36872 8016
rect 38292 7896 38344 7948
rect 36176 7871 36228 7880
rect 36176 7837 36185 7871
rect 36185 7837 36219 7871
rect 36219 7837 36228 7871
rect 36176 7828 36228 7837
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 26424 7692 26476 7744
rect 27620 7692 27672 7744
rect 28448 7735 28500 7744
rect 28448 7701 28457 7735
rect 28457 7701 28491 7735
rect 28491 7701 28500 7735
rect 28448 7692 28500 7701
rect 29736 7735 29788 7744
rect 29736 7701 29745 7735
rect 29745 7701 29779 7735
rect 29779 7701 29788 7735
rect 29736 7692 29788 7701
rect 36268 7760 36320 7812
rect 30012 7692 30064 7744
rect 30748 7692 30800 7744
rect 34796 7692 34848 7744
rect 37280 7760 37332 7812
rect 36912 7692 36964 7744
rect 38844 7871 38896 7880
rect 38844 7837 38853 7871
rect 38853 7837 38887 7871
rect 38887 7837 38896 7871
rect 38844 7828 38896 7837
rect 38660 7760 38712 7812
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 1216 7488 1268 7540
rect 1308 7420 1360 7472
rect 1124 7352 1176 7404
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 7932 7352 7984 7404
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 296 7284 348 7336
rect 7012 7284 7064 7336
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 15568 7531 15620 7540
rect 15568 7497 15577 7531
rect 15577 7497 15611 7531
rect 15611 7497 15620 7531
rect 15568 7488 15620 7497
rect 15752 7488 15804 7540
rect 16396 7488 16448 7540
rect 11520 7352 11572 7404
rect 11612 7352 11664 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 15476 7352 15528 7404
rect 7840 7216 7892 7268
rect 8944 7259 8996 7268
rect 8944 7225 8953 7259
rect 8953 7225 8987 7259
rect 8987 7225 8996 7259
rect 8944 7216 8996 7225
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 7288 7148 7340 7200
rect 9312 7327 9364 7336
rect 9312 7293 9346 7327
rect 9346 7293 9364 7327
rect 9312 7284 9364 7293
rect 9680 7284 9732 7336
rect 11796 7284 11848 7336
rect 12256 7284 12308 7336
rect 12992 7284 13044 7336
rect 14372 7327 14424 7336
rect 14372 7293 14390 7327
rect 14390 7293 14424 7327
rect 14372 7284 14424 7293
rect 15016 7284 15068 7336
rect 19340 7420 19392 7472
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 17776 7352 17828 7404
rect 20352 7488 20404 7540
rect 20536 7488 20588 7540
rect 24216 7488 24268 7540
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 20720 7395 20772 7404
rect 20720 7361 20729 7395
rect 20729 7361 20763 7395
rect 20763 7361 20772 7395
rect 20720 7352 20772 7361
rect 24584 7420 24636 7472
rect 25780 7488 25832 7540
rect 28264 7488 28316 7540
rect 30380 7488 30432 7540
rect 27896 7420 27948 7472
rect 28356 7420 28408 7472
rect 31576 7420 31628 7472
rect 36728 7488 36780 7540
rect 37280 7488 37332 7540
rect 38476 7488 38528 7540
rect 36176 7420 36228 7472
rect 39488 7488 39540 7540
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 19340 7284 19392 7336
rect 19616 7284 19668 7336
rect 21088 7284 21140 7336
rect 21916 7352 21968 7404
rect 22376 7352 22428 7404
rect 25228 7352 25280 7404
rect 25320 7395 25372 7404
rect 25320 7361 25329 7395
rect 25329 7361 25363 7395
rect 25363 7361 25372 7395
rect 25320 7352 25372 7361
rect 26332 7352 26384 7404
rect 27436 7352 27488 7404
rect 27804 7352 27856 7404
rect 21364 7284 21416 7336
rect 22008 7284 22060 7336
rect 24952 7284 25004 7336
rect 25044 7327 25096 7336
rect 25044 7293 25053 7327
rect 25053 7293 25087 7327
rect 25087 7293 25096 7327
rect 25044 7284 25096 7293
rect 9588 7148 9640 7200
rect 9864 7148 9916 7200
rect 10140 7191 10192 7200
rect 10140 7157 10149 7191
rect 10149 7157 10183 7191
rect 10183 7157 10192 7191
rect 10140 7148 10192 7157
rect 10600 7148 10652 7200
rect 13636 7148 13688 7200
rect 14924 7216 14976 7268
rect 14832 7148 14884 7200
rect 19984 7216 20036 7268
rect 24492 7216 24544 7268
rect 19064 7148 19116 7200
rect 19616 7148 19668 7200
rect 20352 7148 20404 7200
rect 24124 7148 24176 7200
rect 24216 7148 24268 7200
rect 26516 7216 26568 7268
rect 28908 7284 28960 7336
rect 31484 7352 31536 7404
rect 34244 7352 34296 7404
rect 34704 7352 34756 7404
rect 36360 7395 36412 7404
rect 36360 7361 36369 7395
rect 36369 7361 36403 7395
rect 36403 7361 36412 7395
rect 36360 7352 36412 7361
rect 36636 7395 36688 7404
rect 36636 7361 36645 7395
rect 36645 7361 36679 7395
rect 36679 7361 36688 7395
rect 36636 7352 36688 7361
rect 39856 7420 39908 7472
rect 37740 7395 37792 7404
rect 37740 7361 37749 7395
rect 37749 7361 37783 7395
rect 37783 7361 37792 7395
rect 37740 7352 37792 7361
rect 38108 7395 38160 7404
rect 38108 7361 38117 7395
rect 38117 7361 38151 7395
rect 38151 7361 38160 7395
rect 38108 7352 38160 7361
rect 38568 7352 38620 7404
rect 38844 7395 38896 7404
rect 38844 7361 38853 7395
rect 38853 7361 38887 7395
rect 38887 7361 38896 7395
rect 38844 7352 38896 7361
rect 39580 7352 39632 7404
rect 27252 7148 27304 7200
rect 32772 7216 32824 7268
rect 38384 7284 38436 7336
rect 39488 7216 39540 7268
rect 34520 7148 34572 7200
rect 35624 7148 35676 7200
rect 39396 7191 39448 7200
rect 39396 7157 39405 7191
rect 39405 7157 39439 7191
rect 39439 7157 39448 7191
rect 39396 7148 39448 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 7748 6944 7800 6996
rect 1216 6876 1268 6928
rect 848 6808 900 6860
rect 7564 6876 7616 6928
rect 756 6740 808 6792
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 8944 6944 8996 6996
rect 9312 6944 9364 6996
rect 8484 6876 8536 6928
rect 1032 6672 1084 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 1768 6604 1820 6656
rect 5540 6740 5592 6792
rect 3516 6604 3568 6656
rect 3700 6672 3752 6724
rect 5448 6715 5500 6724
rect 5448 6681 5457 6715
rect 5457 6681 5491 6715
rect 5491 6681 5500 6715
rect 5448 6672 5500 6681
rect 5724 6604 5776 6656
rect 6276 6740 6328 6792
rect 6460 6672 6512 6724
rect 7656 6740 7708 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8116 6740 8168 6792
rect 7288 6672 7340 6724
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 8300 6604 8352 6656
rect 9496 6808 9548 6860
rect 10048 6851 10100 6860
rect 10048 6817 10066 6851
rect 10066 6817 10100 6851
rect 10048 6808 10100 6817
rect 22560 6944 22612 6996
rect 22652 6944 22704 6996
rect 11428 6919 11480 6928
rect 11428 6885 11437 6919
rect 11437 6885 11471 6919
rect 11471 6885 11480 6919
rect 11428 6876 11480 6885
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 11796 6851 11848 6860
rect 11796 6817 11805 6851
rect 11805 6817 11839 6851
rect 11839 6817 11848 6851
rect 11796 6808 11848 6817
rect 15200 6876 15252 6928
rect 16304 6876 16356 6928
rect 18880 6876 18932 6928
rect 19616 6876 19668 6928
rect 15384 6808 15436 6860
rect 17960 6808 18012 6860
rect 19524 6808 19576 6860
rect 20260 6808 20312 6860
rect 20352 6851 20404 6860
rect 20352 6817 20361 6851
rect 20361 6817 20395 6851
rect 20395 6817 20404 6851
rect 20352 6808 20404 6817
rect 24492 6987 24544 6996
rect 24492 6953 24501 6987
rect 24501 6953 24535 6987
rect 24535 6953 24544 6987
rect 24492 6944 24544 6953
rect 25872 6944 25924 6996
rect 26884 6944 26936 6996
rect 27436 6876 27488 6928
rect 20904 6808 20956 6860
rect 21180 6808 21232 6860
rect 21548 6808 21600 6860
rect 23112 6851 23164 6860
rect 23112 6817 23121 6851
rect 23121 6817 23155 6851
rect 23155 6817 23164 6851
rect 23112 6808 23164 6817
rect 25688 6808 25740 6860
rect 26516 6808 26568 6860
rect 27528 6808 27580 6860
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 11060 6783 11112 6792
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 12900 6783 12952 6792
rect 9404 6604 9456 6656
rect 11796 6672 11848 6724
rect 12900 6749 12912 6783
rect 12912 6749 12946 6783
rect 12946 6749 12952 6783
rect 12900 6740 12952 6749
rect 13268 6740 13320 6792
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 14832 6740 14884 6792
rect 15016 6783 15068 6792
rect 15016 6749 15025 6783
rect 15025 6749 15059 6783
rect 15059 6749 15068 6783
rect 15016 6740 15068 6749
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 28264 6808 28316 6860
rect 36636 6944 36688 6996
rect 39856 6944 39908 6996
rect 37004 6919 37056 6928
rect 37004 6885 37013 6919
rect 37013 6885 37047 6919
rect 37047 6885 37056 6919
rect 37004 6876 37056 6885
rect 37096 6808 37148 6860
rect 37464 6808 37516 6860
rect 37924 6808 37976 6860
rect 38016 6851 38068 6860
rect 38016 6817 38025 6851
rect 38025 6817 38059 6851
rect 38059 6817 38068 6851
rect 38016 6808 38068 6817
rect 38384 6851 38436 6860
rect 38384 6817 38393 6851
rect 38393 6817 38427 6851
rect 38427 6817 38436 6851
rect 38384 6808 38436 6817
rect 16212 6740 16264 6749
rect 14188 6672 14240 6724
rect 17776 6715 17828 6724
rect 17776 6681 17785 6715
rect 17785 6681 17819 6715
rect 17819 6681 17828 6715
rect 17776 6672 17828 6681
rect 17960 6715 18012 6724
rect 17960 6681 17969 6715
rect 17969 6681 18003 6715
rect 18003 6681 18012 6715
rect 17960 6672 18012 6681
rect 18236 6740 18288 6792
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 22008 6740 22060 6792
rect 22100 6783 22152 6792
rect 22100 6749 22109 6783
rect 22109 6749 22143 6783
rect 22143 6749 22152 6783
rect 22100 6740 22152 6749
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 15476 6604 15528 6656
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 18328 6604 18380 6656
rect 19248 6604 19300 6656
rect 20444 6604 20496 6656
rect 20628 6604 20680 6656
rect 21548 6672 21600 6724
rect 22100 6604 22152 6656
rect 25228 6783 25280 6792
rect 25228 6749 25237 6783
rect 25237 6749 25271 6783
rect 25271 6749 25280 6783
rect 25228 6740 25280 6749
rect 25320 6740 25372 6792
rect 23756 6672 23808 6724
rect 26700 6783 26752 6792
rect 26700 6749 26709 6783
rect 26709 6749 26743 6783
rect 26743 6749 26752 6783
rect 26700 6740 26752 6749
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 27804 6740 27856 6792
rect 28172 6783 28224 6792
rect 28172 6749 28181 6783
rect 28181 6749 28215 6783
rect 28215 6749 28224 6783
rect 28172 6740 28224 6749
rect 28356 6740 28408 6792
rect 28816 6740 28868 6792
rect 34612 6740 34664 6792
rect 30104 6672 30156 6724
rect 24032 6604 24084 6656
rect 24124 6647 24176 6656
rect 24124 6613 24133 6647
rect 24133 6613 24167 6647
rect 24167 6613 24176 6647
rect 24124 6604 24176 6613
rect 25688 6604 25740 6656
rect 26608 6604 26660 6656
rect 26700 6604 26752 6656
rect 27804 6604 27856 6656
rect 27896 6647 27948 6656
rect 27896 6613 27905 6647
rect 27905 6613 27939 6647
rect 27939 6613 27948 6647
rect 27896 6604 27948 6613
rect 27988 6604 28040 6656
rect 28632 6604 28684 6656
rect 28724 6604 28776 6656
rect 29000 6604 29052 6656
rect 38752 6740 38804 6792
rect 37556 6672 37608 6724
rect 38476 6604 38528 6656
rect 39672 6604 39724 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 3516 6400 3568 6452
rect 6644 6400 6696 6452
rect 7656 6400 7708 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 5448 6264 5500 6316
rect 8392 6307 8444 6316
rect 8392 6273 8410 6307
rect 8410 6273 8444 6307
rect 8392 6264 8444 6273
rect 572 6196 624 6248
rect 6276 6196 6328 6248
rect 8668 6196 8720 6248
rect 8760 6239 8812 6248
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 8852 6196 8904 6248
rect 9496 6264 9548 6316
rect 10140 6332 10192 6384
rect 10416 6400 10468 6452
rect 11060 6400 11112 6452
rect 11888 6400 11940 6452
rect 12992 6400 13044 6452
rect 14740 6400 14792 6452
rect 10416 6264 10468 6316
rect 11612 6264 11664 6316
rect 12440 6264 12492 6316
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 10508 6196 10560 6248
rect 11704 6196 11756 6248
rect 8116 6060 8168 6112
rect 8668 6060 8720 6112
rect 10692 6060 10744 6112
rect 11060 6060 11112 6112
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 14832 6307 14884 6316
rect 14832 6273 14850 6307
rect 14850 6273 14884 6307
rect 14832 6264 14884 6273
rect 16212 6264 16264 6316
rect 18236 6264 18288 6316
rect 14464 6196 14516 6248
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 18972 6400 19024 6452
rect 19156 6400 19208 6452
rect 15384 6128 15436 6180
rect 18512 6128 18564 6180
rect 12256 6060 12308 6112
rect 13636 6060 13688 6112
rect 14464 6060 14516 6112
rect 14556 6060 14608 6112
rect 16120 6060 16172 6112
rect 16672 6060 16724 6112
rect 18696 6196 18748 6248
rect 19340 6307 19392 6316
rect 19340 6273 19367 6307
rect 19367 6273 19392 6307
rect 19340 6264 19392 6273
rect 19524 6264 19576 6316
rect 20812 6400 20864 6452
rect 21456 6400 21508 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 20260 6375 20312 6384
rect 20260 6341 20269 6375
rect 20269 6341 20303 6375
rect 20303 6341 20312 6375
rect 20260 6332 20312 6341
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 19614 6239 19666 6248
rect 19614 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19666 6239
rect 19614 6196 19666 6205
rect 19800 6196 19852 6248
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 20812 6264 20864 6316
rect 20904 6307 20956 6316
rect 20904 6273 20913 6307
rect 20913 6273 20947 6307
rect 20947 6273 20956 6307
rect 20904 6264 20956 6273
rect 20628 6060 20680 6112
rect 26240 6375 26292 6384
rect 26240 6341 26249 6375
rect 26249 6341 26283 6375
rect 26283 6341 26292 6375
rect 26240 6332 26292 6341
rect 21364 6264 21416 6316
rect 22836 6264 22888 6316
rect 23388 6264 23440 6316
rect 21456 6196 21508 6248
rect 23756 6196 23808 6248
rect 24860 6264 24912 6316
rect 26332 6307 26384 6316
rect 26332 6273 26341 6307
rect 26341 6273 26375 6307
rect 26375 6273 26384 6307
rect 26332 6264 26384 6273
rect 26608 6443 26660 6452
rect 26608 6409 26617 6443
rect 26617 6409 26651 6443
rect 26651 6409 26660 6443
rect 26608 6400 26660 6409
rect 27896 6400 27948 6452
rect 25228 6060 25280 6112
rect 25320 6103 25372 6112
rect 25320 6069 25329 6103
rect 25329 6069 25363 6103
rect 25363 6069 25372 6103
rect 25320 6060 25372 6069
rect 27896 6307 27948 6316
rect 27896 6273 27905 6307
rect 27905 6273 27939 6307
rect 27939 6273 27948 6307
rect 27896 6264 27948 6273
rect 27620 6239 27672 6248
rect 27620 6205 27629 6239
rect 27629 6205 27663 6239
rect 27663 6205 27672 6239
rect 27620 6196 27672 6205
rect 27528 6128 27580 6180
rect 28172 6239 28224 6248
rect 28172 6205 28181 6239
rect 28181 6205 28215 6239
rect 28215 6205 28224 6239
rect 28172 6196 28224 6205
rect 28816 6443 28868 6452
rect 28816 6409 28825 6443
rect 28825 6409 28859 6443
rect 28859 6409 28868 6443
rect 28816 6400 28868 6409
rect 30932 6400 30984 6452
rect 36544 6400 36596 6452
rect 39028 6443 39080 6452
rect 39028 6409 39037 6443
rect 39037 6409 39071 6443
rect 39071 6409 39080 6443
rect 39028 6400 39080 6409
rect 39764 6400 39816 6452
rect 34336 6332 34388 6384
rect 37924 6332 37976 6384
rect 28908 6307 28960 6316
rect 28908 6273 28917 6307
rect 28917 6273 28951 6307
rect 28951 6273 28960 6307
rect 28908 6264 28960 6273
rect 35992 6264 36044 6316
rect 39672 6332 39724 6384
rect 34428 6196 34480 6248
rect 38568 6196 38620 6248
rect 38292 6128 38344 6180
rect 28356 6060 28408 6112
rect 36452 6060 36504 6112
rect 38476 6060 38528 6112
rect 38660 6103 38712 6112
rect 38660 6069 38669 6103
rect 38669 6069 38703 6103
rect 38703 6069 38712 6103
rect 38660 6060 38712 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 1860 5899 1912 5908
rect 1860 5865 1869 5899
rect 1869 5865 1903 5899
rect 1903 5865 1912 5899
rect 1860 5856 1912 5865
rect 2320 5856 2372 5908
rect 6828 5788 6880 5840
rect 7012 5788 7064 5840
rect 8392 5788 8444 5840
rect 848 5720 900 5772
rect 204 5652 256 5704
rect 2504 5720 2556 5772
rect 6920 5720 6972 5772
rect 7564 5720 7616 5772
rect 9680 5856 9732 5908
rect 10692 5856 10744 5908
rect 11060 5788 11112 5840
rect 11152 5788 11204 5840
rect 14648 5856 14700 5908
rect 17960 5788 18012 5840
rect 18696 5788 18748 5840
rect 20352 5856 20404 5908
rect 25228 5856 25280 5908
rect 21916 5788 21968 5840
rect 28172 5788 28224 5840
rect 37832 5856 37884 5908
rect 38200 5899 38252 5908
rect 38200 5865 38209 5899
rect 38209 5865 38243 5899
rect 38243 5865 38252 5899
rect 38200 5856 38252 5865
rect 39580 5856 39632 5908
rect 9680 5720 9732 5772
rect 10784 5720 10836 5772
rect 664 5584 716 5636
rect 3608 5652 3660 5704
rect 7748 5652 7800 5704
rect 8852 5652 8904 5704
rect 11888 5720 11940 5772
rect 12440 5720 12492 5772
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 11704 5652 11756 5704
rect 16764 5720 16816 5772
rect 13176 5652 13228 5704
rect 14740 5652 14792 5704
rect 19156 5720 19208 5772
rect 18604 5652 18656 5704
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 20904 5720 20956 5772
rect 24952 5763 25004 5772
rect 24952 5729 24961 5763
rect 24961 5729 24995 5763
rect 24995 5729 25004 5763
rect 24952 5720 25004 5729
rect 29276 5720 29328 5772
rect 19524 5652 19576 5661
rect 1768 5584 1820 5636
rect 10784 5584 10836 5636
rect 11244 5584 11296 5636
rect 11336 5584 11388 5636
rect 13268 5584 13320 5636
rect 13820 5627 13872 5636
rect 13820 5593 13829 5627
rect 13829 5593 13863 5627
rect 13863 5593 13872 5627
rect 13820 5584 13872 5593
rect 1584 5516 1636 5568
rect 10416 5516 10468 5568
rect 11152 5516 11204 5568
rect 11704 5516 11756 5568
rect 12900 5516 12952 5568
rect 13544 5516 13596 5568
rect 15660 5584 15712 5636
rect 15752 5584 15804 5636
rect 23388 5652 23440 5704
rect 25228 5695 25280 5704
rect 25228 5661 25237 5695
rect 25237 5661 25271 5695
rect 25271 5661 25280 5695
rect 25228 5652 25280 5661
rect 26056 5695 26108 5704
rect 26056 5661 26065 5695
rect 26065 5661 26099 5695
rect 26099 5661 26108 5695
rect 26056 5652 26108 5661
rect 28264 5652 28316 5704
rect 35624 5652 35676 5704
rect 39948 5788 40000 5840
rect 21456 5584 21508 5636
rect 24676 5584 24728 5636
rect 38660 5584 38712 5636
rect 14648 5516 14700 5568
rect 14740 5516 14792 5568
rect 16672 5516 16724 5568
rect 16764 5516 16816 5568
rect 20444 5516 20496 5568
rect 20536 5559 20588 5568
rect 20536 5525 20545 5559
rect 20545 5525 20579 5559
rect 20579 5525 20588 5559
rect 20536 5516 20588 5525
rect 26884 5516 26936 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 5908 5312 5960 5364
rect 6828 5312 6880 5364
rect 13728 5312 13780 5364
rect 20444 5312 20496 5364
rect 20720 5312 20772 5364
rect 23112 5312 23164 5364
rect 28448 5312 28500 5364
rect 28724 5312 28776 5364
rect 34796 5312 34848 5364
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 6644 5244 6696 5296
rect 388 5176 440 5228
rect 848 5108 900 5160
rect 5816 5176 5868 5228
rect 7104 5176 7156 5228
rect 7564 5176 7616 5228
rect 11980 5244 12032 5296
rect 19340 5244 19392 5296
rect 21548 5244 21600 5296
rect 25596 5244 25648 5296
rect 26056 5244 26108 5296
rect 27344 5244 27396 5296
rect 38936 5244 38988 5296
rect 12256 5176 12308 5228
rect 13544 5176 13596 5228
rect 20812 5176 20864 5228
rect 27436 5176 27488 5228
rect 28172 5176 28224 5228
rect 38844 5219 38896 5228
rect 38844 5185 38853 5219
rect 38853 5185 38887 5219
rect 38887 5185 38896 5219
rect 38844 5176 38896 5185
rect 5724 5108 5776 5160
rect 12348 5108 12400 5160
rect 12440 5108 12492 5160
rect 18052 5108 18104 5160
rect 18880 5108 18932 5160
rect 28080 5108 28132 5160
rect 5356 5040 5408 5092
rect 13084 5040 13136 5092
rect 13176 5040 13228 5092
rect 25504 5040 25556 5092
rect 27896 5040 27948 5092
rect 37280 5108 37332 5160
rect 4804 4972 4856 5024
rect 4896 4972 4948 5024
rect 5908 4972 5960 5024
rect 7012 4972 7064 5024
rect 15384 4972 15436 5024
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 28908 4972 28960 5024
rect 29276 5015 29328 5024
rect 29276 4981 29285 5015
rect 29285 4981 29319 5015
rect 29319 4981 29328 5015
rect 29276 4972 29328 4981
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 5080 4768 5132 4820
rect 6276 4768 6328 4820
rect 4988 4632 5040 4684
rect 5816 4675 5868 4684
rect 5816 4641 5834 4675
rect 5834 4641 5868 4675
rect 5816 4632 5868 4641
rect 6644 4675 6696 4684
rect 6644 4641 6653 4675
rect 6653 4641 6687 4675
rect 6687 4641 6696 4675
rect 6644 4632 6696 4641
rect 10508 4768 10560 4820
rect 756 4564 808 4616
rect 848 4496 900 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 4344 4496 4396 4548
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6736 4564 6788 4616
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4896 4428 4948 4480
rect 6644 4496 6696 4548
rect 10232 4632 10284 4684
rect 11520 4768 11572 4820
rect 13176 4768 13228 4820
rect 21456 4700 21508 4752
rect 22284 4768 22336 4820
rect 23848 4768 23900 4820
rect 11428 4632 11480 4684
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 12164 4675 12216 4684
rect 12164 4641 12173 4675
rect 12173 4641 12207 4675
rect 12207 4641 12216 4675
rect 12164 4632 12216 4641
rect 14740 4632 14792 4684
rect 19064 4632 19116 4684
rect 23296 4700 23348 4752
rect 30288 4768 30340 4820
rect 39396 4811 39448 4820
rect 39396 4777 39405 4811
rect 39405 4777 39439 4811
rect 39439 4777 39448 4811
rect 39396 4768 39448 4777
rect 29644 4700 29696 4752
rect 39948 4700 40000 4752
rect 21824 4675 21876 4684
rect 21824 4641 21833 4675
rect 21833 4641 21867 4675
rect 21867 4641 21876 4675
rect 21824 4632 21876 4641
rect 22192 4632 22244 4684
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 14832 4564 14884 4616
rect 16212 4564 16264 4616
rect 7012 4496 7064 4548
rect 7472 4496 7524 4548
rect 8208 4496 8260 4548
rect 16856 4539 16908 4548
rect 16856 4505 16865 4539
rect 16865 4505 16899 4539
rect 16899 4505 16908 4539
rect 16856 4496 16908 4505
rect 17868 4496 17920 4548
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 22560 4607 22612 4616
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 22744 4564 22796 4616
rect 29000 4607 29052 4616
rect 29000 4573 29009 4607
rect 29009 4573 29043 4607
rect 29043 4573 29052 4607
rect 29000 4564 29052 4573
rect 29092 4564 29144 4616
rect 29920 4607 29972 4616
rect 29920 4573 29929 4607
rect 29929 4573 29963 4607
rect 29963 4573 29972 4607
rect 29920 4564 29972 4573
rect 37464 4564 37516 4616
rect 38936 4564 38988 4616
rect 21548 4496 21600 4548
rect 23388 4496 23440 4548
rect 30012 4496 30064 4548
rect 5724 4428 5776 4480
rect 6736 4428 6788 4480
rect 7840 4428 7892 4480
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 10416 4428 10468 4480
rect 11980 4428 12032 4480
rect 15384 4428 15436 4480
rect 18328 4428 18380 4480
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 21824 4428 21876 4480
rect 22468 4428 22520 4480
rect 22560 4428 22612 4480
rect 24584 4428 24636 4480
rect 28264 4471 28316 4480
rect 28264 4437 28273 4471
rect 28273 4437 28307 4471
rect 28307 4437 28316 4471
rect 28264 4428 28316 4437
rect 29552 4428 29604 4480
rect 30656 4428 30708 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 5080 4267 5132 4276
rect 5080 4233 5089 4267
rect 5089 4233 5123 4267
rect 5123 4233 5132 4267
rect 5080 4224 5132 4233
rect 5172 4224 5224 4276
rect 5908 4224 5960 4276
rect 7288 4224 7340 4276
rect 10968 4224 11020 4276
rect 3792 4199 3844 4208
rect 3792 4165 3801 4199
rect 3801 4165 3835 4199
rect 3835 4165 3844 4199
rect 3792 4156 3844 4165
rect 388 4088 440 4140
rect 848 4020 900 4072
rect 3976 4088 4028 4140
rect 5356 4156 5408 4208
rect 10508 4156 10560 4208
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 4896 4088 4948 4140
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7104 4088 7156 4140
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 9404 4088 9456 4140
rect 11704 4156 11756 4208
rect 12532 4224 12584 4276
rect 17684 4224 17736 4276
rect 18604 4224 18656 4276
rect 7656 4020 7708 4072
rect 10508 4020 10560 4072
rect 3700 3884 3752 3936
rect 4068 3884 4120 3936
rect 5540 3884 5592 3936
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 5632 3884 5684 3893
rect 6000 3995 6052 4004
rect 6000 3961 6009 3995
rect 6009 3961 6043 3995
rect 6043 3961 6052 3995
rect 6000 3952 6052 3961
rect 9588 3952 9640 4004
rect 10600 3952 10652 4004
rect 12348 4088 12400 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 19064 4199 19116 4208
rect 19064 4165 19073 4199
rect 19073 4165 19107 4199
rect 19107 4165 19116 4199
rect 19064 4156 19116 4165
rect 18420 4088 18472 4140
rect 21456 4156 21508 4208
rect 10784 4020 10836 4072
rect 11428 4020 11480 4072
rect 16580 4020 16632 4072
rect 16764 4063 16816 4072
rect 16764 4029 16773 4063
rect 16773 4029 16807 4063
rect 16807 4029 16816 4063
rect 16764 4020 16816 4029
rect 17868 4063 17920 4072
rect 17868 4029 17877 4063
rect 17877 4029 17911 4063
rect 17911 4029 17920 4063
rect 17868 4020 17920 4029
rect 19800 4020 19852 4072
rect 20352 4020 20404 4072
rect 21180 4020 21232 4072
rect 21364 4020 21416 4072
rect 22008 4088 22060 4140
rect 22376 4156 22428 4208
rect 22560 4156 22612 4208
rect 23296 4156 23348 4208
rect 22744 4088 22796 4140
rect 23112 4131 23164 4140
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 23388 4131 23440 4140
rect 23388 4097 23397 4131
rect 23397 4097 23431 4131
rect 23431 4097 23440 4131
rect 23388 4088 23440 4097
rect 28356 4224 28408 4276
rect 23572 4088 23624 4140
rect 23848 4156 23900 4208
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 27620 4156 27672 4208
rect 30012 4224 30064 4276
rect 30656 4267 30708 4276
rect 30656 4233 30665 4267
rect 30665 4233 30699 4267
rect 30699 4233 30708 4267
rect 30656 4224 30708 4233
rect 23756 4088 23808 4097
rect 24124 4088 24176 4140
rect 27804 4088 27856 4140
rect 28632 4131 28684 4140
rect 28632 4097 28641 4131
rect 28641 4097 28675 4131
rect 28675 4097 28684 4131
rect 28632 4088 28684 4097
rect 25136 4020 25188 4072
rect 15292 3995 15344 4004
rect 15292 3961 15301 3995
rect 15301 3961 15335 3995
rect 15335 3961 15344 3995
rect 15292 3952 15344 3961
rect 15476 3995 15528 4004
rect 15476 3961 15485 3995
rect 15485 3961 15519 3995
rect 15519 3961 15528 3995
rect 15476 3952 15528 3961
rect 7196 3884 7248 3936
rect 7288 3884 7340 3936
rect 11060 3884 11112 3936
rect 11152 3884 11204 3936
rect 15660 3884 15712 3936
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 20720 3952 20772 4004
rect 21640 3952 21692 4004
rect 21732 3884 21784 3936
rect 22192 3884 22244 3936
rect 23204 3995 23256 4004
rect 23204 3961 23213 3995
rect 23213 3961 23247 3995
rect 23247 3961 23256 3995
rect 23204 3952 23256 3961
rect 23480 3995 23532 4004
rect 23480 3961 23489 3995
rect 23489 3961 23523 3995
rect 23523 3961 23532 3995
rect 23480 3952 23532 3961
rect 26240 3952 26292 4004
rect 27528 4020 27580 4072
rect 28080 4063 28132 4072
rect 28080 4029 28089 4063
rect 28089 4029 28123 4063
rect 28123 4029 28132 4063
rect 28080 4020 28132 4029
rect 27988 3952 28040 4004
rect 28448 4063 28500 4072
rect 28448 4029 28482 4063
rect 28482 4029 28500 4063
rect 30288 4199 30340 4208
rect 30288 4165 30297 4199
rect 30297 4165 30331 4199
rect 30331 4165 30340 4199
rect 30288 4156 30340 4165
rect 29460 4088 29512 4140
rect 29736 4088 29788 4140
rect 28448 4020 28500 4029
rect 29368 4020 29420 4072
rect 39212 4131 39264 4140
rect 39212 4097 39221 4131
rect 39221 4097 39255 4131
rect 39255 4097 39264 4131
rect 39212 4088 39264 4097
rect 40040 4020 40092 4072
rect 39488 3952 39540 4004
rect 22744 3884 22796 3936
rect 23664 3884 23716 3936
rect 26332 3884 26384 3936
rect 28632 3884 28684 3936
rect 29552 3884 29604 3936
rect 30840 3927 30892 3936
rect 30840 3893 30849 3927
rect 30849 3893 30883 3927
rect 30883 3893 30892 3927
rect 30840 3884 30892 3893
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 3792 3680 3844 3732
rect 4988 3723 5040 3732
rect 4988 3689 4997 3723
rect 4997 3689 5031 3723
rect 5031 3689 5040 3723
rect 4988 3680 5040 3689
rect 2412 3612 2464 3664
rect 5540 3655 5592 3664
rect 5540 3621 5549 3655
rect 5549 3621 5583 3655
rect 5583 3621 5592 3655
rect 5540 3612 5592 3621
rect 1032 3544 1084 3596
rect 204 3476 256 3528
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 5172 3544 5224 3596
rect 6736 3680 6788 3732
rect 7012 3680 7064 3732
rect 9496 3680 9548 3732
rect 9588 3723 9640 3732
rect 9588 3689 9597 3723
rect 9597 3689 9631 3723
rect 9631 3689 9640 3723
rect 9588 3680 9640 3689
rect 9772 3680 9824 3732
rect 6920 3612 6972 3664
rect 7840 3612 7892 3664
rect 12440 3680 12492 3732
rect 13636 3680 13688 3732
rect 7564 3587 7616 3596
rect 7564 3553 7582 3587
rect 7582 3553 7616 3587
rect 7564 3544 7616 3553
rect 10784 3612 10836 3664
rect 848 3408 900 3460
rect 3792 3476 3844 3528
rect 4804 3476 4856 3528
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 16580 3680 16632 3732
rect 15568 3612 15620 3664
rect 8392 3476 8444 3485
rect 9772 3476 9824 3528
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 11336 3476 11388 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 16028 3544 16080 3596
rect 17684 3680 17736 3732
rect 17592 3544 17644 3596
rect 18052 3612 18104 3664
rect 20720 3612 20772 3664
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 21180 3544 21232 3553
rect 22100 3544 22152 3596
rect 22284 3587 22336 3596
rect 22284 3553 22293 3587
rect 22293 3553 22327 3587
rect 22327 3553 22336 3587
rect 22284 3544 22336 3553
rect 22560 3544 22612 3596
rect 10048 3408 10100 3460
rect 11980 3408 12032 3460
rect 15292 3451 15344 3460
rect 15292 3417 15301 3451
rect 15301 3417 15335 3451
rect 15335 3417 15344 3451
rect 15292 3408 15344 3417
rect 6644 3340 6696 3392
rect 7472 3340 7524 3392
rect 8852 3340 8904 3392
rect 9588 3340 9640 3392
rect 10140 3383 10192 3392
rect 10140 3349 10149 3383
rect 10149 3349 10183 3383
rect 10183 3349 10192 3383
rect 10140 3340 10192 3349
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 13728 3340 13780 3392
rect 15660 3383 15712 3392
rect 15660 3349 15669 3383
rect 15669 3349 15703 3383
rect 15703 3349 15712 3383
rect 15660 3340 15712 3349
rect 16948 3519 17000 3528
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 17132 3476 17184 3528
rect 17868 3476 17920 3528
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 21916 3476 21968 3528
rect 23020 3544 23072 3596
rect 23296 3587 23348 3596
rect 23296 3553 23330 3587
rect 23330 3553 23348 3587
rect 23296 3544 23348 3553
rect 24124 3723 24176 3732
rect 24124 3689 24133 3723
rect 24133 3689 24167 3723
rect 24167 3689 24176 3723
rect 24124 3680 24176 3689
rect 24400 3723 24452 3732
rect 24400 3689 24409 3723
rect 24409 3689 24443 3723
rect 24443 3689 24452 3723
rect 24400 3680 24452 3689
rect 25872 3680 25924 3732
rect 25780 3612 25832 3664
rect 18144 3408 18196 3460
rect 21548 3408 21600 3460
rect 17776 3340 17828 3392
rect 21456 3340 21508 3392
rect 21640 3340 21692 3392
rect 22100 3340 22152 3392
rect 23204 3519 23256 3528
rect 23204 3485 23213 3519
rect 23213 3485 23247 3519
rect 23247 3485 23256 3519
rect 23204 3476 23256 3485
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 26424 3476 26476 3528
rect 27436 3519 27488 3528
rect 27436 3485 27445 3519
rect 27445 3485 27479 3519
rect 27479 3485 27488 3519
rect 27436 3476 27488 3485
rect 27528 3519 27580 3528
rect 27528 3485 27537 3519
rect 27537 3485 27571 3519
rect 27571 3485 27580 3519
rect 27988 3612 28040 3664
rect 28264 3612 28316 3664
rect 29920 3680 29972 3732
rect 30196 3680 30248 3732
rect 30288 3723 30340 3732
rect 30288 3689 30297 3723
rect 30297 3689 30331 3723
rect 30331 3689 30340 3723
rect 30288 3680 30340 3689
rect 32864 3680 32916 3732
rect 33692 3680 33744 3732
rect 34060 3680 34112 3732
rect 35808 3680 35860 3732
rect 29460 3612 29512 3664
rect 29644 3612 29696 3664
rect 30840 3612 30892 3664
rect 31668 3612 31720 3664
rect 35348 3612 35400 3664
rect 37648 3680 37700 3732
rect 39396 3723 39448 3732
rect 39396 3689 39405 3723
rect 39405 3689 39439 3723
rect 39439 3689 39448 3723
rect 39396 3680 39448 3689
rect 37004 3612 37056 3664
rect 39948 3612 40000 3664
rect 28448 3587 28500 3596
rect 28448 3553 28457 3587
rect 28457 3553 28491 3587
rect 28491 3553 28500 3587
rect 28448 3544 28500 3553
rect 28540 3587 28592 3596
rect 28540 3553 28574 3587
rect 28574 3553 28592 3587
rect 28540 3544 28592 3553
rect 29276 3544 29328 3596
rect 27528 3476 27580 3485
rect 22284 3340 22336 3392
rect 29552 3476 29604 3528
rect 29828 3476 29880 3528
rect 30564 3519 30616 3528
rect 30564 3485 30573 3519
rect 30573 3485 30607 3519
rect 30607 3485 30616 3519
rect 30564 3476 30616 3485
rect 31576 3476 31628 3528
rect 32864 3476 32916 3528
rect 33876 3519 33928 3528
rect 33876 3485 33885 3519
rect 33885 3485 33919 3519
rect 33919 3485 33928 3519
rect 33876 3476 33928 3485
rect 34152 3519 34204 3528
rect 34152 3485 34161 3519
rect 34161 3485 34195 3519
rect 34195 3485 34204 3519
rect 34152 3476 34204 3485
rect 35164 3476 35216 3528
rect 35532 3476 35584 3528
rect 35716 3476 35768 3528
rect 38844 3519 38896 3528
rect 38844 3485 38853 3519
rect 38853 3485 38887 3519
rect 38887 3485 38896 3519
rect 38844 3476 38896 3485
rect 30012 3408 30064 3460
rect 29920 3340 29972 3392
rect 36544 3408 36596 3460
rect 36820 3408 36872 3460
rect 35440 3340 35492 3392
rect 35532 3340 35584 3392
rect 37096 3340 37148 3392
rect 37648 3340 37700 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 4344 3136 4396 3188
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 3884 3068 3936 3120
rect 7380 3136 7432 3188
rect 7840 3136 7892 3188
rect 9864 3136 9916 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 1216 3000 1268 3052
rect 756 2932 808 2984
rect 2504 2932 2556 2984
rect 388 2864 440 2916
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5356 3000 5408 3052
rect 6828 3068 6880 3120
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 8484 3068 8536 3120
rect 11428 3068 11480 3120
rect 17408 3136 17460 3188
rect 12164 3068 12216 3120
rect 21640 3179 21692 3188
rect 21640 3145 21649 3179
rect 21649 3145 21683 3179
rect 21683 3145 21692 3179
rect 21640 3136 21692 3145
rect 8392 3000 8444 3052
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 11980 3000 12032 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 6736 2975 6788 2984
rect 6736 2941 6745 2975
rect 6745 2941 6779 2975
rect 6779 2941 6788 2975
rect 6736 2932 6788 2941
rect 8208 2932 8260 2984
rect 2780 2907 2832 2916
rect 2780 2873 2789 2907
rect 2789 2873 2823 2907
rect 2823 2873 2832 2907
rect 2780 2864 2832 2873
rect 9588 2975 9640 2984
rect 9588 2941 9597 2975
rect 9597 2941 9631 2975
rect 9631 2941 9640 2975
rect 9588 2932 9640 2941
rect 10232 2975 10284 2984
rect 10232 2941 10241 2975
rect 10241 2941 10275 2975
rect 10275 2941 10284 2975
rect 10232 2932 10284 2941
rect 10508 2932 10560 2984
rect 9772 2864 9824 2916
rect 6644 2796 6696 2848
rect 9312 2796 9364 2848
rect 12532 2975 12584 2984
rect 12532 2941 12541 2975
rect 12541 2941 12575 2975
rect 12575 2941 12584 2975
rect 12532 2932 12584 2941
rect 13728 2932 13780 2984
rect 15752 2932 15804 2984
rect 15844 2975 15896 2984
rect 15844 2941 15853 2975
rect 15853 2941 15887 2975
rect 15887 2941 15896 2975
rect 15844 2932 15896 2941
rect 16028 3000 16080 3052
rect 17316 3000 17368 3052
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 17868 3000 17920 3052
rect 22468 3111 22520 3120
rect 22468 3077 22477 3111
rect 22477 3077 22511 3111
rect 22511 3077 22520 3111
rect 22468 3068 22520 3077
rect 22836 3111 22888 3120
rect 22836 3077 22845 3111
rect 22845 3077 22879 3111
rect 22879 3077 22888 3111
rect 22836 3068 22888 3077
rect 22928 3068 22980 3120
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 21916 3043 21968 3052
rect 21916 3009 21925 3043
rect 21925 3009 21959 3043
rect 21959 3009 21968 3043
rect 21916 3000 21968 3009
rect 23112 3000 23164 3052
rect 28356 3136 28408 3188
rect 28448 3136 28500 3188
rect 30748 3136 30800 3188
rect 36268 3136 36320 3188
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 23572 3111 23624 3120
rect 23572 3077 23581 3111
rect 23581 3077 23615 3111
rect 23615 3077 23624 3111
rect 23572 3068 23624 3077
rect 27712 3068 27764 3120
rect 37464 3068 37516 3120
rect 27620 3000 27672 3052
rect 29000 3000 29052 3052
rect 29460 3043 29512 3052
rect 29460 3009 29469 3043
rect 29469 3009 29503 3043
rect 29503 3009 29512 3043
rect 29460 3000 29512 3009
rect 29552 3000 29604 3052
rect 32864 3000 32916 3052
rect 37740 3043 37792 3052
rect 37740 3009 37749 3043
rect 37749 3009 37783 3043
rect 37783 3009 37792 3043
rect 37740 3000 37792 3009
rect 37832 3000 37884 3052
rect 38752 3043 38804 3052
rect 38752 3009 38761 3043
rect 38761 3009 38795 3043
rect 38795 3009 38804 3043
rect 38752 3000 38804 3009
rect 38936 3000 38988 3052
rect 17040 2932 17092 2984
rect 15384 2839 15436 2848
rect 15384 2805 15393 2839
rect 15393 2805 15427 2839
rect 15427 2805 15436 2839
rect 15384 2796 15436 2805
rect 15568 2864 15620 2916
rect 16488 2864 16540 2916
rect 17960 2839 18012 2848
rect 17960 2805 17969 2839
rect 17969 2805 18003 2839
rect 18003 2805 18012 2839
rect 17960 2796 18012 2805
rect 22376 2932 22428 2984
rect 22744 2932 22796 2984
rect 25596 2932 25648 2984
rect 20904 2864 20956 2916
rect 26516 2864 26568 2916
rect 22192 2796 22244 2848
rect 22376 2796 22428 2848
rect 27896 2932 27948 2984
rect 29368 2907 29420 2916
rect 29368 2873 29377 2907
rect 29377 2873 29411 2907
rect 29411 2873 29420 2907
rect 29368 2864 29420 2873
rect 28172 2796 28224 2848
rect 30564 2864 30616 2916
rect 33140 2796 33192 2848
rect 38476 2839 38528 2848
rect 38476 2805 38485 2839
rect 38485 2805 38519 2839
rect 38519 2805 38528 2839
rect 38476 2796 38528 2805
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 1124 2524 1176 2576
rect 7012 2592 7064 2644
rect 14188 2592 14240 2644
rect 14280 2592 14332 2644
rect 14556 2592 14608 2644
rect 14648 2592 14700 2644
rect 23020 2567 23072 2576
rect 23020 2533 23029 2567
rect 23029 2533 23063 2567
rect 23063 2533 23072 2567
rect 23020 2524 23072 2533
rect 204 2388 256 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 1216 2320 1268 2372
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 7012 2431 7064 2440
rect 7012 2397 7021 2431
rect 7021 2397 7055 2431
rect 7055 2397 7064 2431
rect 7012 2388 7064 2397
rect 7472 2388 7524 2440
rect 8300 2388 8352 2440
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 18236 2456 18288 2508
rect 22008 2499 22060 2508
rect 22008 2465 22017 2499
rect 22017 2465 22051 2499
rect 22051 2465 22060 2499
rect 22008 2456 22060 2465
rect 33140 2456 33192 2508
rect 19524 2388 19576 2440
rect 22192 2320 22244 2372
rect 2596 2252 2648 2304
rect 3884 2252 3936 2304
rect 5264 2252 5316 2304
rect 6644 2252 6696 2304
rect 8024 2252 8076 2304
rect 9404 2252 9456 2304
rect 10784 2252 10836 2304
rect 21456 2252 21508 2304
rect 22376 2388 22428 2440
rect 27712 2388 27764 2440
rect 28448 2388 28500 2440
rect 36544 2388 36596 2440
rect 38108 2431 38160 2440
rect 38108 2397 38117 2431
rect 38117 2397 38151 2431
rect 38151 2397 38160 2431
rect 38108 2388 38160 2397
rect 38476 2431 38528 2440
rect 38476 2397 38485 2431
rect 38485 2397 38519 2431
rect 38519 2397 38528 2431
rect 38476 2388 38528 2397
rect 39396 2635 39448 2644
rect 39396 2601 39405 2635
rect 39405 2601 39439 2635
rect 39439 2601 39448 2635
rect 39396 2592 39448 2601
rect 25964 2320 26016 2372
rect 34152 2320 34204 2372
rect 28356 2295 28408 2304
rect 28356 2261 28365 2295
rect 28365 2261 28399 2295
rect 28399 2261 28408 2295
rect 28356 2252 28408 2261
rect 37924 2295 37976 2304
rect 37924 2261 37933 2295
rect 37933 2261 37967 2295
rect 37967 2261 37976 2295
rect 37924 2252 37976 2261
rect 38292 2295 38344 2304
rect 38292 2261 38301 2295
rect 38301 2261 38335 2295
rect 38335 2261 38344 2295
rect 38292 2252 38344 2261
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2252 40000 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 2872 2048 2924 2100
rect 10324 2048 10376 2100
rect 14556 2048 14608 2100
rect 28356 2048 28408 2100
rect 19064 1980 19116 2032
rect 31668 1980 31720 2032
rect 1676 1912 1728 1964
rect 29460 1912 29512 1964
rect 18512 1844 18564 1896
rect 38476 1912 38528 1964
rect 18696 1776 18748 1828
rect 38108 1776 38160 1828
rect 9772 1708 9824 1760
rect 29644 1708 29696 1760
rect 5724 1640 5776 1692
rect 21456 1640 21508 1692
rect 4252 1300 4304 1352
rect 38752 1300 38804 1352
rect 2504 1232 2556 1284
rect 28172 1232 28224 1284
rect 13820 1164 13872 1216
rect 38844 1164 38896 1216
rect 1584 1096 1636 1148
rect 21824 1096 21876 1148
rect 12256 8 12308 60
rect 37740 8 37792 60
<< metal2 >>
rect 3238 11194 3294 11250
rect 3514 11194 3570 11250
rect 3790 11194 3846 11250
rect 4066 11194 4122 11250
rect 4342 11194 4398 11250
rect 4618 11194 4674 11250
rect 4894 11194 4950 11250
rect 5170 11194 5226 11250
rect 5446 11194 5502 11250
rect 5722 11194 5778 11250
rect 5998 11194 6054 11250
rect 6274 11194 6330 11250
rect 6550 11194 6606 11250
rect 6826 11194 6882 11250
rect 7102 11194 7158 11250
rect 7378 11194 7434 11250
rect 7654 11194 7710 11250
rect 7930 11194 7986 11250
rect 8206 11194 8262 11250
rect 8482 11194 8538 11250
rect 8758 11194 8814 11250
rect 9034 11194 9090 11250
rect 9310 11194 9366 11250
rect 9586 11194 9642 11250
rect 9862 11194 9918 11250
rect 10138 11194 10194 11250
rect 10414 11194 10470 11250
rect 10690 11194 10746 11250
rect 10966 11194 11022 11250
rect 11242 11194 11298 11250
rect 11518 11194 11574 11250
rect 11794 11194 11850 11250
rect 12070 11194 12126 11250
rect 12346 11194 12402 11250
rect 12622 11194 12678 11250
rect 12898 11194 12954 11250
rect 13174 11194 13230 11250
rect 13450 11194 13506 11250
rect 13726 11194 13782 11250
rect 14002 11194 14058 11250
rect 14278 11194 14334 11250
rect 14554 11194 14610 11250
rect 14830 11194 14886 11250
rect 15106 11194 15162 11250
rect 15382 11194 15438 11250
rect 15658 11194 15714 11250
rect 15934 11194 15990 11250
rect 16210 11194 16266 11250
rect 16486 11194 16542 11250
rect 16762 11194 16818 11250
rect 17038 11194 17094 11250
rect 17314 11194 17370 11250
rect 17590 11194 17646 11250
rect 17866 11194 17922 11250
rect 18142 11194 18198 11250
rect 18418 11194 18474 11250
rect 18694 11194 18750 11250
rect 18970 11194 19026 11250
rect 19246 11194 19302 11250
rect 19522 11194 19578 11250
rect 19798 11194 19854 11250
rect 20074 11194 20130 11250
rect 20350 11194 20406 11250
rect 20626 11194 20682 11250
rect 20902 11194 20958 11250
rect 21178 11194 21234 11250
rect 21454 11194 21510 11250
rect 21730 11194 21786 11250
rect 22006 11194 22062 11250
rect 22282 11194 22338 11250
rect 22558 11194 22614 11250
rect 22834 11194 22890 11250
rect 23110 11194 23166 11250
rect 23386 11194 23442 11250
rect 23662 11194 23718 11250
rect 23938 11194 23994 11250
rect 24214 11194 24270 11250
rect 24490 11194 24546 11250
rect 24766 11194 24822 11250
rect 25042 11194 25098 11250
rect 25318 11194 25374 11250
rect 25594 11194 25650 11250
rect 25870 11194 25926 11250
rect 26146 11194 26202 11250
rect 26422 11194 26478 11250
rect 26698 11194 26754 11250
rect 26974 11212 27030 11250
rect 26974 11194 26976 11212
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 754 9616 810 9625
rect 754 9551 810 9560
rect 768 8498 796 9551
rect 938 9344 994 9353
rect 938 9279 994 9288
rect 756 8492 808 8498
rect 756 8434 808 8440
rect 570 8256 626 8265
rect 570 8191 626 8200
rect 584 7954 612 8191
rect 572 7948 624 7954
rect 572 7890 624 7896
rect 952 7818 980 9279
rect 1122 8528 1178 8537
rect 1122 8463 1178 8472
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 754 7440 810 7449
rect 1136 7410 1164 8463
rect 1214 7984 1270 7993
rect 1214 7919 1270 7928
rect 1228 7546 1256 7919
rect 1412 7886 1440 9823
rect 3252 9466 3280 11194
rect 3252 9438 3464 9466
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2608 8401 2636 8434
rect 2594 8392 2650 8401
rect 2594 8327 2650 8336
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1674 7984 1730 7993
rect 1674 7919 1730 7928
rect 1688 7886 1716 7919
rect 2792 7886 2820 9007
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 2884 7886 2912 8735
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 3436 8090 3464 9438
rect 3528 8634 3556 11194
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1216 7540 1268 7546
rect 1216 7482 1268 7488
rect 1320 7478 1348 7647
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 1308 7472 1360 7478
rect 1308 7414 1360 7420
rect 754 7375 810 7384
rect 1124 7404 1176 7410
rect 296 7336 348 7342
rect 296 7278 348 7284
rect 308 6905 336 7278
rect 294 6896 350 6905
rect 294 6831 350 6840
rect 768 6798 796 7375
rect 1124 7346 1176 7352
rect 2504 7200 2556 7206
rect 846 7168 902 7177
rect 2504 7142 2556 7148
rect 846 7103 902 7112
rect 860 6866 888 7103
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1216 6928 1268 6934
rect 1216 6870 1268 6876
rect 2318 6896 2374 6905
rect 848 6860 900 6866
rect 848 6802 900 6808
rect 756 6792 808 6798
rect 756 6734 808 6740
rect 1032 6724 1084 6730
rect 1032 6666 1084 6672
rect 1044 6633 1072 6666
rect 1030 6624 1086 6633
rect 1030 6559 1086 6568
rect 1228 6361 1256 6870
rect 2318 6831 2374 6840
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1214 6352 1270 6361
rect 1214 6287 1270 6296
rect 572 6248 624 6254
rect 572 6190 624 6196
rect 584 6089 612 6190
rect 570 6080 626 6089
rect 570 6015 626 6024
rect 202 5808 258 5817
rect 202 5743 258 5752
rect 848 5772 900 5778
rect 216 5710 244 5743
rect 848 5714 900 5720
rect 204 5704 256 5710
rect 204 5646 256 5652
rect 664 5636 716 5642
rect 664 5578 716 5584
rect 676 5545 704 5578
rect 662 5536 718 5545
rect 662 5471 718 5480
rect 860 5273 888 5714
rect 1596 5574 1624 6598
rect 1674 6352 1730 6361
rect 1674 6287 1676 6296
rect 1728 6287 1730 6296
rect 1676 6258 1728 6264
rect 1780 5642 1808 6598
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5914 2360 6831
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1872 5817 1900 5850
rect 1858 5808 1914 5817
rect 2516 5778 2544 7142
rect 3528 6746 3556 8434
rect 3620 7886 3648 8842
rect 3804 8362 3832 11194
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 4080 8090 4108 11194
rect 4356 8362 4384 11194
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4540 8498 4568 8978
rect 4632 8634 4660 11194
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4724 8498 4752 9386
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4908 8090 4936 11194
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 8498 5120 8774
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5184 8294 5212 11194
rect 5460 8634 5488 11194
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5552 8498 5580 10202
rect 5630 8936 5686 8945
rect 5630 8871 5686 8880
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3528 6718 3648 6746
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 3528 6458 3556 6598
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 1858 5743 1914 5752
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 3620 5710 3648 6718
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 1768 5636 1820 5642
rect 1768 5578 1820 5584
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 846 5264 902 5273
rect 388 5228 440 5234
rect 846 5199 902 5208
rect 388 5170 440 5176
rect 400 5001 428 5170
rect 848 5160 900 5166
rect 848 5102 900 5108
rect 2778 5128 2834 5137
rect 386 4992 442 5001
rect 386 4927 442 4936
rect 860 4729 888 5102
rect 2778 5063 2834 5072
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 846 4720 902 4729
rect 846 4655 902 4664
rect 756 4616 808 4622
rect 756 4558 808 4564
rect 768 4457 796 4558
rect 848 4548 900 4554
rect 848 4490 900 4496
rect 754 4448 810 4457
rect 754 4383 810 4392
rect 860 4185 888 4490
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 846 4176 902 4185
rect 388 4140 440 4146
rect 846 4111 902 4120
rect 388 4082 440 4088
rect 400 3913 428 4082
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 386 3904 442 3913
rect 386 3839 442 3848
rect 860 3641 888 4014
rect 846 3632 902 3641
rect 846 3567 902 3576
rect 1032 3596 1084 3602
rect 1032 3538 1084 3544
rect 204 3528 256 3534
rect 204 3470 256 3476
rect 216 3369 244 3470
rect 848 3460 900 3466
rect 848 3402 900 3408
rect 202 3360 258 3369
rect 202 3295 258 3304
rect 860 3097 888 3402
rect 846 3088 902 3097
rect 846 3023 902 3032
rect 756 2984 808 2990
rect 756 2926 808 2932
rect 388 2916 440 2922
rect 388 2858 440 2864
rect 204 2440 256 2446
rect 204 2382 256 2388
rect 216 2281 244 2382
rect 202 2272 258 2281
rect 202 2207 258 2216
rect 400 1737 428 2858
rect 768 2009 796 2926
rect 1044 2553 1072 3538
rect 1216 3052 1268 3058
rect 1216 2994 1268 3000
rect 1228 2825 1256 2994
rect 1214 2816 1270 2825
rect 1214 2751 1270 2760
rect 1124 2576 1176 2582
rect 1030 2544 1086 2553
rect 1124 2518 1176 2524
rect 1030 2479 1086 2488
rect 754 2000 810 2009
rect 754 1935 810 1944
rect 386 1728 442 1737
rect 386 1663 442 1672
rect 1136 56 1164 2518
rect 1216 2372 1268 2378
rect 1216 2314 1268 2320
rect 1228 1465 1256 2314
rect 1214 1456 1270 1465
rect 1214 1391 1270 1400
rect 1596 1154 1624 4422
rect 2410 3904 2466 3913
rect 1950 3836 2258 3845
rect 2410 3839 2466 3848
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2424 3670 2452 3839
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 1970 1716 2382
rect 1676 1964 1728 1970
rect 1676 1906 1728 1912
rect 2516 1290 2544 2926
rect 2792 2922 2820 5063
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3712 3942 3740 6666
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3804 3738 3832 4150
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3804 3534 3832 3674
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3896 3126 3924 7686
rect 5644 6866 5672 8871
rect 5736 8634 5764 11194
rect 5814 9480 5870 9489
rect 5814 9415 5870 9424
rect 5828 8634 5856 9415
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5460 6322 5488 6666
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3602 4016 4082
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 3238 2544 3294 2553
rect 3238 2479 3294 2488
rect 3252 2446 3280 2479
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2504 1284 2556 1290
rect 2504 1226 2556 1232
rect 2608 1170 2636 2246
rect 2884 2106 2912 2382
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 1584 1148 1636 1154
rect 1584 1090 1636 1096
rect 2516 1142 2636 1170
rect 2516 56 2544 1142
rect 3896 56 3924 2246
rect 4080 1737 4108 3878
rect 4066 1728 4122 1737
rect 4066 1663 4122 1672
rect 4264 1358 4292 4422
rect 4356 4146 4384 4490
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4356 3194 4384 4082
rect 4816 3534 4844 4966
rect 4908 4826 4936 4966
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4908 4146 4936 4422
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5000 3738 5028 4626
rect 5092 4282 5120 4762
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5184 3602 5212 4218
rect 5368 4214 5396 5034
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 5184 3058 5212 3538
rect 5368 3058 5396 4150
rect 5552 3942 5580 6734
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 5166 5764 6598
rect 5920 5370 5948 8910
rect 6012 8090 6040 11194
rect 6288 8634 6316 11194
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6564 8090 6592 11194
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6748 8498 6776 9930
rect 6840 8634 6868 11194
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 7116 8090 7144 11194
rect 7288 9240 7340 9246
rect 7288 9182 7340 9188
rect 7300 8498 7328 9182
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7392 8362 7420 11194
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5828 4690 5856 5170
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5920 4622 5948 4966
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5552 3505 5580 3606
rect 5538 3496 5594 3505
rect 5538 3431 5594 3440
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5644 2961 5672 3878
rect 5630 2952 5686 2961
rect 5630 2887 5686 2896
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 5276 56 5304 2246
rect 5736 1698 5764 4422
rect 5920 4282 5948 4558
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6012 4010 6040 7822
rect 6196 4049 6224 7890
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6254 6316 6734
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6288 4826 6316 6190
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6380 4593 6408 7958
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 6920 7880 6972 7886
rect 6918 7848 6920 7857
rect 7196 7880 7248 7886
rect 6972 7848 6974 7857
rect 7196 7822 7248 7828
rect 6918 7783 6974 7792
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6366 4584 6422 4593
rect 6366 4519 6422 4528
rect 6182 4040 6238 4049
rect 6000 4004 6052 4010
rect 6182 3975 6238 3984
rect 6000 3946 6052 3952
rect 6366 3224 6422 3233
rect 6184 3188 6236 3194
rect 6366 3159 6422 3168
rect 6184 3130 6236 3136
rect 6196 3097 6224 3130
rect 6182 3088 6238 3097
rect 6380 3058 6408 3159
rect 6182 3023 6238 3032
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5724 1692 5776 1698
rect 5724 1634 5776 1640
rect 6472 1601 6500 6666
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6656 5302 6684 6394
rect 7024 5846 7052 7278
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 6497 7144 6598
rect 7102 6488 7158 6497
rect 7102 6423 7158 6432
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6840 5681 6868 5782
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6826 5672 6882 5681
rect 6826 5607 6882 5616
rect 6828 5364 6880 5370
rect 6932 5352 6960 5714
rect 6932 5324 7052 5352
rect 6828 5306 6880 5312
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6642 4720 6698 4729
rect 6642 4655 6644 4664
rect 6696 4655 6698 4664
rect 6644 4626 6696 4632
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6656 4298 6684 4490
rect 6748 4486 6776 4558
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6656 4270 6776 4298
rect 6748 3738 6776 4270
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6656 2854 6684 3334
rect 6748 2990 6776 3674
rect 6840 3126 6868 5306
rect 7024 5030 7052 5324
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4554 7052 4966
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7116 4146 7144 5170
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7024 3738 7052 4082
rect 7208 3942 7236 7822
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7300 6730 7328 7142
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 4146 7328 4218
rect 7392 4185 7420 7890
rect 7484 4554 7512 9590
rect 7668 8650 7696 11194
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7576 8634 7696 8650
rect 7564 8628 7696 8634
rect 7616 8622 7696 8628
rect 7564 8570 7616 8576
rect 7852 8498 7880 10066
rect 7944 8634 7972 11194
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8128 8498 8156 9998
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7760 7002 7788 8434
rect 8220 8378 8248 11194
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8312 8566 8340 9046
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8404 8498 8432 9658
rect 8496 8634 8524 11194
rect 8666 9752 8722 9761
rect 8666 9687 8722 9696
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 7840 8356 7892 8362
rect 8220 8350 8340 8378
rect 7840 8298 7892 8304
rect 7852 7274 7880 8298
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8312 8090 8340 8350
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7546 7972 7958
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7930 7440 7986 7449
rect 7930 7375 7932 7384
rect 7984 7375 7986 7384
rect 7932 7346 7984 7352
rect 8220 7313 8248 7754
rect 8404 7426 8432 8230
rect 8312 7410 8432 7426
rect 8300 7404 8432 7410
rect 8352 7398 8432 7404
rect 8300 7346 8352 7352
rect 8206 7304 8262 7313
rect 7840 7268 7892 7274
rect 8206 7239 8262 7248
rect 7840 7210 7892 7216
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7564 6928 7616 6934
rect 8484 6928 8536 6934
rect 7564 6870 7616 6876
rect 7668 6876 8484 6882
rect 7668 6870 8536 6876
rect 7576 5778 7604 6870
rect 7668 6854 8524 6870
rect 7668 6798 7696 6854
rect 7656 6792 7708 6798
rect 8024 6792 8076 6798
rect 7656 6734 7708 6740
rect 8022 6760 8024 6769
rect 8116 6792 8168 6798
rect 8076 6760 8078 6769
rect 8116 6734 8168 6740
rect 8022 6695 8078 6704
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6458 7696 6598
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 8128 6118 8156 6734
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7562 5264 7618 5273
rect 7562 5199 7564 5208
rect 7616 5199 7618 5208
rect 7564 5170 7616 5176
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7378 4176 7434 4185
rect 7288 4140 7340 4146
rect 7378 4111 7434 4120
rect 7288 4082 7340 4088
rect 7196 3936 7248 3942
rect 7288 3936 7340 3942
rect 7196 3878 7248 3884
rect 7286 3904 7288 3913
rect 7340 3904 7342 3913
rect 7286 3839 7342 3848
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6932 3369 6960 3606
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7484 3482 7512 4490
rect 7576 3602 7604 5170
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7668 3641 7696 4014
rect 7654 3632 7710 3641
rect 7564 3596 7616 3602
rect 7654 3567 7710 3576
rect 7564 3538 7616 3544
rect 7656 3528 7708 3534
rect 7484 3476 7656 3482
rect 7484 3470 7708 3476
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 7392 3194 7420 3470
rect 7484 3454 7696 3470
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7024 2446 7052 2586
rect 7484 2446 7512 3334
rect 7576 3233 7604 3454
rect 7562 3224 7618 3233
rect 7562 3159 7618 3168
rect 7760 3176 7788 5646
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 3670 7880 4422
rect 8220 4146 8248 4490
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7840 3188 7892 3194
rect 7760 3148 7840 3176
rect 7840 3130 7892 3136
rect 8206 3088 8262 3097
rect 8206 3023 8262 3032
rect 8220 2990 8248 3023
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8312 2446 8340 6598
rect 8392 6316 8444 6322
rect 8496 6304 8524 6854
rect 8444 6276 8524 6304
rect 8392 6258 8444 6264
rect 8588 6066 8616 8774
rect 8680 7954 8708 9687
rect 8772 8090 8800 11194
rect 9048 9500 9076 11194
rect 8864 9472 9076 9500
rect 8864 8634 8892 9472
rect 9324 8922 9352 11194
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9324 8894 9444 8922
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9416 8090 9444 8894
rect 9508 8498 9536 9862
rect 9600 8634 9628 11194
rect 9680 9784 9732 9790
rect 9680 9726 9732 9732
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8666 7440 8722 7449
rect 8666 7375 8722 7384
rect 8680 6254 8708 7375
rect 8758 6488 8814 6497
rect 8758 6423 8814 6432
rect 8772 6254 8800 6423
rect 8864 6254 8892 7686
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9600 7562 9628 8434
rect 9692 8430 9720 9726
rect 9772 9104 9824 9110
rect 9770 9072 9772 9081
rect 9824 9072 9826 9081
rect 9770 9007 9826 9016
rect 9876 8634 9904 11194
rect 9956 10328 10008 10334
rect 9956 10270 10008 10276
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9508 7534 9628 7562
rect 9218 7440 9274 7449
rect 9218 7375 9220 7384
rect 9272 7375 9274 7384
rect 9220 7346 9272 7352
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8956 7002 8984 7210
rect 9324 7002 9352 7278
rect 9508 7018 9536 7534
rect 9692 7426 9720 7890
rect 9968 7886 9996 10270
rect 10048 9852 10100 9858
rect 10048 9794 10100 9800
rect 10060 8634 10088 9794
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9600 7398 9720 7426
rect 9600 7206 9628 7398
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9312 6996 9364 7002
rect 9508 6990 9628 7018
rect 9312 6938 9364 6944
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9402 6760 9458 6769
rect 9402 6695 9458 6704
rect 9416 6662 9444 6695
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9010 6556 9318 6565
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9508 6322 9536 6802
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8668 6112 8720 6118
rect 8588 6060 8668 6066
rect 8588 6054 8720 6060
rect 8588 6038 8708 6054
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8404 4865 8432 5782
rect 8864 5710 8892 6190
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 8390 4856 8446 4865
rect 8390 4791 8446 4800
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 9600 4162 9628 6990
rect 9692 5914 9720 7278
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9508 4134 9628 4162
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8404 3058 8432 3470
rect 8852 3392 8904 3398
rect 8850 3360 8852 3369
rect 8904 3360 8906 3369
rect 8850 3295 8906 3304
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 9010 3227 9318 3236
rect 8484 3120 8536 3126
rect 8482 3088 8484 3097
rect 8536 3088 8538 3097
rect 8392 3052 8444 3058
rect 8482 3023 8538 3032
rect 9312 3052 9364 3058
rect 8392 2994 8444 3000
rect 9416 3040 9444 4082
rect 9508 3890 9536 4134
rect 9586 4040 9642 4049
rect 9586 3975 9588 3984
rect 9640 3975 9642 3984
rect 9588 3946 9640 3952
rect 9508 3862 9628 3890
rect 9600 3738 9628 3862
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9508 3233 9536 3674
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9494 3224 9550 3233
rect 9494 3159 9550 3168
rect 9364 3012 9444 3040
rect 9312 2994 9364 3000
rect 9600 2990 9628 3334
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9312 2848 9364 2854
rect 9692 2802 9720 5714
rect 9784 3738 9812 7686
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6798 9904 7142
rect 10060 6866 10088 8230
rect 10152 8090 10180 11194
rect 10230 9888 10286 9897
rect 10230 9823 10286 9832
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10244 7886 10272 9823
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10336 8566 10364 9046
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10428 8090 10456 11194
rect 10506 9344 10562 9353
rect 10506 9279 10562 9288
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 10152 6390 10180 7142
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10244 5658 10272 7686
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 6458 10456 6802
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10152 5630 10272 5658
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9784 2922 9812 3470
rect 9876 3194 9904 3470
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10060 3058 10088 3402
rect 10152 3398 10180 5630
rect 10428 5574 10456 6258
rect 10520 6254 10548 9279
rect 10704 8634 10732 11194
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10796 7886 10824 10134
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 7954 10916 9454
rect 10980 8634 11008 11194
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11072 8498 11100 8910
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10244 3602 10272 4626
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10244 2990 10272 3538
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9364 2796 9720 2802
rect 9312 2790 9720 2796
rect 9324 2774 9720 2790
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 6458 1592 6514 1601
rect 6458 1527 6514 1536
rect 6656 56 6684 2246
rect 8036 56 8064 2246
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9416 56 9444 2246
rect 9784 1766 9812 2382
rect 10336 2106 10364 4422
rect 10428 3602 10456 4422
rect 10520 4214 10548 4762
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10520 2990 10548 4014
rect 10612 4010 10640 7142
rect 10888 6866 10916 7890
rect 10980 7721 11008 8434
rect 11256 8090 11284 11194
rect 11426 9208 11482 9217
rect 11426 9143 11482 9152
rect 11440 9042 11468 9143
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11532 8634 11560 11194
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11426 8392 11482 8401
rect 11426 8327 11482 8336
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 10966 7712 11022 7721
rect 10966 7647 11022 7656
rect 11440 6934 11468 8327
rect 11808 8090 11836 11194
rect 12084 8634 12112 11194
rect 12360 8634 12388 11194
rect 12532 9308 12584 9314
rect 12532 9250 12584 9256
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12544 8566 12572 9250
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12636 8090 12664 11194
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12728 8498 12756 9454
rect 12912 8634 12940 11194
rect 13188 8634 13216 11194
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13280 8514 13308 8774
rect 13188 8498 13308 8514
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 13176 8492 13308 8498
rect 13228 8486 13308 8492
rect 13176 8434 13228 8440
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11900 7449 11928 7482
rect 11886 7440 11942 7449
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11612 7404 11664 7410
rect 11886 7375 11942 7384
rect 11612 7346 11664 7352
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 11532 6798 11560 7346
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11072 6458 11100 6734
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11624 6322 11652 7346
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 11808 6866 11836 7278
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11702 6760 11758 6769
rect 11808 6730 11836 6802
rect 11702 6695 11758 6704
rect 11796 6724 11848 6730
rect 11716 6662 11744 6695
rect 11796 6666 11848 6672
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11704 6248 11756 6254
rect 11808 6236 11836 6666
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11756 6208 11836 6236
rect 11704 6190 11756 6196
rect 10692 6112 10744 6118
rect 11060 6112 11112 6118
rect 10692 6054 10744 6060
rect 10782 6080 10838 6089
rect 10704 5914 10732 6054
rect 11060 6054 11112 6060
rect 10782 6015 10838 6024
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5778 10824 6015
rect 11072 5846 11100 6054
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11152 5840 11204 5846
rect 11204 5800 11284 5828
rect 11152 5782 11204 5788
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5409 10824 5578
rect 11164 5574 11192 5646
rect 11256 5642 11284 5800
rect 11900 5778 11928 6394
rect 12268 6118 12296 7278
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12256 6112 12308 6118
rect 12452 6089 12480 6258
rect 12820 6225 12848 6598
rect 12912 6254 12940 6734
rect 13004 6458 13032 7278
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12900 6248 12952 6254
rect 12806 6216 12862 6225
rect 12900 6190 12952 6196
rect 12806 6151 12862 6160
rect 12256 6054 12308 6060
rect 12438 6080 12494 6089
rect 12438 6015 12494 6024
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10782 5400 10838 5409
rect 10782 5335 10838 5344
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10980 4282 11008 4558
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 10784 4072 10836 4078
rect 11348 4060 11376 5578
rect 11716 5574 11744 5646
rect 11704 5568 11756 5574
rect 12452 5545 12480 5714
rect 12912 5574 12940 6190
rect 12900 5568 12952 5574
rect 11704 5510 11756 5516
rect 12438 5536 12494 5545
rect 11520 4820 11572 4826
rect 11440 4780 11520 4808
rect 11440 4690 11468 4780
rect 11520 4762 11572 4768
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11440 4078 11468 4626
rect 10784 4014 10836 4020
rect 11072 4032 11376 4060
rect 11428 4072 11480 4078
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10796 3670 10824 4014
rect 11072 3942 11100 4032
rect 11428 4014 11480 4020
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 11164 3534 11192 3878
rect 11440 3618 11468 4014
rect 11348 3590 11468 3618
rect 11348 3534 11376 3590
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11440 3126 11468 3470
rect 11532 3194 11560 4626
rect 11716 4214 11744 5510
rect 12900 5510 12952 5516
rect 12438 5471 12494 5480
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11992 4690 12020 5238
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12162 4720 12218 4729
rect 11980 4684 12032 4690
rect 12162 4655 12164 4664
rect 11980 4626 12032 4632
rect 12216 4655 12218 4664
rect 12164 4626 12216 4632
rect 11992 4486 12020 4626
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 12162 4176 12218 4185
rect 12162 4111 12218 4120
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11992 3058 12020 3402
rect 12176 3398 12204 4111
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12164 3120 12216 3126
rect 12162 3088 12164 3097
rect 12216 3088 12218 3097
rect 11980 3052 12032 3058
rect 12268 3058 12296 5170
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12360 4146 12388 5102
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12346 3904 12402 3913
rect 12346 3839 12402 3848
rect 12360 3097 12388 3839
rect 12452 3738 12480 5102
rect 13096 5098 13124 8366
rect 13464 8090 13492 11194
rect 13740 8634 13768 11194
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 14016 8362 14044 11194
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 14292 8090 14320 11194
rect 14568 8634 14596 11194
rect 14738 10024 14794 10033
rect 14738 9959 14794 9968
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14660 8498 14688 9046
rect 14752 8566 14780 9959
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5710 13216 6258
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13280 5642 13308 6734
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13556 5574 13584 7686
rect 13648 7206 13676 7686
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4826 13216 5034
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12544 4146 12572 4218
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12346 3088 12402 3097
rect 12162 3023 12218 3032
rect 12256 3052 12308 3058
rect 11980 2994 12032 3000
rect 12346 3023 12402 3032
rect 12256 2994 12308 3000
rect 12544 2990 12572 4082
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 10796 56 10824 2246
rect 12176 66 12296 82
rect 12176 60 12308 66
rect 12176 56 12256 60
rect 1122 0 1178 56
rect 2502 0 2558 56
rect 3882 0 3938 56
rect 5262 0 5318 56
rect 6642 0 6698 56
rect 8022 0 8078 56
rect 9402 0 9458 56
rect 10782 0 10838 56
rect 12162 54 12256 56
rect 12162 0 12218 54
rect 13556 56 13584 5170
rect 13648 3738 13676 6054
rect 13740 5370 13768 8026
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14200 7970 14228 8026
rect 14464 8016 14516 8022
rect 14200 7964 14464 7970
rect 14200 7958 14516 7964
rect 14108 7886 14136 7958
rect 14200 7942 14504 7958
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14280 7880 14332 7886
rect 14332 7840 14412 7868
rect 14280 7822 14332 7828
rect 13832 5794 13860 7822
rect 14384 7342 14412 7840
rect 14372 7336 14424 7342
rect 14424 7296 14504 7324
rect 14372 7278 14424 7284
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14370 7032 14426 7041
rect 14370 6967 14426 6976
rect 14188 6724 14240 6730
rect 14384 6712 14412 6967
rect 14240 6684 14412 6712
rect 14188 6666 14240 6672
rect 14476 6633 14504 7296
rect 14462 6624 14518 6633
rect 14462 6559 14518 6568
rect 14660 6338 14688 8298
rect 14844 8090 14872 11194
rect 15120 8922 15148 11194
rect 14936 8894 15148 8922
rect 14936 8634 14964 8894
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 15396 8634 15424 11194
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14752 7721 14780 7890
rect 14738 7712 14794 7721
rect 14738 7647 14794 7656
rect 14936 7274 14964 8366
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15396 7410 15424 7686
rect 15580 7546 15608 9114
rect 15672 8634 15700 11194
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15764 7546 15792 9318
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 8090 15884 8434
rect 15948 8090 15976 11194
rect 16224 8634 16252 11194
rect 16304 9308 16356 9314
rect 16304 9250 16356 9256
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14844 6798 14872 7142
rect 15028 6798 15056 7278
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 15016 6792 15068 6798
rect 15212 6746 15240 6870
rect 15396 6866 15424 7346
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15068 6740 15240 6746
rect 15016 6734 15240 6740
rect 14752 6458 14780 6734
rect 14844 6633 14872 6734
rect 15028 6718 15240 6734
rect 14830 6624 14886 6633
rect 14830 6559 14886 6568
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14660 6310 14780 6338
rect 14844 6322 14872 6559
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 14464 6248 14516 6254
rect 14648 6248 14700 6254
rect 14516 6196 14596 6202
rect 14464 6190 14596 6196
rect 14648 6190 14700 6196
rect 14476 6174 14596 6190
rect 14568 6118 14596 6174
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 13832 5766 14320 5794
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13726 4856 13782 4865
rect 13726 4791 13782 4800
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3398 13768 4791
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13728 2984 13780 2990
rect 13726 2952 13728 2961
rect 13780 2952 13782 2961
rect 13726 2887 13782 2896
rect 13832 1222 13860 5578
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 14292 2650 14320 5766
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14200 2530 14228 2586
rect 14476 2530 14504 6054
rect 14660 5914 14688 6190
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14752 5710 14780 6310
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 15200 6248 15252 6254
rect 15198 6216 15200 6225
rect 15252 6216 15254 6225
rect 15396 6186 15424 6802
rect 15488 6662 15516 7346
rect 16026 7168 16082 7177
rect 16026 7103 16082 7112
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15658 6216 15714 6225
rect 15198 6151 15254 6160
rect 15384 6180 15436 6186
rect 15658 6151 15714 6160
rect 15384 6122 15436 6128
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 15672 5642 15700 6151
rect 15764 5642 15792 6734
rect 16040 6662 16068 7103
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16132 6118 16160 8434
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16224 7750 16252 7890
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16316 7410 16344 9250
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 7546 16436 8774
rect 16500 8634 16528 11194
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16592 8514 16620 8774
rect 16776 8634 16804 11194
rect 17052 9246 17080 11194
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17040 9240 17092 9246
rect 17040 9182 17092 9188
rect 17236 9178 17264 9590
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17328 8634 17356 11194
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 16500 8486 16620 8514
rect 17132 8492 17184 8498
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6934 16344 7346
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6322 16252 6734
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 14648 5568 14700 5574
rect 14740 5568 14792 5574
rect 14648 5510 14700 5516
rect 14738 5536 14740 5545
rect 14792 5536 14794 5545
rect 14660 2650 14688 5510
rect 14738 5471 14794 5480
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 14830 5400 14886 5409
rect 15010 5403 15318 5412
rect 14830 5335 14886 5344
rect 15566 5400 15622 5409
rect 15566 5335 15622 5344
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14752 2774 14780 4626
rect 14844 4622 14872 5335
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 15396 4486 15424 4966
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 14830 4176 14886 4185
rect 14830 4111 14886 4120
rect 14844 3534 14872 4111
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15304 3641 15332 3946
rect 15290 3632 15346 3641
rect 15290 3567 15346 3576
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 15292 3460 15344 3466
rect 15396 3448 15424 4422
rect 15474 4040 15530 4049
rect 15474 3975 15476 3984
rect 15528 3975 15530 3984
rect 15476 3946 15528 3952
rect 15580 3670 15608 5335
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 15658 4312 15714 4321
rect 15658 4247 15714 4256
rect 15672 3942 15700 4247
rect 16224 4146 16252 4558
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15344 3420 15424 3448
rect 15292 3402 15344 3408
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 15672 3097 15700 3334
rect 15658 3088 15714 3097
rect 15842 3088 15898 3097
rect 15658 3023 15714 3032
rect 15764 3046 15842 3074
rect 15764 2990 15792 3046
rect 16040 3058 16068 3538
rect 15842 3023 15898 3032
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15752 2984 15804 2990
rect 15396 2922 15608 2938
rect 15844 2984 15896 2990
rect 15752 2926 15804 2932
rect 15842 2952 15844 2961
rect 15896 2952 15898 2961
rect 15396 2916 15620 2922
rect 15396 2910 15568 2916
rect 15396 2854 15424 2910
rect 16500 2922 16528 8486
rect 17132 8434 17184 8440
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16684 5574 16712 6054
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16776 5574 16804 5714
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 4078 16804 5510
rect 16854 4584 16910 4593
rect 16854 4519 16856 4528
rect 16908 4519 16910 4528
rect 16856 4490 16908 4496
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16592 3738 16620 4014
rect 17144 3913 17172 8434
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17236 8022 17264 8230
rect 17604 8090 17632 11194
rect 17880 9602 17908 11194
rect 18156 9602 18184 11194
rect 17880 9574 18000 9602
rect 18156 9574 18276 9602
rect 17868 9240 17920 9246
rect 17868 9182 17920 9188
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17788 8498 17816 8978
rect 17880 8634 17908 9182
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17972 7886 18000 9574
rect 18248 7886 18276 9574
rect 18432 8498 18460 11194
rect 18602 9208 18658 9217
rect 18602 9143 18658 9152
rect 18616 9042 18644 9143
rect 18604 9036 18656 9042
rect 18604 8978 18656 8984
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18524 8634 18552 8910
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18708 8498 18736 11194
rect 18880 9784 18932 9790
rect 18880 9726 18932 9732
rect 18788 9240 18840 9246
rect 18788 9182 18840 9188
rect 18800 8566 18828 9182
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18708 8090 18736 8298
rect 18788 8288 18840 8294
rect 18786 8256 18788 8265
rect 18840 8256 18842 8265
rect 18786 8191 18842 8200
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 17960 7744 18012 7750
rect 17222 7712 17278 7721
rect 17960 7686 18012 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17222 7647 17278 7656
rect 17236 7313 17264 7647
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17222 7304 17278 7313
rect 17222 7239 17278 7248
rect 17788 6730 17816 7346
rect 17972 6866 18000 7686
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17788 5137 17816 6666
rect 17972 5846 18000 6666
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18064 5166 18092 7686
rect 18328 7336 18380 7342
rect 18326 7304 18328 7313
rect 18380 7304 18382 7313
rect 18326 7239 18382 7248
rect 18340 7041 18368 7239
rect 18326 7032 18382 7041
rect 18326 6967 18382 6976
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 6322 18276 6734
rect 18340 6662 18368 6967
rect 18892 6934 18920 9726
rect 18984 8498 19012 11194
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18880 6928 18932 6934
rect 18880 6870 18932 6876
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18694 6624 18750 6633
rect 18694 6559 18750 6568
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18052 5160 18104 5166
rect 17774 5128 17830 5137
rect 18052 5102 18104 5108
rect 17774 5063 17830 5072
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17130 3904 17186 3913
rect 17130 3839 17186 3848
rect 17696 3738 17724 4218
rect 17880 4078 17908 4490
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17958 4040 18014 4049
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17592 3596 17644 3602
rect 17328 3556 17592 3584
rect 16948 3528 17000 3534
rect 17132 3528 17184 3534
rect 16948 3470 17000 3476
rect 17052 3488 17132 3516
rect 16960 3369 16988 3470
rect 16946 3360 17002 3369
rect 16946 3295 17002 3304
rect 17052 2990 17080 3488
rect 17132 3470 17184 3476
rect 17328 3058 17356 3556
rect 17592 3538 17644 3544
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17420 3058 17448 3130
rect 17696 3058 17724 3674
rect 17880 3534 17908 4014
rect 17958 3975 18014 3984
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17776 3392 17828 3398
rect 17880 3369 17908 3470
rect 17776 3334 17828 3340
rect 17866 3360 17922 3369
rect 17788 3058 17816 3334
rect 17866 3295 17922 3304
rect 17880 3058 17908 3295
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 15842 2887 15898 2896
rect 16488 2916 16540 2922
rect 15568 2858 15620 2864
rect 16488 2858 16540 2864
rect 15384 2848 15436 2854
rect 17420 2825 17448 2994
rect 17972 2854 18000 3975
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 18064 3448 18092 3606
rect 18144 3460 18196 3466
rect 18064 3420 18144 3448
rect 18144 3402 18196 3408
rect 17960 2848 18012 2854
rect 15384 2790 15436 2796
rect 17406 2816 17462 2825
rect 14752 2746 14964 2774
rect 17960 2790 18012 2796
rect 17406 2751 17462 2760
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14200 2502 14504 2530
rect 14568 2106 14596 2586
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 13820 1216 13872 1222
rect 13820 1158 13872 1164
rect 14936 56 14964 2746
rect 18248 2514 18276 6258
rect 18708 6254 18736 6559
rect 18970 6488 19026 6497
rect 18970 6423 18972 6432
rect 19024 6423 19026 6432
rect 18972 6394 19024 6400
rect 19076 6254 19104 7142
rect 19168 6458 19196 8570
rect 19260 8522 19288 11194
rect 19536 10418 19564 11194
rect 19432 10396 19484 10402
rect 19536 10390 19656 10418
rect 19432 10338 19484 10344
rect 19338 10160 19394 10169
rect 19338 10095 19394 10104
rect 19352 9926 19380 10095
rect 19444 9994 19472 10338
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19248 8516 19300 8522
rect 19248 8458 19300 8464
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19260 8265 19288 8366
rect 19246 8256 19302 8265
rect 19246 8191 19302 8200
rect 19352 7478 19380 8570
rect 19628 8498 19656 10390
rect 19812 8498 19840 11194
rect 19890 10160 19946 10169
rect 19890 10095 19946 10104
rect 19904 9926 19932 10095
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 20088 9874 20116 11194
rect 20364 9874 20392 11194
rect 20088 9846 20208 9874
rect 20364 9846 20484 9874
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19904 8294 19932 9386
rect 20180 8498 20208 9846
rect 20258 8664 20314 8673
rect 20258 8599 20260 8608
rect 20312 8599 20314 8608
rect 20260 8570 20312 8576
rect 20456 8498 20484 9846
rect 20640 8634 20668 11194
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20824 8566 20852 8842
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20916 8498 20944 11194
rect 21192 9874 21220 11194
rect 21192 9846 21404 9874
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 21376 8498 21404 9846
rect 21468 8498 21496 11194
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20812 8356 20864 8362
rect 20996 8356 21048 8362
rect 20812 8298 20864 8304
rect 20916 8316 20996 8344
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19892 8288 19944 8294
rect 20364 8265 20392 8298
rect 19892 8230 19944 8236
rect 20350 8256 20406 8265
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19260 6202 19288 6598
rect 19352 6322 19380 7278
rect 19444 7041 19472 8230
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19628 7342 19656 7822
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19628 7041 19656 7142
rect 19430 7032 19486 7041
rect 19430 6967 19486 6976
rect 19614 7032 19670 7041
rect 19614 6967 19670 6976
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19536 6322 19564 6802
rect 19628 6372 19656 6870
rect 19720 6474 19748 7686
rect 19812 7585 19840 8230
rect 19950 8188 20258 8197
rect 20350 8191 20406 8200
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20824 8129 20852 8298
rect 20810 8120 20866 8129
rect 20260 8084 20312 8090
rect 20810 8055 20866 8064
rect 20260 8026 20312 8032
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19798 7576 19854 7585
rect 19798 7511 19854 7520
rect 19996 7274 20024 7890
rect 20272 7818 20300 8026
rect 20456 7908 20852 7936
rect 20352 7880 20404 7886
rect 20456 7868 20484 7908
rect 20404 7840 20484 7868
rect 20718 7848 20774 7857
rect 20352 7822 20404 7828
rect 20260 7812 20312 7818
rect 20718 7783 20774 7792
rect 20260 7754 20312 7760
rect 20732 7750 20760 7783
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 20364 7206 20392 7482
rect 20444 7404 20496 7410
rect 20548 7392 20576 7482
rect 20496 7364 20576 7392
rect 20720 7404 20772 7410
rect 20444 7346 20496 7352
rect 20824 7392 20852 7908
rect 20772 7364 20852 7392
rect 20720 7346 20772 7352
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19950 7035 20258 7044
rect 20364 6866 20392 7142
rect 20732 7041 20760 7346
rect 20810 7304 20866 7313
rect 20810 7239 20866 7248
rect 20718 7032 20774 7041
rect 20718 6967 20774 6976
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20076 6792 20128 6798
rect 20128 6752 20208 6780
rect 20076 6734 20128 6740
rect 20180 6474 20208 6752
rect 20272 6746 20300 6802
rect 20824 6746 20852 7239
rect 20916 6866 20944 8316
rect 20996 8298 21048 8304
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21010 7644 21318 7653
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21376 7342 21404 8230
rect 21088 7336 21140 7342
rect 21086 7304 21088 7313
rect 21364 7336 21416 7342
rect 21140 7304 21142 7313
rect 21364 7278 21416 7284
rect 21086 7239 21142 7248
rect 21270 7032 21326 7041
rect 21270 6967 21326 6976
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21192 6746 21220 6802
rect 21284 6798 21312 6967
rect 20272 6718 20852 6746
rect 20916 6718 21220 6746
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 20444 6656 20496 6662
rect 20628 6656 20680 6662
rect 20496 6616 20576 6644
rect 20444 6598 20496 6604
rect 19720 6446 19932 6474
rect 20180 6446 20392 6474
rect 19628 6344 19840 6372
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19812 6254 19840 6344
rect 19614 6248 19666 6254
rect 19260 6196 19614 6202
rect 19260 6190 19666 6196
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 18512 6180 18564 6186
rect 19260 6174 19654 6190
rect 18512 6122 18564 6128
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 3534 18368 4422
rect 18418 4312 18474 4321
rect 18418 4247 18474 4256
rect 18432 4146 18460 4247
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 18524 1902 18552 6122
rect 19904 6100 19932 6446
rect 20260 6384 20312 6390
rect 20088 6344 20260 6372
rect 20088 6100 20116 6344
rect 20260 6326 20312 6332
rect 19904 6072 20116 6100
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19338 5944 19394 5953
rect 19950 5947 20258 5956
rect 20364 5914 20392 6446
rect 20548 6322 20576 6616
rect 20628 6598 20680 6604
rect 20810 6624 20866 6633
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20640 6118 20668 6598
rect 20916 6610 20944 6718
rect 20866 6582 20944 6610
rect 20810 6559 20866 6568
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 20810 6488 20866 6497
rect 21010 6491 21318 6500
rect 20810 6423 20812 6432
rect 20864 6423 20866 6432
rect 20812 6394 20864 6400
rect 21376 6322 21404 7278
rect 21468 6458 21496 8298
rect 21560 6866 21588 8366
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 20824 6202 20852 6258
rect 20732 6174 20852 6202
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 19338 5879 19394 5888
rect 20352 5908 20404 5914
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18616 4622 18644 5646
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18616 4282 18644 4558
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18512 1896 18564 1902
rect 18512 1838 18564 1844
rect 18708 1834 18736 5782
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19168 5545 19196 5714
rect 19154 5536 19210 5545
rect 19154 5471 19210 5480
rect 19352 5302 19380 5879
rect 20352 5850 20404 5856
rect 19524 5704 19576 5710
rect 19522 5672 19524 5681
rect 19576 5672 19578 5681
rect 19522 5607 19578 5616
rect 20534 5672 20590 5681
rect 20534 5607 20590 5616
rect 20548 5574 20576 5607
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20456 5370 20484 5510
rect 20732 5370 20760 6174
rect 20916 5778 20944 6258
rect 21468 6254 21496 6394
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 20810 5536 20866 5545
rect 20810 5471 20866 5480
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 20350 5264 20406 5273
rect 20824 5234 20852 5471
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 20350 5199 20406 5208
rect 20812 5228 20864 5234
rect 18880 5160 18932 5166
rect 18786 5128 18842 5137
rect 18880 5102 18932 5108
rect 18786 5063 18842 5072
rect 18800 4486 18828 5063
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18892 3942 18920 5102
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 20364 4865 20392 5199
rect 20812 5170 20864 5176
rect 21364 5024 21416 5030
rect 20902 4992 20958 5001
rect 21364 4966 21416 4972
rect 20902 4927 20958 4936
rect 20350 4856 20406 4865
rect 20350 4791 20406 4800
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 19076 4214 19104 4626
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 18880 3936 18932 3942
rect 19812 3913 19840 4014
rect 20364 3913 20392 4014
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 18880 3878 18932 3884
rect 19798 3904 19854 3913
rect 19798 3839 19854 3848
rect 20350 3904 20406 3913
rect 19950 3836 20258 3845
rect 20350 3839 20406 3848
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20732 3670 20760 3946
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20916 2922 20944 4927
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 21376 4078 21404 4966
rect 21468 4758 21496 5578
rect 21560 5302 21588 6666
rect 21652 5953 21680 9318
rect 21744 8566 21772 11194
rect 22020 8634 22048 11194
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21638 5944 21694 5953
rect 21638 5879 21694 5888
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 21560 4554 21588 5238
rect 21744 4842 21772 8298
rect 21836 6458 21864 8570
rect 22296 8566 22324 11194
rect 22572 8634 22600 11194
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22848 8566 22876 11194
rect 23124 8634 23152 11194
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 22284 8560 22336 8566
rect 22284 8502 22336 8508
rect 22836 8560 22888 8566
rect 22836 8502 22888 8508
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22836 8288 22888 8294
rect 22836 8230 22888 8236
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21928 7750 21956 7958
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21822 6080 21878 6089
rect 21822 6015 21878 6024
rect 21652 4814 21772 4842
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21192 3602 21220 4014
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 21468 3398 21496 4150
rect 21652 4010 21680 4814
rect 21836 4690 21864 6015
rect 21928 5846 21956 7346
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22020 6798 22048 7278
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22112 6662 22140 6734
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 6361 22140 6598
rect 22098 6352 22154 6361
rect 22098 6287 22154 6296
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 22296 5250 22324 8230
rect 22388 7410 22416 8230
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22558 7304 22614 7313
rect 22558 7239 22614 7248
rect 22572 7002 22600 7239
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22296 5222 22416 5250
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 21824 4684 21876 4690
rect 22192 4684 22244 4690
rect 21824 4626 21876 4632
rect 22112 4644 22192 4672
rect 21836 4486 21864 4626
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21640 4004 21692 4010
rect 21640 3946 21692 3952
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21548 3460 21600 3466
rect 21548 3402 21600 3408
rect 21456 3392 21508 3398
rect 21560 3369 21588 3402
rect 21640 3392 21692 3398
rect 21456 3334 21508 3340
rect 21546 3360 21602 3369
rect 21640 3334 21692 3340
rect 21010 3292 21318 3301
rect 21546 3295 21602 3304
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 21652 3194 21680 3334
rect 21744 3233 21772 3878
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 21730 3224 21786 3233
rect 21640 3188 21692 3194
rect 21730 3159 21786 3168
rect 21640 3130 21692 3136
rect 21928 3058 21956 3470
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19522 2680 19578 2689
rect 19950 2683 20258 2692
rect 19522 2615 19578 2624
rect 19536 2446 19564 2615
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 21468 2310 21496 2994
rect 21928 2774 21956 2994
rect 22020 2825 22048 4082
rect 22112 3602 22140 4644
rect 22192 4626 22244 4632
rect 22192 3936 22244 3942
rect 22190 3904 22192 3913
rect 22244 3904 22246 3913
rect 22190 3839 22246 3848
rect 22296 3602 22324 4762
rect 22388 4214 22416 5222
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22572 4486 22600 4558
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22374 3768 22430 3777
rect 22374 3703 22430 3712
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22100 3392 22152 3398
rect 22284 3392 22336 3398
rect 22152 3352 22284 3380
rect 22100 3334 22152 3340
rect 22284 3334 22336 3340
rect 22388 2990 22416 3703
rect 22480 3126 22508 4422
rect 22560 4208 22612 4214
rect 22560 4150 22612 4156
rect 22572 3602 22600 4150
rect 22664 3777 22692 6938
rect 22848 6322 22876 8230
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22834 4992 22890 5001
rect 22834 4927 22890 4936
rect 22848 4690 22876 4927
rect 22940 4729 22968 8230
rect 22926 4720 22982 4729
rect 22836 4684 22888 4690
rect 22926 4655 22982 4664
rect 22836 4626 22888 4632
rect 22744 4616 22796 4622
rect 23032 4570 23060 8230
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23124 7954 23152 8026
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 23110 7168 23166 7177
rect 23110 7103 23166 7112
rect 23124 6866 23152 7103
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 22744 4558 22796 4564
rect 22756 4146 22784 4558
rect 22848 4542 23060 4570
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22650 3768 22706 3777
rect 22650 3703 22706 3712
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22756 2990 22784 3878
rect 22848 3777 22876 4542
rect 23124 4146 23152 5306
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22834 3768 22890 3777
rect 22834 3703 22890 3712
rect 22848 3126 22876 3703
rect 23124 3618 23152 4082
rect 23216 4010 23244 9046
rect 23400 8566 23428 11194
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23400 5710 23428 6258
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23308 4214 23336 4694
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 23296 4208 23348 4214
rect 23296 4150 23348 4156
rect 23400 4146 23428 4490
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23204 4004 23256 4010
rect 23204 3946 23256 3952
rect 23124 3602 23336 3618
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 23124 3596 23348 3602
rect 23124 3590 23296 3596
rect 22926 3224 22982 3233
rect 22926 3159 22982 3168
rect 22940 3126 22968 3159
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22744 2984 22796 2990
rect 22744 2926 22796 2932
rect 22192 2848 22244 2854
rect 21836 2746 21956 2774
rect 22006 2816 22062 2825
rect 22192 2790 22244 2796
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22006 2751 22062 2760
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 19064 2032 19116 2038
rect 19064 1974 19116 1980
rect 20442 2000 20498 2009
rect 18696 1828 18748 1834
rect 18696 1770 18748 1776
rect 17682 504 17738 513
rect 17682 439 17738 448
rect 16302 96 16358 105
rect 12256 2 12308 8
rect 13542 0 13598 56
rect 14922 0 14978 56
rect 17696 56 17724 439
rect 19076 56 19104 1974
rect 20442 1935 20498 1944
rect 20456 56 20484 1935
rect 21468 1698 21496 2246
rect 21456 1692 21508 1698
rect 21456 1634 21508 1640
rect 21836 1154 21864 2746
rect 22020 2514 22048 2751
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22204 2378 22232 2790
rect 22388 2446 22416 2790
rect 23032 2582 23060 3538
rect 23124 3058 23152 3590
rect 23296 3538 23348 3544
rect 23204 3528 23256 3534
rect 23400 3482 23428 4082
rect 23492 4010 23520 9454
rect 23584 4298 23612 10066
rect 23676 8634 23704 11194
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23952 8498 23980 11194
rect 24124 10396 24176 10402
rect 24124 10338 24176 10344
rect 24136 9994 24164 10338
rect 24124 9988 24176 9994
rect 24124 9930 24176 9936
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 24136 8974 24164 9046
rect 24124 8968 24176 8974
rect 24124 8910 24176 8916
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 23756 6724 23808 6730
rect 23756 6666 23808 6672
rect 23768 6254 23796 6666
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 23860 4826 23888 8230
rect 24136 7206 24164 8230
rect 24228 7886 24256 11194
rect 24400 10260 24452 10266
rect 24400 10202 24452 10208
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24228 7206 24256 7482
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 23584 4270 23704 4298
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23256 3476 23428 3482
rect 23204 3470 23428 3476
rect 23216 3454 23428 3470
rect 23584 3126 23612 4082
rect 23676 3942 23704 4270
rect 23860 4214 23888 4762
rect 24044 4321 24072 6598
rect 24136 6497 24164 6598
rect 24122 6488 24178 6497
rect 24122 6423 24178 6432
rect 24030 4312 24086 4321
rect 24030 4247 24086 4256
rect 23848 4208 23900 4214
rect 23754 4176 23810 4185
rect 23848 4150 23900 4156
rect 23754 4111 23756 4120
rect 23808 4111 23810 4120
rect 24124 4140 24176 4146
rect 23756 4082 23808 4088
rect 24124 4082 24176 4088
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 24136 3738 24164 4082
rect 24412 3738 24440 10202
rect 24504 7750 24532 11194
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24596 7478 24624 8570
rect 24780 8498 24808 11194
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24676 8424 24728 8430
rect 24860 8424 24912 8430
rect 24676 8366 24728 8372
rect 24780 8372 24860 8378
rect 24780 8366 24912 8372
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24492 7268 24544 7274
rect 24492 7210 24544 7216
rect 24504 7002 24532 7210
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24688 5642 24716 8366
rect 24780 8350 24900 8366
rect 24676 5636 24728 5642
rect 24676 5578 24728 5584
rect 24780 4865 24808 8350
rect 25056 7886 25084 11194
rect 25332 9874 25360 11194
rect 25608 10305 25636 11194
rect 25884 11014 25912 11194
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25594 10296 25650 10305
rect 25594 10231 25650 10240
rect 25962 10160 26018 10169
rect 25962 10095 26018 10104
rect 25976 9897 26004 10095
rect 26160 9897 26188 11194
rect 25962 9888 26018 9897
rect 25332 9846 25452 9874
rect 25226 9072 25282 9081
rect 25226 9007 25282 9016
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24964 7342 24992 7754
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 25056 7177 25084 7278
rect 25042 7168 25098 7177
rect 25042 7103 25098 7112
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24872 5817 24900 6258
rect 24858 5808 24914 5817
rect 24858 5743 24914 5752
rect 24952 5772 25004 5778
rect 25056 5760 25084 7103
rect 25004 5732 25084 5760
rect 24952 5714 25004 5720
rect 24766 4856 24822 4865
rect 24766 4791 24822 4800
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24596 3534 24624 4422
rect 25148 4078 25176 8055
rect 25240 7886 25268 9007
rect 25424 8498 25452 9846
rect 25962 9823 26018 9832
rect 26146 9888 26202 9897
rect 26146 9823 26202 9832
rect 26436 9738 26464 11194
rect 26712 11082 26740 11194
rect 27028 11194 27030 11212
rect 27250 11194 27306 11250
rect 27526 11194 27582 11250
rect 27802 11194 27858 11250
rect 28078 11194 28134 11250
rect 28354 11194 28410 11250
rect 28630 11194 28686 11250
rect 28906 11194 28962 11250
rect 29182 11194 29238 11250
rect 29458 11194 29514 11250
rect 29734 11194 29790 11250
rect 30010 11194 30066 11250
rect 30286 11194 30342 11250
rect 30562 11194 30618 11250
rect 30838 11194 30894 11250
rect 31114 11194 31170 11250
rect 31390 11194 31446 11250
rect 31666 11194 31722 11250
rect 31942 11194 31998 11250
rect 32218 11194 32274 11250
rect 32494 11194 32550 11250
rect 32770 11194 32826 11250
rect 33046 11194 33102 11250
rect 33322 11194 33378 11250
rect 33598 11194 33654 11250
rect 33874 11194 33930 11250
rect 34150 11194 34206 11250
rect 34426 11194 34482 11250
rect 34702 11194 34758 11250
rect 34978 11194 35034 11250
rect 35254 11194 35310 11250
rect 35530 11194 35586 11250
rect 35806 11194 35862 11250
rect 36082 11194 36138 11250
rect 36358 11194 36414 11250
rect 36634 11194 36690 11250
rect 36910 11194 36966 11250
rect 37186 11194 37242 11250
rect 37372 11212 37424 11218
rect 26976 11154 27028 11160
rect 27264 11150 27292 11194
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26884 10192 26936 10198
rect 26884 10134 26936 10140
rect 26436 9710 26556 9738
rect 25504 8560 25556 8566
rect 25504 8502 25556 8508
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 25240 7410 25268 7822
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25240 6798 25268 7346
rect 25332 6905 25360 7346
rect 25318 6896 25374 6905
rect 25318 6831 25374 6840
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25320 6792 25372 6798
rect 25372 6752 25452 6780
rect 25320 6734 25372 6740
rect 25228 6112 25280 6118
rect 25228 6054 25280 6060
rect 25320 6112 25372 6118
rect 25320 6054 25372 6060
rect 25240 5914 25268 6054
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25226 5808 25282 5817
rect 25226 5743 25282 5752
rect 25240 5710 25268 5743
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25136 4072 25188 4078
rect 25136 4014 25188 4020
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23020 2576 23072 2582
rect 25332 2553 25360 6054
rect 25424 2972 25452 6752
rect 25516 5098 25544 8502
rect 26528 8430 26556 9710
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25608 5302 25636 7890
rect 25700 6866 25728 8298
rect 25778 8256 25834 8265
rect 25778 8191 25834 8200
rect 25792 7546 25820 8191
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25976 7698 26004 7822
rect 25884 7670 26004 7698
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25884 7002 25912 7670
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25700 6662 25728 6802
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 26238 6488 26294 6497
rect 26238 6423 26294 6432
rect 26252 6390 26280 6423
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26344 6322 26372 7346
rect 26332 6316 26384 6322
rect 26332 6258 26384 6264
rect 25870 6216 25926 6225
rect 25870 6151 25926 6160
rect 25596 5296 25648 5302
rect 25596 5238 25648 5244
rect 25504 5092 25556 5098
rect 25504 5034 25556 5040
rect 25778 3768 25834 3777
rect 25884 3738 25912 6151
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26068 5302 26096 5646
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 26238 4720 26294 4729
rect 26238 4655 26294 4664
rect 26252 4010 26280 4655
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25778 3703 25834 3712
rect 25872 3732 25924 3738
rect 25792 3670 25820 3703
rect 25872 3674 25924 3680
rect 25780 3664 25832 3670
rect 25780 3606 25832 3612
rect 26344 3369 26372 3878
rect 26436 3534 26464 7686
rect 26516 7268 26568 7274
rect 26516 7210 26568 7216
rect 26528 6866 26556 7210
rect 26606 7168 26662 7177
rect 26606 7103 26662 7112
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26620 6746 26648 7103
rect 26896 7002 26924 10134
rect 27264 9042 27476 9058
rect 27540 9042 27568 11194
rect 27252 9036 27476 9042
rect 27304 9030 27476 9036
rect 27252 8978 27304 8984
rect 27448 8974 27476 9030
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 27816 8498 27844 11194
rect 27986 10024 28042 10033
rect 27986 9959 28042 9968
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27528 8356 27580 8362
rect 27528 8298 27580 8304
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 27540 7426 27568 8298
rect 27802 7984 27858 7993
rect 27712 7948 27764 7954
rect 27802 7919 27858 7928
rect 27712 7890 27764 7896
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27448 7410 27568 7426
rect 27436 7404 27568 7410
rect 27488 7398 27568 7404
rect 27436 7346 27488 7352
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 26528 6718 26648 6746
rect 26700 6792 26752 6798
rect 26976 6792 27028 6798
rect 26700 6734 26752 6740
rect 26896 6740 26976 6746
rect 26896 6734 27028 6740
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26330 3360 26386 3369
rect 26330 3295 26386 3304
rect 25596 2984 25648 2990
rect 25424 2944 25596 2972
rect 25596 2926 25648 2932
rect 25608 2825 25636 2926
rect 26528 2922 26556 6718
rect 26712 6662 26740 6734
rect 26896 6718 27016 6734
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26620 6458 26648 6598
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26896 5574 26924 6718
rect 27264 6712 27292 7142
rect 27436 6928 27488 6934
rect 27436 6870 27488 6876
rect 27264 6684 27384 6712
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27356 5302 27384 6684
rect 27344 5296 27396 5302
rect 27344 5238 27396 5244
rect 27448 5234 27476 6870
rect 27540 6866 27568 7398
rect 27528 6860 27580 6866
rect 27528 6802 27580 6808
rect 27540 6186 27568 6802
rect 27632 6254 27660 7686
rect 27724 7449 27752 7890
rect 27710 7440 27766 7449
rect 27816 7410 27844 7919
rect 27896 7472 27948 7478
rect 27894 7440 27896 7449
rect 27948 7440 27950 7449
rect 27710 7375 27766 7384
rect 27804 7404 27856 7410
rect 27894 7375 27950 7384
rect 27804 7346 27856 7352
rect 27816 6798 27844 7346
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 28000 6662 28028 9959
rect 28092 8498 28120 11194
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28172 8016 28224 8022
rect 28172 7958 28224 7964
rect 28184 6798 28212 7958
rect 28368 7886 28396 11194
rect 28644 8498 28672 11194
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28276 7546 28304 7822
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28356 7472 28408 7478
rect 28354 7440 28356 7449
rect 28408 7440 28410 7449
rect 28354 7375 28410 7384
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28172 6792 28224 6798
rect 28092 6752 28172 6780
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 27816 6304 27844 6598
rect 27908 6458 27936 6598
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 27896 6316 27948 6322
rect 27816 6276 27896 6304
rect 28092 6304 28120 6752
rect 28172 6734 28224 6740
rect 27948 6276 28120 6304
rect 27896 6258 27948 6264
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 28172 6248 28224 6254
rect 28172 6190 28224 6196
rect 27528 6180 27580 6186
rect 27528 6122 27580 6128
rect 28184 5846 28212 6190
rect 28172 5840 28224 5846
rect 28172 5782 28224 5788
rect 28276 5710 28304 6802
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28368 6118 28396 6734
rect 28356 6112 28408 6118
rect 28356 6054 28408 6060
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 28460 5370 28488 7686
rect 28552 7313 28580 8366
rect 28538 7304 28594 7313
rect 28538 7239 28594 7248
rect 28736 6984 28764 9998
rect 28816 9240 28868 9246
rect 28816 9182 28868 9188
rect 28828 7041 28856 9182
rect 28920 7886 28948 11194
rect 28998 9888 29054 9897
rect 28998 9823 29054 9832
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 28644 6956 28764 6984
rect 28814 7032 28870 7041
rect 28814 6967 28870 6976
rect 28644 6662 28672 6956
rect 28722 6896 28778 6905
rect 28722 6831 28778 6840
rect 28736 6662 28764 6831
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28632 6656 28684 6662
rect 28632 6598 28684 6604
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28828 6458 28856 6734
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28920 6322 28948 7278
rect 29012 6662 29040 9823
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 29104 8566 29132 9114
rect 29196 8566 29224 11194
rect 29274 10296 29330 10305
rect 29274 10231 29330 10240
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29184 8560 29236 8566
rect 29184 8502 29236 8508
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 29104 8090 29132 8230
rect 29092 8084 29144 8090
rect 29092 8026 29144 8032
rect 29000 6656 29052 6662
rect 29000 6598 29052 6604
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 28448 5364 28500 5370
rect 28448 5306 28500 5312
rect 28724 5364 28776 5370
rect 28724 5306 28776 5312
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 28080 5160 28132 5166
rect 28080 5102 28132 5108
rect 27896 5092 27948 5098
rect 27896 5034 27948 5040
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27802 4312 27858 4321
rect 27802 4247 27858 4256
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27434 3904 27490 3913
rect 27434 3839 27490 3848
rect 27448 3534 27476 3839
rect 27540 3534 27568 4014
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 27632 3058 27660 4150
rect 27816 4146 27844 4247
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 26516 2916 26568 2922
rect 26516 2858 26568 2864
rect 25594 2816 25650 2825
rect 25594 2751 25650 2760
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 23020 2518 23072 2524
rect 25318 2544 25374 2553
rect 25318 2479 25374 2488
rect 27724 2446 27752 3062
rect 27908 2990 27936 5034
rect 28092 4078 28120 5102
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 27988 4004 28040 4010
rect 27988 3946 28040 3952
rect 28000 3670 28028 3946
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 27896 2984 27948 2990
rect 27896 2926 27948 2932
rect 28184 2854 28212 5170
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28276 3670 28304 4422
rect 28356 4276 28408 4282
rect 28356 4218 28408 4224
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 28368 3194 28396 4218
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 28448 4072 28500 4078
rect 28448 4014 28500 4020
rect 28460 3913 28488 4014
rect 28644 3942 28672 4082
rect 28632 3936 28684 3942
rect 28446 3904 28502 3913
rect 28502 3862 28580 3890
rect 28632 3878 28684 3884
rect 28446 3839 28502 3848
rect 28552 3602 28580 3862
rect 28448 3596 28500 3602
rect 28448 3538 28500 3544
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 28460 3194 28488 3538
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 28448 3188 28500 3194
rect 28448 3130 28500 3136
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 22192 2372 22244 2378
rect 22192 2314 22244 2320
rect 25964 2372 26016 2378
rect 25964 2314 26016 2320
rect 24582 1864 24638 1873
rect 24582 1799 24638 1808
rect 21824 1148 21876 1154
rect 21824 1090 21876 1096
rect 23202 368 23258 377
rect 23202 303 23258 312
rect 21822 232 21878 241
rect 21822 167 21878 176
rect 21836 56 21864 167
rect 23216 56 23244 303
rect 24596 56 24624 1799
rect 25976 56 26004 2314
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 28184 1290 28212 2790
rect 28460 2446 28488 3130
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28368 2106 28396 2246
rect 28356 2100 28408 2106
rect 28356 2042 28408 2048
rect 28172 1284 28224 1290
rect 28172 1226 28224 1232
rect 27342 640 27398 649
rect 27342 575 27398 584
rect 27356 56 27384 575
rect 28736 56 28764 5306
rect 28920 5030 28948 6258
rect 29288 5778 29316 10231
rect 29368 8356 29420 8362
rect 29368 8298 29420 8304
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 29276 5024 29328 5030
rect 29276 4966 29328 4972
rect 28920 4706 28948 4966
rect 28920 4678 29132 4706
rect 29104 4622 29132 4678
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29092 4616 29144 4622
rect 29092 4558 29144 4564
rect 29012 3058 29040 4558
rect 29288 3602 29316 4966
rect 29380 4321 29408 8298
rect 29472 7886 29500 11194
rect 29644 9988 29696 9994
rect 29644 9930 29696 9936
rect 29552 9104 29604 9110
rect 29552 9046 29604 9052
rect 29460 7880 29512 7886
rect 29460 7822 29512 7828
rect 29564 4486 29592 9046
rect 29656 4758 29684 9930
rect 29748 7886 29776 11194
rect 30024 9602 30052 11194
rect 30024 9574 30144 9602
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29736 7744 29788 7750
rect 29736 7686 29788 7692
rect 29644 4752 29696 4758
rect 29644 4694 29696 4700
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 29366 4312 29422 4321
rect 29366 4247 29422 4256
rect 29748 4146 29776 7686
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29276 3596 29328 3602
rect 29276 3538 29328 3544
rect 29000 3052 29052 3058
rect 29000 2994 29052 3000
rect 29380 2922 29408 4014
rect 29472 3670 29500 4082
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29460 3664 29512 3670
rect 29460 3606 29512 3612
rect 29564 3534 29592 3878
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 29552 3528 29604 3534
rect 29552 3470 29604 3476
rect 29460 3052 29512 3058
rect 29460 2994 29512 3000
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 29368 2916 29420 2922
rect 29368 2858 29420 2864
rect 29472 1970 29500 2994
rect 29460 1964 29512 1970
rect 29460 1906 29512 1912
rect 29564 513 29592 2994
rect 29656 1766 29684 3606
rect 29748 3516 29776 4082
rect 29840 3618 29868 8910
rect 30116 7886 30144 9574
rect 30194 8528 30250 8537
rect 30300 8498 30328 11194
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30194 8463 30250 8472
rect 30288 8492 30340 8498
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30012 7744 30064 7750
rect 30012 7686 30064 7692
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 29932 3738 29960 4558
rect 30024 4554 30052 7686
rect 30104 6724 30156 6730
rect 30104 6666 30156 6672
rect 30012 4548 30064 4554
rect 30012 4490 30064 4496
rect 30012 4276 30064 4282
rect 30012 4218 30064 4224
rect 29920 3732 29972 3738
rect 29920 3674 29972 3680
rect 29840 3590 29960 3618
rect 29828 3528 29880 3534
rect 29748 3488 29828 3516
rect 29828 3470 29880 3476
rect 29932 3398 29960 3590
rect 30024 3466 30052 4218
rect 30012 3460 30064 3466
rect 30012 3402 30064 3408
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29644 1760 29696 1766
rect 29644 1702 29696 1708
rect 29550 504 29606 513
rect 29550 439 29606 448
rect 30116 56 30144 6666
rect 30208 3738 30236 8463
rect 30288 8434 30340 8440
rect 30392 7546 30420 8570
rect 30576 7886 30604 11194
rect 30852 8022 30880 11194
rect 31128 8498 31156 11194
rect 31404 8566 31432 11194
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31392 8560 31444 8566
rect 31392 8502 31444 8508
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 30932 8424 30984 8430
rect 30932 8366 30984 8372
rect 30840 8016 30892 8022
rect 30840 7958 30892 7964
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30748 7744 30800 7750
rect 30748 7686 30800 7692
rect 30380 7540 30432 7546
rect 30380 7482 30432 7488
rect 30286 7032 30342 7041
rect 30286 6967 30342 6976
rect 30300 4978 30328 6967
rect 30300 4950 30420 4978
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 30300 4214 30328 4762
rect 30288 4208 30340 4214
rect 30288 4150 30340 4156
rect 30392 4026 30420 4950
rect 30656 4480 30708 4486
rect 30656 4422 30708 4428
rect 30668 4282 30696 4422
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 30300 3998 30420 4026
rect 30300 3738 30328 3998
rect 30196 3732 30248 3738
rect 30196 3674 30248 3680
rect 30288 3732 30340 3738
rect 30288 3674 30340 3680
rect 30564 3528 30616 3534
rect 30564 3470 30616 3476
rect 30576 2922 30604 3470
rect 30760 3194 30788 7686
rect 30944 6458 30972 8366
rect 31588 7478 31616 8910
rect 31680 7886 31708 11194
rect 31956 9602 31984 11194
rect 31864 9574 31984 9602
rect 31864 7954 31892 9574
rect 32128 9308 32180 9314
rect 32128 9250 32180 9256
rect 32140 8634 32168 9250
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 32232 8378 32260 11194
rect 32508 8634 32536 11194
rect 32784 8650 32812 11194
rect 33060 8838 33088 11194
rect 33336 9602 33364 11194
rect 33336 9574 33456 9602
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 32784 8634 32904 8650
rect 32496 8628 32548 8634
rect 32784 8628 32916 8634
rect 32784 8622 32864 8628
rect 32496 8570 32548 8576
rect 32864 8570 32916 8576
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32232 8350 32352 8378
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 32324 8090 32352 8350
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31576 7472 31628 7478
rect 31576 7414 31628 7420
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 30932 6452 30984 6458
rect 30932 6394 30984 6400
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30852 3670 30880 3878
rect 30840 3664 30892 3670
rect 30840 3606 30892 3612
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30564 2916 30616 2922
rect 30564 2858 30616 2864
rect 31496 56 31524 7346
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32692 5137 32720 8434
rect 32864 8424 32916 8430
rect 32864 8366 32916 8372
rect 32772 7268 32824 7274
rect 32772 7210 32824 7216
rect 32678 5128 32734 5137
rect 32678 5063 32734 5072
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 31668 3664 31720 3670
rect 31668 3606 31720 3612
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 31588 105 31616 3470
rect 31680 2038 31708 3606
rect 32784 2938 32812 7210
rect 32876 3738 32904 8366
rect 33428 8362 33456 9574
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 33520 8634 33548 8774
rect 33612 8634 33640 11194
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33888 8566 33916 11194
rect 33876 8560 33928 8566
rect 33876 8502 33928 8508
rect 33692 8492 33744 8498
rect 33692 8434 33744 8440
rect 34060 8492 34112 8498
rect 34060 8434 34112 8440
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33704 3738 33732 8434
rect 34072 3738 34100 8434
rect 34164 8362 34192 11194
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34152 8356 34204 8362
rect 34152 8298 34204 8304
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 33692 3732 33744 3738
rect 33692 3674 33744 3680
rect 34060 3732 34112 3738
rect 34060 3674 34112 3680
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 34152 3528 34204 3534
rect 34152 3470 34204 3476
rect 32876 3058 32904 3470
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32784 2910 32904 2938
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 31668 2032 31720 2038
rect 31668 1974 31720 1980
rect 31574 96 31630 105
rect 16302 0 16358 40
rect 17682 0 17738 56
rect 19062 0 19118 56
rect 20442 0 20498 56
rect 21822 0 21878 56
rect 23202 0 23258 56
rect 24582 0 24638 56
rect 25962 0 26018 56
rect 27342 0 27398 56
rect 28722 0 28778 56
rect 30102 0 30158 56
rect 31482 0 31538 56
rect 32876 56 32904 2910
rect 33140 2848 33192 2854
rect 33140 2790 33192 2796
rect 33152 2514 33180 2790
rect 33140 2508 33192 2514
rect 33140 2450 33192 2456
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 33888 1873 33916 3470
rect 34164 2378 34192 3470
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 33874 1864 33930 1873
rect 33874 1799 33930 1808
rect 34256 56 34284 7346
rect 34348 6390 34376 9862
rect 34440 8090 34468 11194
rect 34612 11008 34664 11014
rect 34612 10950 34664 10956
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34532 7206 34560 8774
rect 34520 7200 34572 7206
rect 34520 7142 34572 7148
rect 34624 6798 34652 10950
rect 34716 8650 34744 11194
rect 34716 8634 34928 8650
rect 34716 8628 34940 8634
rect 34716 8622 34888 8628
rect 34888 8570 34940 8576
rect 34992 8514 35020 11194
rect 35268 9110 35296 11194
rect 35256 9104 35308 9110
rect 35256 9046 35308 9052
rect 34992 8486 35112 8514
rect 35084 8430 35112 8486
rect 35164 8492 35216 8498
rect 35164 8434 35216 8440
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35072 8424 35124 8430
rect 35072 8366 35124 8372
rect 34704 8288 34756 8294
rect 34704 8230 34756 8236
rect 34716 7410 34744 8230
rect 34796 7744 34848 7750
rect 34796 7686 34848 7692
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 34612 6792 34664 6798
rect 34612 6734 34664 6740
rect 34336 6384 34388 6390
rect 34336 6326 34388 6332
rect 34428 6248 34480 6254
rect 34428 6190 34480 6196
rect 34440 5681 34468 6190
rect 34426 5672 34482 5681
rect 34426 5607 34482 5616
rect 34808 5370 34836 7686
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 35176 3534 35204 8434
rect 35360 3670 35388 8434
rect 35348 3664 35400 3670
rect 35348 3606 35400 3612
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 35452 3398 35480 8434
rect 35544 8090 35572 11194
rect 35624 9852 35676 9858
rect 35624 9794 35676 9800
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35636 7206 35664 9794
rect 35820 8634 35848 11194
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 35624 5704 35676 5710
rect 35624 5646 35676 5652
rect 35532 3528 35584 3534
rect 35532 3470 35584 3476
rect 35544 3398 35572 3470
rect 35440 3392 35492 3398
rect 35440 3334 35492 3340
rect 35532 3392 35584 3398
rect 35532 3334 35584 3340
rect 35636 56 35664 5646
rect 35820 3738 35848 8434
rect 36004 6322 36032 11018
rect 36096 8090 36124 11194
rect 36268 9104 36320 9110
rect 36268 9046 36320 9052
rect 36280 8362 36308 9046
rect 36372 8362 36400 11194
rect 36544 10260 36596 10266
rect 36544 10202 36596 10208
rect 36452 9036 36504 9042
rect 36452 8978 36504 8984
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 36188 7478 36216 7822
rect 36268 7812 36320 7818
rect 36268 7754 36320 7760
rect 36176 7472 36228 7478
rect 36176 7414 36228 7420
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 35808 3732 35860 3738
rect 35808 3674 35860 3680
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 35728 2009 35756 3470
rect 36280 3194 36308 7754
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 35714 2000 35770 2009
rect 35714 1935 35770 1944
rect 36372 1329 36400 7346
rect 36464 6118 36492 8978
rect 36556 6458 36584 10202
rect 36648 8090 36676 11194
rect 36924 8634 36952 11194
rect 37096 9716 37148 9722
rect 37096 9658 37148 9664
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 37004 8492 37056 8498
rect 37004 8434 37056 8440
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36820 8016 36872 8022
rect 36820 7958 36872 7964
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36740 7546 36768 7822
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 36636 7404 36688 7410
rect 36636 7346 36688 7352
rect 36648 7002 36676 7346
rect 36636 6996 36688 7002
rect 36636 6938 36688 6944
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 36452 6112 36504 6118
rect 36452 6054 36504 6060
rect 36832 3466 36860 7958
rect 36912 7744 36964 7750
rect 36912 7686 36964 7692
rect 36544 3460 36596 3466
rect 36544 3402 36596 3408
rect 36820 3460 36872 3466
rect 36820 3402 36872 3408
rect 36556 2446 36584 3402
rect 36924 2774 36952 7686
rect 37016 6934 37044 8434
rect 37004 6928 37056 6934
rect 37004 6870 37056 6876
rect 37108 6866 37136 9658
rect 37200 8362 37228 11194
rect 37462 11194 37518 11250
rect 37738 11194 37794 11250
rect 37372 11154 37424 11160
rect 37280 8832 37332 8838
rect 37280 8774 37332 8780
rect 37292 8498 37320 8774
rect 37384 8650 37412 11154
rect 37476 9654 37504 11194
rect 37556 11144 37608 11150
rect 37556 11086 37608 11092
rect 37464 9648 37516 9654
rect 37464 9590 37516 9596
rect 37384 8622 37504 8650
rect 37280 8492 37332 8498
rect 37280 8434 37332 8440
rect 37188 8356 37240 8362
rect 37188 8298 37240 8304
rect 37280 7812 37332 7818
rect 37280 7754 37332 7760
rect 37292 7546 37320 7754
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 37476 6866 37504 8622
rect 37096 6860 37148 6866
rect 37096 6802 37148 6808
rect 37464 6860 37516 6866
rect 37464 6802 37516 6808
rect 37568 6730 37596 11086
rect 37648 8424 37700 8430
rect 37648 8366 37700 8372
rect 37556 6724 37608 6730
rect 37556 6666 37608 6672
rect 37280 5160 37332 5166
rect 37280 5102 37332 5108
rect 37292 4185 37320 5102
rect 37464 4616 37516 4622
rect 37464 4558 37516 4564
rect 37278 4176 37334 4185
rect 37278 4111 37334 4120
rect 37004 3664 37056 3670
rect 37004 3606 37056 3612
rect 37016 2938 37044 3606
rect 37096 3392 37148 3398
rect 37096 3334 37148 3340
rect 37108 3074 37136 3334
rect 37476 3126 37504 4558
rect 37660 3738 37688 8366
rect 37752 8090 37780 11194
rect 38658 9888 38714 9897
rect 38658 9823 38714 9832
rect 38384 9648 38436 9654
rect 38384 9590 38436 9596
rect 38396 8634 38424 9590
rect 38474 9344 38530 9353
rect 38474 9279 38530 9288
rect 38384 8628 38436 8634
rect 38384 8570 38436 8576
rect 37832 8492 37884 8498
rect 37832 8434 37884 8440
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38384 8492 38436 8498
rect 38384 8434 38436 8440
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37740 7404 37792 7410
rect 37740 7346 37792 7352
rect 37752 4049 37780 7346
rect 37844 5914 37872 8434
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38304 8090 38332 8434
rect 38292 8084 38344 8090
rect 38292 8026 38344 8032
rect 38292 7948 38344 7954
rect 38292 7890 38344 7896
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38120 7313 38148 7346
rect 38106 7304 38162 7313
rect 38106 7239 38162 7248
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38014 6896 38070 6905
rect 37924 6860 37976 6866
rect 38014 6831 38016 6840
rect 37924 6802 37976 6808
rect 38068 6831 38070 6840
rect 38016 6802 38068 6808
rect 37936 6390 37964 6802
rect 37924 6384 37976 6390
rect 37924 6326 37976 6332
rect 38304 6186 38332 7890
rect 38396 7342 38424 8434
rect 38488 7546 38516 9279
rect 38568 8900 38620 8906
rect 38568 8842 38620 8848
rect 38476 7540 38528 7546
rect 38476 7482 38528 7488
rect 38580 7410 38608 8842
rect 38672 8090 38700 9823
rect 39578 9616 39634 9625
rect 39578 9551 39634 9560
rect 38844 8968 38896 8974
rect 38844 8910 38896 8916
rect 38856 8498 38884 8910
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39592 8634 39620 9551
rect 39670 9072 39726 9081
rect 39670 9007 39726 9016
rect 39580 8628 39632 8634
rect 39580 8570 39632 8576
rect 38844 8492 38896 8498
rect 38844 8434 38896 8440
rect 39212 8492 39264 8498
rect 39212 8434 39264 8440
rect 39224 8401 39252 8434
rect 39210 8392 39266 8401
rect 39210 8327 39266 8336
rect 39396 8356 39448 8362
rect 39396 8298 39448 8304
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 39408 7993 39436 8298
rect 39486 8256 39542 8265
rect 39486 8191 39542 8200
rect 39394 7984 39450 7993
rect 39394 7919 39450 7928
rect 38844 7880 38896 7886
rect 38842 7848 38844 7857
rect 38896 7848 38898 7857
rect 38660 7812 38712 7818
rect 38842 7783 38898 7792
rect 38660 7754 38712 7760
rect 38568 7404 38620 7410
rect 38568 7346 38620 7352
rect 38384 7336 38436 7342
rect 38384 7278 38436 7284
rect 38382 6896 38438 6905
rect 38382 6831 38384 6840
rect 38436 6831 38438 6840
rect 38384 6802 38436 6808
rect 38672 6769 38700 7754
rect 38936 7744 38988 7750
rect 38842 7712 38898 7721
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38842 7647 38898 7656
rect 38856 7410 38884 7647
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 39500 7546 39528 8191
rect 39488 7540 39540 7546
rect 39488 7482 39540 7488
rect 38934 7440 38990 7449
rect 38844 7404 38896 7410
rect 38934 7375 38990 7384
rect 39580 7404 39632 7410
rect 38844 7346 38896 7352
rect 39580 7346 39632 7352
rect 39488 7268 39540 7274
rect 39488 7210 39540 7216
rect 39396 7200 39448 7206
rect 39394 7168 39396 7177
rect 39448 7168 39450 7177
rect 39394 7103 39450 7112
rect 39500 6905 39528 7210
rect 39486 6896 39542 6905
rect 39486 6831 39542 6840
rect 38752 6792 38804 6798
rect 38658 6760 38714 6769
rect 39592 6746 39620 7346
rect 38752 6734 38804 6740
rect 38658 6695 38714 6704
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 38292 6180 38344 6186
rect 38292 6122 38344 6128
rect 38488 6118 38516 6598
rect 38568 6248 38620 6254
rect 38568 6190 38620 6196
rect 38476 6112 38528 6118
rect 38476 6054 38528 6060
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37832 5908 37884 5914
rect 37832 5850 37884 5856
rect 38200 5908 38252 5914
rect 38200 5850 38252 5856
rect 38212 5817 38240 5850
rect 38198 5808 38254 5817
rect 38198 5743 38254 5752
rect 38580 5273 38608 6190
rect 38660 6112 38712 6118
rect 38660 6054 38712 6060
rect 38672 5817 38700 6054
rect 38658 5808 38714 5817
rect 38658 5743 38714 5752
rect 38660 5636 38712 5642
rect 38660 5578 38712 5584
rect 38566 5264 38622 5273
rect 38566 5199 38622 5208
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 37738 4040 37794 4049
rect 37738 3975 37794 3984
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 37648 3732 37700 3738
rect 37648 3674 37700 3680
rect 38672 3641 38700 5578
rect 38764 4729 38792 6734
rect 39500 6718 39620 6746
rect 39010 6556 39318 6565
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39028 6452 39080 6458
rect 39028 6394 39080 6400
rect 39040 6361 39068 6394
rect 39026 6352 39082 6361
rect 39026 6287 39082 6296
rect 39394 6080 39450 6089
rect 39394 6015 39450 6024
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39408 5370 39436 6015
rect 39396 5364 39448 5370
rect 39396 5306 39448 5312
rect 38936 5296 38988 5302
rect 38936 5238 38988 5244
rect 39394 5264 39450 5273
rect 38844 5228 38896 5234
rect 38844 5170 38896 5176
rect 38750 4720 38806 4729
rect 38750 4655 38806 4664
rect 38658 3632 38714 3641
rect 38856 3618 38884 5170
rect 38948 4622 38976 5238
rect 39394 5199 39450 5208
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39408 4826 39436 5199
rect 39500 4842 39528 6718
rect 39684 6662 39712 9007
rect 40038 8936 40094 8945
rect 40038 8871 40094 8880
rect 39854 8800 39910 8809
rect 39854 8735 39910 8744
rect 39762 8528 39818 8537
rect 39762 8463 39818 8472
rect 39672 6656 39724 6662
rect 39578 6624 39634 6633
rect 39672 6598 39724 6604
rect 39578 6559 39634 6568
rect 39592 5914 39620 6559
rect 39776 6458 39804 8463
rect 39868 7478 39896 8735
rect 39856 7472 39908 7478
rect 39856 7414 39908 7420
rect 39856 6996 39908 7002
rect 39856 6938 39908 6944
rect 39764 6452 39816 6458
rect 39764 6394 39816 6400
rect 39672 6384 39724 6390
rect 39672 6326 39724 6332
rect 39580 5908 39632 5914
rect 39580 5850 39632 5856
rect 39396 4820 39448 4826
rect 39500 4814 39620 4842
rect 39396 4762 39448 4768
rect 39486 4720 39542 4729
rect 39486 4655 39542 4664
rect 38936 4616 38988 4622
rect 38936 4558 38988 4564
rect 39010 4380 39318 4389
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 39394 4176 39450 4185
rect 39212 4140 39264 4146
rect 39394 4111 39450 4120
rect 39212 4082 39264 4088
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 39026 3839 39082 3848
rect 38658 3567 38714 3576
rect 38764 3590 38884 3618
rect 37648 3392 37700 3398
rect 37648 3334 37700 3340
rect 37464 3120 37516 3126
rect 37108 3046 37228 3074
rect 37464 3062 37516 3068
rect 37016 2910 37136 2938
rect 36924 2746 37044 2774
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36358 1320 36414 1329
rect 36358 1255 36414 1264
rect 37016 56 37044 2746
rect 37108 377 37136 2910
rect 37094 368 37150 377
rect 37094 303 37150 312
rect 37200 241 37228 3046
rect 37660 649 37688 3334
rect 38764 3210 38792 3590
rect 38844 3528 38896 3534
rect 39224 3505 39252 4082
rect 39408 3738 39436 4111
rect 39500 4010 39528 4655
rect 39592 4593 39620 4814
rect 39578 4584 39634 4593
rect 39578 4519 39634 4528
rect 39488 4004 39540 4010
rect 39488 3946 39540 3952
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39394 3632 39450 3641
rect 39394 3567 39450 3576
rect 38844 3470 38896 3476
rect 39210 3496 39266 3505
rect 38672 3182 38792 3210
rect 38672 3097 38700 3182
rect 38658 3088 38714 3097
rect 37740 3052 37792 3058
rect 37740 2994 37792 3000
rect 37832 3052 37884 3058
rect 38658 3023 38714 3032
rect 38752 3052 38804 3058
rect 37832 2994 37884 3000
rect 38752 2994 38804 3000
rect 37646 640 37702 649
rect 37646 575 37702 584
rect 37186 232 37242 241
rect 37186 167 37242 176
rect 37752 66 37780 2994
rect 37844 1737 37872 2994
rect 38476 2848 38528 2854
rect 38476 2790 38528 2796
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38488 2553 38516 2790
rect 38474 2544 38530 2553
rect 38474 2479 38530 2488
rect 38108 2440 38160 2446
rect 38108 2382 38160 2388
rect 38476 2440 38528 2446
rect 38476 2382 38528 2388
rect 37924 2304 37976 2310
rect 37924 2246 37976 2252
rect 37936 2009 37964 2246
rect 37922 2000 37978 2009
rect 37922 1935 37978 1944
rect 38120 1834 38148 2382
rect 38292 2304 38344 2310
rect 38292 2246 38344 2252
rect 38108 1828 38160 1834
rect 38108 1770 38160 1776
rect 38304 1737 38332 2246
rect 38488 1970 38516 2382
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38476 1964 38528 1970
rect 38476 1906 38528 1912
rect 37830 1728 37886 1737
rect 37830 1663 37886 1672
rect 38290 1728 38346 1737
rect 38290 1663 38346 1672
rect 38672 1465 38700 2246
rect 38658 1456 38714 1465
rect 38658 1391 38714 1400
rect 38764 1358 38792 2994
rect 38752 1352 38804 1358
rect 38382 1320 38438 1329
rect 38752 1294 38804 1300
rect 38382 1255 38438 1264
rect 37740 60 37792 66
rect 31574 31 31630 40
rect 32862 0 32918 56
rect 34242 0 34298 56
rect 35622 0 35678 56
rect 37002 0 37058 56
rect 38396 56 38424 1255
rect 38856 1222 38884 3470
rect 39210 3431 39266 3440
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39408 3194 39436 3567
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39394 3088 39450 3097
rect 38936 3052 38988 3058
rect 39394 3023 39450 3032
rect 38936 2994 38988 3000
rect 38948 1601 38976 2994
rect 39028 2848 39080 2854
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 39026 2751 39082 2760
rect 39408 2650 39436 3023
rect 39684 2961 39712 6326
rect 39670 2952 39726 2961
rect 39670 2887 39726 2896
rect 39868 2774 39896 6938
rect 39948 5840 40000 5846
rect 39948 5782 40000 5788
rect 39960 5545 39988 5782
rect 39946 5536 40002 5545
rect 39946 5471 40002 5480
rect 39948 4752 40000 4758
rect 39948 4694 40000 4700
rect 39960 4457 39988 4694
rect 39946 4448 40002 4457
rect 39946 4383 40002 4392
rect 40052 4078 40080 8871
rect 40040 4072 40092 4078
rect 40040 4014 40092 4020
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 39960 3369 39988 3606
rect 39946 3360 40002 3369
rect 39946 3295 40002 3304
rect 39776 2746 39896 2774
rect 39396 2644 39448 2650
rect 39396 2586 39448 2592
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 38934 1592 38990 1601
rect 38934 1527 38990 1536
rect 38844 1216 38896 1222
rect 38844 1158 38896 1164
rect 39776 56 39804 2746
rect 39948 2304 40000 2310
rect 39946 2272 39948 2281
rect 40000 2272 40002 2281
rect 39946 2207 40002 2216
rect 37740 2 37792 8
rect 38382 0 38438 56
rect 39762 0 39818 56
<< via2 >>
rect 1398 9832 1454 9888
rect 754 9560 810 9616
rect 938 9288 994 9344
rect 570 8200 626 8256
rect 1122 8472 1178 8528
rect 754 7384 810 7440
rect 1214 7928 1270 7984
rect 2778 9016 2834 9072
rect 2594 8336 2650 8392
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1674 7928 1730 7984
rect 2870 8744 2926 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1306 7656 1362 7712
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 294 6840 350 6896
rect 846 7112 902 7168
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1030 6568 1086 6624
rect 2318 6840 2374 6896
rect 1214 6296 1270 6352
rect 570 6024 626 6080
rect 202 5752 258 5808
rect 662 5480 718 5536
rect 1674 6316 1730 6352
rect 1674 6296 1676 6316
rect 1676 6296 1728 6316
rect 1728 6296 1730 6316
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1858 5752 1914 5808
rect 5630 8880 5686 8936
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 846 5208 902 5264
rect 386 4936 442 4992
rect 2778 5072 2834 5128
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 846 4664 902 4720
rect 754 4392 810 4448
rect 846 4120 902 4176
rect 386 3848 442 3904
rect 846 3576 902 3632
rect 202 3304 258 3360
rect 846 3032 902 3088
rect 202 2216 258 2272
rect 1214 2760 1270 2816
rect 1030 2488 1086 2544
rect 754 1944 810 2000
rect 386 1672 442 1728
rect 1214 1400 1270 1456
rect 2410 3848 2466 3904
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 5814 9424 5870 9480
rect 3238 2488 3294 2544
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 4066 1672 4122 1728
rect 5538 3440 5594 3496
rect 5630 2896 5686 2952
rect 6918 7828 6920 7848
rect 6920 7828 6972 7848
rect 6972 7828 6974 7848
rect 6918 7792 6974 7828
rect 6366 4528 6422 4584
rect 6182 3984 6238 4040
rect 6366 3168 6422 3224
rect 6182 3032 6238 3088
rect 7102 6432 7158 6488
rect 6826 5616 6882 5672
rect 6642 4684 6698 4720
rect 6642 4664 6644 4684
rect 6644 4664 6696 4684
rect 6696 4664 6698 4684
rect 8666 9696 8722 9752
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7930 7404 7986 7440
rect 7930 7384 7932 7404
rect 7932 7384 7984 7404
rect 7984 7384 7986 7404
rect 8206 7248 8262 7304
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 8022 6740 8024 6760
rect 8024 6740 8076 6760
rect 8076 6740 8078 6760
rect 8022 6704 8078 6740
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 7562 5228 7618 5264
rect 7562 5208 7564 5228
rect 7564 5208 7616 5228
rect 7616 5208 7618 5228
rect 7378 4120 7434 4176
rect 7286 3884 7288 3904
rect 7288 3884 7340 3904
rect 7340 3884 7342 3904
rect 7286 3848 7342 3884
rect 7654 3576 7710 3632
rect 6918 3304 6974 3360
rect 7562 3168 7618 3224
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 8206 3032 8262 3088
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 8666 7384 8722 7440
rect 8758 6432 8814 6488
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 9770 9052 9772 9072
rect 9772 9052 9824 9072
rect 9824 9052 9826 9072
rect 9770 9016 9826 9052
rect 9218 7404 9274 7440
rect 9218 7384 9220 7404
rect 9220 7384 9272 7404
rect 9272 7384 9274 7404
rect 9402 6704 9458 6760
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 8390 4800 8446 4856
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 8850 3340 8852 3360
rect 8852 3340 8904 3360
rect 8904 3340 8906 3360
rect 8850 3304 8906 3340
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 8482 3068 8484 3088
rect 8484 3068 8536 3088
rect 8536 3068 8538 3088
rect 8482 3032 8538 3068
rect 9586 4004 9642 4040
rect 9586 3984 9588 4004
rect 9588 3984 9640 4004
rect 9640 3984 9642 4004
rect 9494 3168 9550 3224
rect 10230 9832 10286 9888
rect 10506 9288 10562 9344
rect 6458 1536 6514 1592
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 11426 9152 11482 9208
rect 11426 8336 11482 8392
rect 10966 7656 11022 7712
rect 11886 7384 11942 7440
rect 11702 6704 11758 6760
rect 10782 6024 10838 6080
rect 12806 6160 12862 6216
rect 12438 6024 12494 6080
rect 10782 5344 10838 5400
rect 12438 5480 12494 5536
rect 12162 4684 12218 4720
rect 12162 4664 12164 4684
rect 12164 4664 12216 4684
rect 12216 4664 12218 4684
rect 12162 4120 12218 4176
rect 12162 3068 12164 3088
rect 12164 3068 12216 3088
rect 12216 3068 12218 3088
rect 12162 3032 12218 3068
rect 12346 3848 12402 3904
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 14738 9968 14794 10024
rect 12346 3032 12402 3088
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 14370 6976 14426 7032
rect 14462 6568 14518 6624
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14738 7656 14794 7712
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 14830 6568 14886 6624
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 13726 4800 13782 4856
rect 13726 2932 13728 2952
rect 13728 2932 13780 2952
rect 13780 2932 13782 2952
rect 13726 2896 13782 2932
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 15198 6196 15200 6216
rect 15200 6196 15252 6216
rect 15252 6196 15254 6216
rect 15198 6160 15254 6196
rect 16026 7112 16082 7168
rect 15658 6160 15714 6216
rect 14738 5516 14740 5536
rect 14740 5516 14792 5536
rect 14792 5516 14794 5536
rect 14738 5480 14794 5516
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 14830 5344 14886 5400
rect 15566 5344 15622 5400
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 14830 4120 14886 4176
rect 15290 3576 15346 3632
rect 15474 4004 15530 4040
rect 15474 3984 15476 4004
rect 15476 3984 15528 4004
rect 15528 3984 15530 4004
rect 15658 4256 15714 4312
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15658 3032 15714 3088
rect 15842 3032 15898 3088
rect 15842 2932 15844 2952
rect 15844 2932 15896 2952
rect 15896 2932 15898 2952
rect 15842 2896 15898 2932
rect 16854 4548 16910 4584
rect 16854 4528 16856 4548
rect 16856 4528 16908 4548
rect 16908 4528 16910 4548
rect 18602 9152 18658 9208
rect 18786 8236 18788 8256
rect 18788 8236 18840 8256
rect 18840 8236 18842 8256
rect 18786 8200 18842 8236
rect 17222 7656 17278 7712
rect 17222 7248 17278 7304
rect 18326 7284 18328 7304
rect 18328 7284 18380 7304
rect 18380 7284 18382 7304
rect 18326 7248 18382 7284
rect 18326 6976 18382 7032
rect 18694 6568 18750 6624
rect 17774 5072 17830 5128
rect 17130 3848 17186 3904
rect 16946 3304 17002 3360
rect 17958 3984 18014 4040
rect 17866 3304 17922 3360
rect 17406 2760 17462 2816
rect 18970 6452 19026 6488
rect 18970 6432 18972 6452
rect 18972 6432 19024 6452
rect 19024 6432 19026 6452
rect 19338 10104 19394 10160
rect 19246 8200 19302 8256
rect 19890 10104 19946 10160
rect 20258 8628 20314 8664
rect 20258 8608 20260 8628
rect 20260 8608 20312 8628
rect 20312 8608 20314 8628
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 19430 6976 19486 7032
rect 19614 6976 19670 7032
rect 20350 8200 20406 8256
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 20810 8064 20866 8120
rect 19798 7520 19854 7576
rect 20718 7792 20774 7848
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 20810 7248 20866 7304
rect 20718 6976 20774 7032
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21086 7284 21088 7304
rect 21088 7284 21140 7304
rect 21140 7284 21142 7304
rect 21086 7248 21142 7284
rect 21270 6976 21326 7032
rect 18418 4256 18474 4312
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19338 5888 19394 5944
rect 20810 6568 20866 6624
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 20810 6452 20866 6488
rect 20810 6432 20812 6452
rect 20812 6432 20864 6452
rect 20864 6432 20866 6452
rect 19154 5480 19210 5536
rect 19522 5652 19524 5672
rect 19524 5652 19576 5672
rect 19576 5652 19578 5672
rect 19522 5616 19578 5652
rect 20534 5616 20590 5672
rect 20810 5480 20866 5536
rect 20350 5208 20406 5264
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 18786 5072 18842 5128
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 20902 4936 20958 4992
rect 20350 4800 20406 4856
rect 19798 3848 19854 3904
rect 20350 3848 20406 3904
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 21638 5888 21694 5944
rect 21822 6024 21878 6080
rect 22098 6296 22154 6352
rect 22558 7248 22614 7304
rect 21546 3304 21602 3360
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 21730 3168 21786 3224
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 19522 2624 19578 2680
rect 22190 3884 22192 3904
rect 22192 3884 22244 3904
rect 22244 3884 22246 3904
rect 22190 3848 22246 3884
rect 22374 3712 22430 3768
rect 22834 4936 22890 4992
rect 22926 4664 22982 4720
rect 23110 7112 23166 7168
rect 22650 3712 22706 3768
rect 22834 3712 22890 3768
rect 22926 3168 22982 3224
rect 22006 2760 22062 2816
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 17682 448 17738 504
rect 16302 40 16358 96
rect 20442 1944 20498 2000
rect 24122 6432 24178 6488
rect 24030 4256 24086 4312
rect 23754 4140 23810 4176
rect 23754 4120 23756 4140
rect 23756 4120 23808 4140
rect 23808 4120 23810 4140
rect 25594 10240 25650 10296
rect 25962 10104 26018 10160
rect 25226 9016 25282 9072
rect 25134 8064 25190 8120
rect 25042 7112 25098 7168
rect 24858 5752 24914 5808
rect 24766 4800 24822 4856
rect 25962 9832 26018 9888
rect 26146 9832 26202 9888
rect 25318 6840 25374 6896
rect 25226 5752 25282 5808
rect 25778 8200 25834 8256
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 26238 6432 26294 6488
rect 25870 6160 25926 6216
rect 25778 3712 25834 3768
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 26238 4664 26294 4720
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 26606 7112 26662 7168
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 27986 9968 28042 10024
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27802 7928 27858 7984
rect 26330 3304 26386 3360
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27710 7384 27766 7440
rect 27894 7420 27896 7440
rect 27896 7420 27948 7440
rect 27948 7420 27950 7440
rect 27894 7384 27950 7420
rect 28354 7420 28356 7440
rect 28356 7420 28408 7440
rect 28408 7420 28410 7440
rect 28354 7384 28410 7420
rect 28538 7248 28594 7304
rect 28998 9832 29054 9888
rect 28814 6976 28870 7032
rect 28722 6840 28778 6896
rect 29274 10240 29330 10296
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27802 4256 27858 4312
rect 27434 3848 27490 3904
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 25594 2760 25650 2816
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 25318 2488 25374 2544
rect 28446 3848 28502 3904
rect 24582 1808 24638 1864
rect 23202 312 23258 368
rect 21822 176 21878 232
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 27342 584 27398 640
rect 29366 4256 29422 4312
rect 30194 8472 30250 8528
rect 29550 448 29606 504
rect 30286 6976 30342 7032
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 32678 5072 32734 5128
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 31574 40 31630 96
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 33874 1808 33930 1864
rect 34426 5616 34482 5672
rect 35714 1944 35770 2000
rect 37278 4120 37334 4176
rect 38658 9832 38714 9888
rect 38474 9288 38530 9344
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 38106 7248 38162 7304
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 38014 6860 38070 6896
rect 38014 6840 38016 6860
rect 38016 6840 38068 6860
rect 38068 6840 38070 6860
rect 39578 9560 39634 9616
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 39670 9016 39726 9072
rect 39210 8336 39266 8392
rect 39486 8200 39542 8256
rect 39394 7928 39450 7984
rect 38842 7828 38844 7848
rect 38844 7828 38896 7848
rect 38896 7828 38898 7848
rect 38842 7792 38898 7828
rect 38382 6860 38438 6896
rect 38382 6840 38384 6860
rect 38384 6840 38436 6860
rect 38436 6840 38438 6860
rect 38842 7656 38898 7712
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 39394 7148 39396 7168
rect 39396 7148 39448 7168
rect 39448 7148 39450 7168
rect 39394 7112 39450 7148
rect 39486 6840 39542 6896
rect 38658 6704 38714 6760
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 38198 5752 38254 5808
rect 38658 5752 38714 5808
rect 38566 5208 38622 5264
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 37738 3984 37794 4040
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39026 6296 39082 6352
rect 39394 6024 39450 6080
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 38750 4664 38806 4720
rect 38658 3576 38714 3632
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 40038 8880 40094 8936
rect 39854 8744 39910 8800
rect 39762 8472 39818 8528
rect 39578 6568 39634 6624
rect 39486 4664 39542 4720
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 36358 1264 36414 1320
rect 37094 312 37150 368
rect 39578 4528 39634 4584
rect 39394 3576 39450 3632
rect 38658 3032 38714 3088
rect 37646 584 37702 640
rect 37186 176 37242 232
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38474 2488 38530 2544
rect 37922 1944 37978 2000
rect 37830 1672 37886 1728
rect 38290 1672 38346 1728
rect 38658 1400 38714 1456
rect 38382 1264 38438 1320
rect 39210 3440 39266 3496
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39394 3032 39450 3088
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 39670 2896 39726 2952
rect 39946 5480 40002 5536
rect 39946 4392 40002 4448
rect 39946 3304 40002 3360
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 38934 1536 38990 1592
rect 39946 2252 39948 2272
rect 39948 2252 40000 2272
rect 40000 2252 40002 2272
rect 39946 2216 40002 2252
<< metal3 >>
rect 25589 10298 25655 10301
rect 29269 10298 29335 10301
rect 25589 10296 29335 10298
rect 25589 10240 25594 10296
rect 25650 10240 29274 10296
rect 29330 10240 29335 10296
rect 25589 10238 29335 10240
rect 25589 10235 25655 10238
rect 29269 10235 29335 10238
rect 19333 10162 19399 10165
rect 19885 10162 19951 10165
rect 19333 10160 19951 10162
rect 19333 10104 19338 10160
rect 19394 10104 19890 10160
rect 19946 10104 19951 10160
rect 19333 10102 19951 10104
rect 19333 10099 19399 10102
rect 19885 10099 19951 10102
rect 25957 10162 26023 10165
rect 28942 10162 28948 10164
rect 25957 10160 28948 10162
rect 25957 10104 25962 10160
rect 26018 10104 28948 10160
rect 25957 10102 28948 10104
rect 25957 10099 26023 10102
rect 28942 10100 28948 10102
rect 29012 10100 29018 10164
rect 14733 10026 14799 10029
rect 27981 10026 28047 10029
rect 14733 10024 28047 10026
rect 14733 9968 14738 10024
rect 14794 9968 27986 10024
rect 28042 9968 28047 10024
rect 14733 9966 28047 9968
rect 14733 9963 14799 9966
rect 27981 9963 28047 9966
rect 0 9890 120 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 120 9830
rect 1393 9827 1459 9830
rect 10225 9890 10291 9893
rect 25957 9890 26023 9893
rect 10225 9888 26023 9890
rect 10225 9832 10230 9888
rect 10286 9832 25962 9888
rect 26018 9832 26023 9888
rect 10225 9830 26023 9832
rect 10225 9827 10291 9830
rect 25957 9827 26023 9830
rect 26141 9890 26207 9893
rect 28993 9890 29059 9893
rect 26141 9888 29059 9890
rect 26141 9832 26146 9888
rect 26202 9832 28998 9888
rect 29054 9832 29059 9888
rect 26141 9830 29059 9832
rect 26141 9827 26207 9830
rect 28993 9827 29059 9830
rect 38653 9890 38719 9893
rect 40880 9890 41000 9920
rect 38653 9888 41000 9890
rect 38653 9832 38658 9888
rect 38714 9832 41000 9888
rect 38653 9830 41000 9832
rect 38653 9827 38719 9830
rect 40880 9800 41000 9830
rect 8661 9754 8727 9757
rect 38326 9754 38332 9756
rect 8661 9752 38332 9754
rect 8661 9696 8666 9752
rect 8722 9696 38332 9752
rect 8661 9694 38332 9696
rect 8661 9691 8727 9694
rect 38326 9692 38332 9694
rect 38396 9692 38402 9756
rect 0 9618 120 9648
rect 749 9618 815 9621
rect 0 9616 815 9618
rect 0 9560 754 9616
rect 810 9560 815 9616
rect 0 9558 815 9560
rect 0 9528 120 9558
rect 749 9555 815 9558
rect 39573 9618 39639 9621
rect 40880 9618 41000 9648
rect 39573 9616 41000 9618
rect 39573 9560 39578 9616
rect 39634 9560 41000 9616
rect 39573 9558 41000 9560
rect 39573 9555 39639 9558
rect 40880 9528 41000 9558
rect 5809 9482 5875 9485
rect 28574 9482 28580 9484
rect 5809 9480 28580 9482
rect 5809 9424 5814 9480
rect 5870 9424 28580 9480
rect 5809 9422 28580 9424
rect 5809 9419 5875 9422
rect 28574 9420 28580 9422
rect 28644 9420 28650 9484
rect 0 9346 120 9376
rect 933 9346 999 9349
rect 0 9344 999 9346
rect 0 9288 938 9344
rect 994 9288 999 9344
rect 0 9286 999 9288
rect 0 9256 120 9286
rect 933 9283 999 9286
rect 10501 9346 10567 9349
rect 37222 9346 37228 9348
rect 10501 9344 37228 9346
rect 10501 9288 10506 9344
rect 10562 9288 37228 9344
rect 10501 9286 37228 9288
rect 10501 9283 10567 9286
rect 37222 9284 37228 9286
rect 37292 9284 37298 9348
rect 38469 9346 38535 9349
rect 40880 9346 41000 9376
rect 38469 9344 41000 9346
rect 38469 9288 38474 9344
rect 38530 9288 41000 9344
rect 38469 9286 41000 9288
rect 38469 9283 38535 9286
rect 40880 9256 41000 9286
rect 11421 9210 11487 9213
rect 18597 9210 18663 9213
rect 11421 9208 18663 9210
rect 11421 9152 11426 9208
rect 11482 9152 18602 9208
rect 18658 9152 18663 9208
rect 11421 9150 18663 9152
rect 11421 9147 11487 9150
rect 18597 9147 18663 9150
rect 0 9074 120 9104
rect 2773 9074 2839 9077
rect 0 9072 2839 9074
rect 0 9016 2778 9072
rect 2834 9016 2839 9072
rect 0 9014 2839 9016
rect 0 8984 120 9014
rect 2773 9011 2839 9014
rect 9765 9074 9831 9077
rect 25221 9074 25287 9077
rect 9765 9072 25287 9074
rect 9765 9016 9770 9072
rect 9826 9016 25226 9072
rect 25282 9016 25287 9072
rect 9765 9014 25287 9016
rect 9765 9011 9831 9014
rect 25221 9011 25287 9014
rect 39665 9074 39731 9077
rect 40880 9074 41000 9104
rect 39665 9072 41000 9074
rect 39665 9016 39670 9072
rect 39726 9016 41000 9072
rect 39665 9014 41000 9016
rect 39665 9011 39731 9014
rect 40880 8984 41000 9014
rect 5625 8938 5691 8941
rect 40033 8938 40099 8941
rect 5625 8936 40099 8938
rect 5625 8880 5630 8936
rect 5686 8880 40038 8936
rect 40094 8880 40099 8936
rect 5625 8878 40099 8880
rect 5625 8875 5691 8878
rect 40033 8875 40099 8878
rect 0 8802 120 8832
rect 2865 8802 2931 8805
rect 0 8800 2931 8802
rect 0 8744 2870 8800
rect 2926 8744 2931 8800
rect 0 8742 2931 8744
rect 0 8712 120 8742
rect 2865 8739 2931 8742
rect 39849 8802 39915 8805
rect 40880 8802 41000 8832
rect 39849 8800 41000 8802
rect 39849 8744 39854 8800
rect 39910 8744 41000 8800
rect 39849 8742 41000 8744
rect 39849 8739 39915 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 19742 8604 19748 8668
rect 19812 8666 19818 8668
rect 20253 8666 20319 8669
rect 19812 8664 20319 8666
rect 19812 8608 20258 8664
rect 20314 8608 20319 8664
rect 19812 8606 20319 8608
rect 19812 8604 19818 8606
rect 20253 8603 20319 8606
rect 0 8530 120 8560
rect 1117 8530 1183 8533
rect 30189 8530 30255 8533
rect 0 8528 1183 8530
rect 0 8472 1122 8528
rect 1178 8472 1183 8528
rect 0 8470 1183 8472
rect 0 8440 120 8470
rect 1117 8467 1183 8470
rect 2730 8528 30255 8530
rect 2730 8472 30194 8528
rect 30250 8472 30255 8528
rect 2730 8470 30255 8472
rect 2589 8394 2655 8397
rect 2730 8394 2790 8470
rect 30189 8467 30255 8470
rect 39757 8530 39823 8533
rect 40880 8530 41000 8560
rect 39757 8528 41000 8530
rect 39757 8472 39762 8528
rect 39818 8472 41000 8528
rect 39757 8470 41000 8472
rect 39757 8467 39823 8470
rect 40880 8440 41000 8470
rect 2589 8392 2790 8394
rect 2589 8336 2594 8392
rect 2650 8336 2790 8392
rect 2589 8334 2790 8336
rect 11421 8394 11487 8397
rect 39205 8394 39271 8397
rect 11421 8392 39271 8394
rect 11421 8336 11426 8392
rect 11482 8336 39210 8392
rect 39266 8336 39271 8392
rect 11421 8334 39271 8336
rect 2589 8331 2655 8334
rect 11421 8331 11487 8334
rect 39205 8331 39271 8334
rect 0 8258 120 8288
rect 565 8258 631 8261
rect 0 8256 631 8258
rect 0 8200 570 8256
rect 626 8200 631 8256
rect 0 8198 631 8200
rect 0 8168 120 8198
rect 565 8195 631 8198
rect 18781 8258 18847 8261
rect 19241 8258 19307 8261
rect 18781 8256 19307 8258
rect 18781 8200 18786 8256
rect 18842 8200 19246 8256
rect 19302 8200 19307 8256
rect 18781 8198 19307 8200
rect 18781 8195 18847 8198
rect 19241 8195 19307 8198
rect 20345 8258 20411 8261
rect 25773 8258 25839 8261
rect 20345 8256 25839 8258
rect 20345 8200 20350 8256
rect 20406 8200 25778 8256
rect 25834 8200 25839 8256
rect 20345 8198 25839 8200
rect 20345 8195 20411 8198
rect 25773 8195 25839 8198
rect 39481 8258 39547 8261
rect 40880 8258 41000 8288
rect 39481 8256 41000 8258
rect 39481 8200 39486 8256
rect 39542 8200 41000 8256
rect 39481 8198 41000 8200
rect 39481 8195 39547 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 20805 8122 20871 8125
rect 25129 8122 25195 8125
rect 20805 8120 25195 8122
rect 20805 8064 20810 8120
rect 20866 8064 25134 8120
rect 25190 8064 25195 8120
rect 20805 8062 25195 8064
rect 20805 8059 20871 8062
rect 25129 8059 25195 8062
rect 0 7986 120 8016
rect 1209 7986 1275 7989
rect 0 7984 1275 7986
rect 0 7928 1214 7984
rect 1270 7928 1275 7984
rect 0 7926 1275 7928
rect 0 7896 120 7926
rect 1209 7923 1275 7926
rect 1669 7986 1735 7989
rect 27797 7986 27863 7989
rect 1669 7984 27863 7986
rect 1669 7928 1674 7984
rect 1730 7928 27802 7984
rect 27858 7928 27863 7984
rect 1669 7926 27863 7928
rect 1669 7923 1735 7926
rect 27797 7923 27863 7926
rect 39389 7986 39455 7989
rect 40880 7986 41000 8016
rect 39389 7984 41000 7986
rect 39389 7928 39394 7984
rect 39450 7928 41000 7984
rect 39389 7926 41000 7928
rect 39389 7923 39455 7926
rect 40880 7896 41000 7926
rect 6913 7850 6979 7853
rect 20713 7850 20779 7853
rect 38837 7850 38903 7853
rect 6913 7848 20779 7850
rect 6913 7792 6918 7848
rect 6974 7792 20718 7848
rect 20774 7792 20779 7848
rect 6913 7790 20779 7792
rect 6913 7787 6979 7790
rect 20713 7787 20779 7790
rect 20854 7848 38903 7850
rect 20854 7792 38842 7848
rect 38898 7792 38903 7848
rect 20854 7790 38903 7792
rect 0 7714 120 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 120 7654
rect 1301 7651 1367 7654
rect 10961 7714 11027 7717
rect 14733 7714 14799 7717
rect 10961 7712 14799 7714
rect 10961 7656 10966 7712
rect 11022 7656 14738 7712
rect 14794 7656 14799 7712
rect 10961 7654 14799 7656
rect 10961 7651 11027 7654
rect 14733 7651 14799 7654
rect 17217 7714 17283 7717
rect 20854 7714 20914 7790
rect 38837 7787 38903 7790
rect 17217 7712 20914 7714
rect 17217 7656 17222 7712
rect 17278 7656 20914 7712
rect 17217 7654 20914 7656
rect 17217 7651 17283 7654
rect 37222 7652 37228 7716
rect 37292 7714 37298 7716
rect 38837 7714 38903 7717
rect 37292 7712 38903 7714
rect 37292 7656 38842 7712
rect 38898 7656 38903 7712
rect 37292 7654 38903 7656
rect 37292 7652 37298 7654
rect 38837 7651 38903 7654
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 19793 7578 19859 7581
rect 20846 7578 20852 7580
rect 9446 7518 14842 7578
rect 0 7442 120 7472
rect 749 7442 815 7445
rect 0 7440 815 7442
rect 0 7384 754 7440
rect 810 7384 815 7440
rect 0 7382 815 7384
rect 0 7352 120 7382
rect 749 7379 815 7382
rect 7925 7442 7991 7445
rect 8661 7442 8727 7445
rect 9213 7442 9279 7445
rect 9446 7442 9506 7518
rect 7925 7440 9506 7442
rect 7925 7384 7930 7440
rect 7986 7384 8666 7440
rect 8722 7384 9218 7440
rect 9274 7384 9506 7440
rect 7925 7382 9506 7384
rect 11881 7442 11947 7445
rect 14782 7442 14842 7518
rect 19793 7576 20852 7578
rect 19793 7520 19798 7576
rect 19854 7520 20852 7576
rect 19793 7518 20852 7520
rect 19793 7515 19859 7518
rect 20846 7516 20852 7518
rect 20916 7516 20922 7580
rect 27705 7442 27771 7445
rect 11881 7440 14658 7442
rect 11881 7384 11886 7440
rect 11942 7384 14658 7440
rect 11881 7382 14658 7384
rect 14782 7440 27771 7442
rect 14782 7384 27710 7440
rect 27766 7384 27771 7440
rect 14782 7382 27771 7384
rect 7925 7379 7991 7382
rect 8661 7379 8727 7382
rect 9213 7379 9279 7382
rect 11881 7379 11947 7382
rect 8201 7306 8267 7309
rect 14598 7306 14658 7382
rect 27705 7379 27771 7382
rect 27889 7442 27955 7445
rect 28349 7442 28415 7445
rect 27889 7440 28415 7442
rect 27889 7384 27894 7440
rect 27950 7384 28354 7440
rect 28410 7384 28415 7440
rect 27889 7382 28415 7384
rect 27889 7379 27955 7382
rect 28349 7379 28415 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 17217 7306 17283 7309
rect 8201 7304 14474 7306
rect 8201 7248 8206 7304
rect 8262 7248 14474 7304
rect 8201 7246 14474 7248
rect 14598 7304 17283 7306
rect 14598 7248 17222 7304
rect 17278 7248 17283 7304
rect 14598 7246 17283 7248
rect 8201 7243 8267 7246
rect 0 7170 120 7200
rect 841 7170 907 7173
rect 0 7168 907 7170
rect 0 7112 846 7168
rect 902 7112 907 7168
rect 0 7110 907 7112
rect 14414 7170 14474 7246
rect 17217 7243 17283 7246
rect 18321 7306 18387 7309
rect 20805 7306 20871 7309
rect 21081 7306 21147 7309
rect 18321 7304 20362 7306
rect 18321 7248 18326 7304
rect 18382 7272 20362 7304
rect 20805 7304 21147 7306
rect 18382 7248 20408 7272
rect 18321 7246 20408 7248
rect 18321 7243 18387 7246
rect 20302 7212 20408 7246
rect 20805 7248 20810 7304
rect 20866 7248 21086 7304
rect 21142 7248 21147 7304
rect 20805 7246 21147 7248
rect 20805 7243 20871 7246
rect 21081 7243 21147 7246
rect 22553 7306 22619 7309
rect 28533 7306 28599 7309
rect 38101 7306 38167 7309
rect 22553 7304 28599 7306
rect 22553 7248 22558 7304
rect 22614 7248 28538 7304
rect 28594 7248 28599 7304
rect 22553 7246 28599 7248
rect 22553 7243 22619 7246
rect 28533 7243 28599 7246
rect 31710 7304 38167 7306
rect 31710 7248 38106 7304
rect 38162 7248 38167 7304
rect 31710 7246 38167 7248
rect 16021 7170 16087 7173
rect 14414 7168 16087 7170
rect 14414 7112 16026 7168
rect 16082 7112 16087 7168
rect 14414 7110 16087 7112
rect 20348 7170 20408 7212
rect 23105 7170 23171 7173
rect 25037 7170 25103 7173
rect 20348 7168 25103 7170
rect 20348 7112 23110 7168
rect 23166 7112 25042 7168
rect 25098 7112 25103 7168
rect 20348 7110 25103 7112
rect 0 7080 120 7110
rect 841 7107 907 7110
rect 16021 7107 16087 7110
rect 23105 7107 23171 7110
rect 25037 7107 25103 7110
rect 26601 7170 26667 7173
rect 31710 7170 31770 7246
rect 38101 7243 38167 7246
rect 26601 7168 31770 7170
rect 26601 7112 26606 7168
rect 26662 7112 31770 7168
rect 26601 7110 31770 7112
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 26601 7107 26667 7110
rect 39389 7107 39455 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 14365 7034 14431 7037
rect 18321 7034 18387 7037
rect 19425 7036 19491 7037
rect 19609 7036 19675 7037
rect 19374 7034 19380 7036
rect 14365 7032 18387 7034
rect 14365 6976 14370 7032
rect 14426 6976 18326 7032
rect 18382 6976 18387 7032
rect 14365 6974 18387 6976
rect 19334 6974 19380 7034
rect 19444 7032 19491 7036
rect 19486 6976 19491 7032
rect 14365 6971 14431 6974
rect 18321 6971 18387 6974
rect 19374 6972 19380 6974
rect 19444 6972 19491 6976
rect 19558 6972 19564 7036
rect 19628 7034 19675 7036
rect 20713 7034 20779 7037
rect 21265 7034 21331 7037
rect 19628 7032 19720 7034
rect 19670 6976 19720 7032
rect 19628 6974 19720 6976
rect 20713 7032 21331 7034
rect 20713 6976 20718 7032
rect 20774 6976 21270 7032
rect 21326 6976 21331 7032
rect 20713 6974 21331 6976
rect 19628 6972 19675 6974
rect 19425 6971 19491 6972
rect 19609 6971 19675 6972
rect 20713 6971 20779 6974
rect 21265 6971 21331 6974
rect 28809 7034 28875 7037
rect 30281 7034 30347 7037
rect 28809 7032 30347 7034
rect 28809 6976 28814 7032
rect 28870 6976 30286 7032
rect 30342 6976 30347 7032
rect 28809 6974 30347 6976
rect 28809 6971 28875 6974
rect 30281 6971 30347 6974
rect 0 6898 120 6928
rect 289 6898 355 6901
rect 0 6896 355 6898
rect 0 6840 294 6896
rect 350 6840 355 6896
rect 0 6838 355 6840
rect 0 6808 120 6838
rect 289 6835 355 6838
rect 2313 6898 2379 6901
rect 25313 6898 25379 6901
rect 2313 6896 25379 6898
rect 2313 6840 2318 6896
rect 2374 6840 25318 6896
rect 25374 6840 25379 6896
rect 2313 6838 25379 6840
rect 2313 6835 2379 6838
rect 25313 6835 25379 6838
rect 28574 6836 28580 6900
rect 28644 6898 28650 6900
rect 28717 6898 28783 6901
rect 28644 6896 28783 6898
rect 28644 6840 28722 6896
rect 28778 6840 28783 6896
rect 28644 6838 28783 6840
rect 28644 6836 28650 6838
rect 28717 6835 28783 6838
rect 28942 6836 28948 6900
rect 29012 6898 29018 6900
rect 38009 6898 38075 6901
rect 38377 6900 38443 6901
rect 29012 6896 38075 6898
rect 29012 6840 38014 6896
rect 38070 6840 38075 6896
rect 29012 6838 38075 6840
rect 29012 6836 29018 6838
rect 38009 6835 38075 6838
rect 38326 6836 38332 6900
rect 38396 6898 38443 6900
rect 39481 6898 39547 6901
rect 40880 6898 41000 6928
rect 38396 6896 38488 6898
rect 38438 6840 38488 6896
rect 38396 6838 38488 6840
rect 39481 6896 41000 6898
rect 39481 6840 39486 6896
rect 39542 6840 41000 6896
rect 39481 6838 41000 6840
rect 38396 6836 38443 6838
rect 38377 6835 38443 6836
rect 39481 6835 39547 6838
rect 40880 6808 41000 6838
rect 8017 6762 8083 6765
rect 9397 6762 9463 6765
rect 8017 6760 9463 6762
rect 8017 6704 8022 6760
rect 8078 6704 9402 6760
rect 9458 6704 9463 6760
rect 8017 6702 9463 6704
rect 8017 6699 8083 6702
rect 9397 6699 9463 6702
rect 11697 6762 11763 6765
rect 38653 6762 38719 6765
rect 11697 6760 38719 6762
rect 11697 6704 11702 6760
rect 11758 6704 38658 6760
rect 38714 6704 38719 6760
rect 11697 6702 38719 6704
rect 11697 6699 11763 6702
rect 38653 6699 38719 6702
rect 0 6626 120 6656
rect 1025 6626 1091 6629
rect 0 6624 1091 6626
rect 0 6568 1030 6624
rect 1086 6568 1091 6624
rect 0 6566 1091 6568
rect 0 6536 120 6566
rect 1025 6563 1091 6566
rect 14457 6626 14523 6629
rect 14825 6626 14891 6629
rect 14457 6624 14891 6626
rect 14457 6568 14462 6624
rect 14518 6568 14830 6624
rect 14886 6568 14891 6624
rect 14457 6566 14891 6568
rect 14457 6563 14523 6566
rect 14825 6563 14891 6566
rect 18689 6626 18755 6629
rect 20805 6626 20871 6629
rect 18689 6624 20871 6626
rect 18689 6568 18694 6624
rect 18750 6568 20810 6624
rect 20866 6568 20871 6624
rect 18689 6566 20871 6568
rect 18689 6563 18755 6566
rect 20805 6563 20871 6566
rect 39573 6626 39639 6629
rect 40880 6626 41000 6656
rect 39573 6624 41000 6626
rect 39573 6568 39578 6624
rect 39634 6568 41000 6624
rect 39573 6566 41000 6568
rect 39573 6563 39639 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 7097 6490 7163 6493
rect 8753 6490 8819 6493
rect 7097 6488 8819 6490
rect 7097 6432 7102 6488
rect 7158 6432 8758 6488
rect 8814 6432 8819 6488
rect 7097 6430 8819 6432
rect 7097 6427 7163 6430
rect 8753 6427 8819 6430
rect 18965 6490 19031 6493
rect 20805 6490 20871 6493
rect 18965 6488 20871 6490
rect 18965 6432 18970 6488
rect 19026 6432 20810 6488
rect 20866 6432 20871 6488
rect 18965 6430 20871 6432
rect 18965 6427 19031 6430
rect 20805 6427 20871 6430
rect 24117 6490 24183 6493
rect 26233 6490 26299 6493
rect 24117 6488 26299 6490
rect 24117 6432 24122 6488
rect 24178 6432 26238 6488
rect 26294 6432 26299 6488
rect 24117 6430 26299 6432
rect 24117 6427 24183 6430
rect 26233 6427 26299 6430
rect 0 6354 120 6384
rect 1209 6354 1275 6357
rect 0 6352 1275 6354
rect 0 6296 1214 6352
rect 1270 6296 1275 6352
rect 0 6294 1275 6296
rect 0 6264 120 6294
rect 1209 6291 1275 6294
rect 1669 6354 1735 6357
rect 22093 6354 22159 6357
rect 1669 6352 22159 6354
rect 1669 6296 1674 6352
rect 1730 6296 22098 6352
rect 22154 6296 22159 6352
rect 1669 6294 22159 6296
rect 1669 6291 1735 6294
rect 22093 6291 22159 6294
rect 39021 6354 39087 6357
rect 40880 6354 41000 6384
rect 39021 6352 41000 6354
rect 39021 6296 39026 6352
rect 39082 6296 41000 6352
rect 39021 6294 41000 6296
rect 39021 6291 39087 6294
rect 40880 6264 41000 6294
rect 12801 6218 12867 6221
rect 15193 6218 15259 6221
rect 12801 6216 15259 6218
rect 12801 6160 12806 6216
rect 12862 6160 15198 6216
rect 15254 6160 15259 6216
rect 12801 6158 15259 6160
rect 12801 6155 12867 6158
rect 15193 6155 15259 6158
rect 15653 6218 15719 6221
rect 25865 6218 25931 6221
rect 15653 6216 25931 6218
rect 15653 6160 15658 6216
rect 15714 6160 25870 6216
rect 25926 6160 25931 6216
rect 15653 6158 25931 6160
rect 15653 6155 15719 6158
rect 25865 6155 25931 6158
rect 0 6082 120 6112
rect 565 6082 631 6085
rect 0 6080 631 6082
rect 0 6024 570 6080
rect 626 6024 631 6080
rect 0 6022 631 6024
rect 0 5992 120 6022
rect 565 6019 631 6022
rect 10777 6082 10843 6085
rect 12433 6082 12499 6085
rect 10777 6080 12499 6082
rect 10777 6024 10782 6080
rect 10838 6024 12438 6080
rect 12494 6024 12499 6080
rect 10777 6022 12499 6024
rect 10777 6019 10843 6022
rect 12433 6019 12499 6022
rect 20846 6020 20852 6084
rect 20916 6082 20922 6084
rect 21817 6082 21883 6085
rect 20916 6080 21883 6082
rect 20916 6024 21822 6080
rect 21878 6024 21883 6080
rect 20916 6022 21883 6024
rect 20916 6020 20922 6022
rect 21817 6019 21883 6022
rect 39389 6082 39455 6085
rect 40880 6082 41000 6112
rect 39389 6080 41000 6082
rect 39389 6024 39394 6080
rect 39450 6024 41000 6080
rect 39389 6022 41000 6024
rect 39389 6019 39455 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 19333 5948 19399 5949
rect 19333 5944 19380 5948
rect 19444 5946 19450 5948
rect 21633 5946 21699 5949
rect 19333 5888 19338 5944
rect 19333 5884 19380 5888
rect 19444 5886 19490 5946
rect 21633 5944 25882 5946
rect 21633 5888 21638 5944
rect 21694 5888 25882 5944
rect 21633 5886 25882 5888
rect 19444 5884 19450 5886
rect 19333 5883 19399 5884
rect 21633 5883 21699 5886
rect 0 5810 120 5840
rect 197 5810 263 5813
rect 0 5808 263 5810
rect 0 5752 202 5808
rect 258 5752 263 5808
rect 0 5750 263 5752
rect 0 5720 120 5750
rect 197 5747 263 5750
rect 1853 5810 1919 5813
rect 24853 5810 24919 5813
rect 25221 5810 25287 5813
rect 1853 5808 25287 5810
rect 1853 5752 1858 5808
rect 1914 5752 24858 5808
rect 24914 5752 25226 5808
rect 25282 5752 25287 5808
rect 1853 5750 25287 5752
rect 25822 5810 25882 5886
rect 38193 5810 38259 5813
rect 25822 5808 38259 5810
rect 25822 5752 38198 5808
rect 38254 5752 38259 5808
rect 25822 5750 38259 5752
rect 1853 5747 1919 5750
rect 24853 5747 24919 5750
rect 25221 5747 25287 5750
rect 38193 5747 38259 5750
rect 38653 5810 38719 5813
rect 40880 5810 41000 5840
rect 38653 5808 41000 5810
rect 38653 5752 38658 5808
rect 38714 5752 41000 5808
rect 38653 5750 41000 5752
rect 38653 5747 38719 5750
rect 40880 5720 41000 5750
rect 6821 5674 6887 5677
rect 19517 5674 19583 5677
rect 6821 5672 19583 5674
rect 6821 5616 6826 5672
rect 6882 5616 19522 5672
rect 19578 5616 19583 5672
rect 6821 5614 19583 5616
rect 6821 5611 6887 5614
rect 19517 5611 19583 5614
rect 20529 5674 20595 5677
rect 34421 5674 34487 5677
rect 20529 5672 34487 5674
rect 20529 5616 20534 5672
rect 20590 5616 34426 5672
rect 34482 5616 34487 5672
rect 20529 5614 34487 5616
rect 20529 5611 20595 5614
rect 34421 5611 34487 5614
rect 0 5538 120 5568
rect 657 5538 723 5541
rect 0 5536 723 5538
rect 0 5480 662 5536
rect 718 5480 723 5536
rect 0 5478 723 5480
rect 0 5448 120 5478
rect 657 5475 723 5478
rect 12433 5538 12499 5541
rect 14733 5538 14799 5541
rect 12433 5536 14799 5538
rect 12433 5480 12438 5536
rect 12494 5480 14738 5536
rect 14794 5480 14799 5536
rect 12433 5478 14799 5480
rect 12433 5475 12499 5478
rect 14733 5475 14799 5478
rect 19149 5538 19215 5541
rect 20805 5538 20871 5541
rect 19149 5536 20871 5538
rect 19149 5480 19154 5536
rect 19210 5480 20810 5536
rect 20866 5480 20871 5536
rect 19149 5478 20871 5480
rect 19149 5475 19215 5478
rect 20805 5475 20871 5478
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 39941 5475 40007 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 10777 5402 10843 5405
rect 14825 5402 14891 5405
rect 10777 5400 14891 5402
rect 10777 5344 10782 5400
rect 10838 5344 14830 5400
rect 14886 5344 14891 5400
rect 10777 5342 14891 5344
rect 10777 5339 10843 5342
rect 14825 5339 14891 5342
rect 15561 5402 15627 5405
rect 15561 5400 20546 5402
rect 15561 5344 15566 5400
rect 15622 5344 20546 5400
rect 15561 5342 20546 5344
rect 15561 5339 15627 5342
rect 0 5266 120 5296
rect 841 5266 907 5269
rect 0 5264 907 5266
rect 0 5208 846 5264
rect 902 5208 907 5264
rect 0 5206 907 5208
rect 0 5176 120 5206
rect 841 5203 907 5206
rect 7557 5266 7623 5269
rect 20345 5266 20411 5269
rect 7557 5264 20411 5266
rect 7557 5208 7562 5264
rect 7618 5208 20350 5264
rect 20406 5208 20411 5264
rect 7557 5206 20411 5208
rect 20486 5266 20546 5342
rect 38561 5266 38627 5269
rect 20486 5264 38627 5266
rect 20486 5208 38566 5264
rect 38622 5208 38627 5264
rect 20486 5206 38627 5208
rect 7557 5203 7623 5206
rect 20345 5203 20411 5206
rect 38561 5203 38627 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 2773 5130 2839 5133
rect 17769 5130 17835 5133
rect 2773 5128 17835 5130
rect 2773 5072 2778 5128
rect 2834 5072 17774 5128
rect 17830 5072 17835 5128
rect 2773 5070 17835 5072
rect 2773 5067 2839 5070
rect 17769 5067 17835 5070
rect 18781 5130 18847 5133
rect 32673 5130 32739 5133
rect 18781 5128 32739 5130
rect 18781 5072 18786 5128
rect 18842 5072 32678 5128
rect 32734 5072 32739 5128
rect 18781 5070 32739 5072
rect 18781 5067 18847 5070
rect 32673 5067 32739 5070
rect 0 4994 120 5024
rect 381 4994 447 4997
rect 0 4992 447 4994
rect 0 4936 386 4992
rect 442 4936 447 4992
rect 0 4934 447 4936
rect 0 4904 120 4934
rect 381 4931 447 4934
rect 20897 4994 20963 4997
rect 22829 4994 22895 4997
rect 20897 4992 22895 4994
rect 20897 4936 20902 4992
rect 20958 4936 22834 4992
rect 22890 4936 22895 4992
rect 20897 4934 22895 4936
rect 20897 4931 20963 4934
rect 22829 4931 22895 4934
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 8385 4858 8451 4861
rect 13721 4858 13787 4861
rect 8385 4856 13787 4858
rect 8385 4800 8390 4856
rect 8446 4800 13726 4856
rect 13782 4800 13787 4856
rect 8385 4798 13787 4800
rect 8385 4795 8451 4798
rect 13721 4795 13787 4798
rect 20345 4858 20411 4861
rect 24761 4858 24827 4861
rect 20345 4856 24827 4858
rect 20345 4800 20350 4856
rect 20406 4800 24766 4856
rect 24822 4800 24827 4856
rect 20345 4798 24827 4800
rect 20345 4795 20411 4798
rect 24761 4795 24827 4798
rect 0 4722 120 4752
rect 841 4722 907 4725
rect 0 4720 907 4722
rect 0 4664 846 4720
rect 902 4664 907 4720
rect 0 4662 907 4664
rect 0 4632 120 4662
rect 841 4659 907 4662
rect 6637 4722 6703 4725
rect 12157 4722 12223 4725
rect 22921 4722 22987 4725
rect 6637 4720 22987 4722
rect 6637 4664 6642 4720
rect 6698 4664 12162 4720
rect 12218 4664 22926 4720
rect 22982 4664 22987 4720
rect 6637 4662 22987 4664
rect 6637 4659 6703 4662
rect 12157 4659 12223 4662
rect 22921 4659 22987 4662
rect 26233 4722 26299 4725
rect 38745 4722 38811 4725
rect 26233 4720 38811 4722
rect 26233 4664 26238 4720
rect 26294 4664 38750 4720
rect 38806 4664 38811 4720
rect 26233 4662 38811 4664
rect 26233 4659 26299 4662
rect 38745 4659 38811 4662
rect 39481 4722 39547 4725
rect 40880 4722 41000 4752
rect 39481 4720 41000 4722
rect 39481 4664 39486 4720
rect 39542 4664 41000 4720
rect 39481 4662 41000 4664
rect 39481 4659 39547 4662
rect 40880 4632 41000 4662
rect 6361 4586 6427 4589
rect 16849 4586 16915 4589
rect 39573 4586 39639 4589
rect 6361 4584 12450 4586
rect 6361 4528 6366 4584
rect 6422 4528 12450 4584
rect 6361 4526 12450 4528
rect 6361 4523 6427 4526
rect 0 4450 120 4480
rect 749 4450 815 4453
rect 0 4448 815 4450
rect 0 4392 754 4448
rect 810 4392 815 4448
rect 0 4390 815 4392
rect 0 4360 120 4390
rect 749 4387 815 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 0 4178 120 4208
rect 841 4178 907 4181
rect 0 4176 907 4178
rect 0 4120 846 4176
rect 902 4120 907 4176
rect 0 4118 907 4120
rect 0 4088 120 4118
rect 841 4115 907 4118
rect 7373 4178 7439 4181
rect 12157 4178 12223 4181
rect 7373 4176 12223 4178
rect 7373 4120 7378 4176
rect 7434 4120 12162 4176
rect 12218 4120 12223 4176
rect 7373 4118 12223 4120
rect 12390 4178 12450 4526
rect 16849 4584 39639 4586
rect 16849 4528 16854 4584
rect 16910 4528 39578 4584
rect 39634 4528 39639 4584
rect 16849 4526 39639 4528
rect 16849 4523 16915 4526
rect 39573 4523 39639 4526
rect 39941 4450 40007 4453
rect 40880 4450 41000 4480
rect 39941 4448 41000 4450
rect 39941 4392 39946 4448
rect 40002 4392 41000 4448
rect 39941 4390 41000 4392
rect 39941 4387 40007 4390
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 15653 4314 15719 4317
rect 18413 4314 18479 4317
rect 15653 4312 18479 4314
rect 15653 4256 15658 4312
rect 15714 4256 18418 4312
rect 18474 4256 18479 4312
rect 15653 4254 18479 4256
rect 15653 4251 15719 4254
rect 18413 4251 18479 4254
rect 24025 4314 24091 4317
rect 27797 4314 27863 4317
rect 29361 4314 29427 4317
rect 24025 4312 26802 4314
rect 24025 4256 24030 4312
rect 24086 4256 26802 4312
rect 24025 4254 26802 4256
rect 24025 4251 24091 4254
rect 14825 4178 14891 4181
rect 23749 4178 23815 4181
rect 12390 4176 23815 4178
rect 12390 4120 14830 4176
rect 14886 4120 23754 4176
rect 23810 4120 23815 4176
rect 12390 4118 23815 4120
rect 26742 4178 26802 4254
rect 27797 4312 29427 4314
rect 27797 4256 27802 4312
rect 27858 4256 29366 4312
rect 29422 4256 29427 4312
rect 27797 4254 29427 4256
rect 27797 4251 27863 4254
rect 29361 4251 29427 4254
rect 37273 4178 37339 4181
rect 26742 4176 37339 4178
rect 26742 4120 37278 4176
rect 37334 4120 37339 4176
rect 26742 4118 37339 4120
rect 7373 4115 7439 4118
rect 12157 4115 12223 4118
rect 14825 4115 14891 4118
rect 23749 4115 23815 4118
rect 37273 4115 37339 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 6177 4042 6243 4045
rect 9581 4042 9647 4045
rect 15469 4042 15535 4045
rect 6177 4040 8402 4042
rect 6177 3984 6182 4040
rect 6238 3984 8402 4040
rect 6177 3982 8402 3984
rect 6177 3979 6243 3982
rect 0 3906 120 3936
rect 381 3906 447 3909
rect 0 3904 447 3906
rect 0 3848 386 3904
rect 442 3848 447 3904
rect 0 3846 447 3848
rect 0 3816 120 3846
rect 381 3843 447 3846
rect 2405 3906 2471 3909
rect 7281 3906 7347 3909
rect 2405 3904 7347 3906
rect 2405 3848 2410 3904
rect 2466 3848 7286 3904
rect 7342 3848 7347 3904
rect 2405 3846 7347 3848
rect 8342 3906 8402 3982
rect 9581 4040 15535 4042
rect 9581 3984 9586 4040
rect 9642 3984 15474 4040
rect 15530 3984 15535 4040
rect 9581 3982 15535 3984
rect 9581 3979 9647 3982
rect 15469 3979 15535 3982
rect 17953 4042 18019 4045
rect 37733 4042 37799 4045
rect 17953 4040 37799 4042
rect 17953 3984 17958 4040
rect 18014 3984 37738 4040
rect 37794 3984 37799 4040
rect 17953 3982 37799 3984
rect 17953 3979 18019 3982
rect 37733 3979 37799 3982
rect 12341 3906 12407 3909
rect 8342 3904 12407 3906
rect 8342 3848 12346 3904
rect 12402 3848 12407 3904
rect 8342 3846 12407 3848
rect 2405 3843 2471 3846
rect 7281 3843 7347 3846
rect 12341 3843 12407 3846
rect 17125 3906 17191 3909
rect 19793 3906 19859 3909
rect 17125 3904 19859 3906
rect 17125 3848 17130 3904
rect 17186 3848 19798 3904
rect 19854 3848 19859 3904
rect 17125 3846 19859 3848
rect 17125 3843 17191 3846
rect 19793 3843 19859 3846
rect 20345 3906 20411 3909
rect 22185 3906 22251 3909
rect 20345 3904 22251 3906
rect 20345 3848 20350 3904
rect 20406 3848 22190 3904
rect 22246 3848 22251 3904
rect 20345 3846 22251 3848
rect 20345 3843 20411 3846
rect 22185 3843 22251 3846
rect 27429 3906 27495 3909
rect 28441 3906 28507 3909
rect 27429 3904 28507 3906
rect 27429 3848 27434 3904
rect 27490 3848 28446 3904
rect 28502 3848 28507 3904
rect 27429 3846 28507 3848
rect 27429 3843 27495 3846
rect 28441 3843 28507 3846
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 39021 3843 39087 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 19742 3770 19748 3772
rect 15150 3710 19748 3770
rect 0 3634 120 3664
rect 841 3634 907 3637
rect 0 3632 907 3634
rect 0 3576 846 3632
rect 902 3576 907 3632
rect 0 3574 907 3576
rect 0 3544 120 3574
rect 841 3571 907 3574
rect 7649 3634 7715 3637
rect 15150 3634 15210 3710
rect 19742 3708 19748 3710
rect 19812 3708 19818 3772
rect 22369 3770 22435 3773
rect 22645 3770 22711 3773
rect 22369 3768 22711 3770
rect 22369 3712 22374 3768
rect 22430 3712 22650 3768
rect 22706 3712 22711 3768
rect 22369 3710 22711 3712
rect 22369 3707 22435 3710
rect 22645 3707 22711 3710
rect 22829 3770 22895 3773
rect 25773 3770 25839 3773
rect 22829 3768 25839 3770
rect 22829 3712 22834 3768
rect 22890 3712 25778 3768
rect 25834 3712 25839 3768
rect 22829 3710 25839 3712
rect 22829 3707 22895 3710
rect 25773 3707 25839 3710
rect 7649 3632 15210 3634
rect 7649 3576 7654 3632
rect 7710 3576 15210 3632
rect 7649 3574 15210 3576
rect 15285 3634 15351 3637
rect 38653 3634 38719 3637
rect 15285 3632 38719 3634
rect 15285 3576 15290 3632
rect 15346 3576 38658 3632
rect 38714 3576 38719 3632
rect 15285 3574 38719 3576
rect 7649 3571 7715 3574
rect 15285 3571 15351 3574
rect 38653 3571 38719 3574
rect 39389 3634 39455 3637
rect 40880 3634 41000 3664
rect 39389 3632 41000 3634
rect 39389 3576 39394 3632
rect 39450 3576 41000 3632
rect 39389 3574 41000 3576
rect 39389 3571 39455 3574
rect 40880 3544 41000 3574
rect 5533 3498 5599 3501
rect 39205 3498 39271 3501
rect 5533 3496 39271 3498
rect 5533 3440 5538 3496
rect 5594 3440 39210 3496
rect 39266 3440 39271 3496
rect 5533 3438 39271 3440
rect 5533 3435 5599 3438
rect 39205 3435 39271 3438
rect 0 3362 120 3392
rect 197 3362 263 3365
rect 0 3360 263 3362
rect 0 3304 202 3360
rect 258 3304 263 3360
rect 0 3302 263 3304
rect 0 3272 120 3302
rect 197 3299 263 3302
rect 6913 3362 6979 3365
rect 8845 3362 8911 3365
rect 6913 3360 8911 3362
rect 6913 3304 6918 3360
rect 6974 3304 8850 3360
rect 8906 3304 8911 3360
rect 6913 3302 8911 3304
rect 6913 3299 6979 3302
rect 8845 3299 8911 3302
rect 16941 3362 17007 3365
rect 17861 3362 17927 3365
rect 16941 3360 17927 3362
rect 16941 3304 16946 3360
rect 17002 3304 17866 3360
rect 17922 3304 17927 3360
rect 16941 3302 17927 3304
rect 16941 3299 17007 3302
rect 17861 3299 17927 3302
rect 21541 3362 21607 3365
rect 26325 3362 26391 3365
rect 21541 3360 26391 3362
rect 21541 3304 21546 3360
rect 21602 3304 26330 3360
rect 26386 3304 26391 3360
rect 21541 3302 26391 3304
rect 21541 3299 21607 3302
rect 26325 3299 26391 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 6361 3226 6427 3229
rect 7557 3226 7623 3229
rect 6361 3224 7623 3226
rect 6361 3168 6366 3224
rect 6422 3168 7562 3224
rect 7618 3168 7623 3224
rect 6361 3166 7623 3168
rect 6361 3163 6427 3166
rect 7557 3163 7623 3166
rect 9489 3226 9555 3229
rect 21725 3226 21791 3229
rect 22921 3226 22987 3229
rect 9489 3224 14106 3226
rect 9489 3168 9494 3224
rect 9550 3168 14106 3224
rect 9489 3166 14106 3168
rect 9489 3163 9555 3166
rect 0 3090 120 3120
rect 841 3090 907 3093
rect 0 3088 907 3090
rect 0 3032 846 3088
rect 902 3032 907 3088
rect 0 3030 907 3032
rect 0 3000 120 3030
rect 841 3027 907 3030
rect 6177 3090 6243 3093
rect 8201 3090 8267 3093
rect 6177 3088 8267 3090
rect 6177 3032 6182 3088
rect 6238 3032 8206 3088
rect 8262 3032 8267 3088
rect 6177 3030 8267 3032
rect 6177 3027 6243 3030
rect 8201 3027 8267 3030
rect 8477 3090 8543 3093
rect 12157 3090 12223 3093
rect 8477 3088 12223 3090
rect 8477 3032 8482 3088
rect 8538 3032 12162 3088
rect 12218 3032 12223 3088
rect 8477 3030 12223 3032
rect 8477 3027 8543 3030
rect 12157 3027 12223 3030
rect 12341 3090 12407 3093
rect 14046 3090 14106 3166
rect 21725 3224 22987 3226
rect 21725 3168 21730 3224
rect 21786 3168 22926 3224
rect 22982 3168 22987 3224
rect 21725 3166 22987 3168
rect 21725 3163 21791 3166
rect 22921 3163 22987 3166
rect 15653 3090 15719 3093
rect 12341 3088 13922 3090
rect 12341 3032 12346 3088
rect 12402 3032 13922 3088
rect 12341 3030 13922 3032
rect 14046 3088 15719 3090
rect 14046 3032 15658 3088
rect 15714 3032 15719 3088
rect 14046 3030 15719 3032
rect 12341 3027 12407 3030
rect 5625 2954 5691 2957
rect 13721 2954 13787 2957
rect 5625 2952 13787 2954
rect 5625 2896 5630 2952
rect 5686 2896 13726 2952
rect 13782 2896 13787 2952
rect 5625 2894 13787 2896
rect 13862 2954 13922 3030
rect 15653 3027 15719 3030
rect 15837 3090 15903 3093
rect 38653 3090 38719 3093
rect 15837 3088 38719 3090
rect 15837 3032 15842 3088
rect 15898 3032 38658 3088
rect 38714 3032 38719 3088
rect 15837 3030 38719 3032
rect 15837 3027 15903 3030
rect 38653 3027 38719 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 15837 2954 15903 2957
rect 39665 2954 39731 2957
rect 13862 2894 15762 2954
rect 5625 2891 5691 2894
rect 13721 2891 13787 2894
rect 0 2818 120 2848
rect 1209 2818 1275 2821
rect 0 2816 1275 2818
rect 0 2760 1214 2816
rect 1270 2760 1275 2816
rect 0 2758 1275 2760
rect 15702 2818 15762 2894
rect 15837 2952 39731 2954
rect 15837 2896 15842 2952
rect 15898 2896 39670 2952
rect 39726 2896 39731 2952
rect 15837 2894 39731 2896
rect 15837 2891 15903 2894
rect 39665 2891 39731 2894
rect 17401 2818 17467 2821
rect 15702 2816 17467 2818
rect 15702 2760 17406 2816
rect 17462 2760 17467 2816
rect 15702 2758 17467 2760
rect 0 2728 120 2758
rect 1209 2755 1275 2758
rect 17401 2755 17467 2758
rect 22001 2818 22067 2821
rect 25589 2818 25655 2821
rect 22001 2816 25655 2818
rect 22001 2760 22006 2816
rect 22062 2760 25594 2816
rect 25650 2760 25655 2816
rect 22001 2758 25655 2760
rect 22001 2755 22067 2758
rect 25589 2755 25655 2758
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 39021 2755 39087 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 19517 2684 19583 2685
rect 19517 2682 19564 2684
rect 19472 2680 19564 2682
rect 19472 2624 19522 2680
rect 19472 2622 19564 2624
rect 19517 2620 19564 2622
rect 19628 2620 19634 2684
rect 19517 2619 19583 2620
rect 0 2546 120 2576
rect 1025 2546 1091 2549
rect 0 2544 1091 2546
rect 0 2488 1030 2544
rect 1086 2488 1091 2544
rect 0 2486 1091 2488
rect 0 2456 120 2486
rect 1025 2483 1091 2486
rect 3233 2546 3299 2549
rect 25313 2546 25379 2549
rect 3233 2544 25379 2546
rect 3233 2488 3238 2544
rect 3294 2488 25318 2544
rect 25374 2488 25379 2544
rect 3233 2486 25379 2488
rect 3233 2483 3299 2486
rect 25313 2483 25379 2486
rect 38469 2546 38535 2549
rect 40880 2546 41000 2576
rect 38469 2544 41000 2546
rect 38469 2488 38474 2544
rect 38530 2488 41000 2544
rect 38469 2486 41000 2488
rect 38469 2483 38535 2486
rect 40880 2456 41000 2486
rect 0 2274 120 2304
rect 197 2274 263 2277
rect 0 2272 263 2274
rect 0 2216 202 2272
rect 258 2216 263 2272
rect 0 2214 263 2216
rect 0 2184 120 2214
rect 197 2211 263 2214
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 0 2002 120 2032
rect 749 2002 815 2005
rect 0 2000 815 2002
rect 0 1944 754 2000
rect 810 1944 815 2000
rect 0 1942 815 1944
rect 0 1912 120 1942
rect 749 1939 815 1942
rect 20437 2002 20503 2005
rect 35709 2002 35775 2005
rect 20437 2000 35775 2002
rect 20437 1944 20442 2000
rect 20498 1944 35714 2000
rect 35770 1944 35775 2000
rect 20437 1942 35775 1944
rect 20437 1939 20503 1942
rect 35709 1939 35775 1942
rect 37917 2002 37983 2005
rect 40880 2002 41000 2032
rect 37917 2000 41000 2002
rect 37917 1944 37922 2000
rect 37978 1944 41000 2000
rect 37917 1942 41000 1944
rect 37917 1939 37983 1942
rect 40880 1912 41000 1942
rect 24577 1866 24643 1869
rect 33869 1866 33935 1869
rect 24577 1864 33935 1866
rect 24577 1808 24582 1864
rect 24638 1808 33874 1864
rect 33930 1808 33935 1864
rect 24577 1806 33935 1808
rect 24577 1803 24643 1806
rect 33869 1803 33935 1806
rect 0 1730 120 1760
rect 381 1730 447 1733
rect 0 1728 447 1730
rect 0 1672 386 1728
rect 442 1672 447 1728
rect 0 1670 447 1672
rect 0 1640 120 1670
rect 381 1667 447 1670
rect 4061 1730 4127 1733
rect 37825 1730 37891 1733
rect 4061 1728 37891 1730
rect 4061 1672 4066 1728
rect 4122 1672 37830 1728
rect 37886 1672 37891 1728
rect 4061 1670 37891 1672
rect 4061 1667 4127 1670
rect 37825 1667 37891 1670
rect 38285 1730 38351 1733
rect 40880 1730 41000 1760
rect 38285 1728 41000 1730
rect 38285 1672 38290 1728
rect 38346 1672 41000 1728
rect 38285 1670 41000 1672
rect 38285 1667 38351 1670
rect 40880 1640 41000 1670
rect 6453 1594 6519 1597
rect 38929 1594 38995 1597
rect 6453 1592 38995 1594
rect 6453 1536 6458 1592
rect 6514 1536 38934 1592
rect 38990 1536 38995 1592
rect 6453 1534 38995 1536
rect 6453 1531 6519 1534
rect 38929 1531 38995 1534
rect 0 1458 120 1488
rect 1209 1458 1275 1461
rect 0 1456 1275 1458
rect 0 1400 1214 1456
rect 1270 1400 1275 1456
rect 0 1398 1275 1400
rect 0 1368 120 1398
rect 1209 1395 1275 1398
rect 38653 1458 38719 1461
rect 40880 1458 41000 1488
rect 38653 1456 41000 1458
rect 38653 1400 38658 1456
rect 38714 1400 41000 1456
rect 38653 1398 41000 1400
rect 38653 1395 38719 1398
rect 40880 1368 41000 1398
rect 36353 1322 36419 1325
rect 38377 1322 38443 1325
rect 36353 1320 38443 1322
rect 36353 1264 36358 1320
rect 36414 1264 38382 1320
rect 38438 1264 38443 1320
rect 36353 1262 38443 1264
rect 36353 1259 36419 1262
rect 38377 1259 38443 1262
rect 27337 642 27403 645
rect 37641 642 37707 645
rect 27337 640 37707 642
rect 27337 584 27342 640
rect 27398 584 37646 640
rect 37702 584 37707 640
rect 27337 582 37707 584
rect 27337 579 27403 582
rect 37641 579 37707 582
rect 17677 506 17743 509
rect 29545 506 29611 509
rect 17677 504 29611 506
rect 17677 448 17682 504
rect 17738 448 29550 504
rect 29606 448 29611 504
rect 17677 446 29611 448
rect 17677 443 17743 446
rect 29545 443 29611 446
rect 23197 370 23263 373
rect 37089 370 37155 373
rect 23197 368 37155 370
rect 23197 312 23202 368
rect 23258 312 37094 368
rect 37150 312 37155 368
rect 23197 310 37155 312
rect 23197 307 23263 310
rect 37089 307 37155 310
rect 21817 234 21883 237
rect 37181 234 37247 237
rect 21817 232 37247 234
rect 21817 176 21822 232
rect 21878 176 37186 232
rect 37242 176 37247 232
rect 21817 174 37247 176
rect 21817 171 21883 174
rect 37181 171 37247 174
rect 16297 98 16363 101
rect 31569 98 31635 101
rect 16297 96 31635 98
rect 16297 40 16302 96
rect 16358 40 31574 96
rect 31630 40 31635 96
rect 16297 38 31635 40
rect 16297 35 16363 38
rect 31569 35 31635 38
<< via3 >>
rect 28948 10100 29012 10164
rect 38332 9692 38396 9756
rect 28580 9420 28644 9484
rect 37228 9284 37292 9348
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 19748 8604 19812 8668
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 37228 7652 37292 7716
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 20852 7516 20916 7580
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 19380 7032 19444 7036
rect 19380 6976 19430 7032
rect 19430 6976 19444 7032
rect 19380 6972 19444 6976
rect 19564 7032 19628 7036
rect 19564 6976 19614 7032
rect 19614 6976 19628 7032
rect 19564 6972 19628 6976
rect 28580 6836 28644 6900
rect 28948 6836 29012 6900
rect 38332 6896 38396 6900
rect 38332 6840 38382 6896
rect 38382 6840 38396 6896
rect 38332 6836 38396 6840
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 20852 6020 20916 6084
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 19380 5944 19444 5948
rect 19380 5888 19394 5944
rect 19394 5888 19444 5944
rect 19380 5884 19444 5888
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 19748 3708 19812 3772
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 19564 2680 19628 2684
rect 19564 2624 19578 2680
rect 19578 2624 19628 2680
rect 19564 2620 19628 2624
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 0 3324 2144
rect 7944 8192 8264 11250
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 7944 6016 8264 7040
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 0 8264 2688
rect 9004 8736 9324 11250
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 9004 6560 9324 7584
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 9004 5472 9324 6496
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 9004 4384 9324 5408
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 9004 3296 9324 4320
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13944 3840 14264 4864
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13944 0 14264 2688
rect 15004 8736 15324 11250
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 15004 7648 15324 8672
rect 19747 8668 19813 8669
rect 19747 8604 19748 8668
rect 19812 8604 19813 8668
rect 19747 8603 19813 8604
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 19379 7036 19445 7037
rect 19379 6972 19380 7036
rect 19444 6972 19445 7036
rect 19379 6971 19445 6972
rect 19563 7036 19629 7037
rect 19563 6972 19564 7036
rect 19628 6972 19629 7036
rect 19563 6971 19629 6972
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 19382 5949 19442 6971
rect 19379 5948 19445 5949
rect 19379 5884 19380 5948
rect 19444 5884 19445 5948
rect 19379 5883 19445 5884
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 19566 2685 19626 6971
rect 19750 3773 19810 8603
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 20851 7580 20917 7581
rect 20851 7516 20852 7580
rect 20916 7516 20917 7580
rect 20851 7515 20917 7516
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 20854 6085 20914 7515
rect 21004 6560 21324 7584
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 20851 6084 20917 6085
rect 20851 6020 20852 6084
rect 20916 6020 20917 6084
rect 20851 6019 20917 6020
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19747 3772 19813 3773
rect 19747 3708 19748 3772
rect 19812 3708 19813 3772
rect 19747 3707 19813 3708
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19563 2684 19629 2685
rect 19563 2620 19564 2684
rect 19628 2620 19629 2684
rect 19563 2619 19629 2620
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 19944 0 20264 2688
rect 21004 5472 21324 6496
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 21004 0 21324 2144
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 28947 10164 29013 10165
rect 28947 10100 28948 10164
rect 29012 10100 29013 10164
rect 28947 10099 29013 10100
rect 28579 9484 28645 9485
rect 28579 9420 28580 9484
rect 28644 9420 28645 9484
rect 28579 9419 28645 9420
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 28582 6901 28642 9419
rect 28950 6901 29010 10099
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 28579 6900 28645 6901
rect 28579 6836 28580 6900
rect 28644 6836 28645 6900
rect 28579 6835 28645 6836
rect 28947 6900 29013 6901
rect 28947 6836 28948 6900
rect 29012 6836 29013 6900
rect 28947 6835 29013 6836
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 37227 9348 37293 9349
rect 37227 9284 37228 9348
rect 37292 9284 37293 9348
rect 37227 9283 37293 9284
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 37230 7717 37290 9283
rect 37944 8192 38264 11250
rect 38331 9756 38397 9757
rect 38331 9692 38332 9756
rect 38396 9692 38397 9756
rect 38331 9691 38397 9692
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37227 7716 37293 7717
rect 37227 7652 37228 7716
rect 37292 7652 37293 7716
rect 37227 7651 37293 7652
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 38334 6901 38394 9691
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 38331 6900 38397 6901
rect 38331 6836 38332 6900
rect 38396 6836 38397 6900
rect 38331 6835 38397 6836
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__mux4_1  _000_
timestamp -3599
transform -1 0 21712 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  _001_
timestamp -3599
transform 1 0 29348 0 -1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  _002_
timestamp -3599
transform -1 0 8648 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _003_
timestamp -3599
transform -1 0 15916 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _004_
timestamp -3599
transform -1 0 11132 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  _005_
timestamp -3599
transform -1 0 23828 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  _006_
timestamp -3599
transform -1 0 12236 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  _007_
timestamp -3599
transform -1 0 26864 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  _008_
timestamp -3599
transform 1 0 25760 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _009_
timestamp -3599
transform -1 0 10304 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _010_
timestamp -3599
transform 1 0 22264 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _011_
timestamp -3599
transform -1 0 9476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _012_
timestamp -3599
transform -1 0 16008 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _013_
timestamp -3599
transform -1 0 6900 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _014_
timestamp -3599
transform 1 0 27508 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _015_
timestamp -3599
transform 1 0 18400 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _016_
timestamp -3599
transform 1 0 26956 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _017_
timestamp -3599
transform 1 0 10212 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _018_
timestamp -3599
transform 1 0 21620 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _019_
timestamp -3599
transform 1 0 8280 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _020_
timestamp -3599
transform -1 0 15456 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _021_
timestamp -3599
transform -1 0 8280 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _022_
timestamp -3599
transform 1 0 27416 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _023_
timestamp -3599
transform -1 0 21344 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  _024_
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _025_
timestamp -3599
transform -1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _026_
timestamp -3599
transform 1 0 16928 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _027_
timestamp -3599
transform 1 0 17848 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _028_
timestamp -3599
transform -1 0 16744 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _029_
timestamp -3599
transform -1 0 16560 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _030_
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _031_
timestamp -3599
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _032_
timestamp -3599
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _033_
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _034_
timestamp -3599
transform 1 0 18032 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _035_
timestamp -3599
transform 1 0 18032 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _036_
timestamp -3599
transform -1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _037_
timestamp -3599
transform -1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _038_
timestamp -3599
transform 1 0 25576 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _039_
timestamp -3599
transform 1 0 26036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _040_
timestamp -3599
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _041_
timestamp -3599
transform 1 0 18308 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _042_
timestamp -3599
transform 1 0 28244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _043_
timestamp -3599
transform -1 0 29348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _044_
timestamp -3599
transform 1 0 3956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _045_
timestamp -3599
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _046_
timestamp -3599
transform 1 0 12880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _047_
timestamp -3599
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _048_
timestamp -3599
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _049_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _050_
timestamp -3599
transform 1 0 21988 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _051_
timestamp -3599
transform 1 0 21160 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _052_
timestamp -3599
transform 1 0 5612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _053_
timestamp -3599
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _054_
timestamp -3599
transform 1 0 25024 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _055_
timestamp -3599
transform 1 0 24932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _056_
timestamp -3599
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _057_
timestamp -3599
transform 1 0 23092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _058_
timestamp -3599
transform -1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _059_
timestamp -3599
transform -1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _060_
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _061_
timestamp -3599
transform 1 0 16744 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _062_
timestamp -3599
transform -1 0 11408 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _063_
timestamp -3599
transform -1 0 11408 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _064_
timestamp -3599
transform 1 0 11776 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _065_
timestamp -3599
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _066_
timestamp -3599
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _067_
timestamp -3599
transform 1 0 6716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _068_
timestamp -3599
transform 1 0 28336 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _069_
timestamp -3599
transform 1 0 27232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _070_
timestamp -3599
transform -1 0 25576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _071_
timestamp -3599
transform -1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp -3599
transform 1 0 18032 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp -3599
transform 1 0 17664 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp -3599
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp -3599
transform -1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _077_
timestamp -3599
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _078_
timestamp -3599
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp -3599
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp -3599
transform 1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp -3599
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _083_
timestamp -3599
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _084_
timestamp -3599
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp -3599
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _086_
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp -3599
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _088_
timestamp -3599
transform 1 0 24932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _089_
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _090_
timestamp -3599
transform 1 0 22448 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp -3599
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _092_
timestamp -3599
transform 1 0 14996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _093_
timestamp -3599
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _094_
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _095_
timestamp -3599
transform 1 0 11684 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _096_
timestamp -3599
transform 1 0 11500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp -3599
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp -3599
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _100_
timestamp -3599
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp -3599
transform 1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp -3599
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_
timestamp -3599
transform 1 0 24748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp -3599
transform 1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp -3599
transform -1 0 29164 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _106_
timestamp -3599
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp -3599
transform -1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp -3599
transform -1 0 33304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp -3599
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp -3599
transform 1 0 36984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp -3599
transform 1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp -3599
transform 1 0 38364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp -3599
transform -1 0 34132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp -3599
transform -1 0 34408 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp -3599
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp -3599
transform 1 0 37536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp -3599
transform 1 0 36984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp -3599
transform -1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp -3599
transform -1 0 30636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp -3599
transform -1 0 34408 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp -3599
transform 1 0 37904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp -3599
transform 1 0 38180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp -3599
transform -1 0 36616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp -3599
transform -1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp -3599
transform -1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp -3599
transform -1 0 30268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp -3599
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp -3599
transform -1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _129_
timestamp -3599
transform -1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp -3599
transform -1 0 29900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp -3599
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp -3599
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp -3599
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _134_
timestamp -3599
transform -1 0 24656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp -3599
transform 1 0 12144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _137_
timestamp -3599
transform -1 0 20976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp -3599
transform -1 0 29992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp -3599
transform -1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp -3599
transform 1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _142_
timestamp -3599
transform -1 0 24288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp -3599
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp -3599
transform -1 0 28796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp -3599
transform -1 0 38732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp -3599
transform -1 0 37628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp -3599
transform -1 0 38364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp -3599
transform -1 0 37996 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp -3599
transform -1 0 37720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp -3599
transform -1 0 38364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp -3599
transform -1 0 36984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp -3599
transform -1 0 38456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp -3599
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _154_
timestamp -3599
transform -1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp -3599
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp -3599
transform -1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp -3599
transform -1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp -3599
transform -1 0 10212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _160_
timestamp -3599
transform -1 0 28520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp -3599
transform 1 0 19504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp -3599
transform -1 0 28612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp -3599
transform 1 0 5244 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp -3599
transform -1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _166_
timestamp -3599
transform -1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp -3599
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp -3599
transform -1 0 28244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp -3599
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _170_
timestamp -3599
transform -1 0 30544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp -3599
transform -1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp -3599
transform -1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _174_
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp -3599
transform -1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _177_
timestamp -3599
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 38824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 38088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 32752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform -1 0 33580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 37444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform -1 0 38824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 2576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform -1 0 9476 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform -1 0 9200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 37812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp -3599
transform -1 0 38916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp -3599
transform -1 0 9476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp -3599
transform -1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp -3599
transform -1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp -3599
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp -3599
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp -3599
transform 1 0 18952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout14
timestamp -3599
transform -1 0 18584 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp -3599
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp -3599
transform -1 0 11408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp -3599
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp -3599
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35
timestamp -3599
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43
timestamp -3599
transform 1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50
timestamp -3599
transform 1 0 5704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65
timestamp -3599
transform 1 0 7084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73
timestamp -3599
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp -3599
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95
timestamp -3599
transform 1 0 9844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_103
timestamp -3599
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp -3599
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636964856
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636964856
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp -3599
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636964856
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_239
timestamp 1636964856
transform 1 0 23092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp -3599
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636964856
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636964856
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp -3599
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636964856
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_293
timestamp -3599
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp -3599
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp -3599
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636964856
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636964856
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp -3599
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636964856
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636964856
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp -3599
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636964856
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636964856
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp -3599
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1636964856
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1636964856
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_43
timestamp -3599
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp -3599
transform 1 0 6624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp -3599
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp -3599
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_100
timestamp 1636964856
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636964856
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp -3599
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_196
timestamp 1636964856
transform 1 0 19136 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_208
timestamp 1636964856
transform 1 0 20240 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_220
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_250
timestamp 1636964856
transform 1 0 24104 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_262
timestamp 1636964856
transform 1 0 25208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp -3599
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_281
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_311
timestamp 1636964856
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_323
timestamp 1636964856
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636964856
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636964856
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636964856
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636964856
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp -3599
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp -3599
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp -3599
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_402
timestamp -3599
transform 1 0 38088 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_12
timestamp 1636964856
transform 1 0 2208 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp -3599
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp -3599
transform 1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp -3599
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp -3599
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_123
timestamp 1636964856
transform 1 0 12420 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp -3599
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_157
timestamp -3599
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp -3599
transform 1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636964856
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp -3599
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp -3599
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_256
timestamp 1636964856
transform 1 0 24656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_268
timestamp 1636964856
transform 1 0 25760 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp -3599
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_323
timestamp 1636964856
transform 1 0 30820 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_335
timestamp -3599
transform 1 0 31924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_341
timestamp -3599
transform 1 0 32476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_350
timestamp -3599
transform 1 0 33304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp -3599
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636964856
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636964856
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_389
timestamp -3599
transform 1 0 36892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_398
timestamp -3599
transform 1 0 37720 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_9
timestamp 1636964856
transform 1 0 1932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp -3599
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_80
timestamp 1636964856
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp -3599
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_97
timestamp -3599
transform 1 0 10028 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp -3599
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp -3599
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_198
timestamp 1636964856
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_210
timestamp 1636964856
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp -3599
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_252
timestamp 1636964856
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_264
timestamp 1636964856
transform 1 0 25392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp -3599
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp -3599
transform 1 0 27324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp -3599
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp -3599
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636964856
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636964856
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636964856
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636964856
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp -3599
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp -3599
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp -3599
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_9
timestamp 1636964856
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp -3599
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp -3599
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636964856
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp -3599
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636964856
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636964856
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp -3599
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_172
timestamp -3599
transform 1 0 16928 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp -3599
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636964856
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp -3599
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp -3599
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636964856
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636964856
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636964856
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_289
timestamp -3599
transform 1 0 27692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_314
timestamp 1636964856
transform 1 0 29992 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_326
timestamp 1636964856
transform 1 0 31096 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_338
timestamp 1636964856
transform 1 0 32200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_350
timestamp 1636964856
transform 1 0 33304 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp -3599
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636964856
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636964856
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636964856
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_401
timestamp -3599
transform 1 0 37996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_409
timestamp -3599
transform 1 0 38732 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1636964856
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1636964856
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_33
timestamp -3599
transform 1 0 4140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp -3599
transform 1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636964856
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636964856
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636964856
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636964856
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp -3599
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -3599
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636964856
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636964856
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636964856
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636964856
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp -3599
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636964856
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636964856
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636964856
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_205
timestamp -3599
transform 1 0 19964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_211
timestamp -3599
transform 1 0 20516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp -3599
transform 1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp -3599
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636964856
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636964856
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636964856
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636964856
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp -3599
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp -3599
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_307
timestamp 1636964856
transform 1 0 29348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 1636964856
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp -3599
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp -3599
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636964856
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636964856
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636964856
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636964856
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp -3599
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp -3599
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp -3599
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_12
timestamp 1636964856
transform 1 0 2208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp -3599
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636964856
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636964856
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636964856
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636964856
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp -3599
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636964856
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_121
timestamp -3599
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp -3599
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp -3599
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_144
timestamp 1636964856
transform 1 0 14352 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_156
timestamp 1636964856
transform 1 0 15456 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_168
timestamp 1636964856
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_180
timestamp 1636964856
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp -3599
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_212
timestamp 1636964856
transform 1 0 20608 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_224
timestamp 1636964856
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_236
timestamp 1636964856
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp -3599
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp -3599
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_283
timestamp 1636964856
transform 1 0 27140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_295
timestamp 1636964856
transform 1 0 28244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636964856
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636964856
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636964856
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636964856
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp -3599
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp -3599
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636964856
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636964856
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp -3599
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_397
timestamp -3599
transform 1 0 37628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_406
timestamp -3599
transform 1 0 38456 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_13
timestamp 1636964856
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_25
timestamp 1636964856
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_37
timestamp 1636964856
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp -3599
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp -3599
transform 1 0 7452 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_91
timestamp -3599
transform 1 0 9476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp -3599
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp -3599
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636964856
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp -3599
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_228
timestamp 1636964856
transform 1 0 22080 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_240
timestamp 1636964856
transform 1 0 23184 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_252
timestamp -3599
transform 1 0 24288 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_258
timestamp -3599
transform 1 0 24840 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636964856
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636964856
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp -3599
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636964856
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636964856
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636964856
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636964856
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp -3599
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_405
timestamp -3599
transform 1 0 38364 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636964856
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -3599
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636964856
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp -3599
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp -3599
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_66
timestamp -3599
transform 1 0 7176 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636964856
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_235
timestamp -3599
transform 1 0 22724 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_266
timestamp -3599
transform 1 0 25576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp -3599
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636964856
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636964856
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636964856
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636964856
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp -3599
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636964856
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp -3599
transform 1 0 35788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_385
timestamp -3599
transform 1 0 36524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_397
timestamp -3599
transform 1 0 37628 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_415
timestamp -3599
transform 1 0 39284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_16
timestamp -3599
transform 1 0 2576 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1636964856
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1636964856
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp -3599
transform 1 0 10212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp -3599
transform 1 0 11960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_134
timestamp -3599
transform 1 0 13432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_156
timestamp -3599
transform 1 0 15456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp -3599
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636964856
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_181
timestamp -3599
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_199
timestamp -3599
transform 1 0 19412 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636964856
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636964856
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp -3599
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp -3599
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636964856
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_317
timestamp -3599
transform 1 0 30268 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_324
timestamp 1636964856
transform 1 0 30912 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636964856
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp -3599
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_357
timestamp -3599
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_362
timestamp 1636964856
transform 1 0 34408 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_374
timestamp -3599
transform 1 0 35512 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_382
timestamp -3599
transform 1 0 36248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp -3599
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp -3599
transform 1 0 4048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_46
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_58
timestamp -3599
transform 1 0 6440 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp -3599
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp -3599
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_95
timestamp -3599
transform 1 0 9844 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp -3599
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_106
timestamp -3599
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp -3599
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp -3599
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp -3599
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp -3599
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp -3599
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_134
timestamp -3599
transform 1 0 13432 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp -3599
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_148
timestamp -3599
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp -3599
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp -3599
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_166
timestamp 1636964856
transform 1 0 16376 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp -3599
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp -3599
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp -3599
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_202
timestamp -3599
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_206
timestamp -3599
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_210
timestamp -3599
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_216
timestamp 1636964856
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_228
timestamp 1636964856
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1636964856
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_259
timestamp -3599
transform 1 0 24932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_264
timestamp -3599
transform 1 0 25392 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_278
timestamp 1636964856
transform 1 0 26680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_290
timestamp -3599
transform 1 0 27784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_296
timestamp -3599
transform 1 0 28336 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_300
timestamp -3599
transform 1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp -3599
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_318
timestamp -3599
transform 1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_343
timestamp 1636964856
transform 1 0 32660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp -3599
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp -3599
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_369
timestamp -3599
transform 1 0 35052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_379
timestamp -3599
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_391
timestamp -3599
transform 1 0 37076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_395
timestamp -3599
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_13
timestamp -3599
transform 1 0 2300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_85
timestamp -3599
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp -3599
transform 1 0 10120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp -3599
transform 1 0 17204 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp -3599
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp -3599
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp -3599
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp -3599
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_329
timestamp -3599
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp -3599
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_340
timestamp -3599
transform 1 0 32384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp -3599
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp -3599
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_409
timestamp -3599
transform 1 0 38732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -3599
transform 1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -3599
transform -1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -3599
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -3599
transform 1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -3599
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -3599
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp -3599
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -3599
transform 1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp -3599
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp -3599
transform 1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -3599
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -3599
transform 1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -3599
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp -3599
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp -3599
transform -1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp -3599
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -3599
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp -3599
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp -3599
transform -1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp -3599
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp -3599
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp -3599
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp -3599
transform -1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp -3599
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp -3599
transform -1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp -3599
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp -3599
transform -1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp -3599
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp -3599
transform -1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp -3599
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp -3599
transform -1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp -3599
transform 1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp -3599
transform -1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp -3599
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp -3599
transform -1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp -3599
transform -1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp -3599
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp -3599
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp -3599
transform 1 0 24380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input55
timestamp -3599
transform -1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp -3599
transform -1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp -3599
transform -1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp -3599
transform 1 0 25300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input59
timestamp -3599
transform 1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp -3599
transform -1 0 26496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp -3599
transform 1 0 27876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp -3599
transform -1 0 30912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input64
timestamp -3599
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp -3599
transform -1 0 31832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66
timestamp -3599
transform -1 0 32108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp -3599
transform -1 0 32384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp -3599
transform 1 0 28152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input69
timestamp -3599
transform -1 0 28704 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp -3599
transform 1 0 29532 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input71
timestamp -3599
transform -1 0 29256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp -3599
transform -1 0 29440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input73
timestamp -3599
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp -3599
transform -1 0 30084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp -3599
transform -1 0 30360 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp -3599
transform 1 0 30452 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output77
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp -3599
transform 1 0 38456 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform 1 0 38916 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 38456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 38272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform -1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform -1 0 35972 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform -1 0 36892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform 1 0 36156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform 1 0 36708 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform -1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform -1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform 1 0 38364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 32936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform 1 0 33304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform 1 0 33672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform 1 0 34040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform -1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform -1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform -1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform 1 0 35420 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform 1 0 35788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform -1 0 3680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 2576 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform -1 0 3312 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform -1 0 4508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform -1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 5336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 5152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform -1 0 6440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform -1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform -1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform 1 0 7176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform -1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform -1 0 7912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform -1 0 8648 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform -1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform -1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform -1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform -1 0 9936 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform -1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform -1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform -1 0 10672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp -3599
transform -1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp -3599
transform -1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp -3599
transform -1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp -3599
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp -3599
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp -3599
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp -3599
transform -1 0 17204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp -3599
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp -3599
transform -1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp -3599
transform -1 0 13892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp -3599
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp -3599
transform -1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp -3599
transform 1 0 14352 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp -3599
transform -1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp -3599
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp -3599
transform -1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp -3599
transform -1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp -3599
transform -1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output181
timestamp -3599
transform -1 0 32660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output182
timestamp -3599
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp -3599
transform -1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp -3599
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp -3599
transform -1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp -3599
transform -1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp -3599
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp -3599
transform -1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp -3599
transform -1 0 11224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_EF_DAC8_190
timestamp -3599
transform -1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 17590 11194 17646 11250 0 FreeSans 224 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 13542 0 13598 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 27342 0 27398 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 28722 0 28778 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 30102 0 30158 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 31482 0 31538 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 32862 0 32918 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 34242 0 34298 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 35622 0 35678 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 37002 0 37058 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 38382 0 38438 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 39762 0 39818 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 14922 0 14978 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 16302 0 16358 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 17682 0 17738 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 19062 0 19118 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 20442 0 20498 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 21822 0 21878 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 23202 0 23258 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 24582 0 24638 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 25962 0 26018 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 32494 11194 32550 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 35254 11194 35310 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 35530 11194 35586 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 35806 11194 35862 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 36082 11194 36138 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 36358 11194 36414 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 36634 11194 36690 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 36910 11194 36966 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 37186 11194 37242 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 37462 11194 37518 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 37738 11194 37794 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 32770 11194 32826 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 33046 11194 33102 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 33322 11194 33378 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 33598 11194 33654 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 33874 11194 33930 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 34150 11194 34206 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 34426 11194 34482 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 34702 11194 34758 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 34978 11194 35034 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 3238 11194 3294 11250 0 FreeSans 224 0 0 0 N1BEG[0]
port 105 nsew signal output
flabel metal2 s 3514 11194 3570 11250 0 FreeSans 224 0 0 0 N1BEG[1]
port 106 nsew signal output
flabel metal2 s 3790 11194 3846 11250 0 FreeSans 224 0 0 0 N1BEG[2]
port 107 nsew signal output
flabel metal2 s 4066 11194 4122 11250 0 FreeSans 224 0 0 0 N1BEG[3]
port 108 nsew signal output
flabel metal2 s 4342 11194 4398 11250 0 FreeSans 224 0 0 0 N2BEG[0]
port 109 nsew signal output
flabel metal2 s 4618 11194 4674 11250 0 FreeSans 224 0 0 0 N2BEG[1]
port 110 nsew signal output
flabel metal2 s 4894 11194 4950 11250 0 FreeSans 224 0 0 0 N2BEG[2]
port 111 nsew signal output
flabel metal2 s 5170 11194 5226 11250 0 FreeSans 224 0 0 0 N2BEG[3]
port 112 nsew signal output
flabel metal2 s 5446 11194 5502 11250 0 FreeSans 224 0 0 0 N2BEG[4]
port 113 nsew signal output
flabel metal2 s 5722 11194 5778 11250 0 FreeSans 224 0 0 0 N2BEG[5]
port 114 nsew signal output
flabel metal2 s 5998 11194 6054 11250 0 FreeSans 224 0 0 0 N2BEG[6]
port 115 nsew signal output
flabel metal2 s 6274 11194 6330 11250 0 FreeSans 224 0 0 0 N2BEG[7]
port 116 nsew signal output
flabel metal2 s 6550 11194 6606 11250 0 FreeSans 224 0 0 0 N2BEGb[0]
port 117 nsew signal output
flabel metal2 s 6826 11194 6882 11250 0 FreeSans 224 0 0 0 N2BEGb[1]
port 118 nsew signal output
flabel metal2 s 7102 11194 7158 11250 0 FreeSans 224 0 0 0 N2BEGb[2]
port 119 nsew signal output
flabel metal2 s 7378 11194 7434 11250 0 FreeSans 224 0 0 0 N2BEGb[3]
port 120 nsew signal output
flabel metal2 s 7654 11194 7710 11250 0 FreeSans 224 0 0 0 N2BEGb[4]
port 121 nsew signal output
flabel metal2 s 7930 11194 7986 11250 0 FreeSans 224 0 0 0 N2BEGb[5]
port 122 nsew signal output
flabel metal2 s 8206 11194 8262 11250 0 FreeSans 224 0 0 0 N2BEGb[6]
port 123 nsew signal output
flabel metal2 s 8482 11194 8538 11250 0 FreeSans 224 0 0 0 N2BEGb[7]
port 124 nsew signal output
flabel metal2 s 8758 11194 8814 11250 0 FreeSans 224 0 0 0 N4BEG[0]
port 125 nsew signal output
flabel metal2 s 11518 11194 11574 11250 0 FreeSans 224 0 0 0 N4BEG[10]
port 126 nsew signal output
flabel metal2 s 11794 11194 11850 11250 0 FreeSans 224 0 0 0 N4BEG[11]
port 127 nsew signal output
flabel metal2 s 12070 11194 12126 11250 0 FreeSans 224 0 0 0 N4BEG[12]
port 128 nsew signal output
flabel metal2 s 12346 11194 12402 11250 0 FreeSans 224 0 0 0 N4BEG[13]
port 129 nsew signal output
flabel metal2 s 12622 11194 12678 11250 0 FreeSans 224 0 0 0 N4BEG[14]
port 130 nsew signal output
flabel metal2 s 12898 11194 12954 11250 0 FreeSans 224 0 0 0 N4BEG[15]
port 131 nsew signal output
flabel metal2 s 9034 11194 9090 11250 0 FreeSans 224 0 0 0 N4BEG[1]
port 132 nsew signal output
flabel metal2 s 9310 11194 9366 11250 0 FreeSans 224 0 0 0 N4BEG[2]
port 133 nsew signal output
flabel metal2 s 9586 11194 9642 11250 0 FreeSans 224 0 0 0 N4BEG[3]
port 134 nsew signal output
flabel metal2 s 9862 11194 9918 11250 0 FreeSans 224 0 0 0 N4BEG[4]
port 135 nsew signal output
flabel metal2 s 10138 11194 10194 11250 0 FreeSans 224 0 0 0 N4BEG[5]
port 136 nsew signal output
flabel metal2 s 10414 11194 10470 11250 0 FreeSans 224 0 0 0 N4BEG[6]
port 137 nsew signal output
flabel metal2 s 10690 11194 10746 11250 0 FreeSans 224 0 0 0 N4BEG[7]
port 138 nsew signal output
flabel metal2 s 10966 11194 11022 11250 0 FreeSans 224 0 0 0 N4BEG[8]
port 139 nsew signal output
flabel metal2 s 11242 11194 11298 11250 0 FreeSans 224 0 0 0 N4BEG[9]
port 140 nsew signal output
flabel metal2 s 13174 11194 13230 11250 0 FreeSans 224 0 0 0 NN4BEG[0]
port 141 nsew signal output
flabel metal2 s 15934 11194 15990 11250 0 FreeSans 224 0 0 0 NN4BEG[10]
port 142 nsew signal output
flabel metal2 s 16210 11194 16266 11250 0 FreeSans 224 0 0 0 NN4BEG[11]
port 143 nsew signal output
flabel metal2 s 16486 11194 16542 11250 0 FreeSans 224 0 0 0 NN4BEG[12]
port 144 nsew signal output
flabel metal2 s 16762 11194 16818 11250 0 FreeSans 224 0 0 0 NN4BEG[13]
port 145 nsew signal output
flabel metal2 s 17038 11194 17094 11250 0 FreeSans 224 0 0 0 NN4BEG[14]
port 146 nsew signal output
flabel metal2 s 17314 11194 17370 11250 0 FreeSans 224 0 0 0 NN4BEG[15]
port 147 nsew signal output
flabel metal2 s 13450 11194 13506 11250 0 FreeSans 224 0 0 0 NN4BEG[1]
port 148 nsew signal output
flabel metal2 s 13726 11194 13782 11250 0 FreeSans 224 0 0 0 NN4BEG[2]
port 149 nsew signal output
flabel metal2 s 14002 11194 14058 11250 0 FreeSans 224 0 0 0 NN4BEG[3]
port 150 nsew signal output
flabel metal2 s 14278 11194 14334 11250 0 FreeSans 224 0 0 0 NN4BEG[4]
port 151 nsew signal output
flabel metal2 s 14554 11194 14610 11250 0 FreeSans 224 0 0 0 NN4BEG[5]
port 152 nsew signal output
flabel metal2 s 14830 11194 14886 11250 0 FreeSans 224 0 0 0 NN4BEG[6]
port 153 nsew signal output
flabel metal2 s 15106 11194 15162 11250 0 FreeSans 224 0 0 0 NN4BEG[7]
port 154 nsew signal output
flabel metal2 s 15382 11194 15438 11250 0 FreeSans 224 0 0 0 NN4BEG[8]
port 155 nsew signal output
flabel metal2 s 15658 11194 15714 11250 0 FreeSans 224 0 0 0 NN4BEG[9]
port 156 nsew signal output
flabel metal2 s 17866 11194 17922 11250 0 FreeSans 224 0 0 0 S1END[0]
port 157 nsew signal input
flabel metal2 s 18142 11194 18198 11250 0 FreeSans 224 0 0 0 S1END[1]
port 158 nsew signal input
flabel metal2 s 18418 11194 18474 11250 0 FreeSans 224 0 0 0 S1END[2]
port 159 nsew signal input
flabel metal2 s 18694 11194 18750 11250 0 FreeSans 224 0 0 0 S1END[3]
port 160 nsew signal input
flabel metal2 s 21178 11194 21234 11250 0 FreeSans 224 0 0 0 S2END[0]
port 161 nsew signal input
flabel metal2 s 21454 11194 21510 11250 0 FreeSans 224 0 0 0 S2END[1]
port 162 nsew signal input
flabel metal2 s 21730 11194 21786 11250 0 FreeSans 224 0 0 0 S2END[2]
port 163 nsew signal input
flabel metal2 s 22006 11194 22062 11250 0 FreeSans 224 0 0 0 S2END[3]
port 164 nsew signal input
flabel metal2 s 22282 11194 22338 11250 0 FreeSans 224 0 0 0 S2END[4]
port 165 nsew signal input
flabel metal2 s 22558 11194 22614 11250 0 FreeSans 224 0 0 0 S2END[5]
port 166 nsew signal input
flabel metal2 s 22834 11194 22890 11250 0 FreeSans 224 0 0 0 S2END[6]
port 167 nsew signal input
flabel metal2 s 23110 11194 23166 11250 0 FreeSans 224 0 0 0 S2END[7]
port 168 nsew signal input
flabel metal2 s 18970 11194 19026 11250 0 FreeSans 224 0 0 0 S2MID[0]
port 169 nsew signal input
flabel metal2 s 19246 11194 19302 11250 0 FreeSans 224 0 0 0 S2MID[1]
port 170 nsew signal input
flabel metal2 s 19522 11194 19578 11250 0 FreeSans 224 0 0 0 S2MID[2]
port 171 nsew signal input
flabel metal2 s 19798 11194 19854 11250 0 FreeSans 224 0 0 0 S2MID[3]
port 172 nsew signal input
flabel metal2 s 20074 11194 20130 11250 0 FreeSans 224 0 0 0 S2MID[4]
port 173 nsew signal input
flabel metal2 s 20350 11194 20406 11250 0 FreeSans 224 0 0 0 S2MID[5]
port 174 nsew signal input
flabel metal2 s 20626 11194 20682 11250 0 FreeSans 224 0 0 0 S2MID[6]
port 175 nsew signal input
flabel metal2 s 20902 11194 20958 11250 0 FreeSans 224 0 0 0 S2MID[7]
port 176 nsew signal input
flabel metal2 s 23386 11194 23442 11250 0 FreeSans 224 0 0 0 S4END[0]
port 177 nsew signal input
flabel metal2 s 26146 11194 26202 11250 0 FreeSans 224 0 0 0 S4END[10]
port 178 nsew signal input
flabel metal2 s 26422 11194 26478 11250 0 FreeSans 224 0 0 0 S4END[11]
port 179 nsew signal input
flabel metal2 s 26698 11194 26754 11250 0 FreeSans 224 0 0 0 S4END[12]
port 180 nsew signal input
flabel metal2 s 26974 11194 27030 11250 0 FreeSans 224 0 0 0 S4END[13]
port 181 nsew signal input
flabel metal2 s 27250 11194 27306 11250 0 FreeSans 224 0 0 0 S4END[14]
port 182 nsew signal input
flabel metal2 s 27526 11194 27582 11250 0 FreeSans 224 0 0 0 S4END[15]
port 183 nsew signal input
flabel metal2 s 23662 11194 23718 11250 0 FreeSans 224 0 0 0 S4END[1]
port 184 nsew signal input
flabel metal2 s 23938 11194 23994 11250 0 FreeSans 224 0 0 0 S4END[2]
port 185 nsew signal input
flabel metal2 s 24214 11194 24270 11250 0 FreeSans 224 0 0 0 S4END[3]
port 186 nsew signal input
flabel metal2 s 24490 11194 24546 11250 0 FreeSans 224 0 0 0 S4END[4]
port 187 nsew signal input
flabel metal2 s 24766 11194 24822 11250 0 FreeSans 224 0 0 0 S4END[5]
port 188 nsew signal input
flabel metal2 s 25042 11194 25098 11250 0 FreeSans 224 0 0 0 S4END[6]
port 189 nsew signal input
flabel metal2 s 25318 11194 25374 11250 0 FreeSans 224 0 0 0 S4END[7]
port 190 nsew signal input
flabel metal2 s 25594 11194 25650 11250 0 FreeSans 224 0 0 0 S4END[8]
port 191 nsew signal input
flabel metal2 s 25870 11194 25926 11250 0 FreeSans 224 0 0 0 S4END[9]
port 192 nsew signal input
flabel metal2 s 27802 11194 27858 11250 0 FreeSans 224 0 0 0 SS4END[0]
port 193 nsew signal input
flabel metal2 s 30562 11194 30618 11250 0 FreeSans 224 0 0 0 SS4END[10]
port 194 nsew signal input
flabel metal2 s 30838 11194 30894 11250 0 FreeSans 224 0 0 0 SS4END[11]
port 195 nsew signal input
flabel metal2 s 31114 11194 31170 11250 0 FreeSans 224 0 0 0 SS4END[12]
port 196 nsew signal input
flabel metal2 s 31390 11194 31446 11250 0 FreeSans 224 0 0 0 SS4END[13]
port 197 nsew signal input
flabel metal2 s 31666 11194 31722 11250 0 FreeSans 224 0 0 0 SS4END[14]
port 198 nsew signal input
flabel metal2 s 31942 11194 31998 11250 0 FreeSans 224 0 0 0 SS4END[15]
port 199 nsew signal input
flabel metal2 s 28078 11194 28134 11250 0 FreeSans 224 0 0 0 SS4END[1]
port 200 nsew signal input
flabel metal2 s 28354 11194 28410 11250 0 FreeSans 224 0 0 0 SS4END[2]
port 201 nsew signal input
flabel metal2 s 28630 11194 28686 11250 0 FreeSans 224 0 0 0 SS4END[3]
port 202 nsew signal input
flabel metal2 s 28906 11194 28962 11250 0 FreeSans 224 0 0 0 SS4END[4]
port 203 nsew signal input
flabel metal2 s 29182 11194 29238 11250 0 FreeSans 224 0 0 0 SS4END[5]
port 204 nsew signal input
flabel metal2 s 29458 11194 29514 11250 0 FreeSans 224 0 0 0 SS4END[6]
port 205 nsew signal input
flabel metal2 s 29734 11194 29790 11250 0 FreeSans 224 0 0 0 SS4END[7]
port 206 nsew signal input
flabel metal2 s 30010 11194 30066 11250 0 FreeSans 224 0 0 0 SS4END[8]
port 207 nsew signal input
flabel metal2 s 30286 11194 30342 11250 0 FreeSans 224 0 0 0 SS4END[9]
port 208 nsew signal input
flabel metal2 s 12162 0 12218 56 0 FreeSans 224 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 32218 11194 32274 11250 0 FreeSans 224 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal2 s 1122 0 1178 56 0 FreeSans 224 0 0 0 VALUE_top0
port 211 nsew signal output
flabel metal2 s 2502 0 2558 56 0 FreeSans 224 0 0 0 VALUE_top1
port 212 nsew signal output
flabel metal2 s 3882 0 3938 56 0 FreeSans 224 0 0 0 VALUE_top2
port 213 nsew signal output
flabel metal2 s 5262 0 5318 56 0 FreeSans 224 0 0 0 VALUE_top3
port 214 nsew signal output
flabel metal2 s 6642 0 6698 56 0 FreeSans 224 0 0 0 VALUE_top4
port 215 nsew signal output
flabel metal2 s 8022 0 8078 56 0 FreeSans 224 0 0 0 VALUE_top5
port 216 nsew signal output
flabel metal2 s 9402 0 9458 56 0 FreeSans 224 0 0 0 VALUE_top6
port 217 nsew signal output
flabel metal2 s 10782 0 10838 56 0 FreeSans 224 0 0 0 VALUE_top7
port 218 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 219 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 220 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal3 666 1428 666 1428 0 FrameData[0]
rlabel metal3 482 4148 482 4148 0 FrameData[10]
rlabel metal3 436 4420 436 4420 0 FrameData[11]
rlabel metal3 482 4692 482 4692 0 FrameData[12]
rlabel metal3 252 4964 252 4964 0 FrameData[13]
rlabel metal3 482 5236 482 5236 0 FrameData[14]
rlabel metal3 390 5508 390 5508 0 FrameData[15]
rlabel metal3 160 5780 160 5780 0 FrameData[16]
rlabel metal3 344 6052 344 6052 0 FrameData[17]
rlabel metal1 2024 6834 2024 6834 0 FrameData[18]
rlabel metal3 574 6596 574 6596 0 FrameData[19]
rlabel metal3 252 1700 252 1700 0 FrameData[1]
rlabel metal3 206 6868 206 6868 0 FrameData[20]
rlabel metal1 1288 6834 1288 6834 0 FrameData[21]
rlabel metal1 1104 6766 1104 6766 0 FrameData[22]
rlabel metal3 712 7684 712 7684 0 FrameData[23]
rlabel metal3 666 7956 666 7956 0 FrameData[24]
rlabel metal3 344 8228 344 8228 0 FrameData[25]
rlabel metal3 620 8500 620 8500 0 FrameData[26]
rlabel metal2 2898 8313 2898 8313 0 FrameData[27]
rlabel metal2 2806 8449 2806 8449 0 FrameData[28]
rlabel metal3 528 9316 528 9316 0 FrameData[29]
rlabel metal3 436 1972 436 1972 0 FrameData[2]
rlabel metal3 436 9588 436 9588 0 FrameData[30]
rlabel metal3 758 9860 758 9860 0 FrameData[31]
rlabel metal3 160 2244 160 2244 0 FrameData[3]
rlabel metal3 574 2516 574 2516 0 FrameData[4]
rlabel metal3 666 2788 666 2788 0 FrameData[5]
rlabel metal3 482 3060 482 3060 0 FrameData[6]
rlabel metal3 160 3332 160 3332 0 FrameData[7]
rlabel metal3 482 3604 482 3604 0 FrameData[8]
rlabel metal3 252 3876 252 3876 0 FrameData[9]
rlabel metal3 39798 1428 39798 1428 0 FrameData_O[0]
rlabel metal2 39422 3927 39422 3927 0 FrameData_O[10]
rlabel metal3 40442 4420 40442 4420 0 FrameData_O[11]
rlabel metal1 39468 3978 39468 3978 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal2 39422 5015 39422 5015 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal3 39798 5780 39798 5780 0 FrameData_O[16]
rlabel metal2 39422 5695 39422 5695 0 FrameData_O[17]
rlabel metal3 39982 6324 39982 6324 0 FrameData_O[18]
rlabel metal1 39514 5882 39514 5882 0 FrameData_O[19]
rlabel metal3 39614 1700 39614 1700 0 FrameData_O[1]
rlabel metal3 40212 6868 40212 6868 0 FrameData_O[20]
rlabel metal3 40166 7140 40166 7140 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 40166 7956 40166 7956 0 FrameData_O[24]
rlabel metal1 39284 7514 39284 7514 0 FrameData_O[25]
rlabel metal1 39606 6426 39606 6426 0 FrameData_O[26]
rlabel metal1 38686 7480 38686 7480 0 FrameData_O[27]
rlabel metal1 39422 6630 39422 6630 0 FrameData_O[28]
rlabel metal1 38410 7514 38410 7514 0 FrameData_O[29]
rlabel metal3 39430 1972 39430 1972 0 FrameData_O[2]
rlabel metal1 39330 8602 39330 8602 0 FrameData_O[30]
rlabel metal2 38686 8959 38686 8959 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 39706 2516 39706 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal2 39422 3383 39422 3383 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal1 17158 5202 17158 5202 0 FrameStrobe[0]
rlabel metal2 27370 327 27370 327 0 FrameStrobe[10]
rlabel metal2 34822 6528 34822 6528 0 FrameStrobe[11]
rlabel metal1 37214 6732 37214 6732 0 FrameStrobe[12]
rlabel metal1 31096 7378 31096 7378 0 FrameStrobe[13]
rlabel metal2 32890 1483 32890 1483 0 FrameStrobe[14]
rlabel metal1 34224 7378 34224 7378 0 FrameStrobe[15]
rlabel metal1 36892 5678 36892 5678 0 FrameStrobe[16]
rlabel metal2 37030 1401 37030 1401 0 FrameStrobe[17]
rlabel metal2 38410 667 38410 667 0 FrameStrobe[18]
rlabel metal2 39790 1401 39790 1401 0 FrameStrobe[19]
rlabel metal2 14950 1401 14950 1401 0 FrameStrobe[1]
rlabel via2 16330 55 16330 55 0 FrameStrobe[2]
rlabel metal2 17710 259 17710 259 0 FrameStrobe[3]
rlabel metal2 19090 1024 19090 1024 0 FrameStrobe[4]
rlabel metal2 20470 1007 20470 1007 0 FrameStrobe[5]
rlabel metal2 21850 123 21850 123 0 FrameStrobe[6]
rlabel metal2 23230 191 23230 191 0 FrameStrobe[7]
rlabel metal2 24610 939 24610 939 0 FrameStrobe[8]
rlabel metal2 25990 1194 25990 1194 0 FrameStrobe[9]
rlabel metal1 32660 8602 32660 8602 0 FrameStrobe_O[0]
rlabel metal2 36294 8704 36294 8704 0 FrameStrobe_O[10]
rlabel metal1 35650 8058 35650 8058 0 FrameStrobe_O[11]
rlabel metal1 36248 8602 36248 8602 0 FrameStrobe_O[12]
rlabel metal1 36248 8058 36248 8058 0 FrameStrobe_O[13]
rlabel metal1 37306 8262 37306 8262 0 FrameStrobe_O[14]
rlabel metal1 36800 8058 36800 8058 0 FrameStrobe_O[15]
rlabel metal1 37352 8602 37352 8602 0 FrameStrobe_O[16]
rlabel metal1 37674 8330 37674 8330 0 FrameStrobe_O[17]
rlabel metal1 38502 8602 38502 8602 0 FrameStrobe_O[18]
rlabel metal1 37904 8058 37904 8058 0 FrameStrobe_O[19]
rlabel metal1 33028 8602 33028 8602 0 FrameStrobe_O[1]
rlabel metal2 33534 8704 33534 8704 0 FrameStrobe_O[2]
rlabel metal1 33672 8330 33672 8330 0 FrameStrobe_O[3]
rlabel metal1 33948 8602 33948 8602 0 FrameStrobe_O[4]
rlabel metal1 34822 8568 34822 8568 0 FrameStrobe_O[5]
rlabel metal1 34684 8330 34684 8330 0 FrameStrobe_O[6]
rlabel metal1 34638 8058 34638 8058 0 FrameStrobe_O[7]
rlabel metal1 35282 8602 35282 8602 0 FrameStrobe_O[8]
rlabel metal1 36018 8364 36018 8364 0 FrameStrobe_O[9]
rlabel via1 19641 6222 19641 6222 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 19090 6698 19090 6698 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit1.Q
rlabel metal1 23000 3570 23000 3570 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit10.Q
rlabel metal1 23690 3570 23690 3570 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 9614 3162 9614 3162 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit12.Q
rlabel metal1 8648 2958 8648 2958 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit13.Q
rlabel metal1 26496 6834 26496 6834 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 26450 5542 26450 5542 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit15.Q
rlabel metal1 25162 6188 25162 6188 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 26266 6409 26266 6409 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 11546 3910 11546 3910 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit18.Q
rlabel metal1 11270 4250 11270 4250 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit19.Q
rlabel metal1 29026 3570 29026 3570 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit2.Q
rlabel metal1 22816 3910 22816 3910 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit20.Q
rlabel metal1 18814 3944 18814 3944 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 10396 6426 10396 6426 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 9890 6970 9890 6970 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit23.Q
rlabel via2 15226 6205 15226 6205 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 14674 6052 14674 6052 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit25.Q
rlabel metal1 7912 3638 7912 3638 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit26.Q
rlabel metal1 7590 3162 7590 3162 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 29394 3468 29394 3468 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit28.Q
rlabel metal1 28336 3162 28336 3162 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit29.Q
rlabel metal1 28244 3638 28244 3638 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 24518 7106 24518 7106 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 20516 7378 20516 7378 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 5014 4182 5014 4182 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 5106 4522 5106 4522 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit5.Q
rlabel metal1 14352 6426 14352 6426 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit6.Q
rlabel metal1 14628 6834 14628 6834 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 8786 6341 8786 6341 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit8.Q
rlabel metal1 7820 6222 7820 6222 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame0_bit9.Q
rlabel metal1 20332 5882 20332 5882 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit16.Q
rlabel metal1 20746 6834 20746 6834 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 21574 3383 21574 3383 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 18906 4522 18906 4522 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 14076 3128 14076 3128 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit20.Q
rlabel via2 15502 3995 15502 3995 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit21.Q
rlabel metal1 12926 6426 12926 6426 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit22.Q
rlabel metal1 14766 7208 14766 7208 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit23.Q
rlabel metal1 8878 6970 8878 6970 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit24.Q
rlabel metal1 9844 5882 9844 5882 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit25.Q
rlabel metal1 20585 3706 20585 3706 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 20930 3927 20930 3927 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit27.Q
rlabel metal1 11730 3570 11730 3570 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit28.Q
rlabel metal1 11914 3128 11914 3128 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 27646 6970 27646 6970 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit30.Q
rlabel metal1 27646 5814 27646 5814 0 Inst_S_EF_DAC8_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 20562 6460 20562 6460 0 Inst_S_EF_DAC8_switch_matrix.N2BEG0
rlabel metal1 29670 3502 29670 3502 0 Inst_S_EF_DAC8_switch_matrix.N2BEG1
rlabel metal1 6302 4114 6302 4114 0 Inst_S_EF_DAC8_switch_matrix.N2BEG2
rlabel metal1 16054 7412 16054 7412 0 Inst_S_EF_DAC8_switch_matrix.N2BEG3
rlabel metal1 9798 6324 9798 6324 0 Inst_S_EF_DAC8_switch_matrix.N2BEG4
rlabel metal2 24610 3978 24610 3978 0 Inst_S_EF_DAC8_switch_matrix.N2BEG5
rlabel metal1 12236 3502 12236 3502 0 Inst_S_EF_DAC8_switch_matrix.N2BEG6
rlabel metal2 28842 6596 28842 6596 0 Inst_S_EF_DAC8_switch_matrix.N2BEG7
rlabel metal1 20930 7820 20930 7820 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb0
rlabel metal1 29670 3706 29670 3706 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb1
rlabel metal1 5060 4114 5060 4114 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb2
rlabel metal1 14812 6630 14812 6630 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb3
rlabel metal1 7866 6086 7866 6086 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb4
rlabel metal2 24150 3910 24150 3910 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb5
rlabel metal1 9154 3162 9154 3162 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb6
rlabel metal1 28750 6732 28750 6732 0 Inst_S_EF_DAC8_switch_matrix.N2BEGb7
rlabel metal2 3450 8755 3450 8755 0 N1BEG[0]
rlabel metal1 3174 8602 3174 8602 0 N1BEG[1]
rlabel metal1 3450 8330 3450 8330 0 N1BEG[2]
rlabel metal1 4186 8058 4186 8058 0 N1BEG[3]
rlabel metal1 3680 8262 3680 8262 0 N2BEG[0]
rlabel metal1 4416 8602 4416 8602 0 N2BEG[1]
rlabel metal1 5014 8058 5014 8058 0 N2BEG[2]
rlabel metal1 4876 8262 4876 8262 0 N2BEG[3]
rlabel metal1 5198 8602 5198 8602 0 N2BEG[4]
rlabel metal1 5658 8602 5658 8602 0 N2BEG[5]
rlabel metal1 6118 8058 6118 8058 0 N2BEG[6]
rlabel metal1 6210 8602 6210 8602 0 N2BEG[7]
rlabel metal1 6670 8058 6670 8058 0 N2BEGb[0]
rlabel metal1 6716 8602 6716 8602 0 N2BEGb[1]
rlabel metal1 7268 8058 7268 8058 0 N2BEGb[2]
rlabel metal1 7176 8330 7176 8330 0 N2BEGb[3]
rlabel metal1 7452 8602 7452 8602 0 N2BEGb[4]
rlabel metal1 7820 8602 7820 8602 0 N2BEGb[5]
rlabel metal1 8372 8058 8372 8058 0 N2BEGb[6]
rlabel metal1 8280 8602 8280 8602 0 N2BEGb[7]
rlabel metal1 8924 8058 8924 8058 0 N4BEG[0]
rlabel metal1 11408 8602 11408 8602 0 N4BEG[10]
rlabel metal1 11914 8058 11914 8058 0 N4BEG[11]
rlabel metal1 12052 8602 12052 8602 0 N4BEG[12]
rlabel metal1 12328 8602 12328 8602 0 N4BEG[13]
rlabel metal1 12788 8058 12788 8058 0 N4BEG[14]
rlabel metal1 12788 8602 12788 8602 0 N4BEG[15]
rlabel metal1 8786 8602 8786 8602 0 N4BEG[1]
rlabel metal1 9522 8058 9522 8058 0 N4BEG[2]
rlabel metal1 9522 8602 9522 8602 0 N4BEG[3]
rlabel metal1 9798 8602 9798 8602 0 N4BEG[4]
rlabel metal1 10120 8058 10120 8058 0 N4BEG[5]
rlabel metal1 10534 8058 10534 8058 0 N4BEG[6]
rlabel metal1 10580 8602 10580 8602 0 N4BEG[7]
rlabel metal1 10902 8602 10902 8602 0 N4BEG[8]
rlabel metal1 11362 8058 11362 8058 0 N4BEG[9]
rlabel metal1 13110 8602 13110 8602 0 NN4BEG[0]
rlabel metal1 16100 8058 16100 8058 0 NN4BEG[10]
rlabel metal1 16146 8602 16146 8602 0 NN4BEG[11]
rlabel metal1 16468 8602 16468 8602 0 NN4BEG[12]
rlabel metal1 16882 8602 16882 8602 0 NN4BEG[13]
rlabel metal1 17940 8602 17940 8602 0 NN4BEG[14]
rlabel metal1 17434 8602 17434 8602 0 NN4BEG[15]
rlabel metal1 13570 8058 13570 8058 0 NN4BEG[1]
rlabel metal1 13616 8602 13616 8602 0 NN4BEG[2]
rlabel metal1 13892 8330 13892 8330 0 NN4BEG[3]
rlabel metal1 14444 8058 14444 8058 0 NN4BEG[4]
rlabel metal1 14536 8602 14536 8602 0 NN4BEG[5]
rlabel metal1 14996 8058 14996 8058 0 NN4BEG[6]
rlabel metal1 14904 8602 14904 8602 0 NN4BEG[7]
rlabel metal1 15318 8602 15318 8602 0 NN4BEG[8]
rlabel metal1 15640 8602 15640 8602 0 NN4BEG[9]
rlabel metal2 17894 10397 17894 10397 0 S1END[0]
rlabel metal2 18170 10397 18170 10397 0 S1END[1]
rlabel metal2 18446 9836 18446 9836 0 S1END[2]
rlabel metal2 18722 9836 18722 9836 0 S1END[3]
rlabel metal2 21206 10533 21206 10533 0 S2END[0]
rlabel metal2 21482 9836 21482 9836 0 S2END[1]
rlabel metal2 21758 9870 21758 9870 0 S2END[2]
rlabel metal2 22034 9904 22034 9904 0 S2END[3]
rlabel metal2 22310 9870 22310 9870 0 S2END[4]
rlabel metal2 22586 9904 22586 9904 0 S2END[5]
rlabel metal2 22862 9870 22862 9870 0 S2END[6]
rlabel metal2 23138 9904 23138 9904 0 S2END[7]
rlabel metal2 18998 9836 18998 9836 0 S2MID[0]
rlabel metal1 19435 8466 19435 8466 0 S2MID[1]
rlabel metal2 19550 10805 19550 10805 0 S2MID[2]
rlabel metal2 19826 9836 19826 9836 0 S2MID[3]
rlabel metal2 20102 10533 20102 10533 0 S2MID[4]
rlabel metal2 20378 10533 20378 10533 0 S2MID[5]
rlabel metal2 20654 9904 20654 9904 0 S2MID[6]
rlabel metal2 20930 9836 20930 9836 0 S2MID[7]
rlabel metal2 23414 9870 23414 9870 0 S4END[0]
rlabel metal1 37582 6766 37582 6766 0 S4END[10]
rlabel metal2 34730 7820 34730 7820 0 S4END[11]
rlabel metal2 36018 8670 36018 8670 0 S4END[12]
rlabel metal2 37398 9911 37398 9911 0 S4END[13]
rlabel metal2 37582 8908 37582 8908 0 S4END[14]
rlabel metal1 38640 6630 38640 6630 0 S4END[15]
rlabel metal2 23690 9904 23690 9904 0 S4END[1]
rlabel metal2 23966 9836 23966 9836 0 S4END[2]
rlabel metal2 24242 9530 24242 9530 0 S4END[3]
rlabel metal2 24518 9462 24518 9462 0 S4END[4]
rlabel metal2 24794 9836 24794 9836 0 S4END[5]
rlabel metal2 25070 9530 25070 9530 0 S4END[6]
rlabel metal2 25346 10533 25346 10533 0 S4END[7]
rlabel metal1 38410 5712 38410 5712 0 S4END[8]
rlabel metal2 34638 8874 34638 8874 0 S4END[9]
rlabel metal2 27830 9836 27830 9836 0 SS4END[0]
rlabel metal2 30590 9530 30590 9530 0 SS4END[10]
rlabel metal2 30866 9598 30866 9598 0 SS4END[11]
rlabel metal2 31142 9836 31142 9836 0 SS4END[12]
rlabel metal2 31418 9870 31418 9870 0 SS4END[13]
rlabel metal2 31694 9530 31694 9530 0 SS4END[14]
rlabel metal2 31970 10397 31970 10397 0 SS4END[15]
rlabel metal2 28106 9836 28106 9836 0 SS4END[1]
rlabel metal2 28382 9530 28382 9530 0 SS4END[2]
rlabel metal2 28658 9836 28658 9836 0 SS4END[3]
rlabel metal2 28934 9530 28934 9530 0 SS4END[4]
rlabel metal2 29210 9870 29210 9870 0 SS4END[5]
rlabel metal2 29486 9530 29486 9530 0 SS4END[6]
rlabel metal2 29762 9530 29762 9530 0 SS4END[7]
rlabel metal2 30038 10397 30038 10397 0 SS4END[8]
rlabel metal2 30314 9836 30314 9836 0 SS4END[9]
rlabel metal2 12190 55 12190 55 0 UserCLK
rlabel metal1 32384 8058 32384 8058 0 UserCLKo
rlabel metal2 1150 1296 1150 1296 0 VALUE_top0
rlabel metal2 2530 599 2530 599 0 VALUE_top1
rlabel metal2 3910 1160 3910 1160 0 VALUE_top2
rlabel metal2 5290 1160 5290 1160 0 VALUE_top3
rlabel metal2 6670 1160 6670 1160 0 VALUE_top4
rlabel metal2 8050 1160 8050 1160 0 VALUE_top5
rlabel metal2 9430 1160 9430 1160 0 VALUE_top6
rlabel metal2 10810 1160 10810 1160 0 VALUE_top7
rlabel metal1 4715 2618 4715 2618 0 net1
rlabel metal2 6670 5848 6670 5848 0 net10
rlabel metal4 37260 8500 37260 8500 0 net100
rlabel metal1 15548 3638 15548 3638 0 net101
rlabel metal2 15410 2873 15410 2873 0 net102
rlabel metal2 38778 5729 38778 5729 0 net103
rlabel metal2 38134 7327 38134 7327 0 net104
rlabel metal1 37168 2414 37168 2414 0 net105
rlabel metal2 38870 8704 38870 8704 0 net106
rlabel metal2 38318 7038 38318 7038 0 net107
rlabel metal1 36018 2482 36018 2482 0 net108
rlabel metal3 20976 1700 20976 1700 0 net109
rlabel metal1 2254 6630 2254 6630 0 net11
rlabel metal1 21528 1326 21528 1326 0 net110
rlabel metal1 39238 2516 39238 2516 0 net111
rlabel metal1 26358 1190 26358 1190 0 net112
rlabel metal3 22724 1564 22724 1564 0 net113
rlabel metal2 40066 6477 40066 6477 0 net114
rlabel metal1 32614 8432 32614 8432 0 net115
rlabel metal1 37904 3706 37904 3706 0 net116
rlabel metal1 35926 7888 35926 7888 0 net117
rlabel metal2 37030 7684 37030 7684 0 net118
rlabel metal2 36202 7650 36202 7650 0 net119
rlabel metal2 17802 5899 17802 5899 0 net12
rlabel metal2 34546 7990 34546 7990 0 net120
rlabel metal1 35558 7514 35558 7514 0 net121
rlabel metal1 37904 5882 37904 5882 0 net122
rlabel metal1 38272 8058 38272 8058 0 net123
rlabel metal1 36570 7276 36570 7276 0 net124
rlabel metal1 37076 7514 37076 7514 0 net125
rlabel metal2 18814 4777 18814 4777 0 net126
rlabel metal1 32936 3706 32936 3706 0 net127
rlabel metal1 33488 3706 33488 3706 0 net128
rlabel metal1 33948 3706 33948 3706 0 net129
rlabel metal1 8280 5746 8280 5746 0 net13
rlabel metal1 36294 3366 36294 3366 0 net130
rlabel metal1 36984 3706 36984 3706 0 net131
rlabel metal1 38410 3400 38410 3400 0 net132
rlabel metal1 34776 3366 34776 3366 0 net133
rlabel metal1 35098 3706 35098 3706 0 net134
rlabel metal2 21850 7514 21850 7514 0 net135
rlabel metal2 2622 8415 2622 8415 0 net136
rlabel metal1 7912 3162 7912 3162 0 net137
rlabel metal2 16054 6885 16054 6885 0 net138
rlabel metal2 9706 9078 9706 9078 0 net139
rlabel metal1 22402 6732 22402 6732 0 net14
rlabel metal2 4554 8738 4554 8738 0 net140
rlabel metal2 6026 5916 6026 5916 0 net141
rlabel metal1 15824 7514 15824 7514 0 net142
rlabel metal1 9154 6086 9154 6086 0 net143
rlabel metal1 5428 8466 5428 8466 0 net144
rlabel metal2 12190 3757 12190 3757 0 net145
rlabel metal2 5842 9027 5842 9027 0 net146
rlabel metal2 20746 7769 20746 7769 0 net147
rlabel metal2 6762 9214 6762 9214 0 net148
rlabel metal1 5658 3978 5658 3978 0 net149
rlabel metal2 23138 6987 23138 6987 0 net15
rlabel metal2 7314 8840 7314 8840 0 net150
rlabel metal1 9154 6630 9154 6630 0 net151
rlabel metal2 7866 9282 7866 9282 0 net152
rlabel metal1 9752 3706 9752 3706 0 net153
rlabel metal2 8142 9248 8142 9248 0 net154
rlabel via2 38410 6851 38410 6851 0 net155
rlabel metal1 5842 5338 5842 5338 0 net156
rlabel metal1 12190 7820 12190 7820 0 net157
rlabel metal1 8050 7242 8050 7242 0 net158
rlabel metal2 12742 8976 12742 8976 0 net159
rlabel metal1 6946 4726 6946 4726 0 net16
rlabel metal1 12581 7854 12581 7854 0 net160
rlabel metal2 14766 9265 14766 9265 0 net161
rlabel metal1 37214 6834 37214 6834 0 net162
rlabel metal1 37352 6426 37352 6426 0 net163
rlabel metal1 36018 6358 36018 6358 0 net164
rlabel metal1 36570 7174 36570 7174 0 net165
rlabel via2 38042 6851 38042 6851 0 net166
rlabel metal1 36754 6868 36754 6868 0 net167
rlabel metal2 21666 7633 21666 7633 0 net168
rlabel metal1 19458 7752 19458 7752 0 net169
rlabel metal1 29210 4590 29210 4590 0 net17
rlabel metal2 13570 6630 13570 6630 0 net170
rlabel metal1 17986 7514 17986 7514 0 net171
rlabel metal2 13754 6698 13754 6698 0 net172
rlabel metal1 15686 8058 15686 8058 0 net173
rlabel metal1 14122 6290 14122 6290 0 net174
rlabel metal2 20378 3961 20378 3961 0 net175
rlabel metal2 9614 3791 9614 3791 0 net176
rlabel metal2 20378 8279 20378 8279 0 net177
rlabel metal1 14444 2618 14444 2618 0 net178
rlabel metal2 13110 6732 13110 6732 0 net179
rlabel metal1 20654 5338 20654 5338 0 net18
rlabel metal1 15548 7242 15548 7242 0 net180
rlabel metal2 7958 7752 7958 7752 0 net181
rlabel metal2 23230 6528 23230 6528 0 net182
rlabel metal2 13662 7446 13662 7446 0 net183
rlabel metal2 19182 5627 19182 5627 0 net184
rlabel metal1 19458 8058 19458 8058 0 net185
rlabel metal2 18814 8874 18814 8874 0 net186
rlabel metal1 37122 3162 37122 3162 0 net187
rlabel metal2 3266 2465 3266 2465 0 net188
rlabel metal2 2898 2244 2898 2244 0 net189
rlabel metal1 16008 3502 16008 3502 0 net19
rlabel metal1 4278 2448 4278 2448 0 net190
rlabel metal1 6279 2414 6279 2414 0 net191
rlabel metal2 7038 2516 7038 2516 0 net192
rlabel metal1 7820 2414 7820 2414 0 net193
rlabel metal2 9798 2074 9798 2074 0 net194
rlabel metal2 19550 2533 19550 2533 0 net195
rlabel metal1 17664 8058 17664 8058 0 net196
rlabel metal1 22310 2346 22310 2346 0 net2
rlabel metal1 1840 6630 1840 6630 0 net20
rlabel metal2 1610 6086 1610 6086 0 net21
rlabel metal1 12535 7378 12535 7378 0 net22
rlabel metal1 11270 6664 11270 6664 0 net23
rlabel metal1 9062 5678 9062 5678 0 net24
rlabel metal2 15364 3434 15364 3434 0 net25
rlabel metal1 18354 3060 18354 3060 0 net26
rlabel metal2 14858 3825 14858 3825 0 net27
rlabel metal2 17434 2907 17434 2907 0 net28
rlabel metal2 2530 2108 2530 2108 0 net29
rlabel metal2 1610 2788 1610 2788 0 net3
rlabel metal1 2231 8398 2231 8398 0 net30
rlabel metal2 1702 7905 1702 7905 0 net31
rlabel metal2 1702 2176 1702 2176 0 net32
rlabel metal2 3818 3944 3818 3944 0 net33
rlabel metal2 4370 3638 4370 3638 0 net34
rlabel metal1 12834 6290 12834 6290 0 net35
rlabel metal1 2024 3638 2024 3638 0 net36
rlabel metal1 5704 6766 5704 6766 0 net37
rlabel metal1 4600 6698 4600 6698 0 net38
rlabel metal1 17112 6766 17112 6766 0 net39
rlabel metal1 5106 3502 5106 3502 0 net4
rlabel metal1 8464 3502 8464 3502 0 net40
rlabel metal2 18538 8772 18538 8772 0 net41
rlabel metal1 21436 7310 21436 7310 0 net42
rlabel metal2 21482 6324 21482 6324 0 net43
rlabel metal1 14950 3468 14950 3468 0 net44
rlabel metal1 22540 3570 22540 3570 0 net45
rlabel metal1 17250 5848 17250 5848 0 net46
rlabel metal1 20470 5644 20470 5644 0 net47
rlabel via2 12190 4675 12190 4675 0 net48
rlabel metal2 22862 3825 22862 3825 0 net49
rlabel metal1 5474 4182 5474 4182 0 net5
rlabel metal1 18630 6154 18630 6154 0 net50
rlabel metal2 19182 7514 19182 7514 0 net51
rlabel metal2 19366 5593 19366 5593 0 net52
rlabel metal2 21850 5355 21850 5355 0 net53
rlabel metal2 19918 8840 19918 8840 0 net54
rlabel metal1 15732 7310 15732 7310 0 net55
rlabel metal3 15180 3672 15180 3672 0 net56
rlabel metal1 27646 4012 27646 4012 0 net57
rlabel metal1 21022 6834 21022 6834 0 net58
rlabel metal1 25760 6834 25760 6834 0 net59
rlabel metal1 2254 5882 2254 5882 0 net6
rlabel metal1 10879 4658 10879 4658 0 net60
rlabel metal1 21712 4658 21712 4658 0 net61
rlabel metal2 17250 8126 17250 8126 0 net62
rlabel metal2 20010 7582 20010 7582 0 net63
rlabel metal2 20378 5032 20378 5032 0 net64
rlabel metal1 29394 4182 29394 4182 0 net65
rlabel metal1 21298 7344 21298 7344 0 net66
rlabel metal1 27888 6222 27888 6222 0 net67
rlabel metal2 30038 6120 30038 6120 0 net68
rlabel metal3 14812 7480 14812 7480 0 net69
rlabel metal2 1886 5831 1886 5831 0 net7
rlabel metal2 32154 8942 32154 8942 0 net70
rlabel metal1 15318 2856 15318 2856 0 net71
rlabel metal2 30774 5440 30774 5440 0 net72
rlabel metal2 29118 8160 29118 8160 0 net73
rlabel metal1 9371 2958 9371 2958 0 net74
rlabel metal2 23138 4726 23138 4726 0 net75
rlabel metal1 10258 6834 10258 6834 0 net76
rlabel metal1 19550 7854 19550 7854 0 net77
rlabel metal2 17250 9384 17250 9384 0 net78
rlabel metal1 29808 4114 29808 4114 0 net79
rlabel metal2 6854 5729 6854 5729 0 net8
rlabel metal1 18814 6188 18814 6188 0 net80
rlabel metal2 28198 7378 28198 7378 0 net81
rlabel metal1 21390 4182 21390 4182 0 net82
rlabel metal1 18446 6154 18446 6154 0 net83
rlabel metal2 21666 3264 21666 3264 0 net84
rlabel metal2 37490 3842 37490 3842 0 net85
rlabel metal2 39238 3791 39238 3791 0 net86
rlabel via2 13754 2941 13754 2941 0 net87
rlabel metal2 38962 4930 38962 4930 0 net88
rlabel metal1 38870 5746 38870 5746 0 net89
rlabel via2 1702 6307 1702 6307 0 net9
rlabel metal2 20562 5593 20562 5593 0 net90
rlabel metal2 37306 4641 37306 4641 0 net91
rlabel via2 15870 2941 15870 2941 0 net92
rlabel metal2 15318 3791 15318 3791 0 net93
rlabel metal1 18354 5814 18354 5814 0 net94
rlabel metal2 17986 3417 17986 3417 0 net95
rlabel via2 16882 4539 16882 4539 0 net96
rlabel metal3 14628 7344 14628 7344 0 net97
rlabel metal2 38686 7259 38686 7259 0 net98
rlabel metal2 39238 8415 39238 8415 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
