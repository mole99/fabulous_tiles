module RegFile (UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire AD0;
 wire AD1;
 wire AD2;
 wire AD3;
 wire A_ADR0;
 wire BD0;
 wire BD1;
 wire BD2;
 wire BD3;
 wire B_ADR0;
 wire net739;
 wire net736;
 wire net729;
 wire net531;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net724;
 wire net525;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net722;
 wire net737;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire \Inst_RegFile_32x4.AD_comb[0] ;
 wire \Inst_RegFile_32x4.AD_comb[1] ;
 wire \Inst_RegFile_32x4.AD_comb[2] ;
 wire \Inst_RegFile_32x4.AD_comb[3] ;
 wire \Inst_RegFile_32x4.AD_reg[0] ;
 wire \Inst_RegFile_32x4.AD_reg[1] ;
 wire \Inst_RegFile_32x4.AD_reg[2] ;
 wire \Inst_RegFile_32x4.AD_reg[3] ;
 wire \Inst_RegFile_32x4.BD_comb[0] ;
 wire \Inst_RegFile_32x4.BD_comb[1] ;
 wire \Inst_RegFile_32x4.BD_comb[2] ;
 wire \Inst_RegFile_32x4.BD_comb[3] ;
 wire \Inst_RegFile_32x4.BD_reg[0] ;
 wire \Inst_RegFile_32x4.BD_reg[1] ;
 wire \Inst_RegFile_32x4.BD_reg[2] ;
 wire \Inst_RegFile_32x4.BD_reg[3] ;
 wire \Inst_RegFile_32x4.mem[0][0] ;
 wire \Inst_RegFile_32x4.mem[0][1] ;
 wire \Inst_RegFile_32x4.mem[0][2] ;
 wire \Inst_RegFile_32x4.mem[0][3] ;
 wire \Inst_RegFile_32x4.mem[10][0] ;
 wire \Inst_RegFile_32x4.mem[10][1] ;
 wire \Inst_RegFile_32x4.mem[10][2] ;
 wire \Inst_RegFile_32x4.mem[10][3] ;
 wire \Inst_RegFile_32x4.mem[11][0] ;
 wire \Inst_RegFile_32x4.mem[11][1] ;
 wire \Inst_RegFile_32x4.mem[11][2] ;
 wire \Inst_RegFile_32x4.mem[11][3] ;
 wire \Inst_RegFile_32x4.mem[12][0] ;
 wire \Inst_RegFile_32x4.mem[12][1] ;
 wire \Inst_RegFile_32x4.mem[12][2] ;
 wire \Inst_RegFile_32x4.mem[12][3] ;
 wire \Inst_RegFile_32x4.mem[13][0] ;
 wire \Inst_RegFile_32x4.mem[13][1] ;
 wire \Inst_RegFile_32x4.mem[13][2] ;
 wire \Inst_RegFile_32x4.mem[13][3] ;
 wire \Inst_RegFile_32x4.mem[14][0] ;
 wire \Inst_RegFile_32x4.mem[14][1] ;
 wire \Inst_RegFile_32x4.mem[14][2] ;
 wire \Inst_RegFile_32x4.mem[14][3] ;
 wire \Inst_RegFile_32x4.mem[15][0] ;
 wire \Inst_RegFile_32x4.mem[15][1] ;
 wire \Inst_RegFile_32x4.mem[15][2] ;
 wire \Inst_RegFile_32x4.mem[15][3] ;
 wire \Inst_RegFile_32x4.mem[16][0] ;
 wire \Inst_RegFile_32x4.mem[16][1] ;
 wire \Inst_RegFile_32x4.mem[16][2] ;
 wire \Inst_RegFile_32x4.mem[16][3] ;
 wire \Inst_RegFile_32x4.mem[17][0] ;
 wire \Inst_RegFile_32x4.mem[17][1] ;
 wire \Inst_RegFile_32x4.mem[17][2] ;
 wire \Inst_RegFile_32x4.mem[17][3] ;
 wire \Inst_RegFile_32x4.mem[18][0] ;
 wire \Inst_RegFile_32x4.mem[18][1] ;
 wire \Inst_RegFile_32x4.mem[18][2] ;
 wire \Inst_RegFile_32x4.mem[18][3] ;
 wire \Inst_RegFile_32x4.mem[19][0] ;
 wire \Inst_RegFile_32x4.mem[19][1] ;
 wire \Inst_RegFile_32x4.mem[19][2] ;
 wire \Inst_RegFile_32x4.mem[19][3] ;
 wire \Inst_RegFile_32x4.mem[1][0] ;
 wire \Inst_RegFile_32x4.mem[1][1] ;
 wire \Inst_RegFile_32x4.mem[1][2] ;
 wire \Inst_RegFile_32x4.mem[1][3] ;
 wire \Inst_RegFile_32x4.mem[20][0] ;
 wire \Inst_RegFile_32x4.mem[20][1] ;
 wire \Inst_RegFile_32x4.mem[20][2] ;
 wire \Inst_RegFile_32x4.mem[20][3] ;
 wire \Inst_RegFile_32x4.mem[21][0] ;
 wire \Inst_RegFile_32x4.mem[21][1] ;
 wire \Inst_RegFile_32x4.mem[21][2] ;
 wire \Inst_RegFile_32x4.mem[21][3] ;
 wire \Inst_RegFile_32x4.mem[22][0] ;
 wire \Inst_RegFile_32x4.mem[22][1] ;
 wire \Inst_RegFile_32x4.mem[22][2] ;
 wire \Inst_RegFile_32x4.mem[22][3] ;
 wire \Inst_RegFile_32x4.mem[23][0] ;
 wire \Inst_RegFile_32x4.mem[23][1] ;
 wire \Inst_RegFile_32x4.mem[23][2] ;
 wire \Inst_RegFile_32x4.mem[23][3] ;
 wire \Inst_RegFile_32x4.mem[24][0] ;
 wire \Inst_RegFile_32x4.mem[24][1] ;
 wire \Inst_RegFile_32x4.mem[24][2] ;
 wire \Inst_RegFile_32x4.mem[24][3] ;
 wire \Inst_RegFile_32x4.mem[25][0] ;
 wire \Inst_RegFile_32x4.mem[25][1] ;
 wire \Inst_RegFile_32x4.mem[25][2] ;
 wire \Inst_RegFile_32x4.mem[25][3] ;
 wire \Inst_RegFile_32x4.mem[26][0] ;
 wire \Inst_RegFile_32x4.mem[26][1] ;
 wire \Inst_RegFile_32x4.mem[26][2] ;
 wire \Inst_RegFile_32x4.mem[26][3] ;
 wire \Inst_RegFile_32x4.mem[27][0] ;
 wire \Inst_RegFile_32x4.mem[27][1] ;
 wire \Inst_RegFile_32x4.mem[27][2] ;
 wire \Inst_RegFile_32x4.mem[27][3] ;
 wire \Inst_RegFile_32x4.mem[28][0] ;
 wire \Inst_RegFile_32x4.mem[28][1] ;
 wire \Inst_RegFile_32x4.mem[28][2] ;
 wire \Inst_RegFile_32x4.mem[28][3] ;
 wire \Inst_RegFile_32x4.mem[29][0] ;
 wire \Inst_RegFile_32x4.mem[29][1] ;
 wire \Inst_RegFile_32x4.mem[29][2] ;
 wire \Inst_RegFile_32x4.mem[29][3] ;
 wire \Inst_RegFile_32x4.mem[2][0] ;
 wire \Inst_RegFile_32x4.mem[2][1] ;
 wire \Inst_RegFile_32x4.mem[2][2] ;
 wire \Inst_RegFile_32x4.mem[2][3] ;
 wire \Inst_RegFile_32x4.mem[30][0] ;
 wire \Inst_RegFile_32x4.mem[30][1] ;
 wire \Inst_RegFile_32x4.mem[30][2] ;
 wire \Inst_RegFile_32x4.mem[30][3] ;
 wire \Inst_RegFile_32x4.mem[31][0] ;
 wire \Inst_RegFile_32x4.mem[31][1] ;
 wire \Inst_RegFile_32x4.mem[31][2] ;
 wire \Inst_RegFile_32x4.mem[31][3] ;
 wire \Inst_RegFile_32x4.mem[3][0] ;
 wire \Inst_RegFile_32x4.mem[3][1] ;
 wire \Inst_RegFile_32x4.mem[3][2] ;
 wire \Inst_RegFile_32x4.mem[3][3] ;
 wire \Inst_RegFile_32x4.mem[4][0] ;
 wire \Inst_RegFile_32x4.mem[4][1] ;
 wire \Inst_RegFile_32x4.mem[4][2] ;
 wire \Inst_RegFile_32x4.mem[4][3] ;
 wire \Inst_RegFile_32x4.mem[5][0] ;
 wire \Inst_RegFile_32x4.mem[5][1] ;
 wire \Inst_RegFile_32x4.mem[5][2] ;
 wire \Inst_RegFile_32x4.mem[5][3] ;
 wire \Inst_RegFile_32x4.mem[6][0] ;
 wire \Inst_RegFile_32x4.mem[6][1] ;
 wire \Inst_RegFile_32x4.mem[6][2] ;
 wire \Inst_RegFile_32x4.mem[6][3] ;
 wire \Inst_RegFile_32x4.mem[7][0] ;
 wire \Inst_RegFile_32x4.mem[7][1] ;
 wire \Inst_RegFile_32x4.mem[7][2] ;
 wire \Inst_RegFile_32x4.mem[7][3] ;
 wire \Inst_RegFile_32x4.mem[8][0] ;
 wire \Inst_RegFile_32x4.mem[8][1] ;
 wire \Inst_RegFile_32x4.mem[8][2] ;
 wire \Inst_RegFile_32x4.mem[8][3] ;
 wire \Inst_RegFile_32x4.mem[9][0] ;
 wire \Inst_RegFile_32x4.mem[9][1] ;
 wire \Inst_RegFile_32x4.mem[9][2] ;
 wire \Inst_RegFile_32x4.mem[9][3] ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_RegFile_switch_matrix.E1BEG0 ;
 wire \Inst_RegFile_switch_matrix.E1BEG1 ;
 wire \Inst_RegFile_switch_matrix.E1BEG2 ;
 wire \Inst_RegFile_switch_matrix.E1BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG0 ;
 wire \Inst_RegFile_switch_matrix.E2BEG1 ;
 wire \Inst_RegFile_switch_matrix.E2BEG2 ;
 wire \Inst_RegFile_switch_matrix.E2BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG4 ;
 wire \Inst_RegFile_switch_matrix.E2BEG5 ;
 wire \Inst_RegFile_switch_matrix.E2BEG6 ;
 wire \Inst_RegFile_switch_matrix.E2BEG7 ;
 wire \Inst_RegFile_switch_matrix.E6BEG0 ;
 wire \Inst_RegFile_switch_matrix.E6BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG0 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG2 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG7 ;
 wire \Inst_RegFile_switch_matrix.N1BEG0 ;
 wire \Inst_RegFile_switch_matrix.N1BEG1 ;
 wire \Inst_RegFile_switch_matrix.N1BEG2 ;
 wire \Inst_RegFile_switch_matrix.N1BEG3 ;
 wire \Inst_RegFile_switch_matrix.N4BEG0 ;
 wire \Inst_RegFile_switch_matrix.N4BEG1 ;
 wire \Inst_RegFile_switch_matrix.N4BEG2 ;
 wire \Inst_RegFile_switch_matrix.N4BEG3 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG0 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG1 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG2 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG3 ;
 wire \Inst_RegFile_switch_matrix.S1BEG0 ;
 wire \Inst_RegFile_switch_matrix.S1BEG1 ;
 wire \Inst_RegFile_switch_matrix.S1BEG2 ;
 wire \Inst_RegFile_switch_matrix.S1BEG3 ;
 wire \Inst_RegFile_switch_matrix.S4BEG0 ;
 wire \Inst_RegFile_switch_matrix.S4BEG1 ;
 wire \Inst_RegFile_switch_matrix.S4BEG2 ;
 wire \Inst_RegFile_switch_matrix.S4BEG3 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG0 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG1 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG2 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG3 ;
 wire \Inst_RegFile_switch_matrix.W1BEG0 ;
 wire \Inst_RegFile_switch_matrix.W1BEG1 ;
 wire \Inst_RegFile_switch_matrix.W1BEG2 ;
 wire \Inst_RegFile_switch_matrix.W1BEG3 ;
 wire \Inst_RegFile_switch_matrix.W6BEG0 ;
 wire \Inst_RegFile_switch_matrix.W6BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG0 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG2 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG3 ;
 wire net210;
 wire net742;
 wire net734;
 wire net526;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net723;
 wire net728;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net725;
 wire net732;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net741;
 wire net727;
 wire net731;
 wire net527;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net726;
 wire net738;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net740;
 wire net735;
 wire net730;
 wire net528;
 wire net319;
 wire net320;
 wire net321;
 wire net721;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net529;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net733;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net530;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net511;
 wire net965;
 wire net966;
 wire net967;
 wire net503;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net505;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net518;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net504;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net516;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net363;
 wire net500;
 wire net501;
 wire net502;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net517;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net532;
 wire net533;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net563;
 wire net717;
 wire net718;
 wire net719;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;

 sg13g2_inv_1 _1510_ (.Y(_1132_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_inv_1 _1511_ (.Y(_1133_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_inv_1 _1512_ (.Y(_1134_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_inv_1 _1513_ (.Y(_1135_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_inv_1 _1514_ (.Y(_1136_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_inv_1 _1515_ (.Y(_1137_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_inv_1 _1516_ (.Y(_1138_),
    .A(net107));
 sg13g2_inv_1 _1517_ (.Y(_1139_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_inv_1 _1518_ (.Y(_1140_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_inv_1 _1519_ (.Y(_1141_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_inv_1 _1520_ (.Y(_1142_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_inv_1 _1521_ (.Y(_1143_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_inv_1 _1522_ (.Y(_1144_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_inv_1 _1523_ (.Y(_1145_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_inv_1 _1524_ (.Y(_1146_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_inv_1 _1525_ (.Y(_1147_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_inv_1 _1526_ (.Y(_1148_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_inv_1 _1527_ (.Y(_1149_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_inv_1 _1528_ (.Y(_1150_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_inv_1 _1529_ (.Y(_1151_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_inv_1 _1530_ (.Y(_1152_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_inv_1 _1531_ (.Y(_1153_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ));
 sg13g2_inv_1 _1532_ (.Y(_1154_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ));
 sg13g2_inv_1 _1533_ (.Y(_1155_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ));
 sg13g2_inv_1 _1534_ (.Y(_1156_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_inv_1 _1535_ (.Y(_1157_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ));
 sg13g2_inv_1 _1536_ (.Y(_1158_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ));
 sg13g2_inv_1 _1537_ (.Y(_1159_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ));
 sg13g2_inv_1 _1538_ (.Y(_1160_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ));
 sg13g2_inv_1 _1539_ (.Y(_1161_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_inv_1 _1540_ (.Y(_1162_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_inv_1 _1541_ (.Y(_1163_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_inv_16 _1542_ (.A(net1015),
    .Y(_1164_));
 sg13g2_inv_2 _1543_ (.Y(_1165_),
    .A(net1003));
 sg13g2_inv_1 _1544_ (.Y(_1166_),
    .A(net1017));
 sg13g2_inv_2 _1545_ (.Y(_1167_),
    .A(net978));
 sg13g2_o21ai_1 _1546_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_1168_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(net988));
 sg13g2_a21oi_1 _1547_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(_1165_),
    .Y(_1169_),
    .B1(_1168_));
 sg13g2_nand2_1 _1548_ (.Y(_1170_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .B(net1033));
 sg13g2_nand2b_1 _1549_ (.Y(_1171_),
    .B(net974),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_a21oi_2 _1550_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .Y(_1172_),
    .A2(_1170_),
    .A1(_1171_));
 sg13g2_nor3_2 _1551_ (.A(_1172_),
    .B(_1169_),
    .C(_1141_),
    .Y(_1173_));
 sg13g2_mux4_1 _1552_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net88),
    .A1(net1019),
    .A2(AD1),
    .A3(net967),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1174_));
 sg13g2_o21ai_1 _1553_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .Y(_1175_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_1174_));
 sg13g2_mux4_1 _1554_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net23),
    .A1(net58),
    .A2(net60),
    .A3(net68),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1176_));
 sg13g2_mux4_1 _1555_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(net32),
    .A1(net40),
    .A2(net3),
    .A3(net11),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_1177_));
 sg13g2_mux2_1 _1556_ (.A0(_1176_),
    .A1(_1177_),
    .S(_1141_),
    .X(_1178_));
 sg13g2_nand2b_1 _1557_ (.Y(_1179_),
    .B(_1178_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_o21ai_1 _1558_ (.B1(_1179_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .A1(_1175_),
    .A2(_1173_));
 sg13g2_mux4_1 _1559_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ),
    .A0(net44),
    .A1(net72),
    .A2(net15),
    .A3(net723),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_1180_));
 sg13g2_or2_1 _1560_ (.X(_1181_),
    .B(_1180_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_mux4_1 _1561_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(net45),
    .A1(net16),
    .A2(net73),
    .A3(net100),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_1182_));
 sg13g2_inv_1 _1562_ (.Y(_1183_),
    .A(_1182_));
 sg13g2_a21oi_1 _1563_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .A2(_1183_),
    .Y(_1184_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_nand2_1 _1564_ (.Y(_1185_),
    .A(net1048),
    .B(net504));
 sg13g2_o21ai_1 _1565_ (.B1(_1185_),
    .Y(_1186_),
    .A1(net1048),
    .A2(net976));
 sg13g2_or2_1 _1566_ (.X(_1187_),
    .B(net1066),
    .A(net1048));
 sg13g2_a21oi_1 _1567_ (.A1(net1048),
    .A2(net1016),
    .Y(_1188_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_a221oi_1 _1568_ (.B2(_1188_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .B1(_1187_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_1189_),
    .A2(_1186_));
 sg13g2_nand2_2 _1569_ (.Y(_1190_),
    .A(net1048),
    .B(net1012));
 sg13g2_nand2b_1 _1570_ (.Y(_1191_),
    .B(net1030),
    .A_N(net1048));
 sg13g2_a21oi_2 _1571_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_1192_),
    .A2(_1190_),
    .A1(_1191_));
 sg13g2_nor2b_1 _1572_ (.A(net1001),
    .B_N(net1048),
    .Y(_1193_));
 sg13g2_o21ai_1 _1573_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .Y(_1194_),
    .A1(net1048),
    .A2(net985));
 sg13g2_o21ai_1 _1574_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .Y(_1195_),
    .A1(_1193_),
    .A2(_1194_));
 sg13g2_o21ai_1 _1575_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .Y(_1196_),
    .A1(_1195_),
    .A2(_1192_));
 sg13g2_mux4_1 _1576_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net1074),
    .A1(net38),
    .A2(net50),
    .A3(net9),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1197_));
 sg13g2_mux4_1 _1577_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .A0(net1217),
    .A1(net66),
    .A2(net85),
    .A3(net93),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .X(_1198_));
 sg13g2_nand2b_1 _1578_ (.Y(_1199_),
    .B(_1197_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_nand2_1 _1579_ (.Y(_1200_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .B(_1198_));
 sg13g2_a21o_1 _1580_ (.A2(_1200_),
    .A1(_1199_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .X(_1201_));
 sg13g2_o21ai_1 _1581_ (.B1(_1201_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .A1(_1189_),
    .A2(_1196_));
 sg13g2_mux2_1 _1582_ (.A0(net80),
    .A1(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_1202_));
 sg13g2_nor2b_1 _1583_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .B_N(net56),
    .Y(_1203_));
 sg13g2_a21oi_1 _1584_ (.A1(net7),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_o21ai_1 _1585_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .Y(_1205_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_1204_));
 sg13g2_a21o_1 _1586_ (.A2(_1202_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .B1(_1205_),
    .X(_1206_));
 sg13g2_mux4_1 _1587_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(net37),
    .A1(net8),
    .A2(net65),
    .A3(net107),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ),
    .X(_1207_));
 sg13g2_nor2_1 _1588_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_nor2b_1 _1589_ (.A(_1208_),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ),
    .Y(_1209_));
 sg13g2_a22oi_1 _1590_ (.Y(_1210_),
    .B1(_1206_),
    .B2(_1209_),
    .A2(_1184_),
    .A1(_1181_));
 sg13g2_nor2b_1 _1591_ (.A(net929),
    .B_N(\Inst_RegFile_32x4.mem[8][0] ),
    .Y(_1211_));
 sg13g2_a21oi_1 _1592_ (.A1(\Inst_RegFile_32x4.mem[9][0] ),
    .A2(net929),
    .Y(_1212_),
    .B1(_1211_));
 sg13g2_nand2b_1 _1593_ (.Y(_1213_),
    .B(\Inst_RegFile_32x4.mem[10][0] ),
    .A_N(net928));
 sg13g2_a21oi_1 _1594_ (.A1(\Inst_RegFile_32x4.mem[11][0] ),
    .A2(net928),
    .Y(_1214_),
    .B1(net1027));
 sg13g2_mux4_1 _1595_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(net1070),
    .A1(net1019),
    .A2(net980),
    .A3(net967),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1215_));
 sg13g2_nor2_1 _1596_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_nor2_1 _1597_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .B(net975),
    .Y(_1217_));
 sg13g2_nor2b_1 _1598_ (.A(net1033),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .Y(_1218_));
 sg13g2_nor3_1 _1599_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .B(_1217_),
    .C(_1218_),
    .Y(_1219_));
 sg13g2_mux2_1 _1600_ (.A0(net988),
    .A1(BD3),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1220_));
 sg13g2_a21o_1 _1601_ (.A2(_1220_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .B1(_1142_),
    .X(_1221_));
 sg13g2_o21ai_1 _1602_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .Y(_1222_),
    .A1(_1219_),
    .A2(_1221_));
 sg13g2_mux2_1 _1603_ (.A0(net3),
    .A1(net11),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1223_));
 sg13g2_mux2_1 _1604_ (.A0(net1074),
    .A1(net40),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1224_));
 sg13g2_mux2_1 _1605_ (.A0(net84),
    .A1(net1072),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1225_));
 sg13g2_mux2_1 _1606_ (.A0(net60),
    .A1(net68),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_1226_));
 sg13g2_mux4_1 _1607_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(_1224_),
    .A1(_1226_),
    .A2(_1223_),
    .A3(_1225_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .X(_1227_));
 sg13g2_nand2b_1 _1608_ (.Y(_1228_),
    .B(_1227_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_o21ai_1 _1609_ (.B1(_1228_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .A1(_1222_),
    .A2(_1216_));
 sg13g2_mux4_1 _1610_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(net46),
    .A1(net101),
    .A2(net74),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_1229_));
 sg13g2_nand2b_1 _1611_ (.Y(_1230_),
    .B(_1229_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_mux4_1 _1612_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(net47),
    .A1(net18),
    .A2(net75),
    .A3(net102),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ),
    .X(_1231_));
 sg13g2_a21oi_1 _1613_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_1231_),
    .Y(_1232_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_mux4_1 _1614_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(net1067),
    .A1(net1018),
    .A2(net979),
    .A3(net504),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_1233_));
 sg13g2_nor2_2 _1615_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_1233_),
    .Y(_1234_));
 sg13g2_nor2_1 _1616_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .B(net1029),
    .Y(_1235_));
 sg13g2_nor2b_1 _1617_ (.A(net1012),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .Y(_1236_));
 sg13g2_nor3_1 _1618_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .B(_1235_),
    .C(_1236_),
    .Y(_1237_));
 sg13g2_mux2_1 _1619_ (.A0(net985),
    .A1(net1001),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0128_));
 sg13g2_a21o_1 _1620_ (.A2(_0128_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .B1(_1143_),
    .X(_0129_));
 sg13g2_o21ai_1 _1621_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .Y(_0130_),
    .A1(_1237_),
    .A2(_0129_));
 sg13g2_mux2_1 _1622_ (.A0(net9),
    .A1(net24),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0131_));
 sg13g2_mux2_1 _1623_ (.A0(net38),
    .A1(net1219),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0132_));
 sg13g2_mux2_1 _1624_ (.A0(net78),
    .A1(net93),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0133_));
 sg13g2_mux2_1 _1625_ (.A0(net1217),
    .A1(net66),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .X(_0134_));
 sg13g2_mux4_1 _1626_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(_0132_),
    .A1(_0134_),
    .A2(_0131_),
    .A3(_0133_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_0135_));
 sg13g2_nand2b_1 _1627_ (.Y(_0136_),
    .B(_0135_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_o21ai_1 _1628_ (.B1(_0136_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .A1(_0130_),
    .A2(_1234_));
 sg13g2_mux4_1 _1629_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ),
    .A0(net51),
    .A1(net93),
    .A2(net83),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_0137_));
 sg13g2_mux4_1 _1630_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(net39),
    .A1(net10),
    .A2(net83),
    .A3(net94),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_0138_));
 sg13g2_inv_1 _1631_ (.Y(_0139_),
    .A(_0138_));
 sg13g2_o21ai_1 _1632_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ),
    .Y(_0140_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .A2(_0139_));
 sg13g2_a21oi_2 _1633_ (.B1(_0140_),
    .Y(_0141_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .A1(_0137_));
 sg13g2_a21oi_2 _1634_ (.B1(_0141_),
    .Y(_0142_),
    .A2(_1232_),
    .A1(_1230_));
 sg13g2_a21o_2 _1635_ (.A2(_1232_),
    .A1(_1230_),
    .B1(_0141_),
    .X(_0143_));
 sg13g2_a221oi_1 _1636_ (.B2(_1214_),
    .C1(net983),
    .B1(_1213_),
    .A1(net1027),
    .Y(_0144_),
    .A2(_1212_));
 sg13g2_nand2_1 _1637_ (.Y(_0145_),
    .A(net1039),
    .B(net963));
 sg13g2_o21ai_1 _1638_ (.B1(_0145_),
    .Y(_0146_),
    .A1(net1039),
    .A2(net976));
 sg13g2_or2_1 _1639_ (.X(_0147_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .A(net1067));
 sg13g2_a21oi_1 _1640_ (.A1(net1039),
    .A2(net1016),
    .Y(_0148_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_a221oi_1 _1641_ (.B2(_0148_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .B1(_0147_),
    .A1(_0146_),
    .Y(_0149_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_nand2_2 _1642_ (.Y(_0150_),
    .A(net1039),
    .B(net1012));
 sg13g2_nand2b_1 _1643_ (.Y(_0151_),
    .B(net1030),
    .A_N(net1039));
 sg13g2_a21oi_2 _1644_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .Y(_0152_),
    .A2(_0150_),
    .A1(_0151_));
 sg13g2_nor2b_1 _1645_ (.A(net1001),
    .B_N(net1039),
    .Y(_0153_));
 sg13g2_o21ai_1 _1646_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .Y(_0154_),
    .A1(net1039),
    .A2(net985));
 sg13g2_o21ai_1 _1647_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .Y(_0155_),
    .A1(_0153_),
    .A2(_0154_));
 sg13g2_o21ai_1 _1648_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ),
    .Y(_0156_),
    .A1(_0155_),
    .A2(_0152_));
 sg13g2_mux4_1 _1649_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(net1074),
    .A1(net38),
    .A2(net57),
    .A3(net9),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0157_));
 sg13g2_mux4_1 _1650_ (.S0(net1039),
    .A0(net1217),
    .A1(net66),
    .A2(net78),
    .A3(net93),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0158_));
 sg13g2_mux2_1 _1651_ (.A0(_0157_),
    .A1(_0158_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .X(_0159_));
 sg13g2_nand2b_1 _1652_ (.Y(_0160_),
    .B(_0159_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_o21ai_1 _1653_ (.B1(_0160_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .A1(_0156_),
    .A2(_0149_));
 sg13g2_o21ai_1 _1654_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .Y(_0161_),
    .A1(_1138_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_a21oi_2 _1655_ (.B1(_0161_),
    .Y(_0162_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG3 ));
 sg13g2_mux2_1 _1656_ (.A0(net24),
    .A1(net78),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .X(_0163_));
 sg13g2_o21ai_1 _1657_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .Y(_0164_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_0163_));
 sg13g2_mux4_1 _1658_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(net56),
    .A1(net6),
    .A2(net63),
    .A3(net90),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ),
    .X(_0165_));
 sg13g2_a21oi_1 _1659_ (.A1(_1144_),
    .A2(_0165_),
    .Y(_0166_),
    .B1(_1145_));
 sg13g2_o21ai_1 _1660_ (.B1(_0166_),
    .Y(_0167_),
    .A1(_0164_),
    .A2(_0162_));
 sg13g2_mux4_1 _1661_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(net108),
    .A1(net1019),
    .A2(net980),
    .A3(net514),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0168_));
 sg13g2_nand2b_1 _1662_ (.Y(_0169_),
    .B(_0168_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_nand2b_1 _1663_ (.Y(_0170_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .A_N(net1003));
 sg13g2_o21ai_1 _1664_ (.B1(_0170_),
    .Y(_0171_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(net989));
 sg13g2_mux2_1 _1665_ (.A0(net975),
    .A1(net1034),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_0172_));
 sg13g2_o21ai_1 _1666_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .Y(_0173_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_0172_));
 sg13g2_a21o_1 _1667_ (.A2(_0171_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .B1(_0173_),
    .X(_0174_));
 sg13g2_and2_1 _1668_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .B(_0169_),
    .X(_0175_));
 sg13g2_mux4_1 _1669_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(net32),
    .A1(net40),
    .A2(net3),
    .A3(net11),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0176_));
 sg13g2_nand2b_1 _1670_ (.Y(_0177_),
    .B(_0176_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_mux4_1 _1671_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .A0(net58),
    .A1(net68),
    .A2(net60),
    .A3(net1070),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .X(_0178_));
 sg13g2_a21oi_1 _1672_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_0178_),
    .Y(_0179_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_a22oi_1 _1673_ (.Y(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .B1(_0177_),
    .B2(_0179_),
    .A2(_0174_),
    .A1(_0175_));
 sg13g2_mux4_1 _1674_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ),
    .A0(net13),
    .A1(net97),
    .A2(net70),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ),
    .X(_0180_));
 sg13g2_mux4_1 _1675_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(net43),
    .A1(net14),
    .A2(net71),
    .A3(net98),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ),
    .X(_0181_));
 sg13g2_nand2_1 _1676_ (.Y(_0182_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .B(_0181_));
 sg13g2_a21oi_2 _1677_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .Y(_0183_),
    .A2(_0180_),
    .A1(_1144_));
 sg13g2_nand2_2 _1678_ (.Y(_0184_),
    .A(_0182_),
    .B(_0183_));
 sg13g2_and2_1 _1679_ (.A(_0184_),
    .B(_0167_),
    .X(_0185_));
 sg13g2_nand2_2 _1680_ (.Y(_0186_),
    .A(_0184_),
    .B(_0167_));
 sg13g2_mux2_1 _1681_ (.A0(\Inst_RegFile_32x4.mem[14][0] ),
    .A1(\Inst_RegFile_32x4.mem[15][0] ),
    .S(net930),
    .X(_0187_));
 sg13g2_nand2b_1 _1682_ (.Y(_0188_),
    .B(net930),
    .A_N(\Inst_RegFile_32x4.mem[13][0] ));
 sg13g2_o21ai_1 _1683_ (.B1(_0188_),
    .Y(_0189_),
    .A1(\Inst_RegFile_32x4.mem[12][0] ),
    .A2(net930));
 sg13g2_a21oi_1 _1684_ (.A1(net1026),
    .A2(_0189_),
    .Y(_0190_),
    .B1(net956));
 sg13g2_o21ai_1 _1685_ (.B1(_0190_),
    .Y(_0191_),
    .A1(net1026),
    .A2(_0187_));
 sg13g2_nand2b_1 _1686_ (.Y(_0192_),
    .B(_0191_),
    .A_N(_0144_));
 sg13g2_nand2_1 _1687_ (.Y(_0193_),
    .A(net1054),
    .B(net966));
 sg13g2_o21ai_1 _1688_ (.B1(_0193_),
    .Y(_0194_),
    .A1(net1054),
    .A2(net976));
 sg13g2_or2_1 _1689_ (.X(_0195_),
    .B(net1070),
    .A(net1054));
 sg13g2_a21oi_1 _1690_ (.A1(net1054),
    .A2(net1016),
    .Y(_0196_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_a221oi_1 _1691_ (.B2(_0196_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .B1(_0195_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .Y(_0197_),
    .A2(_0194_));
 sg13g2_nand2_1 _1692_ (.Y(_0198_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .B(net1032));
 sg13g2_nand2b_1 _1693_ (.Y(_0199_),
    .B(net973),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_a21oi_2 _1694_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .Y(_0200_),
    .A2(_0198_),
    .A1(_0199_));
 sg13g2_nor2b_1 _1695_ (.A(net1002),
    .B_N(net1054),
    .Y(_0201_));
 sg13g2_o21ai_1 _1696_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .Y(_0202_),
    .A1(net1054),
    .A2(net986));
 sg13g2_o21ai_1 _1697_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .Y(_0203_),
    .A1(_0201_),
    .A2(_0202_));
 sg13g2_o21ai_1 _1698_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ),
    .Y(_0204_),
    .A1(_0203_),
    .A2(_0200_));
 sg13g2_mux4_1 _1699_ (.S0(net1054),
    .A0(net11),
    .A1(net60),
    .A2(net68),
    .A3(net1072),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .X(_0205_));
 sg13g2_mux4_1 _1700_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .A0(net1074),
    .A1(net56),
    .A2(net40),
    .A3(net1219),
    .S1(net1054),
    .X(_0206_));
 sg13g2_mux2_1 _1701_ (.A0(_0206_),
    .A1(_0205_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .X(_0207_));
 sg13g2_nand2b_1 _1702_ (.Y(_0208_),
    .B(_0207_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_o21ai_1 _1703_ (.B1(_0208_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .A1(_0204_),
    .A2(_0197_));
 sg13g2_mux4_1 _1704_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ),
    .A0(net34),
    .A1(net62),
    .A2(net22),
    .A3(net89),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0209_));
 sg13g2_mux4_1 _1705_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .A0(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .A2(_0209_),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .S1(_1146_),
    .X(_0210_));
 sg13g2_nand2_1 _1706_ (.Y(_0211_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .B(_0210_));
 sg13g2_nand2_1 _1707_ (.Y(_0212_),
    .A(net1047),
    .B(net966));
 sg13g2_o21ai_1 _1708_ (.B1(_0212_),
    .Y(_0213_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(net976));
 sg13g2_or2_1 _1709_ (.X(_0214_),
    .B(net1047),
    .A(net1068));
 sg13g2_a21oi_1 _1710_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(net1016),
    .Y(_0215_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_a221oi_1 _1711_ (.B2(_0215_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .B1(_0214_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0216_),
    .A2(_0213_));
 sg13g2_nand2_2 _1712_ (.Y(_0217_),
    .A(net1047),
    .B(net1032));
 sg13g2_nand2b_1 _1713_ (.Y(_0218_),
    .B(net972),
    .A_N(net1047));
 sg13g2_a21oi_2 _1714_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0219_),
    .A2(_0218_),
    .A1(_0217_));
 sg13g2_nor2b_1 _1715_ (.A(net1002),
    .B_N(net1047),
    .Y(_0220_));
 sg13g2_o21ai_1 _1716_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0221_),
    .A1(net1047),
    .A2(net1015));
 sg13g2_o21ai_1 _1717_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .Y(_0222_),
    .A1(_0220_),
    .A2(_0221_));
 sg13g2_o21ai_1 _1718_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .Y(_0223_),
    .A1(_0219_),
    .A2(_0222_));
 sg13g2_mux4_1 _1719_ (.S0(net1047),
    .A0(net1073),
    .A1(net41),
    .A2(net1218),
    .A3(net12),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0224_));
 sg13g2_mux4_1 _1720_ (.S0(net1047),
    .A0(net22),
    .A1(net59),
    .A2(net61),
    .A3(net69),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0225_));
 sg13g2_mux2_1 _1721_ (.A0(_0224_),
    .A1(_0225_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .X(_0226_));
 sg13g2_nand2b_1 _1722_ (.Y(_0227_),
    .B(_0226_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_o21ai_1 _1723_ (.B1(_0227_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG6 ),
    .A1(_0223_),
    .A2(_0216_));
 sg13g2_mux4_1 _1724_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .A0(net44),
    .A1(net72),
    .A2(net99),
    .A3(\Inst_RegFile_switch_matrix.E2BEG6 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .X(_0228_));
 sg13g2_mux4_1 _1725_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ),
    .A0(net47),
    .A1(net18),
    .A2(net75),
    .A3(net102),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ),
    .X(_0229_));
 sg13g2_mux2_1 _1726_ (.A0(_0228_),
    .A1(_0229_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .X(_0230_));
 sg13g2_nand2b_1 _1727_ (.Y(_0231_),
    .B(net35),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_a21oi_1 _1728_ (.A1(net63),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .Y(_0232_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_a21oi_1 _1729_ (.A1(_0231_),
    .A2(_0232_),
    .Y(_0233_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_o21ai_1 _1730_ (.B1(_0233_),
    .Y(_0234_),
    .A1(_1146_),
    .A2(_0230_));
 sg13g2_and2_1 _1731_ (.A(_0211_),
    .B(_0234_),
    .X(_0235_));
 sg13g2_nand2_2 _1732_ (.Y(_0236_),
    .A(_0234_),
    .B(_0211_));
 sg13g2_nor2b_1 _1733_ (.A(net922),
    .B_N(\Inst_RegFile_32x4.mem[0][0] ),
    .Y(_0237_));
 sg13g2_a21oi_1 _1734_ (.A1(\Inst_RegFile_32x4.mem[1][0] ),
    .A2(net921),
    .Y(_0238_),
    .B1(_0237_));
 sg13g2_nand2b_1 _1735_ (.Y(_0239_),
    .B(\Inst_RegFile_32x4.mem[2][0] ),
    .A_N(net921));
 sg13g2_a21oi_1 _1736_ (.A1(\Inst_RegFile_32x4.mem[3][0] ),
    .A2(net921),
    .Y(_0240_),
    .B1(net1022));
 sg13g2_a221oi_1 _1737_ (.B2(_0240_),
    .C1(net982),
    .B1(_0239_),
    .A1(net1022),
    .Y(_0241_),
    .A2(_0238_));
 sg13g2_mux2_1 _1738_ (.A0(\Inst_RegFile_32x4.mem[6][0] ),
    .A1(\Inst_RegFile_32x4.mem[7][0] ),
    .S(net930),
    .X(_0242_));
 sg13g2_nor2b_1 _1739_ (.A(net930),
    .B_N(\Inst_RegFile_32x4.mem[4][0] ),
    .Y(_0243_));
 sg13g2_a21oi_1 _1740_ (.A1(\Inst_RegFile_32x4.mem[5][0] ),
    .A2(net930),
    .Y(_0244_),
    .B1(_0243_));
 sg13g2_a21oi_1 _1741_ (.A1(net1026),
    .A2(_0244_),
    .Y(_0245_),
    .B1(net956));
 sg13g2_o21ai_1 _1742_ (.B1(_0245_),
    .Y(_0246_),
    .A1(net1026),
    .A2(_0242_));
 sg13g2_nand2b_1 _1743_ (.Y(_0247_),
    .B(_0246_),
    .A_N(_0241_));
 sg13g2_mux4_1 _1744_ (.S0(net931),
    .A0(\Inst_RegFile_32x4.mem[26][0] ),
    .A1(\Inst_RegFile_32x4.mem[27][0] ),
    .A2(\Inst_RegFile_32x4.mem[24][0] ),
    .A3(\Inst_RegFile_32x4.mem[25][0] ),
    .S1(net1028),
    .X(_0248_));
 sg13g2_mux4_1 _1745_ (.S0(net922),
    .A0(\Inst_RegFile_32x4.mem[30][0] ),
    .A1(\Inst_RegFile_32x4.mem[31][0] ),
    .A2(\Inst_RegFile_32x4.mem[28][0] ),
    .A3(\Inst_RegFile_32x4.mem[29][0] ),
    .S1(net1025),
    .X(_0249_));
 sg13g2_mux2_1 _1746_ (.A0(_0248_),
    .A1(_0249_),
    .S(net982),
    .X(_0250_));
 sg13g2_nor2b_1 _1747_ (.A(net925),
    .B_N(\Inst_RegFile_32x4.mem[16][0] ),
    .Y(_0251_));
 sg13g2_a21oi_1 _1748_ (.A1(\Inst_RegFile_32x4.mem[17][0] ),
    .A2(net925),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_nand2b_1 _1749_ (.Y(_0253_),
    .B(\Inst_RegFile_32x4.mem[18][0] ),
    .A_N(net925));
 sg13g2_a21oi_1 _1750_ (.A1(\Inst_RegFile_32x4.mem[19][0] ),
    .A2(net925),
    .Y(_0254_),
    .B1(net1023));
 sg13g2_a221oi_1 _1751_ (.B2(_0254_),
    .C1(net982),
    .B1(_0253_),
    .A1(net1023),
    .Y(_0255_),
    .A2(_0252_));
 sg13g2_mux2_1 _1752_ (.A0(\Inst_RegFile_32x4.mem[22][0] ),
    .A1(\Inst_RegFile_32x4.mem[23][0] ),
    .S(net926),
    .X(_0256_));
 sg13g2_nor2b_1 _1753_ (.A(net926),
    .B_N(\Inst_RegFile_32x4.mem[20][0] ),
    .Y(_0257_));
 sg13g2_a21oi_1 _1754_ (.A1(\Inst_RegFile_32x4.mem[21][0] ),
    .A2(net926),
    .Y(_0258_),
    .B1(_0257_));
 sg13g2_a21oi_1 _1755_ (.A1(net1024),
    .A2(_0258_),
    .Y(_0259_),
    .B1(net955));
 sg13g2_o21ai_1 _1756_ (.B1(_0259_),
    .Y(_0260_),
    .A1(net1024),
    .A2(_0256_));
 sg13g2_nand2b_1 _1757_ (.Y(_0261_),
    .B(_0260_),
    .A_N(_0255_));
 sg13g2_mux4_1 _1758_ (.S0(_0186_),
    .A0(_0192_),
    .A1(_0247_),
    .A2(_0250_),
    .A3(_0261_),
    .S1(_0236_),
    .X(\Inst_RegFile_32x4.AD_comb[0] ));
 sg13g2_mux2_2 _1759_ (.A0(\Inst_RegFile_32x4.AD_comb[0] ),
    .A1(\Inst_RegFile_32x4.AD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD0));
 sg13g2_mux4_1 _1760_ (.S0(net929),
    .A0(\Inst_RegFile_32x4.mem[10][1] ),
    .A1(\Inst_RegFile_32x4.mem[11][1] ),
    .A2(\Inst_RegFile_32x4.mem[8][1] ),
    .A3(\Inst_RegFile_32x4.mem[9][1] ),
    .S1(net1027),
    .X(_0262_));
 sg13g2_nand2_1 _1761_ (.Y(_0263_),
    .A(net956),
    .B(_0262_));
 sg13g2_mux4_1 _1762_ (.S0(net926),
    .A0(\Inst_RegFile_32x4.mem[14][1] ),
    .A1(\Inst_RegFile_32x4.mem[15][1] ),
    .A2(\Inst_RegFile_32x4.mem[12][1] ),
    .A3(\Inst_RegFile_32x4.mem[13][1] ),
    .S1(net1024),
    .X(_0264_));
 sg13g2_a21oi_1 _1763_ (.A1(net982),
    .A2(_0264_),
    .Y(_0265_),
    .B1(net969));
 sg13g2_mux4_1 _1764_ (.S0(net921),
    .A0(\Inst_RegFile_32x4.mem[2][1] ),
    .A1(\Inst_RegFile_32x4.mem[3][1] ),
    .A2(\Inst_RegFile_32x4.mem[0][1] ),
    .A3(\Inst_RegFile_32x4.mem[1][1] ),
    .S1(net1022),
    .X(_0266_));
 sg13g2_nand2_2 _1765_ (.Y(_0267_),
    .A(_0143_),
    .B(_0266_));
 sg13g2_mux4_1 _1766_ (.S0(net931),
    .A0(\Inst_RegFile_32x4.mem[6][1] ),
    .A1(\Inst_RegFile_32x4.mem[7][1] ),
    .A2(\Inst_RegFile_32x4.mem[4][1] ),
    .A3(\Inst_RegFile_32x4.mem[5][1] ),
    .S1(net1028),
    .X(_0268_));
 sg13g2_a21oi_1 _1767_ (.A1(net983),
    .A2(_0268_),
    .Y(_0269_),
    .B1(_0185_));
 sg13g2_a221oi_1 _1768_ (.B2(_0269_),
    .C1(_0236_),
    .B1(_0267_),
    .A1(_0263_),
    .Y(_0270_),
    .A2(_0265_));
 sg13g2_nor2b_1 _1769_ (.A(net928),
    .B_N(\Inst_RegFile_32x4.mem[24][1] ),
    .Y(_0271_));
 sg13g2_a21oi_1 _1770_ (.A1(\Inst_RegFile_32x4.mem[25][1] ),
    .A2(net928),
    .Y(_0272_),
    .B1(_0271_));
 sg13g2_mux2_1 _1771_ (.A0(\Inst_RegFile_32x4.mem[26][1] ),
    .A1(\Inst_RegFile_32x4.mem[27][1] ),
    .S(net931),
    .X(_0273_));
 sg13g2_a21oi_1 _1772_ (.A1(net1028),
    .A2(_0272_),
    .Y(_0274_),
    .B1(net983));
 sg13g2_o21ai_1 _1773_ (.B1(_0274_),
    .Y(_0275_),
    .A1(net1028),
    .A2(_0273_));
 sg13g2_mux4_1 _1774_ (.S0(net922),
    .A0(\Inst_RegFile_32x4.mem[30][1] ),
    .A1(\Inst_RegFile_32x4.mem[31][1] ),
    .A2(\Inst_RegFile_32x4.mem[28][1] ),
    .A3(\Inst_RegFile_32x4.mem[29][1] ),
    .S1(net1025),
    .X(_0276_));
 sg13g2_a21oi_1 _1775_ (.A1(net982),
    .A2(_0276_),
    .Y(_0277_),
    .B1(net969));
 sg13g2_mux4_1 _1776_ (.S0(net925),
    .A0(\Inst_RegFile_32x4.mem[18][1] ),
    .A1(\Inst_RegFile_32x4.mem[19][1] ),
    .A2(\Inst_RegFile_32x4.mem[16][1] ),
    .A3(\Inst_RegFile_32x4.mem[17][1] ),
    .S1(net1023),
    .X(_0278_));
 sg13g2_nor2b_1 _1777_ (.A(net923),
    .B_N(\Inst_RegFile_32x4.mem[20][1] ),
    .Y(_0279_));
 sg13g2_a21oi_1 _1778_ (.A1(\Inst_RegFile_32x4.mem[21][1] ),
    .A2(net923),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_nor2b_1 _1779_ (.A(net923),
    .B_N(\Inst_RegFile_32x4.mem[22][1] ),
    .Y(_0281_));
 sg13g2_a21oi_1 _1780_ (.A1(\Inst_RegFile_32x4.mem[23][1] ),
    .A2(net923),
    .Y(_0282_),
    .B1(_0281_));
 sg13g2_nand2b_1 _1781_ (.Y(_0283_),
    .B(_0282_),
    .A_N(net1023));
 sg13g2_a21oi_1 _1782_ (.A1(net1023),
    .A2(_0280_),
    .Y(_0284_),
    .B1(net955));
 sg13g2_a22oi_1 _1783_ (.Y(_0285_),
    .B1(_0283_),
    .B2(_0284_),
    .A2(_0278_),
    .A1(net955));
 sg13g2_a221oi_1 _1784_ (.B2(net969),
    .C1(_0235_),
    .B1(_0285_),
    .A1(_0275_),
    .Y(_0286_),
    .A2(_0277_));
 sg13g2_or2_1 _1785_ (.X(\Inst_RegFile_32x4.AD_comb[1] ),
    .B(_0270_),
    .A(_0286_));
 sg13g2_mux2_2 _1786_ (.A0(\Inst_RegFile_32x4.AD_comb[1] ),
    .A1(\Inst_RegFile_32x4.AD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD1));
 sg13g2_mux4_1 _1787_ (.S0(net929),
    .A0(\Inst_RegFile_32x4.mem[10][2] ),
    .A1(\Inst_RegFile_32x4.mem[11][2] ),
    .A2(\Inst_RegFile_32x4.mem[8][2] ),
    .A3(\Inst_RegFile_32x4.mem[9][2] ),
    .S1(net1027),
    .X(_0287_));
 sg13g2_nand2_1 _1788_ (.Y(_0288_),
    .A(net956),
    .B(_0287_));
 sg13g2_mux4_1 _1789_ (.S0(net927),
    .A0(\Inst_RegFile_32x4.mem[14][2] ),
    .A1(\Inst_RegFile_32x4.mem[15][2] ),
    .A2(\Inst_RegFile_32x4.mem[12][2] ),
    .A3(\Inst_RegFile_32x4.mem[13][2] ),
    .S1(net1026),
    .X(_0289_));
 sg13g2_a21oi_1 _1790_ (.A1(net982),
    .A2(_0289_),
    .Y(_0290_),
    .B1(net969));
 sg13g2_mux4_1 _1791_ (.S0(net921),
    .A0(\Inst_RegFile_32x4.mem[2][2] ),
    .A1(\Inst_RegFile_32x4.mem[3][2] ),
    .A2(\Inst_RegFile_32x4.mem[0][2] ),
    .A3(\Inst_RegFile_32x4.mem[1][2] ),
    .S1(net1022),
    .X(_0291_));
 sg13g2_nor2b_1 _1792_ (.A(net926),
    .B_N(\Inst_RegFile_32x4.mem[4][2] ),
    .Y(_0292_));
 sg13g2_a21oi_1 _1793_ (.A1(\Inst_RegFile_32x4.mem[5][2] ),
    .A2(net926),
    .Y(_0293_),
    .B1(_0292_));
 sg13g2_nor2b_1 _1794_ (.A(net926),
    .B_N(\Inst_RegFile_32x4.mem[6][2] ),
    .Y(_0294_));
 sg13g2_a21oi_1 _1795_ (.A1(\Inst_RegFile_32x4.mem[7][2] ),
    .A2(net926),
    .Y(_0295_),
    .B1(_0294_));
 sg13g2_nand2b_1 _1796_ (.Y(_0296_),
    .B(_0295_),
    .A_N(net1024));
 sg13g2_a21oi_1 _1797_ (.A1(net1024),
    .A2(_0293_),
    .Y(_0297_),
    .B1(net956));
 sg13g2_a22oi_1 _1798_ (.Y(_0298_),
    .B1(_0296_),
    .B2(_0297_),
    .A2(_0291_),
    .A1(net955));
 sg13g2_a221oi_1 _1799_ (.B2(net520),
    .C1(_0236_),
    .B1(_0298_),
    .A1(_0288_),
    .Y(_0299_),
    .A2(_0290_));
 sg13g2_mux4_1 _1800_ (.S0(net928),
    .A0(\Inst_RegFile_32x4.mem[26][2] ),
    .A1(\Inst_RegFile_32x4.mem[27][2] ),
    .A2(\Inst_RegFile_32x4.mem[24][2] ),
    .A3(\Inst_RegFile_32x4.mem[25][2] ),
    .S1(net1027),
    .X(_0300_));
 sg13g2_mux4_1 _1801_ (.S0(net921),
    .A0(\Inst_RegFile_32x4.mem[30][2] ),
    .A1(\Inst_RegFile_32x4.mem[31][2] ),
    .A2(\Inst_RegFile_32x4.mem[28][2] ),
    .A3(\Inst_RegFile_32x4.mem[29][2] ),
    .S1(net1022),
    .X(_0301_));
 sg13g2_nand2_2 _1802_ (.Y(_0302_),
    .A(net982),
    .B(_0301_));
 sg13g2_a21oi_1 _1803_ (.A1(net956),
    .A2(_0300_),
    .Y(_0303_),
    .B1(net969));
 sg13g2_mux4_1 _1804_ (.S0(net925),
    .A0(\Inst_RegFile_32x4.mem[18][2] ),
    .A1(\Inst_RegFile_32x4.mem[19][2] ),
    .A2(\Inst_RegFile_32x4.mem[16][2] ),
    .A3(\Inst_RegFile_32x4.mem[17][2] ),
    .S1(net1023),
    .X(_0304_));
 sg13g2_nor2b_1 _1805_ (.A(net924),
    .B_N(\Inst_RegFile_32x4.mem[20][2] ),
    .Y(_0305_));
 sg13g2_a21oi_1 _1806_ (.A1(\Inst_RegFile_32x4.mem[21][2] ),
    .A2(net924),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_nor2b_1 _1807_ (.A(net923),
    .B_N(\Inst_RegFile_32x4.mem[22][2] ),
    .Y(_0307_));
 sg13g2_a21oi_1 _1808_ (.A1(\Inst_RegFile_32x4.mem[23][2] ),
    .A2(net923),
    .Y(_0308_),
    .B1(_0307_));
 sg13g2_nand2b_1 _1809_ (.Y(_0309_),
    .B(_0308_),
    .A_N(net1024));
 sg13g2_a21oi_1 _1810_ (.A1(net1024),
    .A2(_0306_),
    .Y(_0310_),
    .B1(net955));
 sg13g2_a22oi_1 _1811_ (.Y(_0311_),
    .B1(_0309_),
    .B2(_0310_),
    .A2(_0304_),
    .A1(net955));
 sg13g2_a221oi_1 _1812_ (.B2(net520),
    .C1(_0235_),
    .B1(_0311_),
    .A1(_0303_),
    .Y(_0312_),
    .A2(_0302_));
 sg13g2_or2_1 _1813_ (.X(\Inst_RegFile_32x4.AD_comb[2] ),
    .B(_0299_),
    .A(_0312_));
 sg13g2_mux2_2 _1814_ (.A0(\Inst_RegFile_32x4.AD_comb[2] ),
    .A1(\Inst_RegFile_32x4.AD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD2));
 sg13g2_mux4_1 _1815_ (.S0(net929),
    .A0(\Inst_RegFile_32x4.mem[10][3] ),
    .A1(\Inst_RegFile_32x4.mem[11][3] ),
    .A2(\Inst_RegFile_32x4.mem[8][3] ),
    .A3(\Inst_RegFile_32x4.mem[9][3] ),
    .S1(net1027),
    .X(_0313_));
 sg13g2_mux4_1 _1816_ (.S0(net930),
    .A0(\Inst_RegFile_32x4.mem[14][3] ),
    .A1(\Inst_RegFile_32x4.mem[15][3] ),
    .A2(\Inst_RegFile_32x4.mem[12][3] ),
    .A3(\Inst_RegFile_32x4.mem[13][3] ),
    .S1(net1026),
    .X(_0314_));
 sg13g2_nand2_1 _1817_ (.Y(_0315_),
    .A(net983),
    .B(_0314_));
 sg13g2_a21oi_1 _1818_ (.A1(net956),
    .A2(_0313_),
    .Y(_0316_),
    .B1(net969));
 sg13g2_mux4_1 _1819_ (.S0(net921),
    .A0(\Inst_RegFile_32x4.mem[2][3] ),
    .A1(\Inst_RegFile_32x4.mem[3][3] ),
    .A2(\Inst_RegFile_32x4.mem[0][3] ),
    .A3(\Inst_RegFile_32x4.mem[1][3] ),
    .S1(net1022),
    .X(_0317_));
 sg13g2_nand2_1 _1820_ (.Y(_0318_),
    .A(_0143_),
    .B(_0317_));
 sg13g2_mux4_1 _1821_ (.S0(net927),
    .A0(\Inst_RegFile_32x4.mem[6][3] ),
    .A1(\Inst_RegFile_32x4.mem[7][3] ),
    .A2(\Inst_RegFile_32x4.mem[4][3] ),
    .A3(\Inst_RegFile_32x4.mem[5][3] ),
    .S1(net1026),
    .X(_0319_));
 sg13g2_a21oi_1 _1822_ (.A1(net983),
    .A2(_0319_),
    .Y(_0320_),
    .B1(_0185_));
 sg13g2_a221oi_1 _1823_ (.B2(_0320_),
    .C1(_0236_),
    .B1(_0318_),
    .A1(_0315_),
    .Y(_0321_),
    .A2(_0316_));
 sg13g2_mux2_1 _1824_ (.A0(\Inst_RegFile_32x4.mem[26][3] ),
    .A1(\Inst_RegFile_32x4.mem[27][3] ),
    .S(net928),
    .X(_0322_));
 sg13g2_nor2b_1 _1825_ (.A(net928),
    .B_N(\Inst_RegFile_32x4.mem[24][3] ),
    .Y(_0323_));
 sg13g2_a21oi_1 _1826_ (.A1(\Inst_RegFile_32x4.mem[25][3] ),
    .A2(net928),
    .Y(_0324_),
    .B1(_0323_));
 sg13g2_a21oi_1 _1827_ (.A1(net1027),
    .A2(_0324_),
    .Y(_0325_),
    .B1(net983));
 sg13g2_o21ai_1 _1828_ (.B1(_0325_),
    .Y(_0326_),
    .A1(net1026),
    .A2(_0322_));
 sg13g2_mux4_1 _1829_ (.S0(net922),
    .A0(\Inst_RegFile_32x4.mem[30][3] ),
    .A1(\Inst_RegFile_32x4.mem[31][3] ),
    .A2(\Inst_RegFile_32x4.mem[28][3] ),
    .A3(\Inst_RegFile_32x4.mem[29][3] ),
    .S1(net1022),
    .X(_0327_));
 sg13g2_a21oi_1 _1830_ (.A1(net982),
    .A2(_0327_),
    .Y(_0328_),
    .B1(net969));
 sg13g2_mux4_1 _1831_ (.S0(net921),
    .A0(\Inst_RegFile_32x4.mem[18][3] ),
    .A1(\Inst_RegFile_32x4.mem[19][3] ),
    .A2(\Inst_RegFile_32x4.mem[16][3] ),
    .A3(\Inst_RegFile_32x4.mem[17][3] ),
    .S1(net1022),
    .X(_0329_));
 sg13g2_nor2b_1 _1832_ (.A(net924),
    .B_N(\Inst_RegFile_32x4.mem[20][3] ),
    .Y(_0330_));
 sg13g2_a21oi_1 _1833_ (.A1(\Inst_RegFile_32x4.mem[21][3] ),
    .A2(net923),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_nor2b_1 _1834_ (.A(net924),
    .B_N(\Inst_RegFile_32x4.mem[22][3] ),
    .Y(_0332_));
 sg13g2_a21oi_1 _1835_ (.A1(\Inst_RegFile_32x4.mem[23][3] ),
    .A2(net923),
    .Y(_0333_),
    .B1(_0332_));
 sg13g2_nand2b_1 _1836_ (.Y(_0334_),
    .B(_0333_),
    .A_N(net1023));
 sg13g2_a21oi_1 _1837_ (.A1(net1023),
    .A2(_0331_),
    .Y(_0335_),
    .B1(net955));
 sg13g2_a22oi_1 _1838_ (.Y(_0336_),
    .B1(_0334_),
    .B2(_0335_),
    .A2(_0329_),
    .A1(net955));
 sg13g2_a22oi_1 _1839_ (.Y(_0337_),
    .B1(_0336_),
    .B2(net969),
    .A2(_0328_),
    .A1(_0326_));
 sg13g2_a21o_1 _1840_ (.A2(_0236_),
    .A1(_0337_),
    .B1(_0321_),
    .X(\Inst_RegFile_32x4.AD_comb[3] ));
 sg13g2_mux2_2 _1841_ (.A0(\Inst_RegFile_32x4.AD_comb[3] ),
    .A1(\Inst_RegFile_32x4.AD_reg[3] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .X(AD3));
 sg13g2_mux4_1 _1842_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ),
    .A0(net45),
    .A1(net16),
    .A2(net73),
    .A3(net100),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ),
    .X(_0338_));
 sg13g2_inv_1 _1843_ (.Y(_0339_),
    .A(_0338_));
 sg13g2_a21oi_1 _1844_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_0339_),
    .Y(_0340_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_o21ai_1 _1845_ (.B1(_0340_),
    .Y(_0341_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_0228_));
 sg13g2_mux2_1 _1846_ (.A0(net978),
    .A1(net966),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0342_));
 sg13g2_nand2_1 _1847_ (.Y(_0343_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .B(_0342_));
 sg13g2_mux2_1 _1848_ (.A0(net87),
    .A1(net1017),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0344_));
 sg13g2_a21oi_1 _1849_ (.A1(_1133_),
    .A2(_0344_),
    .Y(_0345_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_mux2_1 _1850_ (.A0(net971),
    .A1(net1013),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .X(_0346_));
 sg13g2_o21ai_1 _1851_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .Y(_0347_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(net987));
 sg13g2_a21o_1 _1852_ (.A2(net999),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .B1(_0347_),
    .X(_0348_));
 sg13g2_a21oi_2 _1853_ (.B1(_1134_),
    .Y(_0349_),
    .A2(_0346_),
    .A1(_1133_));
 sg13g2_a221oi_1 _1854_ (.B2(_0349_),
    .C1(_1135_),
    .B1(_0348_),
    .A1(_0343_),
    .Y(_0350_),
    .A2(_0345_));
 sg13g2_mux4_1 _1855_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net1075),
    .A1(net39),
    .A2(net1220),
    .A3(net10),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0351_));
 sg13g2_nor2_1 _1856_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .B(_0351_),
    .Y(_0352_));
 sg13g2_mux4_1 _1857_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .A0(net24),
    .A1(net59),
    .A2(net61),
    .A3(net67),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .X(_0353_));
 sg13g2_o21ai_1 _1858_ (.B1(_1135_),
    .Y(_0354_),
    .A1(_1134_),
    .A2(_0353_));
 sg13g2_nor2_1 _1859_ (.A(_0352_),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_nor2_2 _1860_ (.A(_0350_),
    .B(_0355_),
    .Y(_0356_));
 sg13g2_inv_4 _1861_ (.A(_0356_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG4 ));
 sg13g2_o21ai_1 _1862_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0357_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(net91));
 sg13g2_a21oi_1 _1863_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0356_),
    .Y(_0358_),
    .B1(_0357_));
 sg13g2_nor2b_1 _1864_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .B_N(net52),
    .Y(_0359_));
 sg13g2_a21oi_1 _1865_ (.A1(net84),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_o21ai_1 _1866_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .Y(_0361_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0360_));
 sg13g2_mux4_1 _1867_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(net37),
    .A1(net8),
    .A2(net82),
    .A3(net92),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ),
    .X(_0362_));
 sg13g2_inv_1 _1868_ (.Y(_0363_),
    .A(_0362_));
 sg13g2_nor2_1 _1869_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .B(_0362_),
    .Y(_0364_));
 sg13g2_nor2b_1 _1870_ (.A(_0364_),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .Y(_0365_));
 sg13g2_o21ai_1 _1871_ (.B1(_0365_),
    .Y(_0366_),
    .A1(_0358_),
    .A2(_0361_));
 sg13g2_and2_1 _1872_ (.A(_0341_),
    .B(_0366_),
    .X(_0367_));
 sg13g2_nand2_1 _1873_ (.Y(_0368_),
    .A(_0341_),
    .B(_0366_));
 sg13g2_nor2b_1 _1874_ (.A(net994),
    .B_N(\Inst_RegFile_32x4.mem[10][0] ),
    .Y(_0369_));
 sg13g2_a21oi_1 _1875_ (.A1(\Inst_RegFile_32x4.mem[11][0] ),
    .A2(net994),
    .Y(_0370_),
    .B1(_0369_));
 sg13g2_nand2_1 _1876_ (.Y(_0371_),
    .A(net948),
    .B(_0370_));
 sg13g2_mux4_1 _1877_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net1068),
    .A1(net1017),
    .A2(net978),
    .A3(net965),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0372_));
 sg13g2_nor2_2 _1878_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_0372_),
    .Y(_0373_));
 sg13g2_nor2_1 _1879_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .B(net972),
    .Y(_0374_));
 sg13g2_nor2b_1 _1880_ (.A(net1032),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .Y(_0375_));
 sg13g2_nor3_2 _1881_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .B(_0374_),
    .C(_0375_),
    .Y(_0376_));
 sg13g2_nand2_1 _1882_ (.Y(_0377_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .B(net1002));
 sg13g2_o21ai_1 _1883_ (.B1(_0377_),
    .Y(_0378_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(net1011));
 sg13g2_a21o_1 _1884_ (.A2(_0378_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .B1(_1136_),
    .X(_0379_));
 sg13g2_o21ai_1 _1885_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .Y(_0380_),
    .A1(_0379_),
    .A2(_0376_));
 sg13g2_mux4_1 _1886_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .A0(net1073),
    .A1(net41),
    .A2(net1218),
    .A3(net12),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .X(_0381_));
 sg13g2_mux2_1 _1887_ (.A0(net83),
    .A1(net1071),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0382_));
 sg13g2_mux2_1 _1888_ (.A0(net61),
    .A1(net69),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .X(_0383_));
 sg13g2_nand2b_1 _1889_ (.Y(_0384_),
    .B(_0383_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_a21oi_1 _1890_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_0382_),
    .Y(_0385_),
    .B1(_1136_));
 sg13g2_a21oi_1 _1891_ (.A1(_0384_),
    .A2(_0385_),
    .Y(_0386_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_o21ai_1 _1892_ (.B1(_0386_),
    .Y(_0387_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_0381_));
 sg13g2_o21ai_1 _1893_ (.B1(_0387_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .A1(_0380_),
    .A2(_0373_));
 sg13g2_mux4_1 _1894_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ),
    .A0(net17),
    .A1(net74),
    .A2(net101),
    .A3(net563),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0388_));
 sg13g2_nand2_1 _1895_ (.Y(_0389_),
    .A(net1043),
    .B(net966));
 sg13g2_o21ai_1 _1896_ (.B1(_0389_),
    .Y(_0390_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(net976));
 sg13g2_nor2_1 _1897_ (.A(net1068),
    .B(net1043),
    .Y(_0391_));
 sg13g2_nor2b_1 _1898_ (.A(net1018),
    .B_N(net1043),
    .Y(_0392_));
 sg13g2_nor3_1 _1899_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0391_),
    .C(_0392_),
    .Y(_0393_));
 sg13g2_a21oi_1 _1900_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_0390_),
    .Y(_0394_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_nor2b_1 _1901_ (.A(_0393_),
    .B_N(_0394_),
    .Y(_0395_));
 sg13g2_nor2b_1 _1902_ (.A(net1003),
    .B_N(net1043),
    .Y(_0396_));
 sg13g2_o21ai_1 _1903_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0397_),
    .A1(net1043),
    .A2(net987));
 sg13g2_nand2_2 _1904_ (.Y(_0398_),
    .A(net1043),
    .B(net1014));
 sg13g2_nand2b_1 _1905_ (.Y(_0399_),
    .B(net972),
    .A_N(net1043));
 sg13g2_a21oi_2 _1906_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0400_),
    .A2(_0399_),
    .A1(_0398_));
 sg13g2_o21ai_1 _1907_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .Y(_0401_),
    .A1(_0396_),
    .A2(_0397_));
 sg13g2_o21ai_1 _1908_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ),
    .Y(_0402_),
    .A1(_0401_),
    .A2(_0400_));
 sg13g2_mux4_1 _1909_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(net1075),
    .A1(net39),
    .A2(net1220),
    .A3(net10),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0403_));
 sg13g2_mux4_1 _1910_ (.S0(net1043),
    .A0(net59),
    .A1(net67),
    .A2(net85),
    .A3(net1071),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0404_));
 sg13g2_mux2_1 _1911_ (.A0(_0403_),
    .A1(_0404_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .X(_0405_));
 sg13g2_nand2b_1 _1912_ (.Y(_0406_),
    .B(_0405_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_o21ai_1 _1913_ (.B1(_0406_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .A1(_0402_),
    .A2(_0395_));
 sg13g2_mux4_1 _1914_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .A0(net1215),
    .A1(net79),
    .A2(net109),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .X(_0407_));
 sg13g2_mux4_1 _1915_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(net55),
    .A1(net10),
    .A2(net67),
    .A3(net94),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ),
    .X(_0408_));
 sg13g2_mux4_1 _1916_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .A0(_0388_),
    .A1(_0408_),
    .A2(_0229_),
    .A3(_0407_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .X(_0409_));
 sg13g2_nor2b_1 _1917_ (.A(net995),
    .B_N(\Inst_RegFile_32x4.mem[8][0] ),
    .Y(_0410_));
 sg13g2_a21oi_1 _1918_ (.A1(\Inst_RegFile_32x4.mem[9][0] ),
    .A2(net995),
    .Y(_0411_),
    .B1(_0410_));
 sg13g2_a21oi_1 _1919_ (.A1(_0367_),
    .A2(_0411_),
    .Y(_0412_),
    .B1(net1009));
 sg13g2_nand2_1 _1920_ (.Y(_0413_),
    .A(net1038),
    .B(net504));
 sg13g2_o21ai_1 _1921_ (.B1(_0413_),
    .Y(_0414_),
    .A1(net1038),
    .A2(net976));
 sg13g2_or2_1 _1922_ (.X(_0415_),
    .B(net1038),
    .A(net109));
 sg13g2_a21oi_1 _1923_ (.A1(net1038),
    .A2(_1166_),
    .Y(_0416_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_a221oi_1 _1924_ (.B2(_0416_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .B1(_0415_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0417_),
    .A2(_0414_));
 sg13g2_nand2_1 _1925_ (.Y(_0418_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .B(net1014));
 sg13g2_nand2b_1 _1926_ (.Y(_0419_),
    .B(net973),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_a21oi_2 _1927_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0420_),
    .A2(_0419_),
    .A1(_0418_));
 sg13g2_nor2b_1 _1928_ (.A(net1002),
    .B_N(net1038),
    .Y(_0421_));
 sg13g2_o21ai_1 _1929_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .Y(_0422_),
    .A1(net1038),
    .A2(net987));
 sg13g2_o21ai_1 _1930_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .Y(_0423_),
    .A1(_0421_),
    .A2(_0422_));
 sg13g2_o21ai_1 _1931_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ),
    .Y(_0424_),
    .A1(_0423_),
    .A2(_0420_));
 sg13g2_mux4_1 _1932_ (.S0(net1038),
    .A0(net1075),
    .A1(net39),
    .A2(net1220),
    .A3(net10),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0425_));
 sg13g2_mux4_1 _1933_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .A0(net59),
    .A1(net67),
    .A2(net61),
    .A3(net1071),
    .S1(net1038),
    .X(_0426_));
 sg13g2_mux2_1 _1934_ (.A0(_0425_),
    .A1(_0426_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .X(_0427_));
 sg13g2_nand2b_1 _1935_ (.Y(_0428_),
    .B(_0427_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_o21ai_1 _1936_ (.B1(_0428_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .A1(_0424_),
    .A2(_0417_));
 sg13g2_mux4_1 _1937_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ),
    .A0(net54),
    .A1(net1216),
    .A2(net89),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ),
    .X(_0429_));
 sg13g2_inv_4 _1938_ (.A(_0429_),
    .Y(_0430_));
 sg13g2_mux4_1 _1939_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(net35),
    .A1(net63),
    .A2(net24),
    .A3(net90),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ),
    .X(_0431_));
 sg13g2_inv_1 _1940_ (.Y(_0432_),
    .A(_0431_));
 sg13g2_o21ai_1 _1941_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .Y(_0433_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .A2(_0431_));
 sg13g2_a21o_1 _1942_ (.A2(_0430_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .B1(_0433_),
    .X(_0434_));
 sg13g2_nor2b_1 _1943_ (.A(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .B_N(net71),
    .Y(_0435_));
 sg13g2_a21oi_1 _1944_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .A2(net98),
    .Y(_0436_),
    .B1(_0435_));
 sg13g2_mux2_1 _1945_ (.A0(net43),
    .A1(net14),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .X(_0437_));
 sg13g2_o21ai_1 _1946_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .Y(_0438_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ),
    .A2(_0437_));
 sg13g2_a21oi_1 _1947_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ),
    .A2(_0436_),
    .Y(_0439_),
    .B1(_0438_));
 sg13g2_mux2_1 _1948_ (.A0(net973),
    .A1(net1033),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0440_));
 sg13g2_or2_1 _1949_ (.X(_0441_),
    .B(_0440_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_nor2b_1 _1950_ (.A(BD3),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .Y(_0442_));
 sg13g2_nor2_2 _1951_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .B(BD1),
    .Y(_0443_));
 sg13g2_o21ai_1 _1952_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .Y(_0444_),
    .A1(_0443_),
    .A2(_0442_));
 sg13g2_nand3_1 _1953_ (.B(_0444_),
    .C(_0441_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .Y(_0445_));
 sg13g2_mux4_1 _1954_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net107),
    .A1(net1017),
    .A2(net515),
    .A3(net967),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0446_));
 sg13g2_nand2b_1 _1955_ (.Y(_0447_),
    .B(_0446_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_and2_1 _1956_ (.A(_0447_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_0448_));
 sg13g2_mux4_1 _1957_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(net33),
    .A1(net41),
    .A2(net4),
    .A3(net12),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0449_));
 sg13g2_nand2b_1 _1958_ (.Y(_0450_),
    .B(_0449_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_mux4_1 _1959_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .A0(net59),
    .A1(net69),
    .A2(net61),
    .A3(net1068),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .X(_0451_));
 sg13g2_a21oi_1 _1960_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_0451_),
    .Y(_0452_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_a22oi_1 _1961_ (.Y(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .B1(_0450_),
    .B2(_0452_),
    .A2(_0448_),
    .A1(_0445_));
 sg13g2_or2_1 _1962_ (.X(_0453_),
    .B(net97),
    .A(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_o21ai_1 _1963_ (.B1(_0453_),
    .Y(_0454_),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .A2(_1137_));
 sg13g2_nand2_1 _1964_ (.Y(_0455_),
    .A(net13),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_a21oi_1 _1965_ (.A1(net42),
    .A2(_1137_),
    .Y(_0456_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_a221oi_1 _1966_ (.B2(_0456_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .B1(_0455_),
    .A1(_0454_),
    .Y(_0457_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_o21ai_1 _1967_ (.B1(_1139_),
    .Y(_0458_),
    .A1(_0457_),
    .A2(_0439_));
 sg13g2_and2_2 _1968_ (.A(_0458_),
    .B(_0434_),
    .X(_0459_));
 sg13g2_nand2_2 _1969_ (.Y(_0460_),
    .A(_0434_),
    .B(net518));
 sg13g2_mux4_1 _1970_ (.S0(net997),
    .A0(\Inst_RegFile_32x4.mem[12][0] ),
    .A1(\Inst_RegFile_32x4.mem[13][0] ),
    .A2(\Inst_RegFile_32x4.mem[14][0] ),
    .A3(\Inst_RegFile_32x4.mem[15][0] ),
    .S1(net947),
    .X(_0461_));
 sg13g2_a22oi_1 _1971_ (.Y(_0462_),
    .B1(_0461_),
    .B2(net1008),
    .A2(_0412_),
    .A1(_0371_));
 sg13g2_nand2_1 _1972_ (.Y(_0463_),
    .A(net1053),
    .B(net966));
 sg13g2_o21ai_1 _1973_ (.B1(_0463_),
    .Y(_0464_),
    .A1(net1052),
    .A2(net977));
 sg13g2_nor2b_1 _1974_ (.A(net1052),
    .B_N(net1069),
    .Y(_0465_));
 sg13g2_a21oi_1 _1975_ (.A1(net1052),
    .A2(net506),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_a21oi_1 _1976_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0464_),
    .Y(_0467_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_o21ai_1 _1977_ (.B1(_0467_),
    .Y(_0468_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0466_));
 sg13g2_nor2b_1 _1978_ (.A(net1052),
    .B_N(net971),
    .Y(_0469_));
 sg13g2_a21oi_1 _1979_ (.A1(net1052),
    .A2(net1032),
    .Y(_0470_),
    .B1(_0469_));
 sg13g2_nand2_1 _1980_ (.Y(_0471_),
    .A(net1053),
    .B(net1002));
 sg13g2_o21ai_1 _1981_ (.B1(_0471_),
    .Y(_0472_),
    .A1(net1052),
    .A2(net1011));
 sg13g2_a21oi_2 _1982_ (.B1(_1132_),
    .Y(_0473_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .A1(_0472_));
 sg13g2_o21ai_1 _1983_ (.B1(_0473_),
    .Y(_0474_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0470_));
 sg13g2_nand3_1 _1984_ (.B(_0468_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ),
    .A(_0474_),
    .Y(_0475_));
 sg13g2_mux4_1 _1985_ (.S0(net1052),
    .A0(net33),
    .A1(net41),
    .A2(net55),
    .A3(net4),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .X(_0476_));
 sg13g2_mux2_1 _1986_ (.A0(net69),
    .A1(net1071),
    .S(net1052),
    .X(_0477_));
 sg13g2_nor2b_1 _1987_ (.A(net1053),
    .B_N(net12),
    .Y(_0478_));
 sg13g2_a21oi_1 _1988_ (.A1(net1053),
    .A2(net61),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_a21oi_1 _1989_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0477_),
    .Y(_0480_),
    .B1(_1132_));
 sg13g2_o21ai_1 _1990_ (.B1(_0480_),
    .Y(_0481_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .A2(_0479_));
 sg13g2_o21ai_1 _1991_ (.B1(_0481_),
    .Y(_0482_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .A2(_0476_));
 sg13g2_o21ai_1 _1992_ (.B1(_0475_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ),
    .A2(_0482_));
 sg13g2_mux4_1 _1993_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .A0(_0165_),
    .A1(net516),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .X(_0483_));
 sg13g2_mux4_1 _1994_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ),
    .A0(net15),
    .A1(net99),
    .A2(net72),
    .A3(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ),
    .X(_0484_));
 sg13g2_nand2b_1 _1995_ (.Y(_0485_),
    .B(_0484_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_mux4_1 _1996_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(net47),
    .A1(net18),
    .A2(net75),
    .A3(net102),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0486_));
 sg13g2_a21oi_1 _1997_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(_0486_),
    .Y(_0487_),
    .B1(_1140_));
 sg13g2_nor2b_1 _1998_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .B_N(net36),
    .Y(_0488_));
 sg13g2_a21oi_1 _1999_ (.A1(net64),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_a221oi_1 _2000_ (.B2(_1140_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .B1(_0489_),
    .A1(_0485_),
    .Y(_0490_),
    .A2(_0487_));
 sg13g2_a21oi_2 _2001_ (.B1(_0490_),
    .Y(_0491_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .A1(_0483_));
 sg13g2_a21o_1 _2002_ (.A2(_0483_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .B1(_0490_),
    .X(_0492_));
 sg13g2_mux4_1 _2003_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[0][0] ),
    .A1(\Inst_RegFile_32x4.mem[1][0] ),
    .A2(\Inst_RegFile_32x4.mem[2][0] ),
    .A3(\Inst_RegFile_32x4.mem[3][0] ),
    .S1(net944),
    .X(_0493_));
 sg13g2_nand2b_1 _2004_ (.Y(_0494_),
    .B(_0493_),
    .A_N(net1004));
 sg13g2_mux4_1 _2005_ (.S0(net997),
    .A0(\Inst_RegFile_32x4.mem[4][0] ),
    .A1(\Inst_RegFile_32x4.mem[5][0] ),
    .A2(\Inst_RegFile_32x4.mem[6][0] ),
    .A3(\Inst_RegFile_32x4.mem[7][0] ),
    .S1(net947),
    .X(_0495_));
 sg13g2_a21oi_1 _2006_ (.A1(net1007),
    .A2(_0495_),
    .Y(_0496_),
    .B1(_0460_));
 sg13g2_a22oi_1 _2007_ (.Y(_0497_),
    .B1(_0494_),
    .B2(_0496_),
    .A2(_0462_),
    .A1(_0460_));
 sg13g2_nor2b_1 _2008_ (.A(net996),
    .B_N(\Inst_RegFile_32x4.mem[24][0] ),
    .Y(_0498_));
 sg13g2_a21oi_1 _2009_ (.A1(\Inst_RegFile_32x4.mem[25][0] ),
    .A2(net993),
    .Y(_0499_),
    .B1(_0498_));
 sg13g2_mux2_1 _2010_ (.A0(\Inst_RegFile_32x4.mem[26][0] ),
    .A1(\Inst_RegFile_32x4.mem[27][0] ),
    .S(net998),
    .X(_0500_));
 sg13g2_a21oi_1 _2011_ (.A1(net1036),
    .A2(_0499_),
    .Y(_0501_),
    .B1(net1009));
 sg13g2_o21ai_1 _2012_ (.B1(_0501_),
    .Y(_0502_),
    .A1(net1036),
    .A2(_0500_));
 sg13g2_mux4_1 _2013_ (.S0(net992),
    .A0(\Inst_RegFile_32x4.mem[28][0] ),
    .A1(\Inst_RegFile_32x4.mem[29][0] ),
    .A2(\Inst_RegFile_32x4.mem[30][0] ),
    .A3(\Inst_RegFile_32x4.mem[31][0] ),
    .S1(net946),
    .X(_0503_));
 sg13g2_a21oi_2 _2014_ (.B1(_0459_),
    .Y(_0504_),
    .A2(_0503_),
    .A1(net1004));
 sg13g2_mux4_1 _2015_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[16][0] ),
    .A1(\Inst_RegFile_32x4.mem[17][0] ),
    .A2(\Inst_RegFile_32x4.mem[18][0] ),
    .A3(\Inst_RegFile_32x4.mem[19][0] ),
    .S1(net945),
    .X(_0505_));
 sg13g2_nand2b_1 _2016_ (.Y(_0506_),
    .B(_0505_),
    .A_N(net1005));
 sg13g2_mux4_1 _2017_ (.S0(net992),
    .A0(\Inst_RegFile_32x4.mem[20][0] ),
    .A1(\Inst_RegFile_32x4.mem[21][0] ),
    .A2(\Inst_RegFile_32x4.mem[22][0] ),
    .A3(\Inst_RegFile_32x4.mem[23][0] ),
    .S1(net945),
    .X(_0507_));
 sg13g2_a21oi_1 _2018_ (.A1(net1005),
    .A2(_0507_),
    .Y(_0508_),
    .B1(net943));
 sg13g2_a221oi_1 _2019_ (.B2(_0508_),
    .C1(_0491_),
    .B1(_0506_),
    .A1(_0502_),
    .Y(_0509_),
    .A2(_0504_));
 sg13g2_a21o_1 _2020_ (.A2(_0497_),
    .A1(_0491_),
    .B1(_0509_),
    .X(\Inst_RegFile_32x4.BD_comb[0] ));
 sg13g2_mux2_2 _2021_ (.A0(\Inst_RegFile_32x4.BD_comb[0] ),
    .A1(\Inst_RegFile_32x4.BD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD0));
 sg13g2_mux2_1 _2022_ (.A0(\Inst_RegFile_32x4.mem[24][1] ),
    .A1(\Inst_RegFile_32x4.mem[25][1] ),
    .S(net993),
    .X(_0510_));
 sg13g2_nand2b_1 _2023_ (.Y(_0511_),
    .B(net998),
    .A_N(\Inst_RegFile_32x4.mem[27][1] ));
 sg13g2_o21ai_1 _2024_ (.B1(_0511_),
    .Y(_0512_),
    .A1(\Inst_RegFile_32x4.mem[26][1] ),
    .A2(net998));
 sg13g2_a21oi_1 _2025_ (.A1(net948),
    .A2(_0512_),
    .Y(_0513_),
    .B1(net1009));
 sg13g2_o21ai_1 _2026_ (.B1(_0513_),
    .Y(_0514_),
    .A1(net948),
    .A2(_0510_));
 sg13g2_mux4_1 _2027_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[28][1] ),
    .A1(\Inst_RegFile_32x4.mem[29][1] ),
    .A2(\Inst_RegFile_32x4.mem[30][1] ),
    .A3(\Inst_RegFile_32x4.mem[31][1] ),
    .S1(net944),
    .X(_0515_));
 sg13g2_a21oi_2 _2028_ (.B1(_0459_),
    .Y(_0516_),
    .A2(_0515_),
    .A1(net1004));
 sg13g2_nand2_2 _2029_ (.Y(_0517_),
    .A(_0514_),
    .B(_0516_));
 sg13g2_mux4_1 _2030_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[16][1] ),
    .A1(\Inst_RegFile_32x4.mem[17][1] ),
    .A2(\Inst_RegFile_32x4.mem[18][1] ),
    .A3(\Inst_RegFile_32x4.mem[19][1] ),
    .S1(net945),
    .X(_0518_));
 sg13g2_nand2b_1 _2031_ (.Y(_0519_),
    .B(_0518_),
    .A_N(net1005));
 sg13g2_mux4_1 _2032_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[20][1] ),
    .A1(\Inst_RegFile_32x4.mem[21][1] ),
    .A2(\Inst_RegFile_32x4.mem[22][1] ),
    .A3(\Inst_RegFile_32x4.mem[23][1] ),
    .S1(net945),
    .X(_0520_));
 sg13g2_a21oi_1 _2033_ (.A1(net1007),
    .A2(_0520_),
    .Y(_0521_),
    .B1(net943));
 sg13g2_a21oi_2 _2034_ (.B1(net532),
    .Y(_0522_),
    .A2(_0521_),
    .A1(_0519_));
 sg13g2_mux4_1 _2035_ (.S0(net995),
    .A0(\Inst_RegFile_32x4.mem[8][1] ),
    .A1(\Inst_RegFile_32x4.mem[9][1] ),
    .A2(\Inst_RegFile_32x4.mem[10][1] ),
    .A3(\Inst_RegFile_32x4.mem[11][1] ),
    .S1(net947),
    .X(_0523_));
 sg13g2_nand2b_1 _2036_ (.Y(_0524_),
    .B(_0523_),
    .A_N(net1008));
 sg13g2_mux4_1 _2037_ (.S0(net992),
    .A0(\Inst_RegFile_32x4.mem[12][1] ),
    .A1(\Inst_RegFile_32x4.mem[13][1] ),
    .A2(\Inst_RegFile_32x4.mem[14][1] ),
    .A3(\Inst_RegFile_32x4.mem[15][1] ),
    .S1(net946),
    .X(_0525_));
 sg13g2_a21oi_1 _2038_ (.A1(net1006),
    .A2(_0525_),
    .Y(_0526_),
    .B1(_0459_));
 sg13g2_mux4_1 _2039_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[0][1] ),
    .A1(\Inst_RegFile_32x4.mem[1][1] ),
    .A2(\Inst_RegFile_32x4.mem[2][1] ),
    .A3(\Inst_RegFile_32x4.mem[3][1] ),
    .S1(net944),
    .X(_0527_));
 sg13g2_nand2b_1 _2040_ (.Y(_0528_),
    .B(_0527_),
    .A_N(net1006));
 sg13g2_mux4_1 _2041_ (.S0(net998),
    .A0(\Inst_RegFile_32x4.mem[4][1] ),
    .A1(\Inst_RegFile_32x4.mem[5][1] ),
    .A2(\Inst_RegFile_32x4.mem[6][1] ),
    .A3(\Inst_RegFile_32x4.mem[7][1] ),
    .S1(net948),
    .X(_0529_));
 sg13g2_a21oi_1 _2042_ (.A1(net1006),
    .A2(_0529_),
    .Y(_0530_),
    .B1(net943));
 sg13g2_a221oi_1 _2043_ (.B2(_0530_),
    .C1(_0492_),
    .B1(_0528_),
    .A1(_0524_),
    .Y(_0531_),
    .A2(_0526_));
 sg13g2_a21o_1 _2044_ (.A2(_0517_),
    .A1(_0522_),
    .B1(_0531_),
    .X(\Inst_RegFile_32x4.BD_comb[1] ));
 sg13g2_mux2_2 _2045_ (.A0(\Inst_RegFile_32x4.BD_comb[1] ),
    .A1(\Inst_RegFile_32x4.BD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD1));
 sg13g2_nor2b_1 _2046_ (.A(net993),
    .B_N(\Inst_RegFile_32x4.mem[24][3] ),
    .Y(_0532_));
 sg13g2_a21oi_1 _2047_ (.A1(\Inst_RegFile_32x4.mem[25][3] ),
    .A2(net993),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_mux2_1 _2048_ (.A0(\Inst_RegFile_32x4.mem[26][3] ),
    .A1(\Inst_RegFile_32x4.mem[27][3] ),
    .S(net993),
    .X(_0534_));
 sg13g2_a21oi_1 _2049_ (.A1(net1036),
    .A2(_0533_),
    .Y(_0535_),
    .B1(net1008));
 sg13g2_o21ai_1 _2050_ (.B1(_0535_),
    .Y(_0536_),
    .A1(net1036),
    .A2(_0534_));
 sg13g2_mux4_1 _2051_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[28][3] ),
    .A1(\Inst_RegFile_32x4.mem[29][3] ),
    .A2(\Inst_RegFile_32x4.mem[30][3] ),
    .A3(\Inst_RegFile_32x4.mem[31][3] ),
    .S1(net944),
    .X(_0537_));
 sg13g2_a21oi_1 _2052_ (.A1(net1004),
    .A2(_0537_),
    .Y(_0538_),
    .B1(_0459_));
 sg13g2_mux4_1 _2053_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[16][3] ),
    .A1(\Inst_RegFile_32x4.mem[17][3] ),
    .A2(\Inst_RegFile_32x4.mem[18][3] ),
    .A3(\Inst_RegFile_32x4.mem[19][3] ),
    .S1(net944),
    .X(_0539_));
 sg13g2_nand2b_1 _2054_ (.Y(_0540_),
    .B(_0539_),
    .A_N(net1005));
 sg13g2_mux4_1 _2055_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[20][3] ),
    .A1(\Inst_RegFile_32x4.mem[21][3] ),
    .A2(\Inst_RegFile_32x4.mem[22][3] ),
    .A3(\Inst_RegFile_32x4.mem[23][3] ),
    .S1(net945),
    .X(_0541_));
 sg13g2_a21oi_2 _2056_ (.B1(net943),
    .Y(_0542_),
    .A2(_0541_),
    .A1(net1005));
 sg13g2_a221oi_1 _2057_ (.B2(_0540_),
    .C1(net519),
    .B1(_0542_),
    .A1(_0536_),
    .Y(_0543_),
    .A2(_0538_));
 sg13g2_nor2b_1 _2058_ (.A(net994),
    .B_N(\Inst_RegFile_32x4.mem[10][3] ),
    .Y(_0544_));
 sg13g2_a21oi_1 _2059_ (.A1(\Inst_RegFile_32x4.mem[11][3] ),
    .A2(net994),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_nand2_1 _2060_ (.Y(_0546_),
    .A(net947),
    .B(_0545_));
 sg13g2_nor2b_1 _2061_ (.A(net995),
    .B_N(\Inst_RegFile_32x4.mem[8][3] ),
    .Y(_0547_));
 sg13g2_a21oi_1 _2062_ (.A1(\Inst_RegFile_32x4.mem[9][3] ),
    .A2(net995),
    .Y(_0548_),
    .B1(_0547_));
 sg13g2_a21oi_1 _2063_ (.A1(net1036),
    .A2(_0548_),
    .Y(_0549_),
    .B1(net1008));
 sg13g2_mux4_1 _2064_ (.S0(net997),
    .A0(\Inst_RegFile_32x4.mem[12][3] ),
    .A1(\Inst_RegFile_32x4.mem[13][3] ),
    .A2(\Inst_RegFile_32x4.mem[14][3] ),
    .A3(\Inst_RegFile_32x4.mem[15][3] ),
    .S1(net947),
    .X(_0550_));
 sg13g2_a22oi_1 _2065_ (.Y(_0551_),
    .B1(_0550_),
    .B2(net1008),
    .A2(_0549_),
    .A1(_0546_));
 sg13g2_mux4_1 _2066_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[0][3] ),
    .A1(\Inst_RegFile_32x4.mem[1][3] ),
    .A2(\Inst_RegFile_32x4.mem[2][3] ),
    .A3(\Inst_RegFile_32x4.mem[3][3] ),
    .S1(net944),
    .X(_0552_));
 sg13g2_nand2b_1 _2067_ (.Y(_0553_),
    .B(_0552_),
    .A_N(net1004));
 sg13g2_mux4_1 _2068_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[4][3] ),
    .A1(\Inst_RegFile_32x4.mem[5][3] ),
    .A2(\Inst_RegFile_32x4.mem[6][3] ),
    .A3(\Inst_RegFile_32x4.mem[7][3] ),
    .S1(net947),
    .X(_0554_));
 sg13g2_a21oi_1 _2069_ (.A1(net1006),
    .A2(_0554_),
    .Y(_0555_),
    .B1(net943));
 sg13g2_a22oi_1 _2070_ (.Y(_0556_),
    .B1(_0553_),
    .B2(_0555_),
    .A2(_0551_),
    .A1(_0460_));
 sg13g2_a21o_1 _2071_ (.A2(_0556_),
    .A1(net519),
    .B1(_0543_),
    .X(\Inst_RegFile_32x4.BD_comb[3] ));
 sg13g2_mux2_2 _2072_ (.A0(\Inst_RegFile_32x4.BD_comb[3] ),
    .A1(\Inst_RegFile_32x4.BD_reg[3] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD3));
 sg13g2_nor2b_1 _2073_ (.A(net993),
    .B_N(\Inst_RegFile_32x4.mem[24][2] ),
    .Y(_0557_));
 sg13g2_a21oi_1 _2074_ (.A1(\Inst_RegFile_32x4.mem[25][2] ),
    .A2(net993),
    .Y(_0558_),
    .B1(_0557_));
 sg13g2_mux2_1 _2075_ (.A0(\Inst_RegFile_32x4.mem[26][2] ),
    .A1(\Inst_RegFile_32x4.mem[27][2] ),
    .S(net993),
    .X(_0559_));
 sg13g2_a21oi_1 _2076_ (.A1(net1036),
    .A2(_0558_),
    .Y(_0560_),
    .B1(net1008));
 sg13g2_o21ai_1 _2077_ (.B1(_0560_),
    .Y(_0561_),
    .A1(net1036),
    .A2(_0559_));
 sg13g2_mux4_1 _2078_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[28][2] ),
    .A1(\Inst_RegFile_32x4.mem[29][2] ),
    .A2(\Inst_RegFile_32x4.mem[30][2] ),
    .A3(\Inst_RegFile_32x4.mem[31][2] ),
    .S1(net944),
    .X(_0562_));
 sg13g2_a21oi_2 _2079_ (.B1(_0459_),
    .Y(_0563_),
    .A2(_0562_),
    .A1(net1004));
 sg13g2_mux4_1 _2080_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[16][2] ),
    .A1(\Inst_RegFile_32x4.mem[17][2] ),
    .A2(\Inst_RegFile_32x4.mem[18][2] ),
    .A3(\Inst_RegFile_32x4.mem[19][2] ),
    .S1(net945),
    .X(_0564_));
 sg13g2_nand2b_1 _2081_ (.Y(_0565_),
    .B(_0564_),
    .A_N(net1005));
 sg13g2_mux4_1 _2082_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[20][2] ),
    .A1(\Inst_RegFile_32x4.mem[21][2] ),
    .A2(\Inst_RegFile_32x4.mem[22][2] ),
    .A3(\Inst_RegFile_32x4.mem[23][2] ),
    .S1(net945),
    .X(_0566_));
 sg13g2_a21oi_1 _2083_ (.A1(net1004),
    .A2(_0566_),
    .Y(_0567_),
    .B1(net943));
 sg13g2_a221oi_1 _2084_ (.B2(_0567_),
    .C1(net532),
    .B1(_0565_),
    .A1(_0561_),
    .Y(_0568_),
    .A2(_0563_));
 sg13g2_nor2b_1 _2085_ (.A(net994),
    .B_N(\Inst_RegFile_32x4.mem[10][2] ),
    .Y(_0569_));
 sg13g2_a21oi_1 _2086_ (.A1(\Inst_RegFile_32x4.mem[11][2] ),
    .A2(net994),
    .Y(_0570_),
    .B1(_0569_));
 sg13g2_nand2_1 _2087_ (.Y(_0571_),
    .A(net947),
    .B(_0570_));
 sg13g2_nor2b_1 _2088_ (.A(net994),
    .B_N(\Inst_RegFile_32x4.mem[8][2] ),
    .Y(_0572_));
 sg13g2_a21oi_1 _2089_ (.A1(\Inst_RegFile_32x4.mem[9][2] ),
    .A2(net994),
    .Y(_0573_),
    .B1(_0572_));
 sg13g2_a21oi_1 _2090_ (.A1(net1036),
    .A2(_0573_),
    .Y(_0574_),
    .B1(net1008));
 sg13g2_mux4_1 _2091_ (.S0(net997),
    .A0(\Inst_RegFile_32x4.mem[12][2] ),
    .A1(\Inst_RegFile_32x4.mem[13][2] ),
    .A2(\Inst_RegFile_32x4.mem[14][2] ),
    .A3(\Inst_RegFile_32x4.mem[15][2] ),
    .S1(net947),
    .X(_0575_));
 sg13g2_a22oi_1 _2092_ (.Y(_0576_),
    .B1(_0575_),
    .B2(net1008),
    .A2(_0574_),
    .A1(_0571_));
 sg13g2_mux4_1 _2093_ (.S0(net990),
    .A0(\Inst_RegFile_32x4.mem[0][2] ),
    .A1(\Inst_RegFile_32x4.mem[1][2] ),
    .A2(\Inst_RegFile_32x4.mem[2][2] ),
    .A3(\Inst_RegFile_32x4.mem[3][2] ),
    .S1(net944),
    .X(_0577_));
 sg13g2_nand2b_1 _2094_ (.Y(_0578_),
    .B(_0577_),
    .A_N(net1004));
 sg13g2_mux4_1 _2095_ (.S0(net991),
    .A0(\Inst_RegFile_32x4.mem[4][2] ),
    .A1(\Inst_RegFile_32x4.mem[5][2] ),
    .A2(\Inst_RegFile_32x4.mem[6][2] ),
    .A3(\Inst_RegFile_32x4.mem[7][2] ),
    .S1(net945),
    .X(_0579_));
 sg13g2_a21oi_1 _2096_ (.A1(net1007),
    .A2(_0579_),
    .Y(_0580_),
    .B1(net943));
 sg13g2_a22oi_1 _2097_ (.Y(_0581_),
    .B1(_0578_),
    .B2(_0580_),
    .A2(_0576_),
    .A1(net943));
 sg13g2_a21o_1 _2098_ (.A2(_0581_),
    .A1(net532),
    .B1(_0568_),
    .X(\Inst_RegFile_32x4.BD_comb[2] ));
 sg13g2_mux2_1 _2099_ (.A0(\Inst_RegFile_32x4.BD_comb[2] ),
    .A1(\Inst_RegFile_32x4.BD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .X(BD2));
 sg13g2_o21ai_1 _2100_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .Y(_0582_),
    .A1(net1055),
    .A2(net986));
 sg13g2_a21o_1 _2101_ (.A2(_1165_),
    .A1(net1055),
    .B1(_0582_),
    .X(_0583_));
 sg13g2_a21oi_1 _2102_ (.A1(net1055),
    .A2(net1011),
    .Y(_0584_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_o21ai_1 _2103_ (.B1(_0584_),
    .Y(_0585_),
    .A1(net1055),
    .A2(net971));
 sg13g2_nand3_1 _2104_ (.B(_0583_),
    .C(_0585_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .Y(_0586_));
 sg13g2_nand2_1 _2105_ (.Y(_0587_),
    .A(net1055),
    .B(net719));
 sg13g2_o21ai_1 _2106_ (.B1(_0587_),
    .Y(_0588_),
    .A1(net1055),
    .A2(net977));
 sg13g2_nor2b_1 _2107_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .B_N(net1068),
    .Y(_0589_));
 sg13g2_a21oi_1 _2108_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(net1017),
    .Y(_0590_),
    .B1(_0589_));
 sg13g2_a21oi_1 _2109_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .A2(_0588_),
    .Y(_0591_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_o21ai_1 _2110_ (.B1(_0591_),
    .Y(_0592_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .A2(_0590_));
 sg13g2_nand3_1 _2111_ (.B(_0586_),
    .C(_0592_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .Y(_0593_));
 sg13g2_mux4_1 _2112_ (.S0(net1055),
    .A0(net10),
    .A1(net59),
    .A2(net67),
    .A3(net1071),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0594_));
 sg13g2_mux4_1 _2113_ (.S0(net1055),
    .A0(net1075),
    .A1(net39),
    .A2(net57),
    .A3(net1220),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .X(_0595_));
 sg13g2_nor2b_1 _2114_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .B_N(_0595_),
    .Y(_0596_));
 sg13g2_a21oi_2 _2115_ (.B1(_0596_),
    .Y(_0597_),
    .A2(_0594_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_o21ai_1 _2116_ (.B1(_0593_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .A1(_0597_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_mux2_1 _2117_ (.A0(net81),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .X(_0598_));
 sg13g2_nor2b_1 _2118_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .B_N(net53),
    .Y(_0599_));
 sg13g2_a21oi_1 _2119_ (.A1(net21),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .Y(_0600_),
    .B1(_0599_));
 sg13g2_o21ai_1 _2120_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_0601_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_0600_));
 sg13g2_a21oi_2 _2121_ (.B1(_0601_),
    .Y(_0602_),
    .A2(_0598_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_mux4_1 _2122_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(net41),
    .A1(net12),
    .A2(net69),
    .A3(net106),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ),
    .X(_0603_));
 sg13g2_o21ai_1 _2123_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .Y(_0604_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0603_));
 sg13g2_mux2_1 _2124_ (.A0(net76),
    .A1(net510),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .X(_0605_));
 sg13g2_nand2b_1 _2125_ (.Y(_0606_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .A_N(net19));
 sg13g2_nor2_1 _2126_ (.A(net48),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0607_));
 sg13g2_nor2_1 _2127_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .B(_0607_),
    .Y(_0608_));
 sg13g2_a221oi_1 _2128_ (.B2(_0608_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .B1(_0606_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .Y(_0609_),
    .A2(_0605_));
 sg13g2_nand2b_1 _2129_ (.Y(_0610_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ),
    .A_N(net20));
 sg13g2_o21ai_1 _2130_ (.B1(_0610_),
    .Y(_0611_),
    .A1(net49),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_mux2_1 _2131_ (.A0(net77),
    .A1(net104),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ),
    .X(_0612_));
 sg13g2_o21ai_1 _2132_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .Y(_0613_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_0611_));
 sg13g2_a21oi_1 _2133_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ),
    .A2(_0612_),
    .Y(_0614_),
    .B1(_0613_));
 sg13g2_or3_1 _2134_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .B(_0609_),
    .C(_0614_),
    .X(_0615_));
 sg13g2_o21ai_1 _2135_ (.B1(_0615_),
    .Y(B_ADR0),
    .A1(_0604_),
    .A2(_0602_));
 sg13g2_nand2_1 _2136_ (.Y(_0616_),
    .A(net1057),
    .B(net963));
 sg13g2_o21ai_1 _2137_ (.B1(_0616_),
    .Y(_0617_),
    .A1(net1056),
    .A2(net976));
 sg13g2_nor2b_1 _2138_ (.A(net1056),
    .B_N(net1066),
    .Y(_0618_));
 sg13g2_a21oi_1 _2139_ (.A1(net1056),
    .A2(net1018),
    .Y(_0619_),
    .B1(_0618_));
 sg13g2_a21oi_1 _2140_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0617_),
    .Y(_0620_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_o21ai_1 _2141_ (.B1(_0620_),
    .Y(_0621_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0619_));
 sg13g2_nor2b_1 _2142_ (.A(net1056),
    .B_N(net1029),
    .Y(_0622_));
 sg13g2_a21oi_1 _2143_ (.A1(net1056),
    .A2(net1012),
    .Y(_0623_),
    .B1(_0622_));
 sg13g2_mux2_1 _2144_ (.A0(net985),
    .A1(net1001),
    .S(net1056),
    .X(_0624_));
 sg13g2_o21ai_1 _2145_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .Y(_0625_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0623_));
 sg13g2_a21oi_2 _2146_ (.B1(_0625_),
    .Y(_0626_),
    .A2(_0624_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_nand2_1 _2147_ (.Y(_0627_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ),
    .B(_0621_));
 sg13g2_nor2b_1 _2148_ (.A(net1056),
    .B_N(net1216),
    .Y(_0628_));
 sg13g2_a21oi_1 _2149_ (.A1(net66),
    .A2(net1057),
    .Y(_0629_),
    .B1(_0628_));
 sg13g2_mux2_1 _2150_ (.A0(net93),
    .A1(net109),
    .S(net1057),
    .X(_0630_));
 sg13g2_o21ai_1 _2151_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .Y(_0631_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0629_));
 sg13g2_a21oi_1 _2152_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .A2(_0630_),
    .Y(_0632_),
    .B1(_0631_));
 sg13g2_mux4_1 _2153_ (.S0(net1056),
    .A0(net38),
    .A1(net50),
    .A2(net1219),
    .A3(net9),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .X(_0633_));
 sg13g2_nor2_1 _2154_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ),
    .B(_0632_),
    .Y(_0634_));
 sg13g2_o21ai_1 _2155_ (.B1(_0634_),
    .Y(_0635_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .A2(_0633_));
 sg13g2_o21ai_1 _2156_ (.B1(_0635_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .A1(_0627_),
    .A2(_0626_));
 sg13g2_mux2_1 _2157_ (.A0(net92),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ),
    .X(_0636_));
 sg13g2_nor2b_1 _2158_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ),
    .B_N(net53),
    .Y(_0637_));
 sg13g2_a21oi_1 _2159_ (.A1(net8),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ),
    .Y(_0638_),
    .B1(_0637_));
 sg13g2_o21ai_1 _2160_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .Y(_0639_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ),
    .A2(_0638_));
 sg13g2_a21o_1 _2161_ (.A2(_0636_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ),
    .B1(_0639_),
    .X(_0640_));
 sg13g2_mux4_1 _2162_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ),
    .A0(net41),
    .A1(net69),
    .A2(net23),
    .A3(net96),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ),
    .X(_0641_));
 sg13g2_o21ai_1 _2163_ (.B1(_0640_),
    .Y(_0642_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_0641_));
 sg13g2_mux4_1 _2164_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(net48),
    .A1(net19),
    .A2(net103),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ),
    .X(_0643_));
 sg13g2_nand2b_1 _2165_ (.Y(_0644_),
    .B(_0643_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_mux4_1 _2166_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ),
    .A0(net49),
    .A1(net20),
    .A2(net77),
    .A3(net104),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_0645_));
 sg13g2_a21oi_1 _2167_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_0645_),
    .Y(_0646_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_a22oi_1 _2168_ (.Y(A_ADR0),
    .B1(_0644_),
    .B2(_0646_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ),
    .A1(_0642_));
 sg13g2_mux4_1 _2169_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(net105),
    .A1(net1017),
    .A2(net978),
    .A3(net971),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0647_));
 sg13g2_nand2b_1 _2170_ (.Y(_0648_),
    .B(_1147_),
    .A_N(_0647_));
 sg13g2_nor2b_1 _2171_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .B_N(net1031),
    .Y(_0649_));
 sg13g2_a21oi_1 _2172_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(net1013),
    .Y(_0650_),
    .B1(_0649_));
 sg13g2_mux2_1 _2173_ (.A0(net986),
    .A1(net1002),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0651_));
 sg13g2_a21oi_1 _2174_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0651_),
    .Y(_0652_),
    .B1(_1147_));
 sg13g2_o21ai_1 _2175_ (.B1(_0652_),
    .Y(_0653_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0650_));
 sg13g2_nand3_1 _2176_ (.B(_0648_),
    .C(_0653_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .Y(_0654_));
 sg13g2_mux4_1 _2177_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(net1075),
    .A1(net37),
    .A2(net56),
    .A3(net8),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0655_));
 sg13g2_mux2_1 _2178_ (.A0(net81),
    .A1(net92),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .X(_0656_));
 sg13g2_nor2b_1 _2179_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .B_N(net1215),
    .Y(_0657_));
 sg13g2_a21oi_1 _2180_ (.A1(net65),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .Y(_0658_),
    .B1(_0657_));
 sg13g2_a21oi_1 _2181_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0656_),
    .Y(_0659_),
    .B1(_1147_));
 sg13g2_o21ai_1 _2182_ (.B1(_0659_),
    .Y(_0660_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .A2(_0658_));
 sg13g2_o21ai_1 _2183_ (.B1(_0660_),
    .Y(_0661_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0655_));
 sg13g2_o21ai_1 _2184_ (.B1(_0654_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0661_));
 sg13g2_nor2b_1 _2185_ (.A(net1002),
    .B_N(net1044),
    .Y(_0662_));
 sg13g2_o21ai_1 _2186_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .Y(_0663_),
    .A1(net1044),
    .A2(net987));
 sg13g2_nand2_1 _2187_ (.Y(_0664_),
    .A(net1044),
    .B(net1013));
 sg13g2_nand2b_1 _2188_ (.Y(_0665_),
    .B(net1031),
    .A_N(net1044));
 sg13g2_a21oi_1 _2189_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_o21ai_1 _2190_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .Y(_0667_),
    .A1(_0662_),
    .A2(_0663_));
 sg13g2_nand2_1 _2191_ (.Y(_0668_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .B(net971));
 sg13g2_o21ai_1 _2192_ (.B1(_0668_),
    .Y(_0669_),
    .A1(net1044),
    .A2(net977));
 sg13g2_or2_1 _2193_ (.X(_0670_),
    .B(net1044),
    .A(net105));
 sg13g2_a21oi_1 _2194_ (.A1(net1044),
    .A2(net1016),
    .Y(_0671_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_a221oi_1 _2195_ (.B2(_0671_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .B1(_0670_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .Y(_0672_),
    .A2(_0669_));
 sg13g2_o21ai_1 _2196_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_0673_),
    .A1(_0666_),
    .A2(_0667_));
 sg13g2_mux4_1 _2197_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .A0(net37),
    .A1(net8),
    .A2(net1220),
    .A3(net23),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0674_));
 sg13g2_mux4_1 _2198_ (.S0(net1044),
    .A0(net1215),
    .A1(net65),
    .A2(net81),
    .A3(net92),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .X(_0675_));
 sg13g2_mux2_1 _2199_ (.A0(_0674_),
    .A1(_0675_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .X(_0676_));
 sg13g2_nand2b_1 _2200_ (.Y(_0677_),
    .B(_0676_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_o21ai_1 _2201_ (.B1(_0677_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .A1(_0673_),
    .A2(_0672_));
 sg13g2_o21ai_1 _2202_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .Y(_0678_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(net988));
 sg13g2_a21oi_1 _2203_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_1165_),
    .Y(_0679_),
    .B1(_0678_));
 sg13g2_nor2b_1 _2204_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .B_N(net1034),
    .Y(_0680_));
 sg13g2_a21oi_2 _2205_ (.B1(_0680_),
    .Y(_0681_),
    .A2(net1015),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_o21ai_1 _2206_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .Y(_0682_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0681_));
 sg13g2_mux4_1 _2207_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(net105),
    .A1(net1019),
    .A2(net980),
    .A3(net974),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0683_));
 sg13g2_nor2_1 _2208_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_o21ai_1 _2209_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .Y(_0685_),
    .A1(_0679_),
    .A2(_0682_));
 sg13g2_or2_1 _2210_ (.X(_0686_),
    .B(_0685_),
    .A(_0684_));
 sg13g2_mux4_1 _2211_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(net31),
    .A1(net37),
    .A2(net53),
    .A3(net8),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0687_));
 sg13g2_mux4_1 _2212_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .A0(net1215),
    .A1(net65),
    .A2(net84),
    .A3(net92),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .X(_0688_));
 sg13g2_nor2b_1 _2213_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .B_N(_0687_),
    .Y(_0689_));
 sg13g2_a21oi_1 _2214_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0688_),
    .Y(_0690_),
    .B1(_0689_));
 sg13g2_o21ai_1 _2215_ (.B1(_0686_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0690_));
 sg13g2_mux2_1 _2216_ (.A0(net988),
    .A1(BD3),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .X(_0691_));
 sg13g2_nor2b_1 _2217_ (.A(net1058),
    .B_N(net1033),
    .Y(_0692_));
 sg13g2_a21oi_2 _2218_ (.B1(_0692_),
    .Y(_0693_),
    .A2(net1015),
    .A1(net1058));
 sg13g2_o21ai_1 _2219_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .Y(_0694_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0693_));
 sg13g2_a21oi_2 _2220_ (.B1(_0694_),
    .Y(_0695_),
    .A2(_0691_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_mux2_1 _2221_ (.A0(net980),
    .A1(net974),
    .S(net1058),
    .X(_0696_));
 sg13g2_nor2b_1 _2222_ (.A(net1058),
    .B_N(net1065),
    .Y(_0697_));
 sg13g2_a21oi_1 _2223_ (.A1(net1058),
    .A2(net1019),
    .Y(_0698_),
    .B1(_0697_));
 sg13g2_a21oi_1 _2224_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0696_),
    .Y(_0699_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_o21ai_1 _2225_ (.B1(_0699_),
    .Y(_0700_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0698_));
 sg13g2_nand2_1 _2226_ (.Y(_0701_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .B(_0700_));
 sg13g2_mux4_1 _2227_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .A0(net37),
    .A1(net1220),
    .A2(net53),
    .A3(net8),
    .S1(net1058),
    .X(_0702_));
 sg13g2_mux2_1 _2228_ (.A0(net92),
    .A1(net108),
    .S(net1058),
    .X(_0703_));
 sg13g2_mux2_1 _2229_ (.A0(net1214),
    .A1(net65),
    .S(net1058),
    .X(_0704_));
 sg13g2_nand2b_1 _2230_ (.Y(_0705_),
    .B(_0704_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_a21oi_1 _2231_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .A2(_0703_),
    .Y(_0706_),
    .B1(_1148_));
 sg13g2_a21oi_1 _2232_ (.A1(_0705_),
    .A2(_0706_),
    .Y(_0707_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_o21ai_1 _2233_ (.B1(_0707_),
    .Y(_0708_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0702_));
 sg13g2_o21ai_1 _2234_ (.B1(_0708_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .A1(_0701_),
    .A2(_0695_));
 sg13g2_mux2_1 _2235_ (.A0(net963),
    .A1(net970),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_0709_));
 sg13g2_nor2b_1 _2236_ (.A(net1040),
    .B_N(net1066),
    .Y(_0710_));
 sg13g2_a21oi_1 _2237_ (.A1(net1040),
    .A2(net1018),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_a21oi_1 _2238_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0709_),
    .Y(_0712_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_o21ai_1 _2239_ (.B1(_0712_),
    .Y(_0713_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0711_));
 sg13g2_o21ai_1 _2240_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0714_),
    .A1(net1040),
    .A2(net984));
 sg13g2_a21o_1 _2241_ (.A2(net999),
    .A1(net1040),
    .B1(_0714_),
    .X(_0715_));
 sg13g2_a21oi_2 _2242_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0716_),
    .A2(net1010),
    .A1(net1040));
 sg13g2_o21ai_1 _2243_ (.B1(_0716_),
    .Y(_0717_),
    .A1(net1040),
    .A2(net1029));
 sg13g2_nand3_1 _2244_ (.B(_0717_),
    .C(_0715_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0718_));
 sg13g2_nand3_1 _2245_ (.B(_0713_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .A(_0718_),
    .Y(_0719_));
 sg13g2_mux4_1 _2246_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .A0(net1076),
    .A1(net7),
    .A2(net36),
    .A3(net1216),
    .S1(net1040),
    .X(_0720_));
 sg13g2_mux4_1 _2247_ (.S0(net1040),
    .A0(net64),
    .A1(net80),
    .A2(net83),
    .A3(net91),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0721_));
 sg13g2_nor2b_1 _2248_ (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .B_N(_0720_),
    .Y(_0722_));
 sg13g2_a21oi_1 _2249_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0721_),
    .Y(_0723_),
    .B1(_0722_));
 sg13g2_o21ai_1 _2250_ (.B1(_0719_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0723_));
 sg13g2_mux2_1 _2251_ (.A0(net963),
    .A1(net970),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .X(_0724_));
 sg13g2_or2_1 _2252_ (.X(_0725_),
    .B(net1045),
    .A(net1066));
 sg13g2_a21oi_1 _2253_ (.A1(net1045),
    .A2(net1016),
    .Y(_0726_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_a221oi_1 _2254_ (.B2(_0726_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .B1(_0725_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .Y(_0727_),
    .A2(_0724_));
 sg13g2_o21ai_1 _2255_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .Y(_0728_),
    .A1(net1045),
    .A2(net984));
 sg13g2_a21oi_1 _2256_ (.A1(net1045),
    .A2(net999),
    .Y(_0729_),
    .B1(_0728_));
 sg13g2_a21oi_2 _2257_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .Y(_0730_),
    .A2(net1010),
    .A1(net1045));
 sg13g2_o21ai_1 _2258_ (.B1(_0730_),
    .Y(_0731_),
    .A1(net1045),
    .A2(net1029));
 sg13g2_nand2_2 _2259_ (.Y(_0732_),
    .A(_0731_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_o21ai_1 _2260_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0733_),
    .A1(_0732_),
    .A2(_0729_));
 sg13g2_mux4_1 _2261_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .A0(net36),
    .A1(net7),
    .A2(net1221),
    .A3(net1216),
    .S1(net1045),
    .X(_0734_));
 sg13g2_mux4_1 _2262_ (.S0(net1045),
    .A0(net64),
    .A1(net80),
    .A2(net91),
    .A3(net107),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0735_));
 sg13g2_inv_1 _2263_ (.Y(_0736_),
    .A(_0735_));
 sg13g2_a21oi_1 _2264_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0736_),
    .Y(_0737_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_o21ai_1 _2265_ (.B1(_0737_),
    .Y(_0738_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0734_));
 sg13g2_o21ai_1 _2266_ (.B1(_0738_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .A1(_0733_),
    .A2(_0727_));
 sg13g2_mux4_1 _2267_ (.S0(net1050),
    .A0(net1066),
    .A1(net1018),
    .A2(net504),
    .A3(net973),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .X(_0739_));
 sg13g2_or2_1 _2268_ (.X(_0740_),
    .B(_0739_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_a21oi_2 _2269_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_0741_),
    .A2(net1010),
    .A1(net1050));
 sg13g2_o21ai_1 _2270_ (.B1(_0741_),
    .Y(_0742_),
    .A1(net1050),
    .A2(net1030));
 sg13g2_o21ai_1 _2271_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .Y(_0743_),
    .A1(net1050),
    .A2(net985));
 sg13g2_a21o_1 _2272_ (.A2(net999),
    .A1(net1050),
    .B1(_0743_),
    .X(_0744_));
 sg13g2_nand3_1 _2273_ (.B(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .C(_0744_),
    .A(_0742_),
    .Y(_0745_));
 sg13g2_nand3_1 _2274_ (.B(_0740_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .A(_0745_),
    .Y(_0746_));
 sg13g2_nor2b_1 _2275_ (.A(net1049),
    .B_N(net7),
    .Y(_0747_));
 sg13g2_a21oi_1 _2276_ (.A1(net1216),
    .A2(net1049),
    .Y(_0748_),
    .B1(_0747_));
 sg13g2_nor2b_1 _2277_ (.A(net1049),
    .B_N(net64),
    .Y(_0749_));
 sg13g2_a21oi_1 _2278_ (.A1(net91),
    .A2(net1049),
    .Y(_0750_),
    .B1(_0749_));
 sg13g2_nor2b_1 _2279_ (.A(net1049),
    .B_N(net52),
    .Y(_0751_));
 sg13g2_a21oi_1 _2280_ (.A1(net55),
    .A2(net1049),
    .Y(_0752_),
    .B1(_0751_));
 sg13g2_nor2b_1 _2281_ (.A(net1049),
    .B_N(net1076),
    .Y(_0753_));
 sg13g2_a21oi_1 _2282_ (.A1(net36),
    .A2(net1049),
    .Y(_0754_),
    .B1(_0753_));
 sg13g2_mux4_1 _2283_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .A0(_0754_),
    .A1(_0752_),
    .A2(_0748_),
    .A3(_0750_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .X(_0755_));
 sg13g2_o21ai_1 _2284_ (.B1(_0746_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_0755_));
 sg13g2_mux2_1 _2285_ (.A0(net718),
    .A1(net970),
    .S(net1059),
    .X(_0756_));
 sg13g2_or2_1 _2286_ (.X(_0757_),
    .B(net1059),
    .A(net1066));
 sg13g2_a21oi_1 _2287_ (.A1(net1059),
    .A2(_1166_),
    .Y(_0758_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_a221oi_1 _2288_ (.B2(_0758_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .B1(_0757_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .Y(_0759_),
    .A2(_0756_));
 sg13g2_a21oi_2 _2289_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .Y(_0760_),
    .A2(net1011),
    .A1(net1059));
 sg13g2_o21ai_1 _2290_ (.B1(_0760_),
    .Y(_0761_),
    .A1(net1059),
    .A2(net1031));
 sg13g2_o21ai_1 _2291_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .Y(_0762_),
    .A1(net1059),
    .A2(net987));
 sg13g2_a21oi_1 _2292_ (.A1(net1059),
    .A2(net999),
    .Y(_0763_),
    .B1(_0762_));
 sg13g2_nand2_2 _2293_ (.Y(_0764_),
    .A(_0761_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_o21ai_1 _2294_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ),
    .Y(_0765_),
    .A1(_0764_),
    .A2(_0763_));
 sg13g2_mux4_1 _2295_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .A0(net36),
    .A1(net1221),
    .A2(net52),
    .A3(net7),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .X(_0766_));
 sg13g2_mux4_1 _2296_ (.S0(net1059),
    .A0(net22),
    .A1(net1217),
    .A2(net64),
    .A3(net91),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .X(_0767_));
 sg13g2_inv_1 _2297_ (.Y(_0768_),
    .A(_0767_));
 sg13g2_a21oi_1 _2298_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0768_),
    .Y(_0769_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_o21ai_1 _2299_ (.B1(_0769_),
    .Y(_0770_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .A2(_0766_));
 sg13g2_o21ai_1 _2300_ (.B1(_0770_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .A1(_0765_),
    .A2(_0759_));
 sg13g2_nand2_1 _2301_ (.Y(_0771_),
    .A(net1037),
    .B(net719));
 sg13g2_o21ai_1 _2302_ (.B1(_0771_),
    .Y(_0772_),
    .A1(net1037),
    .A2(net977));
 sg13g2_or2_1 _2303_ (.X(_0773_),
    .B(net1037),
    .A(net106));
 sg13g2_a21oi_1 _2304_ (.A1(net1037),
    .A2(net1016),
    .Y(_0774_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_a221oi_1 _2305_ (.B2(_0774_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .B1(_0773_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_0775_),
    .A2(_0772_));
 sg13g2_nand2_1 _2306_ (.Y(_0776_),
    .A(net1037),
    .B(net1031));
 sg13g2_nand2b_1 _2307_ (.Y(_0777_),
    .B(net971),
    .A_N(net1037));
 sg13g2_a21oi_1 _2308_ (.A1(_0776_),
    .A2(_0777_),
    .Y(_0778_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_nor2b_1 _2309_ (.A(net986),
    .B_N(net1037),
    .Y(_0779_));
 sg13g2_o21ai_1 _2310_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .Y(_0780_),
    .A1(net1037),
    .A2(net1013));
 sg13g2_o21ai_1 _2311_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .Y(_0781_),
    .A1(_0779_),
    .A2(_0780_));
 sg13g2_o21ai_1 _2312_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ),
    .Y(_0782_),
    .A1(_0778_),
    .A2(_0781_));
 sg13g2_mux4_1 _2313_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .A0(net58),
    .A1(net62),
    .A2(net60),
    .A3(net1072),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_0783_));
 sg13g2_mux4_1 _2314_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .A0(net1076),
    .A1(net1221),
    .A2(net34),
    .A3(net5),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(_0784_));
 sg13g2_mux2_1 _2315_ (.A0(_0784_),
    .A1(_0783_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .X(_0785_));
 sg13g2_nand2b_1 _2316_ (.Y(_0786_),
    .B(_0785_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_o21ai_1 _2317_ (.B1(_0786_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .A1(_0775_),
    .A2(_0782_));
 sg13g2_mux2_1 _2318_ (.A0(net963),
    .A1(net970),
    .S(net1041),
    .X(_0787_));
 sg13g2_or2_1 _2319_ (.X(_0788_),
    .B(net1041),
    .A(net1065));
 sg13g2_a21oi_1 _2320_ (.A1(net1041),
    .A2(net976),
    .Y(_0789_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_a221oi_1 _2321_ (.B2(_0789_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .B1(_0788_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0790_),
    .A2(_0787_));
 sg13g2_a21oi_2 _2322_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0791_),
    .A2(net1010),
    .A1(net1041));
 sg13g2_o21ai_1 _2323_ (.B1(_0791_),
    .Y(_0792_),
    .A1(net1041),
    .A2(net1029));
 sg13g2_o21ai_1 _2324_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .Y(_0793_),
    .A1(net1041),
    .A2(net984));
 sg13g2_a21oi_1 _2325_ (.A1(net1041),
    .A2(net999),
    .Y(_0794_),
    .B1(_0793_));
 sg13g2_nand2_2 _2326_ (.Y(_0795_),
    .A(_0792_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_o21ai_1 _2327_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ),
    .Y(_0796_),
    .A1(_0795_),
    .A2(_0794_));
 sg13g2_mux4_1 _2328_ (.S0(net1041),
    .A0(net1073),
    .A1(net35),
    .A2(net6),
    .A3(net1214),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0797_));
 sg13g2_mux4_1 _2329_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(net63),
    .A1(net79),
    .A2(net82),
    .A3(net90),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .X(_0798_));
 sg13g2_inv_1 _2330_ (.Y(_0799_),
    .A(_0798_));
 sg13g2_a21oi_1 _2331_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_0799_),
    .Y(_0800_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_o21ai_1 _2332_ (.B1(_0800_),
    .Y(_0801_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .A2(_0797_));
 sg13g2_o21ai_1 _2333_ (.B1(_0801_),
    .Y(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .A1(_0796_),
    .A2(_0790_));
 sg13g2_nor2b_1 _2334_ (.A(net1042),
    .B_N(net1014),
    .Y(_0802_));
 sg13g2_a21oi_2 _2335_ (.B1(_0802_),
    .Y(_0803_),
    .A2(net987),
    .A1(net1042));
 sg13g2_mux2_1 _2336_ (.A0(net972),
    .A1(net1032),
    .S(net1042),
    .X(_0804_));
 sg13g2_a21oi_1 _2337_ (.A1(_1149_),
    .A2(_0804_),
    .Y(_0805_),
    .B1(_1150_));
 sg13g2_o21ai_1 _2338_ (.B1(_0805_),
    .Y(_0806_),
    .A1(_0803_),
    .A2(_1149_));
 sg13g2_mux2_1 _2339_ (.A0(net979),
    .A1(net966),
    .S(net1042),
    .X(_0807_));
 sg13g2_nor2b_1 _2340_ (.A(net1042),
    .B_N(net1070),
    .Y(_0808_));
 sg13g2_a21oi_1 _2341_ (.A1(net1042),
    .A2(net506),
    .Y(_0809_),
    .B1(_0808_));
 sg13g2_a21oi_1 _2342_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0807_),
    .Y(_0810_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_o21ai_1 _2343_ (.B1(_0810_),
    .Y(_0811_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0809_));
 sg13g2_nand3_1 _2344_ (.B(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ),
    .C(_0811_),
    .A(_0806_),
    .Y(_0812_));
 sg13g2_mux4_1 _2345_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(net1076),
    .A1(net1221),
    .A2(net34),
    .A3(net5),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0813_));
 sg13g2_mux2_1 _2346_ (.A0(net82),
    .A1(net1072),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_0814_));
 sg13g2_nor2b_1 _2347_ (.A(net1042),
    .B_N(net58),
    .Y(_0815_));
 sg13g2_a21oi_1 _2348_ (.A1(net62),
    .A2(net1042),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_a21oi_1 _2349_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0814_),
    .Y(_0817_),
    .B1(_1150_));
 sg13g2_o21ai_1 _2350_ (.B1(_0817_),
    .Y(_0818_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0816_));
 sg13g2_o21ai_1 _2351_ (.B1(_0818_),
    .Y(_0819_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .A2(_0813_));
 sg13g2_o21ai_1 _2352_ (.B1(_0812_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0819_));
 sg13g2_o21ai_1 _2353_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_0820_),
    .A1(net1046),
    .A2(net984));
 sg13g2_a21oi_1 _2354_ (.A1(net1046),
    .A2(net999),
    .Y(_0821_),
    .B1(_0820_));
 sg13g2_a21oi_2 _2355_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .Y(_0822_),
    .A2(net1010),
    .A1(net1046));
 sg13g2_o21ai_1 _2356_ (.B1(_0822_),
    .Y(_0823_),
    .A1(net1046),
    .A2(net1029));
 sg13g2_nand2_2 _2357_ (.Y(_0824_),
    .A(_0823_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_mux4_1 _2358_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .A0(net1065),
    .A1(net963),
    .A2(net979),
    .A3(net970),
    .S1(net1046),
    .X(_0825_));
 sg13g2_nor2_1 _2359_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_0825_),
    .Y(_0826_));
 sg13g2_o21ai_1 _2360_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .Y(_0827_),
    .A1(_0824_),
    .A2(_0821_));
 sg13g2_mux4_1 _2361_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .A0(net35),
    .A1(net6),
    .A2(net1218),
    .A3(net1214),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(_0828_));
 sg13g2_mux2_1 _2362_ (.A0(net90),
    .A1(net106),
    .S(net1046),
    .X(_0829_));
 sg13g2_nor2b_1 _2363_ (.A(net1046),
    .B_N(net63),
    .Y(_0830_));
 sg13g2_a21oi_1 _2364_ (.A1(net79),
    .A2(net1046),
    .Y(_0831_),
    .B1(_0830_));
 sg13g2_o21ai_1 _2365_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0832_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_0831_));
 sg13g2_a21oi_1 _2366_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_0829_),
    .Y(_0833_),
    .B1(_0832_));
 sg13g2_nor2_1 _2367_ (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .B(_0833_),
    .Y(_0834_));
 sg13g2_o21ai_1 _2368_ (.B1(_0834_),
    .Y(_0835_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0828_));
 sg13g2_o21ai_1 _2369_ (.B1(_0835_),
    .Y(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .A1(_0827_),
    .A2(_0826_));
 sg13g2_mux4_1 _2370_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(net1072),
    .A1(net1019),
    .A2(AD1),
    .A3(net967),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .X(_0836_));
 sg13g2_nand2_1 _2371_ (.Y(_0837_),
    .A(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .B(net988));
 sg13g2_o21ai_1 _2372_ (.B1(_0837_),
    .Y(_0838_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(net1011));
 sg13g2_nor2b_1 _2373_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .B_N(net974),
    .Y(_0839_));
 sg13g2_a21oi_1 _2374_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(net1033),
    .Y(_0840_),
    .B1(_0839_));
 sg13g2_o21ai_1 _2375_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .Y(_0841_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .A2(_0840_));
 sg13g2_a21oi_1 _2376_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .A2(_0838_),
    .Y(_0842_),
    .B1(_0841_));
 sg13g2_o21ai_1 _2377_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_0843_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0836_));
 sg13g2_mux4_1 _2378_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .A0(net30),
    .A1(net1221),
    .A2(net34),
    .A3(net5),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0844_));
 sg13g2_mux4_1 _2379_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .A0(net21),
    .A1(net60),
    .A2(net58),
    .A3(net62),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0845_));
 sg13g2_inv_1 _2380_ (.Y(_0846_),
    .A(_0845_));
 sg13g2_a21oi_1 _2381_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0846_),
    .Y(_0847_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_o21ai_1 _2382_ (.B1(_0847_),
    .Y(_0848_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0844_));
 sg13g2_o21ai_1 _2383_ (.B1(_0848_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG7 ),
    .A1(_0842_),
    .A2(_0843_));
 sg13g2_mux4_1 _2384_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .A0(net1065),
    .A1(net504),
    .A2(net979),
    .A3(net970),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0849_));
 sg13g2_nor2b_1 _2385_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .B_N(net1030),
    .Y(_0850_));
 sg13g2_a21oi_2 _2386_ (.B1(_0850_),
    .Y(_0851_),
    .A2(net1012),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_mux2_1 _2387_ (.A0(net984),
    .A1(net1001),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0852_));
 sg13g2_o21ai_1 _2388_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_0853_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0851_));
 sg13g2_a21oi_2 _2389_ (.B1(_0853_),
    .Y(_0854_),
    .A2(_0852_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_nor2b_1 _2390_ (.A(_0854_),
    .B_N(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .Y(_0855_));
 sg13g2_o21ai_1 _2391_ (.B1(_0855_),
    .Y(_0856_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_0849_));
 sg13g2_nor2b_1 _2392_ (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .B_N(net6),
    .Y(_0857_));
 sg13g2_a21oi_1 _2393_ (.A1(net1214),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .Y(_0858_),
    .B1(_0857_));
 sg13g2_mux2_1 _2394_ (.A0(net63),
    .A1(net90),
    .S(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .X(_0859_));
 sg13g2_o21ai_1 _2395_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .Y(_0860_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0858_));
 sg13g2_a21o_1 _2396_ (.A2(_0859_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .B1(_0860_),
    .X(_0861_));
 sg13g2_mux4_1 _2397_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(net1073),
    .A1(net35),
    .A2(net51),
    .A3(net54),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .X(_0862_));
 sg13g2_o21ai_1 _2398_ (.B1(_0861_),
    .Y(_0863_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_0862_));
 sg13g2_o21ai_1 _2399_ (.B1(_0856_),
    .Y(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0863_));
 sg13g2_nand2_1 _2400_ (.Y(_0864_),
    .A(net1051),
    .B(net986));
 sg13g2_o21ai_1 _2401_ (.B1(_0864_),
    .Y(_0865_),
    .A1(net1051),
    .A2(net1011));
 sg13g2_nor2b_1 _2402_ (.A(net1051),
    .B_N(net972),
    .Y(_0866_));
 sg13g2_a21oi_1 _2403_ (.A1(net1051),
    .A2(net1031),
    .Y(_0867_),
    .B1(_0866_));
 sg13g2_o21ai_1 _2404_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .Y(_0868_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0867_));
 sg13g2_a21oi_2 _2405_ (.B1(_0868_),
    .Y(_0869_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .A1(_0865_));
 sg13g2_mux4_1 _2406_ (.S0(net1051),
    .A0(net1070),
    .A1(net1017),
    .A2(net978),
    .A3(net719),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .X(_0870_));
 sg13g2_o21ai_1 _2407_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ),
    .Y(_0871_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .A2(_0870_));
 sg13g2_mux2_1 _2408_ (.A0(net5),
    .A1(net58),
    .S(net1051),
    .X(_0872_));
 sg13g2_mux2_1 _2409_ (.A0(net62),
    .A1(net1072),
    .S(net1051),
    .X(_0873_));
 sg13g2_mux2_1 _2410_ (.A0(net54),
    .A1(net1221),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .X(_0874_));
 sg13g2_mux2_1 _2411_ (.A0(net1076),
    .A1(net34),
    .S(net1051),
    .X(_0875_));
 sg13g2_mux4_1 _2412_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .A0(_0875_),
    .A1(_0874_),
    .A2(_0872_),
    .A3(_0873_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .X(_0876_));
 sg13g2_nand2b_1 _2413_ (.Y(_0877_),
    .B(_0876_),
    .A_N(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_o21ai_1 _2414_ (.B1(_0877_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .A1(_0871_),
    .A2(_0869_));
 sg13g2_mux2_1 _2415_ (.A0(net963),
    .A1(net970),
    .S(net1060),
    .X(_0878_));
 sg13g2_nor2b_1 _2416_ (.A(net1060),
    .B_N(net1065),
    .Y(_0879_));
 sg13g2_a21oi_1 _2417_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(net979),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_a21oi_1 _2418_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .A2(_0878_),
    .Y(_0881_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_o21ai_1 _2419_ (.B1(_0881_),
    .Y(_0882_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .A2(_0880_));
 sg13g2_a21oi_2 _2420_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_0883_),
    .A2(net1010),
    .A1(net1060));
 sg13g2_o21ai_1 _2421_ (.B1(_0883_),
    .Y(_0884_),
    .A1(net1060),
    .A2(net1029));
 sg13g2_o21ai_1 _2422_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .Y(_0885_),
    .A1(net1060),
    .A2(net984));
 sg13g2_a21o_1 _2423_ (.A2(net999),
    .A1(net1060),
    .B1(_0885_),
    .X(_0886_));
 sg13g2_nand3_1 _2424_ (.B(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .C(_0886_),
    .A(_0884_),
    .Y(_0887_));
 sg13g2_nand3_1 _2425_ (.B(_0882_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ),
    .A(_0887_),
    .Y(_0888_));
 sg13g2_mux4_1 _2426_ (.S0(net1060),
    .A0(net35),
    .A1(net51),
    .A2(net1218),
    .A3(net6),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0889_));
 sg13g2_mux4_1 _2427_ (.S0(net1060),
    .A0(net21),
    .A1(net1214),
    .A2(net63),
    .A3(net90),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .X(_0890_));
 sg13g2_nor2b_1 _2428_ (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .B_N(_0889_),
    .Y(_0891_));
 sg13g2_a21oi_1 _2429_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .A2(_0890_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_o21ai_1 _2430_ (.B1(_0888_),
    .Y(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ),
    .A2(_0892_));
 sg13g2_mux4_1 _2431_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A0(net56),
    .A1(net1219),
    .A2(net84),
    .A3(net1070),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0893_));
 sg13g2_mux4_1 _2432_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .A0(net1017),
    .A1(net718),
    .A2(net979),
    .A3(net971),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0894_));
 sg13g2_mux4_1 _2433_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ),
    .A0(net46),
    .A1(net74),
    .A2(net17),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_0895_));
 sg13g2_mux4_1 _2434_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ),
    .A0(net46),
    .A1(net101),
    .A2(net17),
    .A3(net503),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_0896_));
 sg13g2_mux4_1 _2435_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A0(_0896_),
    .A1(_0895_),
    .A2(net499),
    .A3(net500),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .X(_0897_));
 sg13g2_mux4_1 _2436_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .A0(net1031),
    .A1(net987),
    .A2(net1012),
    .A3(net1001),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .X(_0898_));
 sg13g2_mux4_1 _2437_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .A0(_0893_),
    .A1(_0894_),
    .A2(_0898_),
    .A3(_0897_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.W6BEG1 ));
 sg13g2_nand2b_1 _2438_ (.Y(_0899_),
    .B(net55),
    .A_N(net1062));
 sg13g2_a21oi_1 _2439_ (.A1(net4),
    .A2(net1062),
    .Y(_0900_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_nor2b_1 _2440_ (.A(net1062),
    .B_N(net83),
    .Y(_0901_));
 sg13g2_a21oi_1 _2441_ (.A1(net1068),
    .A2(net1061),
    .Y(_0902_),
    .B1(_0901_));
 sg13g2_a221oi_1 _2442_ (.B2(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .B1(_0902_),
    .A1(_0899_),
    .Y(_0903_),
    .A2(_0900_));
 sg13g2_nor2b_1 _2443_ (.A(net1061),
    .B_N(net719),
    .Y(_0904_));
 sg13g2_a21oi_1 _2444_ (.A1(net1061),
    .A2(net971),
    .Y(_0905_),
    .B1(_0904_));
 sg13g2_a21oi_1 _2445_ (.A1(net1061),
    .A2(net978),
    .Y(_0906_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_o21ai_1 _2446_ (.B1(_0906_),
    .Y(_0907_),
    .A1(net1061),
    .A2(net1016));
 sg13g2_a21oi_1 _2447_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_0905_),
    .Y(_0908_),
    .B1(_1151_));
 sg13g2_a21oi_1 _2448_ (.A1(_0907_),
    .A2(_0908_),
    .Y(_0909_),
    .B1(_0903_));
 sg13g2_mux4_1 _2449_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ),
    .A0(net45),
    .A1(net16),
    .A2(net73),
    .A3(net100),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ),
    .X(_0910_));
 sg13g2_mux4_1 _2450_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(net45),
    .A1(net16),
    .A2(net73),
    .A3(net100),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ),
    .X(_0911_));
 sg13g2_mux2_1 _2451_ (.A0(_0911_),
    .A1(_0910_),
    .S(net1061),
    .X(_0912_));
 sg13g2_o21ai_1 _2452_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .Y(_0913_),
    .A1(net1061),
    .A2(_1183_));
 sg13g2_a21oi_1 _2453_ (.A1(net1062),
    .A2(_0338_),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_nor2_1 _2454_ (.A(_1151_),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_o21ai_1 _2455_ (.B1(_0915_),
    .Y(_0916_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_0912_));
 sg13g2_mux4_1 _2456_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A0(net1031),
    .A1(net986),
    .A2(net1013),
    .A3(net1003),
    .S1(net1061),
    .X(_0917_));
 sg13g2_a21oi_1 _2457_ (.A1(_1151_),
    .A2(_0917_),
    .Y(_0918_),
    .B1(_1152_));
 sg13g2_a22oi_1 _2458_ (.Y(\Inst_RegFile_switch_matrix.W6BEG0 ),
    .B1(_0916_),
    .B2(_0918_),
    .A2(_0909_),
    .A1(_1152_));
 sg13g2_mux4_1 _2459_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(net38),
    .A1(net66),
    .A2(net21),
    .A3(net93),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ),
    .X(_0919_));
 sg13g2_mux4_1 _2460_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .A0(net1030),
    .A1(net499),
    .A2(net500),
    .A3(_0919_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_0920_));
 sg13g2_mux4_1 _2461_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .A0(net1075),
    .A1(net59),
    .A2(net1071),
    .A3(net1018),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .X(_0921_));
 sg13g2_mux2_1 _2462_ (.A0(_0921_),
    .A1(_0920_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG3 ));
 sg13g2_mux4_1 _2463_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(net38),
    .A1(net9),
    .A2(net84),
    .A3(net93),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ),
    .X(_0922_));
 sg13g2_o21ai_1 _2464_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .Y(_0923_),
    .A1(_1153_),
    .A2(_0922_));
 sg13g2_a21oi_1 _2465_ (.A1(_1153_),
    .A2(_0339_),
    .Y(_0924_),
    .B1(_0923_));
 sg13g2_nor2_1 _2466_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .B(_1165_),
    .Y(_0925_));
 sg13g2_a21oi_1 _2467_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_1182_),
    .Y(_0926_),
    .B1(_0925_));
 sg13g2_o21ai_1 _2468_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .Y(_0927_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_0926_));
 sg13g2_nor2_1 _2469_ (.A(_0924_),
    .B(_0927_),
    .Y(_0928_));
 sg13g2_mux4_1 _2470_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .A0(net1076),
    .A1(net58),
    .A2(net1072),
    .A3(net972),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .X(_0929_));
 sg13g2_nor2_1 _2471_ (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .B(_0929_),
    .Y(_0930_));
 sg13g2_nor2_1 _2472_ (.A(_0928_),
    .B(_0930_),
    .Y(\Inst_RegFile_switch_matrix.WW4BEG2 ));
 sg13g2_mux4_1 _2473_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .A0(net984),
    .A1(_0895_),
    .A2(_0896_),
    .A3(_0138_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .X(_0931_));
 sg13g2_mux4_1 _2474_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .A0(net1073),
    .A1(net61),
    .A2(net1069),
    .A3(net504),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .X(_0932_));
 sg13g2_mux2_1 _2475_ (.A0(_0932_),
    .A1(_0931_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG1 ));
 sg13g2_mux4_1 _2476_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .A0(net1013),
    .A1(_0910_),
    .A2(_0911_),
    .A3(_0408_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .X(_0933_));
 sg13g2_mux4_1 _2477_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .A0(net1074),
    .A1(net60),
    .A2(net1070),
    .A3(net978),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .X(_0934_));
 sg13g2_mux2_1 _2478_ (.A0(_0934_),
    .A1(_0933_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ),
    .X(\Inst_RegFile_switch_matrix.WW4BEG0 ));
 sg13g2_mux4_1 _2479_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ),
    .A0(net34),
    .A1(net62),
    .A2(net5),
    .A3(net109),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0935_));
 sg13g2_mux4_1 _2480_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .A0(net1034),
    .A1(net499),
    .A2(net500),
    .A3(_0935_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_0936_));
 sg13g2_mux4_1 _2481_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .A0(net31),
    .A1(net2),
    .A2(net1071),
    .A3(net1020),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .X(_0937_));
 sg13g2_mux2_1 _2482_ (.A0(_0937_),
    .A1(_0936_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG3 ));
 sg13g2_o21ai_1 _2483_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .Y(_0938_),
    .A1(_1154_),
    .A2(_0209_));
 sg13g2_a21oi_1 _2484_ (.A1(_1154_),
    .A2(_0339_),
    .Y(_0939_),
    .B1(_0938_));
 sg13g2_nor2_1 _2485_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .B(_1165_),
    .Y(_0940_));
 sg13g2_a21oi_1 _2486_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_1182_),
    .Y(_0941_),
    .B1(_0940_));
 sg13g2_o21ai_1 _2487_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .Y(_0942_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0941_));
 sg13g2_nor2_1 _2488_ (.A(_0939_),
    .B(_0942_),
    .Y(_0943_));
 sg13g2_mux4_1 _2489_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A0(net30),
    .A1(net1),
    .A2(net86),
    .A3(net974),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .X(_0944_));
 sg13g2_nor2_1 _2490_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .B(_0944_),
    .Y(_0945_));
 sg13g2_nor2_1 _2491_ (.A(_0943_),
    .B(_0945_),
    .Y(\Inst_RegFile_switch_matrix.SS4BEG2 ));
 sg13g2_mux4_1 _2492_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .A0(net985),
    .A1(_0895_),
    .A2(_0896_),
    .A3(_0165_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .X(_0946_));
 sg13g2_mux4_1 _2493_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .A0(net1073),
    .A1(net1218),
    .A2(net1069),
    .A3(net505),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .X(_0947_));
 sg13g2_mux2_2 _2494_ (.A0(_0947_),
    .A1(_0946_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ),
    .X(\Inst_RegFile_switch_matrix.SS4BEG1 ));
 sg13g2_a21oi_1 _2495_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .A2(_0432_),
    .Y(_0948_),
    .B1(_1155_));
 sg13g2_o21ai_1 _2496_ (.B1(_0948_),
    .Y(_0949_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .A2(_0910_));
 sg13g2_nor2_2 _2497_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .B(net1010),
    .Y(_0950_));
 sg13g2_a21oi_2 _2498_ (.B1(_0950_),
    .Y(_0951_),
    .A2(_0911_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ));
 sg13g2_o21ai_1 _2499_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ),
    .Y(_0952_),
    .A1(_0951_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ));
 sg13g2_inv_2 _2500_ (.Y(_0953_),
    .A(_0952_));
 sg13g2_mux4_1 _2501_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .A0(net1074),
    .A1(net1219),
    .A2(net88),
    .A3(net980),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .X(_0954_));
 sg13g2_nor2_1 _2502_ (.A(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ),
    .B(_0954_),
    .Y(_0955_));
 sg13g2_a21oi_2 _2503_ (.B1(_0955_),
    .Y(\Inst_RegFile_switch_matrix.SS4BEG0 ),
    .A2(_0953_),
    .A1(_0949_));
 sg13g2_mux4_1 _2504_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .A0(net57),
    .A1(net85),
    .A2(net1219),
    .A3(net1070),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0956_));
 sg13g2_mux4_1 _2505_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .A0(net1020),
    .A1(net967),
    .A2(net980),
    .A3(net974),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0957_));
 sg13g2_mux4_1 _2506_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .A0(_0896_),
    .A1(_0895_),
    .A2(net499),
    .A3(net500),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .X(_0958_));
 sg13g2_mux4_1 _2507_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .A0(net1034),
    .A1(net989),
    .A2(net1015),
    .A3(net1003),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .X(_0959_));
 sg13g2_mux4_1 _2508_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .A0(_0956_),
    .A1(_0957_),
    .A2(_0959_),
    .A3(_0958_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .X(\Inst_RegFile_switch_matrix.E6BEG1 ));
 sg13g2_nand2b_1 _2509_ (.Y(_0960_),
    .B(net54),
    .A_N(net1063));
 sg13g2_a21oi_1 _2510_ (.A1(net1218),
    .A2(net1064),
    .Y(_0961_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_nor2b_1 _2511_ (.A(net1063),
    .B_N(net82),
    .Y(_0962_));
 sg13g2_a21oi_1 _2512_ (.A1(net1068),
    .A2(net1063),
    .Y(_0963_),
    .B1(_0962_));
 sg13g2_a221oi_1 _2513_ (.B2(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .B1(_0963_),
    .A1(_0960_),
    .Y(_0964_),
    .A2(_0961_));
 sg13g2_nor2b_1 _2514_ (.A(net1064),
    .B_N(net967),
    .Y(_0965_));
 sg13g2_a21oi_1 _2515_ (.A1(net1064),
    .A2(net972),
    .Y(_0966_),
    .B1(_0965_));
 sg13g2_a21oi_1 _2516_ (.A1(net1063),
    .A2(net978),
    .Y(_0967_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_o21ai_1 _2517_ (.B1(_0967_),
    .Y(_0968_),
    .A1(net1063),
    .A2(_1166_));
 sg13g2_a21oi_1 _2518_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0966_),
    .Y(_0969_),
    .B1(_1156_));
 sg13g2_a21oi_1 _2519_ (.A1(_0968_),
    .A2(_0969_),
    .Y(_0970_),
    .B1(_0964_));
 sg13g2_mux2_1 _2520_ (.A0(_0911_),
    .A1(_0910_),
    .S(net1063),
    .X(_0971_));
 sg13g2_o21ai_1 _2521_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .Y(_0972_),
    .A1(net1063),
    .A2(_1183_));
 sg13g2_a21oi_1 _2522_ (.A1(net1063),
    .A2(_0338_),
    .Y(_0973_),
    .B1(_0972_));
 sg13g2_nor2_1 _2523_ (.A(_1156_),
    .B(_0973_),
    .Y(_0974_));
 sg13g2_o21ai_1 _2524_ (.B1(_0974_),
    .Y(_0975_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .A2(_0971_));
 sg13g2_mux4_1 _2525_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .A0(net1033),
    .A1(net988),
    .A2(net1015),
    .A3(net1003),
    .S1(net1064),
    .X(_0976_));
 sg13g2_a21oi_2 _2526_ (.B1(_1157_),
    .Y(_0977_),
    .A2(_1156_),
    .A1(_0976_));
 sg13g2_a22oi_1 _2527_ (.Y(\Inst_RegFile_switch_matrix.E6BEG0 ),
    .B1(_0975_),
    .B2(_0977_),
    .A2(_0970_),
    .A1(_1157_));
 sg13g2_mux4_1 _2528_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ),
    .A0(net40),
    .A1(net11),
    .A2(net85),
    .A3(net95),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ),
    .X(_0978_));
 sg13g2_mux4_1 _2529_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(net1033),
    .A1(net499),
    .A2(net500),
    .A3(_0978_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0979_));
 sg13g2_mux4_1 _2530_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .A0(net1075),
    .A1(net1220),
    .A2(net59),
    .A3(net1019),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .X(_0980_));
 sg13g2_mux2_1 _2531_ (.A0(_0980_),
    .A1(_0979_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.EE4BEG3 ));
 sg13g2_mux4_1 _2532_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(net57),
    .A1(net11),
    .A2(net68),
    .A3(net95),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_0981_));
 sg13g2_o21ai_1 _2533_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .Y(_0982_),
    .A1(_1158_),
    .A2(_0981_));
 sg13g2_a21oi_1 _2534_ (.A1(_1158_),
    .A2(_0339_),
    .Y(_0983_),
    .B1(_0982_));
 sg13g2_nor2_1 _2535_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .B(_1165_),
    .Y(_0984_));
 sg13g2_a21oi_1 _2536_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_1182_),
    .Y(_0985_),
    .B1(_0984_));
 sg13g2_o21ai_1 _2537_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .Y(_0986_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_0985_));
 sg13g2_nor2_1 _2538_ (.A(_0983_),
    .B(_0986_),
    .Y(_0987_));
 sg13g2_mux4_1 _2539_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .A0(net1076),
    .A1(net1221),
    .A2(net58),
    .A3(net974),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .X(_0988_));
 sg13g2_nor2_1 _2540_ (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_nor2_1 _2541_ (.A(_0987_),
    .B(_0989_),
    .Y(\Inst_RegFile_switch_matrix.EE4BEG2 ));
 sg13g2_mux4_1 _2542_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .A0(net988),
    .A1(_0895_),
    .A2(_0896_),
    .A3(_0641_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .X(_0990_));
 sg13g2_mux4_1 _2543_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A0(net1073),
    .A1(net1218),
    .A2(net61),
    .A3(net967),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .X(_0991_));
 sg13g2_mux2_2 _2544_ (.A0(_0991_),
    .A1(_0990_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ),
    .X(\Inst_RegFile_switch_matrix.EE4BEG1 ));
 sg13g2_mux4_1 _2545_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .A0(net1015),
    .A1(_0910_),
    .A2(_0911_),
    .A3(_0603_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .X(_0992_));
 sg13g2_mux4_1 _2546_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .A0(net1074),
    .A1(net1219),
    .A2(net60),
    .A3(net980),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .X(_0993_));
 sg13g2_mux2_1 _2547_ (.A0(_0993_),
    .A1(_0992_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ),
    .X(\Inst_RegFile_switch_matrix.EE4BEG0 ));
 sg13g2_mux4_1 _2548_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(net54),
    .A1(net64),
    .A2(net7),
    .A3(net91),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ),
    .X(_0994_));
 sg13g2_mux4_1 _2549_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .A0(net1033),
    .A1(net499),
    .A2(net500),
    .A3(_0994_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0995_));
 sg13g2_mux4_1 _2550_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .A0(net1075),
    .A1(net1220),
    .A2(net1071),
    .A3(net1019),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .X(_0996_));
 sg13g2_mux2_1 _2551_ (.A0(_0996_),
    .A1(_0995_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG3 ));
 sg13g2_mux4_1 _2552_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ),
    .A0(net36),
    .A1(net64),
    .A2(net7),
    .A3(net108),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ),
    .X(_0997_));
 sg13g2_o21ai_1 _2553_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .Y(_0998_),
    .A1(_1159_),
    .A2(_0997_));
 sg13g2_a21oi_1 _2554_ (.A1(_1159_),
    .A2(_0339_),
    .Y(_0999_),
    .B1(_0998_));
 sg13g2_nor2_1 _2555_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .B(_1165_),
    .Y(_1000_));
 sg13g2_a21oi_1 _2556_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_1182_),
    .Y(_1001_),
    .B1(_1000_));
 sg13g2_o21ai_1 _2557_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .Y(_1002_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_1001_));
 sg13g2_nor2_1 _2558_ (.A(_0999_),
    .B(_1002_),
    .Y(_1003_));
 sg13g2_mux4_1 _2559_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .A0(net1076),
    .A1(net1221),
    .A2(net1072),
    .A3(net974),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .X(_1004_));
 sg13g2_nor2_2 _2560_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_nor2_1 _2561_ (.A(_1003_),
    .B(_1005_),
    .Y(\Inst_RegFile_switch_matrix.NN4BEG2 ));
 sg13g2_mux4_1 _2562_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .A0(net986),
    .A1(_0895_),
    .A2(_0896_),
    .A3(_1207_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .X(_1006_));
 sg13g2_mux4_1 _2563_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .A0(net1073),
    .A1(net1218),
    .A2(net1068),
    .A3(net718),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .X(_1007_));
 sg13g2_mux2_1 _2564_ (.A0(_1007_),
    .A1(_1006_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ),
    .X(\Inst_RegFile_switch_matrix.NN4BEG1 ));
 sg13g2_a21oi_1 _2565_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .A2(_0363_),
    .Y(_1008_),
    .B1(_1160_));
 sg13g2_o21ai_1 _2566_ (.B1(_1008_),
    .Y(_1009_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .A2(_0910_));
 sg13g2_nor2_2 _2567_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .B(net1010),
    .Y(_1010_));
 sg13g2_a21oi_2 _2568_ (.B1(_1010_),
    .Y(_1011_),
    .A2(_0911_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ));
 sg13g2_o21ai_1 _2569_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .Y(_1012_),
    .A1(_1011_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ));
 sg13g2_inv_2 _2570_ (.Y(_1013_),
    .A(_1012_));
 sg13g2_mux4_1 _2571_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .A0(net1074),
    .A1(net1219),
    .A2(net88),
    .A3(net980),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .X(_1014_));
 sg13g2_nor2_1 _2572_ (.A(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_a21oi_2 _2573_ (.B1(_1015_),
    .Y(\Inst_RegFile_switch_matrix.NN4BEG0 ),
    .A2(_1013_),
    .A1(_1009_));
 sg13g2_mux4_1 _2574_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(net57),
    .A1(net81),
    .A2(net106),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_1016_));
 sg13g2_mux4_1 _2575_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .A0(net1018),
    .A1(_0486_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .A3(_1016_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG3 ));
 sg13g2_mux4_1 _2576_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ),
    .A0(net1001),
    .A1(_0338_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .A3(net522),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG2 ));
 sg13g2_mux4_1 _2577_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .A0(net984),
    .A1(_0645_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .A3(net502),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG1 ));
 sg13g2_mux4_1 _2578_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ),
    .A0(net52),
    .A1(net96),
    .A2(net7),
    .A3(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ),
    .X(_1017_));
 sg13g2_mux4_1 _2579_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ),
    .A0(net43),
    .A1(net14),
    .A2(net71),
    .A3(net98),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ),
    .X(_1018_));
 sg13g2_mux4_1 _2580_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ),
    .A0(net1012),
    .A1(net512),
    .A2(_1018_),
    .A3(_1017_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .X(\Inst_RegFile_switch_matrix.W1BEG0 ));
 sg13g2_mux4_1 _2581_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ),
    .A0(net63),
    .A1(net1067),
    .A2(net78),
    .A3(net975),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG3 ));
 sg13g2_mux4_1 _2582_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ),
    .A0(net62),
    .A1(net1065),
    .A2(net81),
    .A3(net967),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG2 ));
 sg13g2_mux4_1 _2583_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ),
    .A0(net1216),
    .A1(net65),
    .A2(net80),
    .A3(net979),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG1 ));
 sg13g2_mux4_1 _2584_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ),
    .A0(net1214),
    .A1(net79),
    .A2(net64),
    .A3(net1020),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ),
    .X(\Inst_RegFile_switch_matrix.S4BEG0 ));
 sg13g2_mux4_1 _2585_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .A0(net1003),
    .A1(_0486_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .A3(_1016_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _2586_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ),
    .A0(net985),
    .A1(_0338_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .A3(net522),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _2587_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .A0(net1015),
    .A1(_0645_),
    .A2(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .A3(_0137_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _2588_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ),
    .A0(net1030),
    .A1(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .A2(_1018_),
    .A3(_1017_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .X(\Inst_RegFile_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _2589_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .A0(net988),
    .A1(_0486_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .A3(_1016_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG3 ));
 sg13g2_mux4_1 _2590_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ),
    .A0(net1012),
    .A1(_0338_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .A3(net522),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG2 ));
 sg13g2_mux4_1 _2591_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .A0(net1034),
    .A1(_0645_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .A3(_0137_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG1 ));
 sg13g2_mux4_1 _2592_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ),
    .A0(net975),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .A2(_1018_),
    .A3(_1017_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .X(\Inst_RegFile_switch_matrix.E1BEG0 ));
 sg13g2_mux4_1 _2593_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ),
    .A0(net35),
    .A1(net50),
    .A2(net1066),
    .A3(net1001),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG3 ));
 sg13g2_mux4_1 _2594_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ),
    .A0(net34),
    .A1(net1065),
    .A2(net53),
    .A3(net986),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG2 ));
 sg13g2_mux4_1 _2595_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ),
    .A0(net37),
    .A1(net52),
    .A2(net1216),
    .A3(net1013),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG1 ));
 sg13g2_mux4_1 _2596_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ),
    .A0(net36),
    .A1(net51),
    .A2(net1214),
    .A3(net1031),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ),
    .X(\Inst_RegFile_switch_matrix.N4BEG0 ));
 sg13g2_mux4_1 _2597_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .A0(net1013),
    .A1(_0486_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .A3(_1016_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _2598_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ),
    .A0(net1029),
    .A1(_0338_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .A3(net521),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG2 ));
 sg13g2_mux4_1 _2599_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .A0(net970),
    .A1(_0645_),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .A3(net502),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG1 ));
 sg13g2_mux4_1 _2600_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ),
    .A0(net963),
    .A1(net509),
    .A2(_1018_),
    .A3(_1017_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .X(\Inst_RegFile_switch_matrix.N1BEG0 ));
 sg13g2_mux4_1 _2601_ (.S0(_1161_),
    .A0(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .A1(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .A2(net721),
    .A3(_0935_),
    .S1(_1162_),
    .X(_1019_));
 sg13g2_nand2b_1 _2602_ (.Y(_1020_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ),
    .A_N(_1019_));
 sg13g2_nor2_1 _2603_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .B(_1180_),
    .Y(_1021_));
 sg13g2_o21ai_1 _2604_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .Y(_1022_),
    .A1(_1161_),
    .A2(_1231_));
 sg13g2_mux2_1 _2605_ (.A0(net34),
    .A1(net62),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .X(_1023_));
 sg13g2_a21oi_1 _2606_ (.A1(_1162_),
    .A2(_1023_),
    .Y(_1024_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_o21ai_1 _2607_ (.B1(_1024_),
    .Y(_1025_),
    .A1(_1021_),
    .A2(_1022_));
 sg13g2_and2_1 _2608_ (.A(_1020_),
    .B(_1025_),
    .X(_1026_));
 sg13g2_mux4_1 _2609_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(net50),
    .A1(net1066),
    .A2(net82),
    .A3(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_1027_));
 sg13g2_mux4_1 _2610_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ),
    .A0(net42),
    .A1(net97),
    .A2(net70),
    .A3(net524),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ),
    .X(_1028_));
 sg13g2_mux4_1 _2611_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .A0(_1028_),
    .A1(_1018_),
    .A2(_0209_),
    .A3(_1027_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_1029_));
 sg13g2_nand2_1 _2612_ (.Y(_1030_),
    .A(_1026_),
    .B(_1029_));
 sg13g2_mux4_1 _2613_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(net47),
    .A1(net18),
    .A2(net75),
    .A3(net102),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_1031_));
 sg13g2_mux4_1 _2614_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(net55),
    .A1(net22),
    .A2(net79),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ),
    .X(_1032_));
 sg13g2_mux4_1 _2615_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .A0(_0895_),
    .A1(_0922_),
    .A2(_1031_),
    .A3(_1032_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_1033_));
 sg13g2_nor2_1 _2616_ (.A(_1030_),
    .B(_1033_),
    .Y(_1034_));
 sg13g2_mux2_1 _2617_ (.A0(net108),
    .A1(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .X(_1035_));
 sg13g2_nor2b_1 _2618_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .B_N(net8),
    .Y(_1036_));
 sg13g2_a21oi_1 _2619_ (.A1(net85),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .Y(_1037_),
    .B1(_1036_));
 sg13g2_o21ai_1 _2620_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_1038_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_1037_));
 sg13g2_a21oi_1 _2621_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(_1035_),
    .Y(_1039_),
    .B1(_1038_));
 sg13g2_o21ai_1 _2622_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .Y(_1040_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0981_));
 sg13g2_or2_1 _2623_ (.X(_1041_),
    .B(_1040_),
    .A(_1039_));
 sg13g2_mux4_1 _2624_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(net19),
    .A1(net76),
    .A2(net103),
    .A3(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_1042_));
 sg13g2_mux4_1 _2625_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ),
    .A0(net49),
    .A1(net20),
    .A2(net77),
    .A3(net104),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_1043_));
 sg13g2_inv_1 _2626_ (.Y(_1044_),
    .A(_1043_));
 sg13g2_a21oi_1 _2627_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1044_),
    .Y(_1045_),
    .B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_o21ai_1 _2628_ (.B1(_1045_),
    .Y(_1046_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_1042_));
 sg13g2_and2_1 _2629_ (.A(_1041_),
    .B(_1046_),
    .X(_1047_));
 sg13g2_nand2_1 _2630_ (.Y(_1048_),
    .A(_1041_),
    .B(_1046_));
 sg13g2_and2_1 _2631_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .B(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .X(_1049_));
 sg13g2_a21oi_1 _2632_ (.A1(_1163_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .Y(_1050_),
    .B1(_1049_));
 sg13g2_nor2_1 _2633_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .B(_0432_),
    .Y(_1051_));
 sg13g2_a21oi_1 _2634_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .Y(_1052_),
    .B1(_1051_));
 sg13g2_mux4_1 _2635_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(net44),
    .A1(net99),
    .A2(net15),
    .A3(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ),
    .X(_1053_));
 sg13g2_and2_1 _2636_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .B(_1031_),
    .X(_1054_));
 sg13g2_a21oi_2 _2637_ (.B1(_1054_),
    .Y(_1055_),
    .A2(_1053_),
    .A1(_1163_));
 sg13g2_nand2b_1 _2638_ (.Y(_1056_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A_N(net65));
 sg13g2_o21ai_1 _2639_ (.B1(_1056_),
    .Y(_1057_),
    .A1(net37),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_mux4_1 _2640_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .A0(_1057_),
    .A1(_1055_),
    .A2(_1052_),
    .A3(_1050_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ),
    .X(_1058_));
 sg13g2_mux4_1 _2641_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .A0(_1053_),
    .A1(_0997_),
    .A2(_0910_),
    .A3(_1017_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ),
    .X(_1059_));
 sg13g2_inv_1 _2642_ (.Y(_1060_),
    .A(_1059_));
 sg13g2_nor3_2 _2643_ (.A(_1058_),
    .B(_1048_),
    .C(_1059_),
    .Y(_1061_));
 sg13g2_nand2_2 _2644_ (.Y(_1062_),
    .A(_1061_),
    .B(_1034_));
 sg13g2_mux4_1 _2645_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(net48),
    .A1(net76),
    .A2(net103),
    .A3(net517),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ),
    .X(_1063_));
 sg13g2_mux4_1 _2646_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ),
    .A0(net49),
    .A1(net20),
    .A2(net77),
    .A3(net104),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ),
    .X(_1064_));
 sg13g2_mux4_1 _2647_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .A0(_1063_),
    .A1(_1064_),
    .A2(_0978_),
    .A3(_1016_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .X(_1065_));
 sg13g2_mux2_1 _2648_ (.A0(net942),
    .A1(net844),
    .S(_1062_),
    .X(_0000_));
 sg13g2_mux4_1 _2649_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ),
    .A0(net23),
    .A1(net96),
    .A2(net80),
    .A3(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ),
    .X(_1066_));
 sg13g2_mux4_1 _2650_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(_0484_),
    .A1(_0911_),
    .A2(_0994_),
    .A3(_1066_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ),
    .X(_1067_));
 sg13g2_mux2_1 _2651_ (.A0(net953),
    .A1(net767),
    .S(_1062_),
    .X(_0001_));
 sg13g2_mux4_1 _2652_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ),
    .A0(net51),
    .A1(net1065),
    .A2(net1214),
    .A3(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ),
    .X(_1068_));
 sg13g2_mux4_1 _2653_ (.S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ),
    .A0(_0896_),
    .A1(_0919_),
    .A2(_0486_),
    .A3(_1068_),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .X(_1069_));
 sg13g2_mux2_1 _2654_ (.A0(net961),
    .A1(net805),
    .S(_1062_),
    .X(_0002_));
 sg13g2_mux2_1 _2655_ (.A0(net78),
    .A1(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .X(_1070_));
 sg13g2_nor2b_1 _2656_ (.A(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .B_N(net50),
    .Y(_1071_));
 sg13g2_a21oi_1 _2657_ (.A1(net1216),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .Y(_1072_),
    .B1(_1071_));
 sg13g2_o21ai_1 _2658_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_1073_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_1072_));
 sg13g2_a21oi_1 _2659_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_1070_),
    .Y(_1074_),
    .B1(_1073_));
 sg13g2_o21ai_1 _2660_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .Y(_1075_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0935_));
 sg13g2_mux2_1 _2661_ (.A0(net70),
    .A1(net508),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .X(_1076_));
 sg13g2_nand2b_1 _2662_ (.Y(_1077_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .A_N(net13));
 sg13g2_nor2_1 _2663_ (.A(net42),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .Y(_1078_));
 sg13g2_nor2_1 _2664_ (.A(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_1078_),
    .Y(_1079_));
 sg13g2_a221oi_1 _2665_ (.B2(_1079_),
    .C1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .B1(_1077_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .Y(_1080_),
    .A2(_1076_));
 sg13g2_nand2b_1 _2666_ (.Y(_1081_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ),
    .A_N(net14));
 sg13g2_o21ai_1 _2667_ (.B1(_1081_),
    .Y(_1082_),
    .A1(net43),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_mux2_1 _2668_ (.A0(net71),
    .A1(net98),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ),
    .X(_1083_));
 sg13g2_o21ai_1 _2669_ (.B1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .Y(_1084_),
    .A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_1082_));
 sg13g2_a21oi_1 _2670_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ),
    .A2(_1083_),
    .Y(_1085_),
    .B1(_1084_));
 sg13g2_or3_1 _2671_ (.A(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .B(_1080_),
    .C(_1085_),
    .X(_1086_));
 sg13g2_o21ai_1 _2672_ (.B1(_1086_),
    .Y(_1087_),
    .A1(_1074_),
    .A2(_1075_));
 sg13g2_mux2_1 _2673_ (.A0(net935),
    .A1(net799),
    .S(_1062_),
    .X(_0003_));
 sg13g2_nor3_2 _2674_ (.A(_1058_),
    .B(_1047_),
    .C(_1059_),
    .Y(_1088_));
 sg13g2_nand2_2 _2675_ (.Y(_1089_),
    .A(_1088_),
    .B(_1034_));
 sg13g2_mux2_1 _2676_ (.A0(net942),
    .A1(net850),
    .S(_1089_),
    .X(_0004_));
 sg13g2_mux2_1 _2677_ (.A0(net952),
    .A1(net810),
    .S(_1089_),
    .X(_0005_));
 sg13g2_mux2_1 _2678_ (.A0(net961),
    .A1(net782),
    .S(_1089_),
    .X(_0006_));
 sg13g2_mux2_1 _2679_ (.A0(net935),
    .A1(net830),
    .S(_1089_),
    .X(_0007_));
 sg13g2_nor3_2 _2680_ (.A(_1048_),
    .B(_1060_),
    .C(_1058_),
    .Y(_1090_));
 sg13g2_nand2_2 _2681_ (.Y(_1091_),
    .A(_1090_),
    .B(_1034_));
 sg13g2_mux2_1 _2682_ (.A0(net942),
    .A1(net757),
    .S(_1091_),
    .X(_0008_));
 sg13g2_mux2_1 _2683_ (.A0(net952),
    .A1(net755),
    .S(_1091_),
    .X(_0009_));
 sg13g2_mux2_1 _2684_ (.A0(net961),
    .A1(net768),
    .S(_1091_),
    .X(_0010_));
 sg13g2_mux2_1 _2685_ (.A0(net935),
    .A1(net744),
    .S(_1091_),
    .X(_0011_));
 sg13g2_nor3_2 _2686_ (.A(_1047_),
    .B(_1060_),
    .C(_1058_),
    .Y(_1092_));
 sg13g2_nand2_2 _2687_ (.Y(_1093_),
    .A(_1092_),
    .B(_1034_));
 sg13g2_mux2_1 _2688_ (.A0(net942),
    .A1(net807),
    .S(_1093_),
    .X(_0012_));
 sg13g2_mux2_1 _2689_ (.A0(net952),
    .A1(net794),
    .S(_1093_),
    .X(_0013_));
 sg13g2_mux2_1 _2690_ (.A0(net960),
    .A1(net819),
    .S(_1093_),
    .X(_0014_));
 sg13g2_mux2_1 _2691_ (.A0(net935),
    .A1(net849),
    .S(_1093_),
    .X(_0015_));
 sg13g2_nor2b_1 _2692_ (.A(_1030_),
    .B_N(_1033_),
    .Y(_1094_));
 sg13g2_nand2_2 _2693_ (.Y(_1095_),
    .A(_1061_),
    .B(_1094_));
 sg13g2_mux2_1 _2694_ (.A0(net937),
    .A1(net812),
    .S(_1095_),
    .X(_0016_));
 sg13g2_mux2_1 _2695_ (.A0(net950),
    .A1(net769),
    .S(_1095_),
    .X(_0017_));
 sg13g2_mux2_1 _2696_ (.A0(net959),
    .A1(net776),
    .S(_1095_),
    .X(_0018_));
 sg13g2_mux2_1 _2697_ (.A0(net933),
    .A1(net789),
    .S(_1095_),
    .X(_0019_));
 sg13g2_nor2_1 _2698_ (.A(_1026_),
    .B(_1029_),
    .Y(_1096_));
 sg13g2_nor3_1 _2699_ (.A(_1026_),
    .B(_1029_),
    .C(_1033_),
    .Y(_1097_));
 sg13g2_and2_2 _2700_ (.A(_1090_),
    .B(_1097_),
    .X(_1098_));
 sg13g2_mux2_1 _2701_ (.A0(net738),
    .A1(net937),
    .S(_1098_),
    .X(_0020_));
 sg13g2_mux2_1 _2702_ (.A0(net728),
    .A1(net949),
    .S(_1098_),
    .X(_0021_));
 sg13g2_mux2_1 _2703_ (.A0(net745),
    .A1(net959),
    .S(_1098_),
    .X(_0022_));
 sg13g2_mux2_1 _2704_ (.A0(net733),
    .A1(net932),
    .S(_1098_),
    .X(_0023_));
 sg13g2_nand2_2 _2705_ (.Y(_1099_),
    .A(_1090_),
    .B(_1094_));
 sg13g2_mux2_1 _2706_ (.A0(net937),
    .A1(net775),
    .S(_1099_),
    .X(_0024_));
 sg13g2_mux2_1 _2707_ (.A0(net950),
    .A1(net820),
    .S(_1099_),
    .X(_0025_));
 sg13g2_mux2_1 _2708_ (.A0(net959),
    .A1(net842),
    .S(_1099_),
    .X(_0026_));
 sg13g2_mux2_1 _2709_ (.A0(net933),
    .A1(net787),
    .S(_1099_),
    .X(_0027_));
 sg13g2_nand2b_1 _2710_ (.Y(_1100_),
    .B(_1029_),
    .A_N(_1026_));
 sg13g2_nor2_1 _2711_ (.A(_1033_),
    .B(_1100_),
    .Y(_1101_));
 sg13g2_nand2_2 _2712_ (.Y(_1102_),
    .A(_1088_),
    .B(_1101_));
 sg13g2_mux2_1 _2713_ (.A0(net941),
    .A1(net821),
    .S(_1102_),
    .X(_0028_));
 sg13g2_mux2_1 _2714_ (.A0(net953),
    .A1(net831),
    .S(_1102_),
    .X(_0029_));
 sg13g2_mux2_1 _2715_ (.A0(net961),
    .A1(net823),
    .S(_1102_),
    .X(_0030_));
 sg13g2_mux2_1 _2716_ (.A0(net935),
    .A1(net811),
    .S(_1102_),
    .X(_0031_));
 sg13g2_nor2b_1 _2717_ (.A(_1100_),
    .B_N(_1033_),
    .Y(_1103_));
 sg13g2_and2_2 _2718_ (.A(_1088_),
    .B(_1103_),
    .X(_1104_));
 sg13g2_mux2_1 _2719_ (.A0(net740),
    .A1(net940),
    .S(_1104_),
    .X(_0032_));
 sg13g2_mux2_1 _2720_ (.A0(net751),
    .A1(net951),
    .S(_1104_),
    .X(_0033_));
 sg13g2_mux2_1 _2721_ (.A0(net753),
    .A1(net960),
    .S(_1104_),
    .X(_0034_));
 sg13g2_mux2_1 _2722_ (.A0(net741),
    .A1(net934),
    .S(_1104_),
    .X(_0035_));
 sg13g2_nand3b_1 _2723_ (.B(_1025_),
    .C(_1020_),
    .Y(_1105_),
    .A_N(_1029_));
 sg13g2_nor2_2 _2724_ (.A(_1033_),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nand2_2 _2725_ (.Y(_1107_),
    .A(_1088_),
    .B(_1106_));
 sg13g2_mux2_1 _2726_ (.A0(net938),
    .A1(net798),
    .S(_1107_),
    .X(_0036_));
 sg13g2_mux2_1 _2727_ (.A0(net949),
    .A1(net834),
    .S(_1107_),
    .X(_0037_));
 sg13g2_mux2_1 _2728_ (.A0(net958),
    .A1(net785),
    .S(_1107_),
    .X(_0038_));
 sg13g2_mux2_1 _2729_ (.A0(net936),
    .A1(net822),
    .S(_1107_),
    .X(_0039_));
 sg13g2_nor2b_2 _2730_ (.A(_1105_),
    .B_N(_1033_),
    .Y(_1108_));
 sg13g2_nand2_2 _2731_ (.Y(_1109_),
    .A(_1090_),
    .B(_1108_));
 sg13g2_mux2_1 _2732_ (.A0(net939),
    .A1(net758),
    .S(_1109_),
    .X(_0040_));
 sg13g2_mux2_1 _2733_ (.A0(net951),
    .A1(net793),
    .S(_1109_),
    .X(_0041_));
 sg13g2_mux2_1 _2734_ (.A0(net958),
    .A1(net840),
    .S(_1109_),
    .X(_0042_));
 sg13g2_mux2_1 _2735_ (.A0(net933),
    .A1(net795),
    .S(_1109_),
    .X(_0043_));
 sg13g2_nand2_2 _2736_ (.Y(_1110_),
    .A(_1092_),
    .B(_1108_));
 sg13g2_mux2_1 _2737_ (.A0(net939),
    .A1(net841),
    .S(_1110_),
    .X(_0044_));
 sg13g2_mux2_1 _2738_ (.A0(net951),
    .A1(net832),
    .S(_1110_),
    .X(_0045_));
 sg13g2_mux2_1 _2739_ (.A0(net958),
    .A1(net847),
    .S(_1110_),
    .X(_0046_));
 sg13g2_mux2_1 _2740_ (.A0(net933),
    .A1(net828),
    .S(_1110_),
    .X(_0047_));
 sg13g2_nand2_2 _2741_ (.Y(_1111_),
    .A(_1090_),
    .B(_1103_));
 sg13g2_mux2_1 _2742_ (.A0(net940),
    .A1(net756),
    .S(_1111_),
    .X(_0048_));
 sg13g2_mux2_1 _2743_ (.A0(net954),
    .A1(net806),
    .S(_1111_),
    .X(_0049_));
 sg13g2_mux2_1 _2744_ (.A0(net960),
    .A1(net766),
    .S(_1111_),
    .X(_0050_));
 sg13g2_mux2_1 _2745_ (.A0(net934),
    .A1(net778),
    .S(_1111_),
    .X(_0051_));
 sg13g2_and2_2 _2746_ (.A(_1092_),
    .B(_1103_),
    .X(_1112_));
 sg13g2_mux2_1 _2747_ (.A0(net760),
    .A1(net940),
    .S(_1112_),
    .X(_0052_));
 sg13g2_mux2_1 _2748_ (.A0(net750),
    .A1(net951),
    .S(_1112_),
    .X(_0053_));
 sg13g2_mux2_1 _2749_ (.A0(net752),
    .A1(net960),
    .S(_1112_),
    .X(_0054_));
 sg13g2_mux2_1 _2750_ (.A0(net736),
    .A1(net934),
    .S(_1112_),
    .X(_0055_));
 sg13g2_nand2_2 _2751_ (.Y(_1113_),
    .A(_1061_),
    .B(_1106_));
 sg13g2_mux2_1 _2752_ (.A0(net938),
    .A1(net774),
    .S(_1113_),
    .X(_0056_));
 sg13g2_mux2_1 _2753_ (.A0(net949),
    .A1(net845),
    .S(_1113_),
    .X(_0057_));
 sg13g2_mux2_1 _2754_ (.A0(net958),
    .A1(net848),
    .S(_1113_),
    .X(_0058_));
 sg13g2_mux2_1 _2755_ (.A0(net932),
    .A1(net818),
    .S(_1113_),
    .X(_0059_));
 sg13g2_nand2_2 _2756_ (.Y(_1114_),
    .A(_1090_),
    .B(_1106_));
 sg13g2_mux2_1 _2757_ (.A0(net938),
    .A1(net779),
    .S(_1114_),
    .X(_0060_));
 sg13g2_mux2_1 _2758_ (.A0(net949),
    .A1(net836),
    .S(_1114_),
    .X(_0061_));
 sg13g2_mux2_1 _2759_ (.A0(net958),
    .A1(net846),
    .S(_1114_),
    .X(_0062_));
 sg13g2_mux2_1 _2760_ (.A0(net932),
    .A1(net837),
    .S(_1114_),
    .X(_0063_));
 sg13g2_nand2_2 _2761_ (.Y(_1115_),
    .A(_1088_),
    .B(_1097_));
 sg13g2_mux2_1 _2762_ (.A0(net937),
    .A1(net843),
    .S(_1115_),
    .X(_0064_));
 sg13g2_mux2_1 _2763_ (.A0(net949),
    .A1(net765),
    .S(_1115_),
    .X(_0065_));
 sg13g2_mux2_1 _2764_ (.A0(net959),
    .A1(net784),
    .S(_1115_),
    .X(_0066_));
 sg13g2_mux2_1 _2765_ (.A0(net932),
    .A1(net773),
    .S(_1115_),
    .X(_0067_));
 sg13g2_nand2_2 _2766_ (.Y(_1116_),
    .A(_1061_),
    .B(_1108_));
 sg13g2_mux2_1 _2767_ (.A0(net939),
    .A1(net762),
    .S(_1116_),
    .X(_0068_));
 sg13g2_mux2_1 _2768_ (.A0(net951),
    .A1(net763),
    .S(_1116_),
    .X(_0069_));
 sg13g2_mux2_1 _2769_ (.A0(net958),
    .A1(net761),
    .S(_1116_),
    .X(_0070_));
 sg13g2_mux2_1 _2770_ (.A0(net933),
    .A1(net817),
    .S(_1116_),
    .X(_0071_));
 sg13g2_nand2_2 _2771_ (.Y(_1117_),
    .A(_1108_),
    .B(_1088_));
 sg13g2_mux2_1 _2772_ (.A0(net939),
    .A1(net815),
    .S(_1117_),
    .X(_0072_));
 sg13g2_mux2_1 _2773_ (.A0(net951),
    .A1(net838),
    .S(_1117_),
    .X(_0073_));
 sg13g2_mux2_1 _2774_ (.A0(net958),
    .A1(net802),
    .S(_1117_),
    .X(_0074_));
 sg13g2_mux2_1 _2775_ (.A0(net933),
    .A1(net814),
    .S(_1117_),
    .X(_0075_));
 sg13g2_nand2_2 _2776_ (.Y(_1118_),
    .A(_1092_),
    .B(_1106_));
 sg13g2_mux2_1 _2777_ (.A0(net939),
    .A1(net781),
    .S(_1118_),
    .X(_0076_));
 sg13g2_mux2_1 _2778_ (.A0(net949),
    .A1(net826),
    .S(_1118_),
    .X(_0077_));
 sg13g2_mux2_1 _2779_ (.A0(net958),
    .A1(net839),
    .S(_1118_),
    .X(_0078_));
 sg13g2_mux2_1 _2780_ (.A0(net933),
    .A1(net783),
    .S(_1118_),
    .X(_0079_));
 sg13g2_nand2_2 _2781_ (.Y(_1119_),
    .A(_1088_),
    .B(_1094_));
 sg13g2_mux2_1 _2782_ (.A0(net937),
    .A1(net772),
    .S(_1119_),
    .X(_0080_));
 sg13g2_mux2_1 _2783_ (.A0(net950),
    .A1(net800),
    .S(_1119_),
    .X(_0081_));
 sg13g2_mux2_1 _2784_ (.A0(net959),
    .A1(net808),
    .S(_1119_),
    .X(_0082_));
 sg13g2_mux2_1 _2785_ (.A0(net932),
    .A1(net809),
    .S(_1119_),
    .X(_0083_));
 sg13g2_nand2_2 _2786_ (.Y(_1120_),
    .A(_1092_),
    .B(_1094_));
 sg13g2_mux2_1 _2787_ (.A0(net937),
    .A1(net824),
    .S(_1120_),
    .X(_0084_));
 sg13g2_mux2_1 _2788_ (.A0(net950),
    .A1(net827),
    .S(_1120_),
    .X(_0085_));
 sg13g2_mux2_1 _2789_ (.A0(net959),
    .A1(net829),
    .S(_1120_),
    .X(_0086_));
 sg13g2_mux2_1 _2790_ (.A0(net932),
    .A1(net851),
    .S(_1120_),
    .X(_0087_));
 sg13g2_nand2_2 _2791_ (.Y(_1121_),
    .A(_1092_),
    .B(_1097_));
 sg13g2_mux2_1 _2792_ (.A0(net937),
    .A1(net792),
    .S(_1121_),
    .X(_0088_));
 sg13g2_mux2_1 _2793_ (.A0(net949),
    .A1(net801),
    .S(_1121_),
    .X(_0089_));
 sg13g2_mux2_1 _2794_ (.A0(net959),
    .A1(net780),
    .S(_1121_),
    .X(_0090_));
 sg13g2_mux2_1 _2795_ (.A0(net932),
    .A1(net791),
    .S(_1121_),
    .X(_0091_));
 sg13g2_and2_1 _2796_ (.A(_1033_),
    .B(_1096_),
    .X(_1122_));
 sg13g2_and2_2 _2797_ (.A(_1061_),
    .B(_1122_),
    .X(_1123_));
 sg13g2_mux2_1 _2798_ (.A0(net726),
    .A1(net940),
    .S(_1123_),
    .X(_0092_));
 sg13g2_mux2_1 _2799_ (.A0(net732),
    .A1(net952),
    .S(_1123_),
    .X(_0093_));
 sg13g2_mux2_1 _2800_ (.A0(net734),
    .A1(net962),
    .S(_1123_),
    .X(_0094_));
 sg13g2_mux2_1 _2801_ (.A0(net727),
    .A1(net934),
    .S(_1123_),
    .X(_0095_));
 sg13g2_nand2_2 _2802_ (.Y(_1124_),
    .A(_1088_),
    .B(_1122_));
 sg13g2_mux2_1 _2803_ (.A0(net940),
    .A1(net777),
    .S(_1124_),
    .X(_0096_));
 sg13g2_mux2_1 _2804_ (.A0(net952),
    .A1(net788),
    .S(_1124_),
    .X(_0097_));
 sg13g2_mux2_1 _2805_ (.A0(net962),
    .A1(net764),
    .S(_1124_),
    .X(_0098_));
 sg13g2_mux2_1 _2806_ (.A0(net934),
    .A1(net797),
    .S(_1124_),
    .X(_0099_));
 sg13g2_and2_1 _2807_ (.A(_1090_),
    .B(_1122_),
    .X(_1125_));
 sg13g2_mux2_1 _2808_ (.A0(net724),
    .A1(net940),
    .S(_1125_),
    .X(_0100_));
 sg13g2_mux2_1 _2809_ (.A0(net746),
    .A1(net952),
    .S(_1125_),
    .X(_0101_));
 sg13g2_mux2_1 _2810_ (.A0(net729),
    .A1(net960),
    .S(_1125_),
    .X(_0102_));
 sg13g2_mux2_1 _2811_ (.A0(net737),
    .A1(net934),
    .S(_1125_),
    .X(_0103_));
 sg13g2_nand2_2 _2812_ (.Y(_1126_),
    .A(_1092_),
    .B(_1122_));
 sg13g2_mux2_1 _2813_ (.A0(net940),
    .A1(net835),
    .S(_1126_),
    .X(_0104_));
 sg13g2_mux2_1 _2814_ (.A0(net952),
    .A1(net770),
    .S(_1126_),
    .X(_0105_));
 sg13g2_mux2_1 _2815_ (.A0(net960),
    .A1(net803),
    .S(_1126_),
    .X(_0106_));
 sg13g2_mux2_1 _2816_ (.A0(net934),
    .A1(net786),
    .S(_1126_),
    .X(_0107_));
 sg13g2_and2_2 _2817_ (.A(_1061_),
    .B(_1101_),
    .X(_1127_));
 sg13g2_mux2_1 _2818_ (.A0(net731),
    .A1(net941),
    .S(_1127_),
    .X(_0108_));
 sg13g2_mux2_1 _2819_ (.A0(net747),
    .A1(net952),
    .S(_1127_),
    .X(_0109_));
 sg13g2_mux2_1 _2820_ (.A0(net730),
    .A1(net960),
    .S(_1127_),
    .X(_0110_));
 sg13g2_mux2_1 _2821_ (.A0(net748),
    .A1(net935),
    .S(_1127_),
    .X(_0111_));
 sg13g2_and2_2 _2822_ (.A(_1061_),
    .B(_1097_),
    .X(_1128_));
 sg13g2_mux2_1 _2823_ (.A0(net739),
    .A1(net937),
    .S(_1128_),
    .X(_0112_));
 sg13g2_mux2_1 _2824_ (.A0(net735),
    .A1(net949),
    .S(_1128_),
    .X(_0113_));
 sg13g2_mux2_1 _2825_ (.A0(net742),
    .A1(net959),
    .S(_1128_),
    .X(_0114_));
 sg13g2_mux2_1 _2826_ (.A0(net749),
    .A1(net932),
    .S(_1128_),
    .X(_0115_));
 sg13g2_and2_2 _2827_ (.A(_1090_),
    .B(_1101_),
    .X(_1129_));
 sg13g2_mux2_1 _2828_ (.A0(net759),
    .A1(net941),
    .S(_1129_),
    .X(_0116_));
 sg13g2_mux2_1 _2829_ (.A0(net754),
    .A1(net953),
    .S(_1129_),
    .X(_0117_));
 sg13g2_mux2_1 _2830_ (.A0(net725),
    .A1(net961),
    .S(_1129_),
    .X(_0118_));
 sg13g2_mux2_1 _2831_ (.A0(net743),
    .A1(net935),
    .S(_1129_),
    .X(_0119_));
 sg13g2_nand2_2 _2832_ (.Y(_1130_),
    .A(_1092_),
    .B(_1101_));
 sg13g2_mux2_1 _2833_ (.A0(net941),
    .A1(net804),
    .S(_1130_),
    .X(_0120_));
 sg13g2_mux2_1 _2834_ (.A0(net953),
    .A1(net796),
    .S(_1130_),
    .X(_0121_));
 sg13g2_mux2_1 _2835_ (.A0(net961),
    .A1(net833),
    .S(_1130_),
    .X(_0122_));
 sg13g2_mux2_1 _2836_ (.A0(net935),
    .A1(net790),
    .S(_1130_),
    .X(_0123_));
 sg13g2_nand2_2 _2837_ (.Y(_1131_),
    .A(_1061_),
    .B(_1103_));
 sg13g2_mux2_1 _2838_ (.A0(net940),
    .A1(net825),
    .S(_1131_),
    .X(_0124_));
 sg13g2_mux2_1 _2839_ (.A0(net954),
    .A1(net771),
    .S(_1131_),
    .X(_0125_));
 sg13g2_mux2_1 _2840_ (.A0(net960),
    .A1(net813),
    .S(_1131_),
    .X(_0126_));
 sg13g2_mux2_1 _2841_ (.A0(net934),
    .A1(net816),
    .S(_1131_),
    .X(_0127_));
 sg13g2_dfrbp_1 _2842_ (.CLK(UserCLK),
    .RESET_B(net439),
    .D(_0000_),
    .Q_N(_1365_),
    .Q(\Inst_RegFile_32x4.mem[24][0] ));
 sg13g2_dfrbp_1 _2843_ (.CLK(UserCLK),
    .RESET_B(net487),
    .D(_0001_),
    .Q_N(_1364_),
    .Q(\Inst_RegFile_32x4.mem[24][1] ));
 sg13g2_dfrbp_1 _2844_ (.CLK(UserCLK),
    .RESET_B(net486),
    .D(_0002_),
    .Q_N(_1363_),
    .Q(\Inst_RegFile_32x4.mem[24][2] ));
 sg13g2_dfrbp_1 _2845_ (.CLK(UserCLK),
    .RESET_B(net485),
    .D(_0003_),
    .Q_N(_1362_),
    .Q(\Inst_RegFile_32x4.mem[24][3] ));
 sg13g2_dfrbp_1 _2846_ (.CLK(UserCLK),
    .RESET_B(net484),
    .D(_0004_),
    .Q_N(_1361_),
    .Q(\Inst_RegFile_32x4.mem[25][0] ));
 sg13g2_dfrbp_1 _2847_ (.CLK(UserCLK),
    .RESET_B(net483),
    .D(_0005_),
    .Q_N(_1360_),
    .Q(\Inst_RegFile_32x4.mem[25][1] ));
 sg13g2_dfrbp_1 _2848_ (.CLK(UserCLK),
    .RESET_B(net482),
    .D(_0006_),
    .Q_N(_1359_),
    .Q(\Inst_RegFile_32x4.mem[25][2] ));
 sg13g2_dfrbp_1 _2849_ (.CLK(UserCLK),
    .RESET_B(net481),
    .D(_0007_),
    .Q_N(_1358_),
    .Q(\Inst_RegFile_32x4.mem[25][3] ));
 sg13g2_dfrbp_1 _2850_ (.CLK(UserCLK),
    .RESET_B(net480),
    .D(_0008_),
    .Q_N(_1357_),
    .Q(\Inst_RegFile_32x4.mem[26][0] ));
 sg13g2_dfrbp_1 _2851_ (.CLK(UserCLK),
    .RESET_B(net479),
    .D(_0009_),
    .Q_N(_1356_),
    .Q(\Inst_RegFile_32x4.mem[26][1] ));
 sg13g2_dfrbp_1 _2852_ (.CLK(UserCLK),
    .RESET_B(net478),
    .D(_0010_),
    .Q_N(_1355_),
    .Q(\Inst_RegFile_32x4.mem[26][2] ));
 sg13g2_dfrbp_1 _2853_ (.CLK(UserCLK),
    .RESET_B(net477),
    .D(_0011_),
    .Q_N(_1354_),
    .Q(\Inst_RegFile_32x4.mem[26][3] ));
 sg13g2_dfrbp_1 _2854_ (.CLK(UserCLK),
    .RESET_B(net476),
    .D(_0012_),
    .Q_N(_1353_),
    .Q(\Inst_RegFile_32x4.mem[27][0] ));
 sg13g2_dfrbp_1 _2855_ (.CLK(UserCLK),
    .RESET_B(net475),
    .D(_0013_),
    .Q_N(_1352_),
    .Q(\Inst_RegFile_32x4.mem[27][1] ));
 sg13g2_dfrbp_1 _2856_ (.CLK(UserCLK),
    .RESET_B(net474),
    .D(_0014_),
    .Q_N(_1351_),
    .Q(\Inst_RegFile_32x4.mem[27][2] ));
 sg13g2_dfrbp_1 _2857_ (.CLK(UserCLK),
    .RESET_B(net473),
    .D(_0015_),
    .Q_N(_1350_),
    .Q(\Inst_RegFile_32x4.mem[27][3] ));
 sg13g2_dfrbp_1 _2858_ (.CLK(UserCLK),
    .RESET_B(net472),
    .D(_0016_),
    .Q_N(_1349_),
    .Q(\Inst_RegFile_32x4.mem[28][0] ));
 sg13g2_dfrbp_1 _2859_ (.CLK(UserCLK),
    .RESET_B(net471),
    .D(_0017_),
    .Q_N(_1348_),
    .Q(\Inst_RegFile_32x4.mem[28][1] ));
 sg13g2_dfrbp_1 _2860_ (.CLK(UserCLK),
    .RESET_B(net470),
    .D(_0018_),
    .Q_N(_1347_),
    .Q(\Inst_RegFile_32x4.mem[28][2] ));
 sg13g2_dfrbp_1 _2861_ (.CLK(UserCLK),
    .RESET_B(net469),
    .D(_0019_),
    .Q_N(_1346_),
    .Q(\Inst_RegFile_32x4.mem[28][3] ));
 sg13g2_dfrbp_1 _2862_ (.CLK(UserCLK),
    .RESET_B(net468),
    .D(_0020_),
    .Q_N(_1345_),
    .Q(\Inst_RegFile_32x4.mem[2][0] ));
 sg13g2_dfrbp_1 _2863_ (.CLK(UserCLK),
    .RESET_B(net467),
    .D(_0021_),
    .Q_N(_1344_),
    .Q(\Inst_RegFile_32x4.mem[2][1] ));
 sg13g2_dfrbp_1 _2864_ (.CLK(UserCLK),
    .RESET_B(net466),
    .D(_0022_),
    .Q_N(_1343_),
    .Q(\Inst_RegFile_32x4.mem[2][2] ));
 sg13g2_dfrbp_1 _2865_ (.CLK(UserCLK),
    .RESET_B(net465),
    .D(_0023_),
    .Q_N(_1342_),
    .Q(\Inst_RegFile_32x4.mem[2][3] ));
 sg13g2_dfrbp_1 _2866_ (.CLK(UserCLK),
    .RESET_B(net464),
    .D(_0024_),
    .Q_N(_1341_),
    .Q(\Inst_RegFile_32x4.mem[30][0] ));
 sg13g2_dfrbp_1 _2867_ (.CLK(UserCLK),
    .RESET_B(net463),
    .D(_0025_),
    .Q_N(_1340_),
    .Q(\Inst_RegFile_32x4.mem[30][1] ));
 sg13g2_dfrbp_1 _2868_ (.CLK(UserCLK),
    .RESET_B(net462),
    .D(_0026_),
    .Q_N(_1339_),
    .Q(\Inst_RegFile_32x4.mem[30][2] ));
 sg13g2_dfrbp_1 _2869_ (.CLK(UserCLK),
    .RESET_B(net461),
    .D(_0027_),
    .Q_N(_1338_),
    .Q(\Inst_RegFile_32x4.mem[30][3] ));
 sg13g2_dfrbp_1 _2870_ (.CLK(UserCLK),
    .RESET_B(net460),
    .D(_0028_),
    .Q_N(_1337_),
    .Q(\Inst_RegFile_32x4.mem[9][0] ));
 sg13g2_dfrbp_1 _2871_ (.CLK(UserCLK),
    .RESET_B(net459),
    .D(_0029_),
    .Q_N(_1336_),
    .Q(\Inst_RegFile_32x4.mem[9][1] ));
 sg13g2_dfrbp_1 _2872_ (.CLK(UserCLK),
    .RESET_B(net458),
    .D(_0030_),
    .Q_N(_1335_),
    .Q(\Inst_RegFile_32x4.mem[9][2] ));
 sg13g2_dfrbp_1 _2873_ (.CLK(UserCLK),
    .RESET_B(net457),
    .D(_0031_),
    .Q_N(_1334_),
    .Q(\Inst_RegFile_32x4.mem[9][3] ));
 sg13g2_dfrbp_1 _2874_ (.CLK(UserCLK),
    .RESET_B(net456),
    .D(_0032_),
    .Q_N(_1333_),
    .Q(\Inst_RegFile_32x4.mem[13][0] ));
 sg13g2_dfrbp_1 _2875_ (.CLK(UserCLK),
    .RESET_B(net455),
    .D(_0033_),
    .Q_N(_1332_),
    .Q(\Inst_RegFile_32x4.mem[13][1] ));
 sg13g2_dfrbp_1 _2876_ (.CLK(UserCLK),
    .RESET_B(net454),
    .D(_0034_),
    .Q_N(_1331_),
    .Q(\Inst_RegFile_32x4.mem[13][2] ));
 sg13g2_dfrbp_1 _2877_ (.CLK(UserCLK),
    .RESET_B(net453),
    .D(_0035_),
    .Q_N(_1330_),
    .Q(\Inst_RegFile_32x4.mem[13][3] ));
 sg13g2_dfrbp_1 _2878_ (.CLK(UserCLK),
    .RESET_B(net452),
    .D(_0036_),
    .Q_N(_1329_),
    .Q(\Inst_RegFile_32x4.mem[17][0] ));
 sg13g2_dfrbp_1 _2879_ (.CLK(UserCLK),
    .RESET_B(net451),
    .D(_0037_),
    .Q_N(_1328_),
    .Q(\Inst_RegFile_32x4.mem[17][1] ));
 sg13g2_dfrbp_1 _2880_ (.CLK(UserCLK),
    .RESET_B(net450),
    .D(_0038_),
    .Q_N(_1327_),
    .Q(\Inst_RegFile_32x4.mem[17][2] ));
 sg13g2_dfrbp_1 _2881_ (.CLK(UserCLK),
    .RESET_B(net449),
    .D(_0039_),
    .Q_N(_1326_),
    .Q(\Inst_RegFile_32x4.mem[17][3] ));
 sg13g2_dfrbp_1 _2882_ (.CLK(UserCLK),
    .RESET_B(net448),
    .D(_0040_),
    .Q_N(_1325_),
    .Q(\Inst_RegFile_32x4.mem[22][0] ));
 sg13g2_dfrbp_1 _2883_ (.CLK(UserCLK),
    .RESET_B(net447),
    .D(_0041_),
    .Q_N(_1324_),
    .Q(\Inst_RegFile_32x4.mem[22][1] ));
 sg13g2_dfrbp_1 _2884_ (.CLK(UserCLK),
    .RESET_B(net438),
    .D(_0042_),
    .Q_N(_1323_),
    .Q(\Inst_RegFile_32x4.mem[22][2] ));
 sg13g2_dfrbp_1 _2885_ (.CLK(UserCLK),
    .RESET_B(net437),
    .D(_0043_),
    .Q_N(_1322_),
    .Q(\Inst_RegFile_32x4.mem[22][3] ));
 sg13g2_dfrbp_1 _2886_ (.CLK(UserCLK),
    .RESET_B(net436),
    .D(_0044_),
    .Q_N(_1321_),
    .Q(\Inst_RegFile_32x4.mem[23][0] ));
 sg13g2_dfrbp_1 _2887_ (.CLK(UserCLK),
    .RESET_B(net435),
    .D(_0045_),
    .Q_N(_1320_),
    .Q(\Inst_RegFile_32x4.mem[23][1] ));
 sg13g2_dfrbp_1 _2888_ (.CLK(UserCLK),
    .RESET_B(net434),
    .D(_0046_),
    .Q_N(_1319_),
    .Q(\Inst_RegFile_32x4.mem[23][2] ));
 sg13g2_dfrbp_1 _2889_ (.CLK(UserCLK),
    .RESET_B(net433),
    .D(_0047_),
    .Q_N(_1318_),
    .Q(\Inst_RegFile_32x4.mem[23][3] ));
 sg13g2_dfrbp_1 _2890_ (.CLK(UserCLK),
    .RESET_B(net432),
    .D(_0048_),
    .Q_N(_1317_),
    .Q(\Inst_RegFile_32x4.mem[14][0] ));
 sg13g2_dfrbp_1 _2891_ (.CLK(UserCLK),
    .RESET_B(net431),
    .D(_0049_),
    .Q_N(_1316_),
    .Q(\Inst_RegFile_32x4.mem[14][1] ));
 sg13g2_dfrbp_1 _2892_ (.CLK(UserCLK),
    .RESET_B(net430),
    .D(_0050_),
    .Q_N(_1315_),
    .Q(\Inst_RegFile_32x4.mem[14][2] ));
 sg13g2_dfrbp_1 _2893_ (.CLK(UserCLK),
    .RESET_B(net429),
    .D(_0051_),
    .Q_N(_1314_),
    .Q(\Inst_RegFile_32x4.mem[14][3] ));
 sg13g2_dfrbp_1 _2894_ (.CLK(UserCLK),
    .RESET_B(net428),
    .D(_0052_),
    .Q_N(_1313_),
    .Q(\Inst_RegFile_32x4.mem[15][0] ));
 sg13g2_dfrbp_1 _2895_ (.CLK(UserCLK),
    .RESET_B(net427),
    .D(_0053_),
    .Q_N(_1312_),
    .Q(\Inst_RegFile_32x4.mem[15][1] ));
 sg13g2_dfrbp_1 _2896_ (.CLK(UserCLK),
    .RESET_B(net426),
    .D(_0054_),
    .Q_N(_1311_),
    .Q(\Inst_RegFile_32x4.mem[15][2] ));
 sg13g2_dfrbp_1 _2897_ (.CLK(UserCLK),
    .RESET_B(net425),
    .D(_0055_),
    .Q_N(_1310_),
    .Q(\Inst_RegFile_32x4.mem[15][3] ));
 sg13g2_dfrbp_1 _2898_ (.CLK(UserCLK),
    .RESET_B(net424),
    .D(_0056_),
    .Q_N(_1309_),
    .Q(\Inst_RegFile_32x4.mem[16][0] ));
 sg13g2_dfrbp_1 _2899_ (.CLK(UserCLK),
    .RESET_B(net423),
    .D(_0057_),
    .Q_N(_1308_),
    .Q(\Inst_RegFile_32x4.mem[16][1] ));
 sg13g2_dfrbp_1 _2900_ (.CLK(UserCLK),
    .RESET_B(net422),
    .D(_0058_),
    .Q_N(_1307_),
    .Q(\Inst_RegFile_32x4.mem[16][2] ));
 sg13g2_dfrbp_1 _2901_ (.CLK(UserCLK),
    .RESET_B(net421),
    .D(_0059_),
    .Q_N(_1306_),
    .Q(\Inst_RegFile_32x4.mem[16][3] ));
 sg13g2_dfrbp_1 _2902_ (.CLK(UserCLK),
    .RESET_B(net420),
    .D(_0060_),
    .Q_N(_1305_),
    .Q(\Inst_RegFile_32x4.mem[18][0] ));
 sg13g2_dfrbp_1 _2903_ (.CLK(UserCLK),
    .RESET_B(net419),
    .D(_0061_),
    .Q_N(_1304_),
    .Q(\Inst_RegFile_32x4.mem[18][1] ));
 sg13g2_dfrbp_1 _2904_ (.CLK(UserCLK),
    .RESET_B(net418),
    .D(_0062_),
    .Q_N(_1303_),
    .Q(\Inst_RegFile_32x4.mem[18][2] ));
 sg13g2_dfrbp_1 _2905_ (.CLK(UserCLK),
    .RESET_B(net417),
    .D(_0063_),
    .Q_N(_1302_),
    .Q(\Inst_RegFile_32x4.mem[18][3] ));
 sg13g2_dfrbp_1 _2906_ (.CLK(UserCLK),
    .RESET_B(net416),
    .D(_0064_),
    .Q_N(_1301_),
    .Q(\Inst_RegFile_32x4.mem[1][0] ));
 sg13g2_dfrbp_1 _2907_ (.CLK(UserCLK),
    .RESET_B(net415),
    .D(_0065_),
    .Q_N(_1300_),
    .Q(\Inst_RegFile_32x4.mem[1][1] ));
 sg13g2_dfrbp_1 _2908_ (.CLK(UserCLK),
    .RESET_B(net414),
    .D(_0066_),
    .Q_N(_1299_),
    .Q(\Inst_RegFile_32x4.mem[1][2] ));
 sg13g2_dfrbp_1 _2909_ (.CLK(UserCLK),
    .RESET_B(net413),
    .D(_0067_),
    .Q_N(_1298_),
    .Q(\Inst_RegFile_32x4.mem[1][3] ));
 sg13g2_dfrbp_1 _2910_ (.CLK(UserCLK),
    .RESET_B(net412),
    .D(_0068_),
    .Q_N(_1297_),
    .Q(\Inst_RegFile_32x4.mem[20][0] ));
 sg13g2_dfrbp_1 _2911_ (.CLK(UserCLK),
    .RESET_B(net411),
    .D(_0069_),
    .Q_N(_1296_),
    .Q(\Inst_RegFile_32x4.mem[20][1] ));
 sg13g2_dfrbp_1 _2912_ (.CLK(UserCLK),
    .RESET_B(net410),
    .D(_0070_),
    .Q_N(_1295_),
    .Q(\Inst_RegFile_32x4.mem[20][2] ));
 sg13g2_dfrbp_1 _2913_ (.CLK(UserCLK),
    .RESET_B(net409),
    .D(_0071_),
    .Q_N(_1294_),
    .Q(\Inst_RegFile_32x4.mem[20][3] ));
 sg13g2_dfrbp_1 _2914_ (.CLK(UserCLK),
    .RESET_B(net408),
    .D(_0072_),
    .Q_N(_1293_),
    .Q(\Inst_RegFile_32x4.mem[21][0] ));
 sg13g2_dfrbp_1 _2915_ (.CLK(UserCLK),
    .RESET_B(net407),
    .D(_0073_),
    .Q_N(_1292_),
    .Q(\Inst_RegFile_32x4.mem[21][1] ));
 sg13g2_dfrbp_1 _2916_ (.CLK(UserCLK),
    .RESET_B(net406),
    .D(_0074_),
    .Q_N(_1291_),
    .Q(\Inst_RegFile_32x4.mem[21][2] ));
 sg13g2_dfrbp_1 _2917_ (.CLK(UserCLK),
    .RESET_B(net440),
    .D(_0075_),
    .Q_N(_1366_),
    .Q(\Inst_RegFile_32x4.mem[21][3] ));
 sg13g2_dlhq_1 _2918_ (.D(net1167),
    .GATE(net1130),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ));
 sg13g2_dlhq_1 _2919_ (.D(net1161),
    .GATE(net1130),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ));
 sg13g2_dlhq_1 _2920_ (.D(net1159),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ));
 sg13g2_dlhq_1 _2921_ (.D(net1157),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ));
 sg13g2_dlhq_1 _2922_ (.D(net1154),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ));
 sg13g2_dlhq_1 _2923_ (.D(net1152),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ));
 sg13g2_dlhq_1 _2924_ (.D(net1151),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ));
 sg13g2_dlhq_1 _2925_ (.D(net1149),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ));
 sg13g2_dlhq_1 _2926_ (.D(net1211),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ));
 sg13g2_dlhq_1 _2927_ (.D(net1208),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ));
 sg13g2_dlhq_1 _2928_ (.D(net1206),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ));
 sg13g2_dlhq_1 _2929_ (.D(net1203),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ));
 sg13g2_dlhq_1 _2930_ (.D(net1202),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ));
 sg13g2_dlhq_1 _2931_ (.D(net1199),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ));
 sg13g2_dlhq_1 _2932_ (.D(net1196),
    .GATE(net1130),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ));
 sg13g2_dlhq_1 _2933_ (.D(net1195),
    .GATE(net1128),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ));
 sg13g2_dlhq_1 _2934_ (.D(net1192),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ));
 sg13g2_dlhq_1 _2935_ (.D(net1190),
    .GATE(net1129),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ));
 sg13g2_dlhq_1 _2936_ (.D(net1186),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ));
 sg13g2_dlhq_1 _2937_ (.D(net1184),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ));
 sg13g2_dlhq_1 _2938_ (.D(net1182),
    .GATE(net1130),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ));
 sg13g2_dlhq_1 _2939_ (.D(net1181),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ));
 sg13g2_dlhq_1 _2940_ (.D(net1178),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ));
 sg13g2_dlhq_1 _2941_ (.D(net1176),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ));
 sg13g2_dlhq_1 _2942_ (.D(net1174),
    .GATE(net27),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ));
 sg13g2_dlhq_1 _2943_ (.D(net1172),
    .GATE(net1130),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ));
 sg13g2_dlhq_1 _2944_ (.D(net1170),
    .GATE(net27),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ));
 sg13g2_dlhq_1 _2945_ (.D(net1168),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ));
 sg13g2_dlhq_1 _2946_ (.D(net1165),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ));
 sg13g2_dlhq_1 _2947_ (.D(net1163),
    .GATE(net1127),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ));
 sg13g2_dlhq_1 _2948_ (.D(net1213),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ));
 sg13g2_dlhq_1 _2949_ (.D(net1189),
    .GATE(net1136),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ));
 sg13g2_dlhq_1 _2950_ (.D(net1167),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ));
 sg13g2_dlhq_1 _2951_ (.D(net1161),
    .GATE(net1136),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ));
 sg13g2_dlhq_1 _2952_ (.D(net1158),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ));
 sg13g2_dlhq_1 _2953_ (.D(net1156),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ));
 sg13g2_dlhq_1 _2954_ (.D(net25),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ));
 sg13g2_dlhq_1 _2955_ (.D(net26),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ));
 sg13g2_dlhq_1 _2956_ (.D(net1150),
    .GATE(net1133),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ));
 sg13g2_dlhq_1 _2957_ (.D(net1148),
    .GATE(net1133),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ));
 sg13g2_dlhq_1 _2958_ (.D(net1210),
    .GATE(net1135),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ));
 sg13g2_dlhq_1 _2959_ (.D(net1208),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ));
 sg13g2_dlhq_1 _2960_ (.D(net1207),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ));
 sg13g2_dlhq_1 _2961_ (.D(net1203),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ));
 sg13g2_dlhq_1 _2962_ (.D(net1202),
    .GATE(net1135),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ));
 sg13g2_dlhq_1 _2963_ (.D(net1200),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ));
 sg13g2_dlhq_1 _2964_ (.D(net1197),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ));
 sg13g2_dlhq_1 _2965_ (.D(net1194),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ));
 sg13g2_dlhq_1 _2966_ (.D(net1193),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ));
 sg13g2_dlhq_1 _2967_ (.D(net1191),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ));
 sg13g2_dlhq_1 _2968_ (.D(net1186),
    .GATE(net1133),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ));
 sg13g2_dlhq_1 _2969_ (.D(net1184),
    .GATE(net1133),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ));
 sg13g2_dlhq_1 _2970_ (.D(net1183),
    .GATE(net1133),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ));
 sg13g2_dlhq_1 _2971_ (.D(net1180),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ));
 sg13g2_dlhq_1 _2972_ (.D(net1179),
    .GATE(net1132),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ));
 sg13g2_dlhq_1 _2973_ (.D(net1176),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ));
 sg13g2_dlhq_1 _2974_ (.D(net1174),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ));
 sg13g2_dlhq_1 _2975_ (.D(net1173),
    .GATE(net1134),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ));
 sg13g2_dlhq_1 _2976_ (.D(net1170),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ));
 sg13g2_dlhq_1 _2977_ (.D(net1168),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ));
 sg13g2_dlhq_1 _2978_ (.D(net1164),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ));
 sg13g2_dlhq_1 _2979_ (.D(net1162),
    .GATE(net1131),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ));
 sg13g2_dlhq_1 _2980_ (.D(net1212),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ));
 sg13g2_dlhq_1 _2981_ (.D(net1188),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ));
 sg13g2_dlhq_1 _2982_ (.D(net1166),
    .GATE(net1141),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ));
 sg13g2_dlhq_1 _2983_ (.D(net1161),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ));
 sg13g2_dlhq_1 _2984_ (.D(net1159),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ));
 sg13g2_dlhq_1 _2985_ (.D(net1157),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ));
 sg13g2_dlhq_1 _2986_ (.D(net1154),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ));
 sg13g2_dlhq_1 _2987_ (.D(net1152),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ));
 sg13g2_dlhq_1 _2988_ (.D(net1150),
    .GATE(net1140),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ));
 sg13g2_dlhq_1 _2989_ (.D(net1148),
    .GATE(net1140),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ));
 sg13g2_dlhq_1 _2990_ (.D(net1210),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ));
 sg13g2_dlhq_1 _2991_ (.D(net1209),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ));
 sg13g2_dlhq_1 _2992_ (.D(net1207),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ));
 sg13g2_dlhq_1 _2993_ (.D(net1205),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ));
 sg13g2_dlhq_1 _2994_ (.D(net1202),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ));
 sg13g2_dlhq_1 _2995_ (.D(net1198),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ));
 sg13g2_dlhq_1 _2996_ (.D(net1196),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ));
 sg13g2_dlhq_1 _2997_ (.D(net1194),
    .GATE(net1137),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ));
 sg13g2_dlhq_1 _2998_ (.D(net1193),
    .GATE(net1141),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ));
 sg13g2_dlhq_1 _2999_ (.D(net1191),
    .GATE(net1140),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ));
 sg13g2_dlhq_1 _3000_ (.D(net1187),
    .GATE(net1140),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ));
 sg13g2_dlhq_1 _3001_ (.D(net1185),
    .GATE(net1140),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ));
 sg13g2_dlhq_1 _3002_ (.D(net1182),
    .GATE(net1140),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ));
 sg13g2_dlhq_1 _3003_ (.D(net1180),
    .GATE(net1139),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ));
 sg13g2_dlhq_1 _3004_ (.D(net1178),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ));
 sg13g2_dlhq_1 _3005_ (.D(net1176),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ));
 sg13g2_dlhq_1 _3006_ (.D(net1175),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ));
 sg13g2_dlhq_1 _3007_ (.D(net1172),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ));
 sg13g2_dlhq_1 _3008_ (.D(net1171),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ));
 sg13g2_dlhq_1 _3009_ (.D(net1168),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ));
 sg13g2_dlhq_1 _3010_ (.D(net1164),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ));
 sg13g2_dlhq_1 _3011_ (.D(net1162),
    .GATE(net1138),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ));
 sg13g2_dlhq_1 _3012_ (.D(net1212),
    .GATE(net1079),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ));
 sg13g2_dlhq_1 _3013_ (.D(net1188),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ));
 sg13g2_dlhq_1 _3014_ (.D(net1166),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ));
 sg13g2_dlhq_1 _3015_ (.D(net1160),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ));
 sg13g2_dlhq_1 _3016_ (.D(net1158),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ));
 sg13g2_dlhq_1 _3017_ (.D(net1156),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ));
 sg13g2_dlhq_1 _3018_ (.D(net1155),
    .GATE(net1079),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ));
 sg13g2_dlhq_1 _3019_ (.D(net1153),
    .GATE(net1079),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ));
 sg13g2_dlhq_1 _3020_ (.D(net1151),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ));
 sg13g2_dlhq_1 _3021_ (.D(net1149),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ));
 sg13g2_dlhq_1 _3022_ (.D(net1211),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ));
 sg13g2_dlhq_1 _3023_ (.D(net1208),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ));
 sg13g2_dlhq_1 _3024_ (.D(net1206),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ));
 sg13g2_dlhq_1 _3025_ (.D(net1203),
    .GATE(net1079),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ));
 sg13g2_dlhq_1 _3026_ (.D(net1201),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ));
 sg13g2_dlhq_1 _3027_ (.D(net1199),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ));
 sg13g2_dlhq_1 _3028_ (.D(net1197),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ));
 sg13g2_dlhq_1 _3029_ (.D(net1194),
    .GATE(net1078),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ));
 sg13g2_dlhq_1 _3030_ (.D(net1192),
    .GATE(net1081),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ));
 sg13g2_dlhq_1 _3031_ (.D(net1190),
    .GATE(net1081),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ));
 sg13g2_dlhq_1 _3032_ (.D(net1187),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ));
 sg13g2_dlhq_1 _3033_ (.D(net1185),
    .GATE(net29),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ));
 sg13g2_dlhq_1 _3034_ (.D(net1182),
    .GATE(net1080),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _3035_ (.D(net1180),
    .GATE(net1080),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _3036_ (.D(net1179),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _3037_ (.D(net1176),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _3038_ (.D(net1175),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _3039_ (.D(net1172),
    .GATE(net1077),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _3040_ (.D(net1170),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _3041_ (.D(net1169),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _3042_ (.D(net1165),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _3043_ (.D(net1163),
    .GATE(net1082),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _3044_ (.D(net1213),
    .GATE(net1087),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _3045_ (.D(net1188),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _3046_ (.D(net1167),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _3047_ (.D(net1161),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _3048_ (.D(net1159),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _3049_ (.D(net1157),
    .GATE(net1085),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _3050_ (.D(net1154),
    .GATE(net1085),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _3051_ (.D(net1153),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _3052_ (.D(net1151),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _3053_ (.D(net1148),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _3054_ (.D(net1210),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _3055_ (.D(net1209),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _3056_ (.D(net1207),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _3057_ (.D(net1204),
    .GATE(net1086),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _3058_ (.D(net1201),
    .GATE(net1085),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _3059_ (.D(net1198),
    .GATE(net1085),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _3060_ (.D(net1196),
    .GATE(net1085),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _3061_ (.D(net1194),
    .GATE(net1085),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _3062_ (.D(net1193),
    .GATE(net1087),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _3063_ (.D(net1191),
    .GATE(net1087),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _3064_ (.D(net1186),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _3065_ (.D(net1184),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _3066_ (.D(net1182),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _3067_ (.D(net1180),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _3068_ (.D(net1178),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _3069_ (.D(net1176),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _3070_ (.D(net1174),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _3071_ (.D(net1173),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _3072_ (.D(net1170),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _3073_ (.D(net1168),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _3074_ (.D(net1164),
    .GATE(net1083),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _3075_ (.D(net1162),
    .GATE(net1084),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _3076_ (.D(net1213),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _3077_ (.D(net1189),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _3078_ (.D(net1166),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _3079_ (.D(net1160),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _3080_ (.D(net1158),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _3081_ (.D(net1156),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _3082_ (.D(net1154),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _3083_ (.D(net1152),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _3084_ (.D(net1150),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _3085_ (.D(net1148),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _3086_ (.D(net1210),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _3087_ (.D(net1208),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _3088_ (.D(net1207),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _3089_ (.D(net1204),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _3090_ (.D(net1201),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _3091_ (.D(net1198),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _3092_ (.D(net1196),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _3093_ (.D(net1195),
    .GATE(net1092),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _3094_ (.D(net1193),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _3095_ (.D(net1190),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _3096_ (.D(net1186),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _3097_ (.D(net1184),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _3098_ (.D(net1182),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _3099_ (.D(net1180),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _3100_ (.D(net1179),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _3101_ (.D(net1177),
    .GATE(net1090),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _3102_ (.D(net1174),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _3103_ (.D(net1173),
    .GATE(net1091),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _3104_ (.D(net1170),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _3105_ (.D(net1169),
    .GATE(net1089),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _3106_ (.D(net1164),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _3107_ (.D(net1162),
    .GATE(net1088),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _3108_ (.D(net1212),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _3109_ (.D(net1189),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _3110_ (.D(net1166),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _3111_ (.D(net1160),
    .GATE(net1097),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _3112_ (.D(net1159),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _3113_ (.D(net1157),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _3114_ (.D(net1155),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _3115_ (.D(net1152),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _3116_ (.D(net1150),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _3117_ (.D(net1148),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _3118_ (.D(net1211),
    .GATE(net1097),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _3119_ (.D(net1208),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _3120_ (.D(net1207),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _3121_ (.D(net1204),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _3122_ (.D(net1201),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _3123_ (.D(net1198),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _3124_ (.D(net1197),
    .GATE(net1097),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _3125_ (.D(net1195),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _3126_ (.D(net1192),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _3127_ (.D(net1190),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _3128_ (.D(net1186),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _3129_ (.D(net1185),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _3130_ (.D(net1182),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _3131_ (.D(net1180),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _3132_ (.D(net1179),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _3133_ (.D(net1177),
    .GATE(net1095),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _3134_ (.D(net1175),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _3135_ (.D(net1172),
    .GATE(net1094),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _3136_ (.D(net1170),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _3137_ (.D(net1169),
    .GATE(net1096),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _3138_ (.D(net1164),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _3139_ (.D(net1162),
    .GATE(net1093),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _3140_ (.D(net1213),
    .GATE(net28),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _3141_ (.D(net1189),
    .GATE(net1102),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _3142_ (.D(net1167),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _3143_ (.D(net1161),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _3144_ (.D(net1158),
    .GATE(net1099),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _3145_ (.D(net1156),
    .GATE(net1099),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _3146_ (.D(net1154),
    .GATE(net1099),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _3147_ (.D(net1152),
    .GATE(net1099),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _3148_ (.D(net1151),
    .GATE(net1102),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _3149_ (.D(net1149),
    .GATE(net1102),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _3150_ (.D(net1210),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _3151_ (.D(net1209),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _3152_ (.D(net1206),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _3153_ (.D(net1203),
    .GATE(net1099),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _3154_ (.D(net1201),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _3155_ (.D(net1198),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _3156_ (.D(net1196),
    .GATE(net1102),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _3157_ (.D(net1194),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _3158_ (.D(net1192),
    .GATE(net1101),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _3159_ (.D(net1190),
    .GATE(net1101),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _3160_ (.D(net1186),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _3161_ (.D(net1184),
    .GATE(net1099),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _3162_ (.D(net1182),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _3163_ (.D(net1180),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _3164_ (.D(net1178),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _3165_ (.D(net1177),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _3166_ (.D(net1174),
    .GATE(net1100),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _3167_ (.D(net1172),
    .GATE(net1101),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _3168_ (.D(net1171),
    .GATE(net1101),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _3169_ (.D(net1168),
    .GATE(net1101),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _3170_ (.D(net1164),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _3171_ (.D(net1162),
    .GATE(net1098),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _3172_ (.D(net1212),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _3173_ (.D(net1188),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _3174_ (.D(net1166),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _3175_ (.D(net1160),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _3176_ (.D(net1159),
    .GATE(net1104),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _3177_ (.D(net1157),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _3178_ (.D(net1155),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _3179_ (.D(net1153),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _3180_ (.D(net1150),
    .GATE(net1108),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _3181_ (.D(net1148),
    .GATE(net1108),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _3182_ (.D(net1210),
    .GATE(net1108),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _3183_ (.D(net1209),
    .GATE(net1108),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _3184_ (.D(net1206),
    .GATE(net1103),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _3185_ (.D(net1203),
    .GATE(net1104),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _3186_ (.D(net1202),
    .GATE(net1104),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _3187_ (.D(net1199),
    .GATE(net1104),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _3188_ (.D(net1196),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _3189_ (.D(net1195),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _3190_ (.D(net1192),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _3191_ (.D(net1190),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _3192_ (.D(net1186),
    .GATE(net1107),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _3193_ (.D(net1184),
    .GATE(net1107),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _3194_ (.D(net1183),
    .GATE(net1107),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _3195_ (.D(net1181),
    .GATE(net1107),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _3196_ (.D(net1178),
    .GATE(net1106),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _3197_ (.D(net1176),
    .GATE(net1106),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _3198_ (.D(net1175),
    .GATE(net1106),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _3199_ (.D(net1172),
    .GATE(net1106),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _3200_ (.D(net1171),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _3201_ (.D(net1168),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _3202_ (.D(net1164),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _3203_ (.D(net1163),
    .GATE(net1105),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _3204_ (.D(net1212),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _3205_ (.D(net1188),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _3206_ (.D(net1166),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _3207_ (.D(net1160),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _3208_ (.D(net1158),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _3209_ (.D(net1156),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _3210_ (.D(net1155),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _3211_ (.D(net1153),
    .GATE(net1109),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _3212_ (.D(net1150),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _3213_ (.D(net1148),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _3214_ (.D(net1211),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _3215_ (.D(net1209),
    .GATE(net1114),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _3216_ (.D(net1206),
    .GATE(net1110),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _3217_ (.D(net1203),
    .GATE(net1110),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _3218_ (.D(net1202),
    .GATE(net1110),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _3219_ (.D(net1199),
    .GATE(net1110),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _3220_ (.D(net1196),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _3221_ (.D(net1194),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _3222_ (.D(net1192),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _3223_ (.D(net1190),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _3224_ (.D(net1187),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _3225_ (.D(net1185),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _3226_ (.D(net1183),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _3227_ (.D(net1181),
    .GATE(net1112),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _3228_ (.D(net1178),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _3229_ (.D(net1176),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _3230_ (.D(net1175),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _3231_ (.D(net1172),
    .GATE(net1111),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _3232_ (.D(net1170),
    .GATE(net1113),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _3233_ (.D(net1169),
    .GATE(net1113),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _3234_ (.D(net1165),
    .GATE(net1113),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _3235_ (.D(net1163),
    .GATE(net1113),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _3236_ (.D(net1212),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _3237_ (.D(net1188),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _3238_ (.D(net1166),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _3239_ (.D(net1160),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _3240_ (.D(net1158),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _3241_ (.D(net1156),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _3242_ (.D(net1154),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _3243_ (.D(net1152),
    .GATE(net1115),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _3244_ (.D(net1151),
    .GATE(net1119),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _3245_ (.D(net1149),
    .GATE(net1119),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _3246_ (.D(net1211),
    .GATE(net1119),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _3247_ (.D(net1208),
    .GATE(net1119),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _3248_ (.D(net1206),
    .GATE(net1116),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _3249_ (.D(net1203),
    .GATE(net1116),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _3250_ (.D(net1201),
    .GATE(net1116),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _3251_ (.D(net1198),
    .GATE(net1116),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _3252_ (.D(net1196),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _3253_ (.D(net1194),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _3254_ (.D(net1193),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _3255_ (.D(net1191),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _3256_ (.D(net1187),
    .GATE(net1120),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _3257_ (.D(net1184),
    .GATE(net1120),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _3258_ (.D(net1183),
    .GATE(net1120),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _3259_ (.D(net1181),
    .GATE(net1120),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _3260_ (.D(net1178),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _3261_ (.D(net1176),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _3262_ (.D(net1174),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _3263_ (.D(net1172),
    .GATE(net1117),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _3264_ (.D(net1171),
    .GATE(net1118),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _3265_ (.D(net1168),
    .GATE(net1118),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _3266_ (.D(net1165),
    .GATE(net1118),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _3267_ (.D(net1163),
    .GATE(net1118),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _3268_ (.D(net1212),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _3269_ (.D(net1188),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _3270_ (.D(net1166),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _3271_ (.D(net1160),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _3272_ (.D(net1158),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _3273_ (.D(net1156),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _3274_ (.D(net1154),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _3275_ (.D(net1152),
    .GATE(net1121),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _3276_ (.D(net1151),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _3277_ (.D(net1149),
    .GATE(net1124),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _3278_ (.D(net1211),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _3279_ (.D(net1208),
    .GATE(net1124),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _3280_ (.D(net1206),
    .GATE(net1122),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _3281_ (.D(net1203),
    .GATE(net1122),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _3282_ (.D(net1201),
    .GATE(net1122),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _3283_ (.D(net1198),
    .GATE(net1122),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _3284_ (.D(net1197),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _3285_ (.D(net1194),
    .GATE(net1122),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _3286_ (.D(net1192),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _3287_ (.D(net1191),
    .GATE(net1125),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _3288_ (.D(net1187),
    .GATE(net1126),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _3289_ (.D(net1185),
    .GATE(net1126),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _3290_ (.D(net1183),
    .GATE(net1126),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _3291_ (.D(net1181),
    .GATE(net1126),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _3292_ (.D(net1178),
    .GATE(net1124),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _3293_ (.D(net1177),
    .GATE(net1124),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _3294_ (.D(net1175),
    .GATE(net1124),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _3295_ (.D(net1173),
    .GATE(net1124),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _3296_ (.D(net1171),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _3297_ (.D(net1168),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _3298_ (.D(net1165),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _3299_ (.D(net1162),
    .GATE(net1123),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _3300_ (.D(net1212),
    .GATE(net1146),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _3301_ (.D(net1188),
    .GATE(net1146),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _3302_ (.D(net1167),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _3303_ (.D(net1160),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _3304_ (.D(net1158),
    .GATE(net1143),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _3305_ (.D(net1156),
    .GATE(net1143),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _3306_ (.D(net1154),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _3307_ (.D(net1152),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _3308_ (.D(net1150),
    .GATE(net1145),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _3309_ (.D(net1149),
    .GATE(net1145),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _3310_ (.D(net1210),
    .GATE(net1147),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _3311_ (.D(net1208),
    .GATE(net1147),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _3312_ (.D(net1206),
    .GATE(net1143),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _3313_ (.D(net1204),
    .GATE(net1143),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _3314_ (.D(net1201),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _3315_ (.D(net1198),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _3316_ (.D(net1197),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _3317_ (.D(net1195),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _3318_ (.D(net1192),
    .GATE(net1146),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _3319_ (.D(net1190),
    .GATE(net1146),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _3320_ (.D(net1186),
    .GATE(net1143),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _3321_ (.D(net1184),
    .GATE(net1143),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _3322_ (.D(net1182),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _3323_ (.D(net1180),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _3324_ (.D(net1179),
    .GATE(net1145),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _3325_ (.D(net1177),
    .GATE(net1145),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _3326_ (.D(net1174),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _3327_ (.D(net1173),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _3328_ (.D(net1170),
    .GATE(net1146),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _3329_ (.D(net1169),
    .GATE(net1144),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _3330_ (.D(net1164),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _3331_ (.D(net1162),
    .GATE(net1142),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_dfrbp_1 _3332_ (.CLK(UserCLK),
    .RESET_B(net441),
    .D(\Inst_RegFile_32x4.BD_comb[0] ),
    .Q_N(_1367_),
    .Q(\Inst_RegFile_32x4.BD_reg[0] ));
 sg13g2_dfrbp_1 _3333_ (.CLK(UserCLK),
    .RESET_B(net442),
    .D(\Inst_RegFile_32x4.BD_comb[1] ),
    .Q_N(_1368_),
    .Q(\Inst_RegFile_32x4.BD_reg[1] ));
 sg13g2_dfrbp_1 _3334_ (.CLK(UserCLK),
    .RESET_B(net443),
    .D(\Inst_RegFile_32x4.BD_comb[2] ),
    .Q_N(_1369_),
    .Q(\Inst_RegFile_32x4.BD_reg[2] ));
 sg13g2_dfrbp_1 _3335_ (.CLK(UserCLK),
    .RESET_B(net444),
    .D(\Inst_RegFile_32x4.BD_comb[3] ),
    .Q_N(_1370_),
    .Q(\Inst_RegFile_32x4.BD_reg[3] ));
 sg13g2_dfrbp_1 _3336_ (.CLK(UserCLK),
    .RESET_B(net445),
    .D(\Inst_RegFile_32x4.AD_comb[0] ),
    .Q_N(_1371_),
    .Q(\Inst_RegFile_32x4.AD_reg[0] ));
 sg13g2_dfrbp_1 _3337_ (.CLK(UserCLK),
    .RESET_B(net446),
    .D(\Inst_RegFile_32x4.AD_comb[1] ),
    .Q_N(_1372_),
    .Q(\Inst_RegFile_32x4.AD_reg[1] ));
 sg13g2_dfrbp_1 _3338_ (.CLK(UserCLK),
    .RESET_B(net488),
    .D(\Inst_RegFile_32x4.AD_comb[2] ),
    .Q_N(_1373_),
    .Q(\Inst_RegFile_32x4.AD_reg[2] ));
 sg13g2_dfrbp_1 _3339_ (.CLK(UserCLK),
    .RESET_B(net405),
    .D(\Inst_RegFile_32x4.AD_comb[3] ),
    .Q_N(_1290_),
    .Q(\Inst_RegFile_32x4.AD_reg[3] ));
 sg13g2_dfrbp_1 _3340_ (.CLK(UserCLK),
    .RESET_B(net404),
    .D(_0076_),
    .Q_N(_1289_),
    .Q(\Inst_RegFile_32x4.mem[19][0] ));
 sg13g2_dfrbp_1 _3341_ (.CLK(UserCLK),
    .RESET_B(net403),
    .D(_0077_),
    .Q_N(_1288_),
    .Q(\Inst_RegFile_32x4.mem[19][1] ));
 sg13g2_dfrbp_1 _3342_ (.CLK(UserCLK),
    .RESET_B(net402),
    .D(_0078_),
    .Q_N(_1287_),
    .Q(\Inst_RegFile_32x4.mem[19][2] ));
 sg13g2_dfrbp_1 _3343_ (.CLK(UserCLK),
    .RESET_B(net401),
    .D(_0079_),
    .Q_N(_1286_),
    .Q(\Inst_RegFile_32x4.mem[19][3] ));
 sg13g2_dfrbp_1 _3344_ (.CLK(UserCLK),
    .RESET_B(net400),
    .D(_0080_),
    .Q_N(_1285_),
    .Q(\Inst_RegFile_32x4.mem[29][0] ));
 sg13g2_dfrbp_1 _3345_ (.CLK(UserCLK),
    .RESET_B(net399),
    .D(_0081_),
    .Q_N(_1284_),
    .Q(\Inst_RegFile_32x4.mem[29][1] ));
 sg13g2_dfrbp_1 _3346_ (.CLK(UserCLK),
    .RESET_B(net398),
    .D(_0082_),
    .Q_N(_1283_),
    .Q(\Inst_RegFile_32x4.mem[29][2] ));
 sg13g2_dfrbp_1 _3347_ (.CLK(UserCLK),
    .RESET_B(net397),
    .D(_0083_),
    .Q_N(_1282_),
    .Q(\Inst_RegFile_32x4.mem[29][3] ));
 sg13g2_dfrbp_1 _3348_ (.CLK(UserCLK),
    .RESET_B(net396),
    .D(_0084_),
    .Q_N(_1281_),
    .Q(\Inst_RegFile_32x4.mem[31][0] ));
 sg13g2_dfrbp_1 _3349_ (.CLK(UserCLK),
    .RESET_B(net395),
    .D(_0085_),
    .Q_N(_1280_),
    .Q(\Inst_RegFile_32x4.mem[31][1] ));
 sg13g2_dfrbp_1 _3350_ (.CLK(UserCLK),
    .RESET_B(net394),
    .D(_0086_),
    .Q_N(_1279_),
    .Q(\Inst_RegFile_32x4.mem[31][2] ));
 sg13g2_dfrbp_1 _3351_ (.CLK(UserCLK),
    .RESET_B(net393),
    .D(_0087_),
    .Q_N(_1278_),
    .Q(\Inst_RegFile_32x4.mem[31][3] ));
 sg13g2_dfrbp_1 _3352_ (.CLK(UserCLK),
    .RESET_B(net392),
    .D(_0088_),
    .Q_N(_1277_),
    .Q(\Inst_RegFile_32x4.mem[3][0] ));
 sg13g2_dfrbp_1 _3353_ (.CLK(UserCLK),
    .RESET_B(net391),
    .D(_0089_),
    .Q_N(_1276_),
    .Q(\Inst_RegFile_32x4.mem[3][1] ));
 sg13g2_dfrbp_1 _3354_ (.CLK(UserCLK),
    .RESET_B(net390),
    .D(_0090_),
    .Q_N(_1275_),
    .Q(\Inst_RegFile_32x4.mem[3][2] ));
 sg13g2_dfrbp_1 _3355_ (.CLK(UserCLK),
    .RESET_B(net389),
    .D(_0091_),
    .Q_N(_1274_),
    .Q(\Inst_RegFile_32x4.mem[3][3] ));
 sg13g2_dfrbp_1 _3356_ (.CLK(UserCLK),
    .RESET_B(net388),
    .D(_0092_),
    .Q_N(_1273_),
    .Q(\Inst_RegFile_32x4.mem[4][0] ));
 sg13g2_dfrbp_1 _3357_ (.CLK(UserCLK),
    .RESET_B(net387),
    .D(_0093_),
    .Q_N(_1272_),
    .Q(\Inst_RegFile_32x4.mem[4][1] ));
 sg13g2_dfrbp_1 _3358_ (.CLK(UserCLK),
    .RESET_B(net386),
    .D(_0094_),
    .Q_N(_1271_),
    .Q(\Inst_RegFile_32x4.mem[4][2] ));
 sg13g2_dfrbp_1 _3359_ (.CLK(UserCLK),
    .RESET_B(net385),
    .D(_0095_),
    .Q_N(_1270_),
    .Q(\Inst_RegFile_32x4.mem[4][3] ));
 sg13g2_dfrbp_1 _3360_ (.CLK(UserCLK),
    .RESET_B(net384),
    .D(_0096_),
    .Q_N(_1269_),
    .Q(\Inst_RegFile_32x4.mem[5][0] ));
 sg13g2_dfrbp_1 _3361_ (.CLK(UserCLK),
    .RESET_B(net383),
    .D(_0097_),
    .Q_N(_1268_),
    .Q(\Inst_RegFile_32x4.mem[5][1] ));
 sg13g2_dfrbp_1 _3362_ (.CLK(UserCLK),
    .RESET_B(net382),
    .D(_0098_),
    .Q_N(_1267_),
    .Q(\Inst_RegFile_32x4.mem[5][2] ));
 sg13g2_dfrbp_1 _3363_ (.CLK(UserCLK),
    .RESET_B(net381),
    .D(_0099_),
    .Q_N(_1266_),
    .Q(\Inst_RegFile_32x4.mem[5][3] ));
 sg13g2_dfrbp_1 _3364_ (.CLK(UserCLK),
    .RESET_B(net380),
    .D(_0100_),
    .Q_N(_1265_),
    .Q(\Inst_RegFile_32x4.mem[6][0] ));
 sg13g2_dfrbp_1 _3365_ (.CLK(UserCLK),
    .RESET_B(net379),
    .D(_0101_),
    .Q_N(_1264_),
    .Q(\Inst_RegFile_32x4.mem[6][1] ));
 sg13g2_dfrbp_1 _3366_ (.CLK(UserCLK),
    .RESET_B(net378),
    .D(_0102_),
    .Q_N(_1263_),
    .Q(\Inst_RegFile_32x4.mem[6][2] ));
 sg13g2_dfrbp_1 _3367_ (.CLK(UserCLK),
    .RESET_B(net377),
    .D(_0103_),
    .Q_N(_1262_),
    .Q(\Inst_RegFile_32x4.mem[6][3] ));
 sg13g2_dfrbp_1 _3368_ (.CLK(UserCLK),
    .RESET_B(net376),
    .D(_0104_),
    .Q_N(_1261_),
    .Q(\Inst_RegFile_32x4.mem[7][0] ));
 sg13g2_dfrbp_1 _3369_ (.CLK(UserCLK),
    .RESET_B(net375),
    .D(_0105_),
    .Q_N(_1260_),
    .Q(\Inst_RegFile_32x4.mem[7][1] ));
 sg13g2_dfrbp_1 _3370_ (.CLK(UserCLK),
    .RESET_B(net374),
    .D(_0106_),
    .Q_N(_1259_),
    .Q(\Inst_RegFile_32x4.mem[7][2] ));
 sg13g2_dfrbp_1 _3371_ (.CLK(UserCLK),
    .RESET_B(net373),
    .D(_0107_),
    .Q_N(_1258_),
    .Q(\Inst_RegFile_32x4.mem[7][3] ));
 sg13g2_dfrbp_1 _3372_ (.CLK(UserCLK),
    .RESET_B(net372),
    .D(_0108_),
    .Q_N(_1257_),
    .Q(\Inst_RegFile_32x4.mem[8][0] ));
 sg13g2_dfrbp_1 _3373_ (.CLK(UserCLK),
    .RESET_B(net371),
    .D(_0109_),
    .Q_N(_1256_),
    .Q(\Inst_RegFile_32x4.mem[8][1] ));
 sg13g2_dfrbp_1 _3374_ (.CLK(UserCLK),
    .RESET_B(net370),
    .D(_0110_),
    .Q_N(_1255_),
    .Q(\Inst_RegFile_32x4.mem[8][2] ));
 sg13g2_dfrbp_1 _3375_ (.CLK(UserCLK),
    .RESET_B(net369),
    .D(_0111_),
    .Q_N(_1254_),
    .Q(\Inst_RegFile_32x4.mem[8][3] ));
 sg13g2_dfrbp_1 _3376_ (.CLK(UserCLK),
    .RESET_B(net368),
    .D(_0112_),
    .Q_N(_1253_),
    .Q(\Inst_RegFile_32x4.mem[0][0] ));
 sg13g2_dfrbp_1 _3377_ (.CLK(UserCLK),
    .RESET_B(net367),
    .D(_0113_),
    .Q_N(_1252_),
    .Q(\Inst_RegFile_32x4.mem[0][1] ));
 sg13g2_dfrbp_1 _3378_ (.CLK(UserCLK),
    .RESET_B(net366),
    .D(_0114_),
    .Q_N(_1251_),
    .Q(\Inst_RegFile_32x4.mem[0][2] ));
 sg13g2_dfrbp_1 _3379_ (.CLK(UserCLK),
    .RESET_B(net365),
    .D(_0115_),
    .Q_N(_1250_),
    .Q(\Inst_RegFile_32x4.mem[0][3] ));
 sg13g2_dfrbp_1 _3380_ (.CLK(UserCLK),
    .RESET_B(net364),
    .D(_0116_),
    .Q_N(_1249_),
    .Q(\Inst_RegFile_32x4.mem[10][0] ));
 sg13g2_dfrbp_1 _3381_ (.CLK(UserCLK),
    .RESET_B(net363),
    .D(_0117_),
    .Q_N(_1248_),
    .Q(\Inst_RegFile_32x4.mem[10][1] ));
 sg13g2_dfrbp_1 _3382_ (.CLK(UserCLK),
    .RESET_B(net498),
    .D(_0118_),
    .Q_N(_1247_),
    .Q(\Inst_RegFile_32x4.mem[10][2] ));
 sg13g2_dfrbp_1 _3383_ (.CLK(UserCLK),
    .RESET_B(net497),
    .D(_0119_),
    .Q_N(_1246_),
    .Q(\Inst_RegFile_32x4.mem[10][3] ));
 sg13g2_dfrbp_1 _3384_ (.CLK(UserCLK),
    .RESET_B(net496),
    .D(_0120_),
    .Q_N(_1245_),
    .Q(\Inst_RegFile_32x4.mem[11][0] ));
 sg13g2_dfrbp_1 _3385_ (.CLK(UserCLK),
    .RESET_B(net495),
    .D(_0121_),
    .Q_N(_1244_),
    .Q(\Inst_RegFile_32x4.mem[11][1] ));
 sg13g2_dfrbp_1 _3386_ (.CLK(UserCLK),
    .RESET_B(net494),
    .D(_0122_),
    .Q_N(_1243_),
    .Q(\Inst_RegFile_32x4.mem[11][2] ));
 sg13g2_dfrbp_1 _3387_ (.CLK(UserCLK),
    .RESET_B(net493),
    .D(_0123_),
    .Q_N(_1242_),
    .Q(\Inst_RegFile_32x4.mem[11][3] ));
 sg13g2_dfrbp_1 _3388_ (.CLK(UserCLK),
    .RESET_B(net492),
    .D(_0124_),
    .Q_N(_1241_),
    .Q(\Inst_RegFile_32x4.mem[12][0] ));
 sg13g2_dfrbp_1 _3389_ (.CLK(UserCLK),
    .RESET_B(net491),
    .D(_0125_),
    .Q_N(_1240_),
    .Q(\Inst_RegFile_32x4.mem[12][1] ));
 sg13g2_dfrbp_1 _3390_ (.CLK(UserCLK),
    .RESET_B(net490),
    .D(_0126_),
    .Q_N(_1239_),
    .Q(\Inst_RegFile_32x4.mem[12][2] ));
 sg13g2_dfrbp_1 _3391_ (.CLK(UserCLK),
    .RESET_B(net489),
    .D(_0127_),
    .Q_N(_1238_),
    .Q(\Inst_RegFile_32x4.mem[12][3] ));
 sg13g2_tiehi _3380__364 (.L_HI(net364));
 sg13g2_tiehi _3379__365 (.L_HI(net365));
 sg13g2_tiehi _3378__366 (.L_HI(net366));
 sg13g2_tiehi _3377__367 (.L_HI(net367));
 sg13g2_tiehi _3376__368 (.L_HI(net368));
 sg13g2_tiehi _3375__369 (.L_HI(net369));
 sg13g2_tiehi _3374__370 (.L_HI(net370));
 sg13g2_tiehi _3373__371 (.L_HI(net371));
 sg13g2_tiehi _3372__372 (.L_HI(net372));
 sg13g2_tiehi _3371__373 (.L_HI(net373));
 sg13g2_tiehi _3370__374 (.L_HI(net374));
 sg13g2_tiehi _3369__375 (.L_HI(net375));
 sg13g2_tiehi _3368__376 (.L_HI(net376));
 sg13g2_tiehi _3367__377 (.L_HI(net377));
 sg13g2_tiehi _3366__378 (.L_HI(net378));
 sg13g2_tiehi _3365__379 (.L_HI(net379));
 sg13g2_tiehi _3364__380 (.L_HI(net380));
 sg13g2_tiehi _3363__381 (.L_HI(net381));
 sg13g2_tiehi _3362__382 (.L_HI(net382));
 sg13g2_tiehi _3361__383 (.L_HI(net383));
 sg13g2_tiehi _3360__384 (.L_HI(net384));
 sg13g2_tiehi _3359__385 (.L_HI(net385));
 sg13g2_tiehi _3358__386 (.L_HI(net386));
 sg13g2_tiehi _3357__387 (.L_HI(net387));
 sg13g2_tiehi _3356__388 (.L_HI(net388));
 sg13g2_tiehi _3355__389 (.L_HI(net389));
 sg13g2_tiehi _3354__390 (.L_HI(net390));
 sg13g2_tiehi _3353__391 (.L_HI(net391));
 sg13g2_tiehi _3352__392 (.L_HI(net392));
 sg13g2_tiehi _3351__393 (.L_HI(net393));
 sg13g2_tiehi _3350__394 (.L_HI(net394));
 sg13g2_tiehi _3349__395 (.L_HI(net395));
 sg13g2_tiehi _3348__396 (.L_HI(net396));
 sg13g2_tiehi _3347__397 (.L_HI(net397));
 sg13g2_tiehi _3346__398 (.L_HI(net398));
 sg13g2_tiehi _3345__399 (.L_HI(net399));
 sg13g2_tiehi _3344__400 (.L_HI(net400));
 sg13g2_tiehi _3343__401 (.L_HI(net401));
 sg13g2_tiehi _3342__402 (.L_HI(net402));
 sg13g2_tiehi _3341__403 (.L_HI(net403));
 sg13g2_tiehi _3340__404 (.L_HI(net404));
 sg13g2_tiehi _3339__405 (.L_HI(net405));
 sg13g2_tiehi _2916__406 (.L_HI(net406));
 sg13g2_tiehi _2915__407 (.L_HI(net407));
 sg13g2_tiehi _2914__408 (.L_HI(net408));
 sg13g2_tiehi _2913__409 (.L_HI(net409));
 sg13g2_tiehi _2912__410 (.L_HI(net410));
 sg13g2_tiehi _2911__411 (.L_HI(net411));
 sg13g2_tiehi _2910__412 (.L_HI(net412));
 sg13g2_tiehi _2909__413 (.L_HI(net413));
 sg13g2_tiehi _2908__414 (.L_HI(net414));
 sg13g2_tiehi _2907__415 (.L_HI(net415));
 sg13g2_tiehi _2906__416 (.L_HI(net416));
 sg13g2_tiehi _2905__417 (.L_HI(net417));
 sg13g2_tiehi _2904__418 (.L_HI(net418));
 sg13g2_tiehi _2903__419 (.L_HI(net419));
 sg13g2_tiehi _2902__420 (.L_HI(net420));
 sg13g2_tiehi _2901__421 (.L_HI(net421));
 sg13g2_tiehi _2900__422 (.L_HI(net422));
 sg13g2_tiehi _2899__423 (.L_HI(net423));
 sg13g2_tiehi _2898__424 (.L_HI(net424));
 sg13g2_tiehi _2897__425 (.L_HI(net425));
 sg13g2_tiehi _2896__426 (.L_HI(net426));
 sg13g2_tiehi _2895__427 (.L_HI(net427));
 sg13g2_tiehi _2894__428 (.L_HI(net428));
 sg13g2_tiehi _2893__429 (.L_HI(net429));
 sg13g2_tiehi _2892__430 (.L_HI(net430));
 sg13g2_tiehi _2891__431 (.L_HI(net431));
 sg13g2_tiehi _2890__432 (.L_HI(net432));
 sg13g2_tiehi _2889__433 (.L_HI(net433));
 sg13g2_tiehi _2888__434 (.L_HI(net434));
 sg13g2_tiehi _2887__435 (.L_HI(net435));
 sg13g2_tiehi _2886__436 (.L_HI(net436));
 sg13g2_tiehi _2885__437 (.L_HI(net437));
 sg13g2_tiehi _2884__438 (.L_HI(net438));
 sg13g2_tiehi _2842__439 (.L_HI(net439));
 sg13g2_tiehi _2917__440 (.L_HI(net440));
 sg13g2_tiehi _3332__441 (.L_HI(net441));
 sg13g2_tiehi _3333__442 (.L_HI(net442));
 sg13g2_tiehi _3334__443 (.L_HI(net443));
 sg13g2_tiehi _3335__444 (.L_HI(net444));
 sg13g2_tiehi _3336__445 (.L_HI(net445));
 sg13g2_tiehi _3337__446 (.L_HI(net446));
 sg13g2_tiehi _2883__447 (.L_HI(net447));
 sg13g2_tiehi _2882__448 (.L_HI(net448));
 sg13g2_tiehi _2881__449 (.L_HI(net449));
 sg13g2_tiehi _2880__450 (.L_HI(net450));
 sg13g2_tiehi _2879__451 (.L_HI(net451));
 sg13g2_tiehi _2878__452 (.L_HI(net452));
 sg13g2_tiehi _2877__453 (.L_HI(net453));
 sg13g2_tiehi _2876__454 (.L_HI(net454));
 sg13g2_tiehi _2875__455 (.L_HI(net455));
 sg13g2_tiehi _2874__456 (.L_HI(net456));
 sg13g2_tiehi _2873__457 (.L_HI(net457));
 sg13g2_tiehi _2872__458 (.L_HI(net458));
 sg13g2_tiehi _2871__459 (.L_HI(net459));
 sg13g2_tiehi _2870__460 (.L_HI(net460));
 sg13g2_tiehi _2869__461 (.L_HI(net461));
 sg13g2_tiehi _2868__462 (.L_HI(net462));
 sg13g2_tiehi _2867__463 (.L_HI(net463));
 sg13g2_tiehi _2866__464 (.L_HI(net464));
 sg13g2_tiehi _2865__465 (.L_HI(net465));
 sg13g2_tiehi _2864__466 (.L_HI(net466));
 sg13g2_tiehi _2863__467 (.L_HI(net467));
 sg13g2_tiehi _2862__468 (.L_HI(net468));
 sg13g2_tiehi _2861__469 (.L_HI(net469));
 sg13g2_tiehi _2860__470 (.L_HI(net470));
 sg13g2_tiehi _2859__471 (.L_HI(net471));
 sg13g2_tiehi _2858__472 (.L_HI(net472));
 sg13g2_tiehi _2857__473 (.L_HI(net473));
 sg13g2_tiehi _2856__474 (.L_HI(net474));
 sg13g2_tiehi _2855__475 (.L_HI(net475));
 sg13g2_tiehi _2854__476 (.L_HI(net476));
 sg13g2_tiehi _2853__477 (.L_HI(net477));
 sg13g2_tiehi _2852__478 (.L_HI(net478));
 sg13g2_tiehi _2851__479 (.L_HI(net479));
 sg13g2_tiehi _2850__480 (.L_HI(net480));
 sg13g2_tiehi _2849__481 (.L_HI(net481));
 sg13g2_tiehi _2848__482 (.L_HI(net482));
 sg13g2_tiehi _2847__483 (.L_HI(net483));
 sg13g2_tiehi _2846__484 (.L_HI(net484));
 sg13g2_tiehi _2845__485 (.L_HI(net485));
 sg13g2_tiehi _2844__486 (.L_HI(net486));
 sg13g2_tiehi _2843__487 (.L_HI(net487));
 sg13g2_tiehi _3338__488 (.L_HI(net488));
 sg13g2_tiehi _3391__489 (.L_HI(net489));
 sg13g2_tiehi _3390__490 (.L_HI(net490));
 sg13g2_tiehi _3389__491 (.L_HI(net491));
 sg13g2_tiehi _3388__492 (.L_HI(net492));
 sg13g2_tiehi _3387__493 (.L_HI(net493));
 sg13g2_tiehi _3386__494 (.L_HI(net494));
 sg13g2_tiehi _3385__495 (.L_HI(net495));
 sg13g2_tiehi _3384__496 (.L_HI(net496));
 sg13g2_tiehi _3383__497 (.L_HI(net497));
 sg13g2_tiehi _3382__498 (.L_HI(net498));
 sg13g2_dlygate4sd1_1 rebuffer1 (.A(_1229_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold241 (.A(\Inst_RegFile_32x4.mem[0][0] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold238 (.A(\Inst_RegFile_32x4.mem[15][3] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold231 (.A(\Inst_RegFile_32x4.mem[6][2] ),
    .X(net729));
 sg13g2_buf_2 rebuffer33 (.A(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .X(net531));
 sg13g2_buf_2 _3532_ (.A(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .X(net114));
 sg13g2_buf_2 _3533_ (.A(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .X(net115));
 sg13g2_buf_2 _3534_ (.A(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .X(net116));
 sg13g2_buf_8 _3535_ (.A(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .X(net117));
 sg13g2_buf_1 _3536_ (.A(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .X(net118));
 sg13g2_buf_8 _3537_ (.A(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .X(net119));
 sg13g2_buf_1 _3538_ (.A(\Inst_RegFile_switch_matrix.E2BEG6 ),
    .X(net120));
 sg13g2_buf_2 _3539_ (.A(\Inst_RegFile_switch_matrix.E2BEG7 ),
    .X(net121));
 sg13g2_buf_1 _3540_ (.A(net13),
    .X(net122));
 sg13g2_buf_1 _3541_ (.A(net14),
    .X(net123));
 sg13g2_buf_1 _3542_ (.A(net15),
    .X(net124));
 sg13g2_buf_1 _3543_ (.A(net16),
    .X(net125));
 sg13g2_buf_1 _3544_ (.A(net17),
    .X(net126));
 sg13g2_buf_1 _3545_ (.A(net18),
    .X(net127));
 sg13g2_buf_1 _3546_ (.A(net19),
    .X(net128));
 sg13g2_buf_1 _3547_ (.A(net20),
    .X(net129));
 sg13g2_buf_1 _3548_ (.A(E6END[2]),
    .X(net130));
 sg13g2_buf_1 _3549_ (.A(E6END[3]),
    .X(net133));
 sg13g2_buf_1 _3550_ (.A(E6END[4]),
    .X(net134));
 sg13g2_buf_1 _3551_ (.A(E6END[5]),
    .X(net135));
 sg13g2_buf_1 _3552_ (.A(E6END[6]),
    .X(net136));
 sg13g2_buf_1 _3553_ (.A(E6END[7]),
    .X(net137));
 sg13g2_buf_1 _3554_ (.A(E6END[8]),
    .X(net138));
 sg13g2_buf_1 _3555_ (.A(E6END[9]),
    .X(net139));
 sg13g2_buf_1 _3556_ (.A(E6END[10]),
    .X(net140));
 sg13g2_buf_1 _3557_ (.A(E6END[11]),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold226 (.A(\Inst_RegFile_32x4.mem[6][0] ),
    .X(net724));
 sg13g2_buf_2 rebuffer27 (.A(AD2),
    .X(net525));
 sg13g2_buf_1 _3560_ (.A(EE4END[4]),
    .X(net142));
 sg13g2_buf_1 _3561_ (.A(EE4END[5]),
    .X(net149));
 sg13g2_buf_1 _3562_ (.A(EE4END[6]),
    .X(net150));
 sg13g2_buf_1 _3563_ (.A(EE4END[7]),
    .X(net151));
 sg13g2_buf_1 _3564_ (.A(EE4END[8]),
    .X(net152));
 sg13g2_buf_1 _3565_ (.A(EE4END[9]),
    .X(net153));
 sg13g2_buf_1 _3566_ (.A(EE4END[10]),
    .X(net154));
 sg13g2_buf_1 _3567_ (.A(EE4END[11]),
    .X(net155));
 sg13g2_buf_1 _3568_ (.A(EE4END[12]),
    .X(net156));
 sg13g2_buf_1 _3569_ (.A(EE4END[13]),
    .X(net157));
 sg13g2_buf_1 _3570_ (.A(EE4END[14]),
    .X(net143));
 sg13g2_buf_1 _3571_ (.A(EE4END[15]),
    .X(net144));
 sg13g2_dlygate4sd1_1 rebuffer224 (.A(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold239 (.A(\Inst_RegFile_32x4.mem[6][3] ),
    .X(net737));
 sg13g2_buf_2 _3574_ (.A(\Inst_RegFile_switch_matrix.EE4BEG2 ),
    .X(net147));
 sg13g2_buf_1 _3575_ (.A(\Inst_RegFile_switch_matrix.EE4BEG3 ),
    .X(net148));
 sg13g2_buf_1 _3576_ (.A(net1213),
    .X(net158));
 sg13g2_buf_1 _3577_ (.A(net1189),
    .X(net169));
 sg13g2_buf_1 _3578_ (.A(net1167),
    .X(net180));
 sg13g2_buf_1 _3579_ (.A(net1161),
    .X(net183));
 sg13g2_buf_1 _3580_ (.A(net1159),
    .X(net184));
 sg13g2_buf_1 _3581_ (.A(net1157),
    .X(net185));
 sg13g2_buf_1 _3582_ (.A(net25),
    .X(net186));
 sg13g2_buf_1 _3583_ (.A(net26),
    .X(net187));
 sg13g2_buf_1 _3584_ (.A(net1150),
    .X(net188));
 sg13g2_buf_1 _3585_ (.A(net1148),
    .X(net189));
 sg13g2_buf_1 _3586_ (.A(net1210),
    .X(net159));
 sg13g2_buf_1 _3587_ (.A(net1209),
    .X(net160));
 sg13g2_buf_1 _3588_ (.A(net1207),
    .X(net161));
 sg13g2_buf_1 _3589_ (.A(net1205),
    .X(net162));
 sg13g2_buf_1 _3590_ (.A(net1202),
    .X(net163));
 sg13g2_buf_1 _3591_ (.A(net1200),
    .X(net164));
 sg13g2_buf_1 _3592_ (.A(net1197),
    .X(net165));
 sg13g2_buf_1 _3593_ (.A(net1195),
    .X(net166));
 sg13g2_buf_1 _3594_ (.A(net1193),
    .X(net167));
 sg13g2_buf_1 _3595_ (.A(net1191),
    .X(net168));
 sg13g2_buf_1 _3596_ (.A(net1187),
    .X(net170));
 sg13g2_buf_1 _3597_ (.A(net1185),
    .X(net171));
 sg13g2_buf_1 _3598_ (.A(net1183),
    .X(net172));
 sg13g2_buf_1 _3599_ (.A(net1181),
    .X(net173));
 sg13g2_buf_1 _3600_ (.A(net1179),
    .X(net174));
 sg13g2_buf_1 _3601_ (.A(net1177),
    .X(net175));
 sg13g2_buf_1 _3602_ (.A(net1174),
    .X(net176));
 sg13g2_buf_1 _3603_ (.A(net1173),
    .X(net177));
 sg13g2_buf_1 _3604_ (.A(net1171),
    .X(net178));
 sg13g2_buf_1 _3605_ (.A(net1169),
    .X(net179));
 sg13g2_buf_1 _3606_ (.A(net1165),
    .X(net181));
 sg13g2_buf_1 _3607_ (.A(net1163),
    .X(net182));
 sg13g2_buf_1 _3608_ (.A(net1144),
    .X(net190));
 sg13g2_buf_1 _3609_ (.A(net1126),
    .X(net201));
 sg13g2_buf_1 _3610_ (.A(net1120),
    .X(net202));
 sg13g2_buf_1 _3611_ (.A(net1112),
    .X(net203));
 sg13g2_buf_1 _3612_ (.A(net1108),
    .X(net204));
 sg13g2_buf_1 _3613_ (.A(net1102),
    .X(net205));
 sg13g2_buf_1 _3614_ (.A(net1095),
    .X(net206));
 sg13g2_buf_1 _3615_ (.A(net1090),
    .X(net207));
 sg13g2_buf_1 _3616_ (.A(net1087),
    .X(net208));
 sg13g2_buf_1 _3617_ (.A(net1082),
    .X(net209));
 sg13g2_buf_1 _3618_ (.A(net1140),
    .X(net191));
 sg13g2_buf_1 _3619_ (.A(net1134),
    .X(net192));
 sg13g2_buf_1 _3620_ (.A(net1130),
    .X(net193));
 sg13g2_buf_1 _3621_ (.A(FrameStrobe[13]),
    .X(net194));
 sg13g2_buf_1 _3622_ (.A(FrameStrobe[14]),
    .X(net195));
 sg13g2_buf_1 _3623_ (.A(FrameStrobe[15]),
    .X(net196));
 sg13g2_buf_1 _3624_ (.A(FrameStrobe[16]),
    .X(net197));
 sg13g2_buf_1 _3625_ (.A(FrameStrobe[17]),
    .X(net198));
 sg13g2_buf_1 _3626_ (.A(FrameStrobe[18]),
    .X(net199));
 sg13g2_buf_1 _3627_ (.A(FrameStrobe[19]),
    .X(net200));
 sg13g2_buf_8 _3628_ (.A(\Inst_RegFile_switch_matrix.N1BEG0 ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold244 (.A(\Inst_RegFile_32x4.mem[0][2] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold236 (.A(\Inst_RegFile_32x4.mem[4][2] ),
    .X(net734));
 sg13g2_dlygate4sd1_1 rebuffer28 (.A(net528),
    .X(net526));
 sg13g2_buf_8 _3632_ (.A(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .X(net214));
 sg13g2_buf_2 _3633_ (.A(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .X(net215));
 sg13g2_buf_8 _3634_ (.A(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .X(net216));
 sg13g2_buf_1 _3635_ (.A(net717),
    .X(net217));
 sg13g2_buf_1 _3636_ (.A(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .X(net218));
 sg13g2_dlygate4sd1_1 rebuffer225 (.A(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold230 (.A(\Inst_RegFile_32x4.mem[2][1] ),
    .X(net728));
 sg13g2_buf_1 _3639_ (.A(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .X(net221));
 sg13g2_buf_1 _3640_ (.A(net42),
    .X(net222));
 sg13g2_buf_1 _3641_ (.A(net43),
    .X(net223));
 sg13g2_buf_1 _3642_ (.A(net44),
    .X(net224));
 sg13g2_buf_1 _3643_ (.A(net45),
    .X(net225));
 sg13g2_buf_1 _3644_ (.A(net46),
    .X(net226));
 sg13g2_buf_1 _3645_ (.A(net47),
    .X(net227));
 sg13g2_buf_1 _3646_ (.A(net48),
    .X(net228));
 sg13g2_buf_1 _3647_ (.A(net49),
    .X(net229));
 sg13g2_buf_1 _3648_ (.A(N4END[4]),
    .X(net230));
 sg13g2_buf_1 _3649_ (.A(N4END[5]),
    .X(net237));
 sg13g2_buf_1 _3650_ (.A(N4END[6]),
    .X(net238));
 sg13g2_buf_1 _3651_ (.A(N4END[7]),
    .X(net239));
 sg13g2_buf_1 _3652_ (.A(N4END[8]),
    .X(net240));
 sg13g2_buf_1 _3653_ (.A(N4END[9]),
    .X(net241));
 sg13g2_buf_1 _3654_ (.A(N4END[10]),
    .X(net242));
 sg13g2_buf_1 _3655_ (.A(N4END[11]),
    .X(net243));
 sg13g2_buf_1 _3656_ (.A(N4END[12]),
    .X(net244));
 sg13g2_buf_1 _3657_ (.A(N4END[13]),
    .X(net245));
 sg13g2_buf_1 _3658_ (.A(N4END[14]),
    .X(net231));
 sg13g2_buf_1 _3659_ (.A(N4END[15]),
    .X(net232));
 sg13g2_buf_1 _3660_ (.A(\Inst_RegFile_switch_matrix.N4BEG0 ),
    .X(net233));
 sg13g2_buf_1 _3661_ (.A(\Inst_RegFile_switch_matrix.N4BEG1 ),
    .X(net234));
 sg13g2_buf_1 _3662_ (.A(\Inst_RegFile_switch_matrix.N4BEG2 ),
    .X(net235));
 sg13g2_buf_1 _3663_ (.A(\Inst_RegFile_switch_matrix.N4BEG3 ),
    .X(net236));
 sg13g2_buf_1 _3664_ (.A(NN4END[4]),
    .X(net246));
 sg13g2_buf_1 _3665_ (.A(NN4END[5]),
    .X(net253));
 sg13g2_buf_1 _3666_ (.A(NN4END[6]),
    .X(net254));
 sg13g2_buf_1 _3667_ (.A(NN4END[7]),
    .X(net255));
 sg13g2_buf_1 _3668_ (.A(NN4END[8]),
    .X(net256));
 sg13g2_buf_1 _3669_ (.A(NN4END[9]),
    .X(net257));
 sg13g2_buf_1 _3670_ (.A(NN4END[10]),
    .X(net258));
 sg13g2_buf_1 _3671_ (.A(NN4END[11]),
    .X(net259));
 sg13g2_buf_1 _3672_ (.A(NN4END[12]),
    .X(net260));
 sg13g2_buf_1 _3673_ (.A(NN4END[13]),
    .X(net261));
 sg13g2_buf_1 _3674_ (.A(NN4END[14]),
    .X(net247));
 sg13g2_buf_1 _3675_ (.A(NN4END[15]),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold227 (.A(\Inst_RegFile_32x4.mem[10][2] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold234 (.A(\Inst_RegFile_32x4.mem[4][1] ),
    .X(net732));
 sg13g2_buf_1 _3678_ (.A(\Inst_RegFile_switch_matrix.NN4BEG2 ),
    .X(net251));
 sg13g2_buf_1 _3679_ (.A(\Inst_RegFile_switch_matrix.NN4BEG3 ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold243 (.A(\Inst_RegFile_32x4.mem[13][3] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold229 (.A(\Inst_RegFile_32x4.mem[4][3] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold233 (.A(\Inst_RegFile_32x4.mem[8][0] ),
    .X(net731));
 sg13g2_dlygate4sd1_1 rebuffer29 (.A(net529),
    .X(net527));
 sg13g2_buf_1 _3684_ (.A(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .X(net266));
 sg13g2_buf_1 _3685_ (.A(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .X(net267));
 sg13g2_buf_2 _3686_ (.A(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .X(net268));
 sg13g2_buf_1 _3687_ (.A(net511),
    .X(net269));
 sg13g2_buf_1 _3688_ (.A(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .X(net270));
 sg13g2_buf_1 _3689_ (.A(net501),
    .X(net271));
 sg13g2_buf_1 _3690_ (.A(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .X(net272));
 sg13g2_buf_8 _3691_ (.A(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .X(net273));
 sg13g2_buf_1 _3692_ (.A(net70),
    .X(net274));
 sg13g2_buf_1 _3693_ (.A(net71),
    .X(net275));
 sg13g2_buf_1 _3694_ (.A(net72),
    .X(net276));
 sg13g2_buf_1 _3695_ (.A(net73),
    .X(net277));
 sg13g2_buf_1 _3696_ (.A(net74),
    .X(net278));
 sg13g2_buf_1 _3697_ (.A(net75),
    .X(net279));
 sg13g2_buf_1 _3698_ (.A(net76),
    .X(net280));
 sg13g2_buf_1 _3699_ (.A(net77),
    .X(net281));
 sg13g2_buf_1 _3700_ (.A(S4END[4]),
    .X(net282));
 sg13g2_buf_1 _3701_ (.A(S4END[5]),
    .X(net289));
 sg13g2_buf_1 _3702_ (.A(S4END[6]),
    .X(net290));
 sg13g2_buf_1 _3703_ (.A(S4END[7]),
    .X(net291));
 sg13g2_buf_1 _3704_ (.A(S4END[8]),
    .X(net292));
 sg13g2_buf_1 _3705_ (.A(S4END[9]),
    .X(net293));
 sg13g2_buf_1 _3706_ (.A(S4END[10]),
    .X(net294));
 sg13g2_buf_1 _3707_ (.A(S4END[11]),
    .X(net295));
 sg13g2_buf_1 _3708_ (.A(S4END[12]),
    .X(net296));
 sg13g2_buf_1 _3709_ (.A(S4END[13]),
    .X(net297));
 sg13g2_buf_1 _3710_ (.A(S4END[14]),
    .X(net283));
 sg13g2_buf_1 _3711_ (.A(S4END[15]),
    .X(net284));
 sg13g2_buf_1 _3712_ (.A(\Inst_RegFile_switch_matrix.S4BEG0 ),
    .X(net285));
 sg13g2_buf_1 _3713_ (.A(\Inst_RegFile_switch_matrix.S4BEG1 ),
    .X(net286));
 sg13g2_buf_1 _3714_ (.A(\Inst_RegFile_switch_matrix.S4BEG2 ),
    .X(net287));
 sg13g2_buf_1 _3715_ (.A(\Inst_RegFile_switch_matrix.S4BEG3 ),
    .X(net288));
 sg13g2_buf_1 _3716_ (.A(SS4END[4]),
    .X(net298));
 sg13g2_buf_1 _3717_ (.A(SS4END[5]),
    .X(net305));
 sg13g2_buf_1 _3718_ (.A(SS4END[6]),
    .X(net306));
 sg13g2_buf_1 _3719_ (.A(SS4END[7]),
    .X(net307));
 sg13g2_buf_1 _3720_ (.A(SS4END[8]),
    .X(net308));
 sg13g2_buf_1 _3721_ (.A(SS4END[9]),
    .X(net309));
 sg13g2_buf_1 _3722_ (.A(SS4END[10]),
    .X(net310));
 sg13g2_buf_1 _3723_ (.A(SS4END[11]),
    .X(net311));
 sg13g2_buf_1 _3724_ (.A(SS4END[12]),
    .X(net312));
 sg13g2_buf_1 _3725_ (.A(SS4END[13]),
    .X(net313));
 sg13g2_buf_1 _3726_ (.A(SS4END[14]),
    .X(net299));
 sg13g2_buf_1 _3727_ (.A(SS4END[15]),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold228 (.A(\Inst_RegFile_32x4.mem[4][0] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold240 (.A(\Inst_RegFile_32x4.mem[2][0] ),
    .X(net738));
 sg13g2_buf_8 _3730_ (.A(\Inst_RegFile_switch_matrix.SS4BEG2 ),
    .X(net303));
 sg13g2_buf_1 _3731_ (.A(\Inst_RegFile_switch_matrix.SS4BEG3 ),
    .X(net304));
 sg13g2_buf_1 _3732_ (.A(UserCLK),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold242 (.A(\Inst_RegFile_32x4.mem[13][0] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold237 (.A(\Inst_RegFile_32x4.mem[0][1] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold232 (.A(\Inst_RegFile_32x4.mem[8][2] ),
    .X(net730));
 sg13g2_dlygate4sd1_1 rebuffer30 (.A(net530),
    .X(net528));
 sg13g2_buf_1 _3737_ (.A(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .X(net319));
 sg13g2_buf_1 _3738_ (.A(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .X(net320));
 sg13g2_buf_1 _3739_ (.A(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .X(net321));
 sg13g2_dlygate4sd1_1 rebuffer223 (.A(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .X(net721));
 sg13g2_buf_1 _3741_ (.A(net523),
    .X(net323));
 sg13g2_buf_2 _3742_ (.A(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .X(net324));
 sg13g2_buf_8 _3743_ (.A(net722),
    .X(net325));
 sg13g2_buf_2 _3744_ (.A(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .X(net326));
 sg13g2_buf_1 _3745_ (.A(net97),
    .X(net327));
 sg13g2_buf_1 _3746_ (.A(net98),
    .X(net328));
 sg13g2_buf_1 _3747_ (.A(net99),
    .X(net329));
 sg13g2_buf_1 _3748_ (.A(net100),
    .X(net330));
 sg13g2_buf_1 _3749_ (.A(net101),
    .X(net331));
 sg13g2_buf_1 _3750_ (.A(net102),
    .X(net332));
 sg13g2_buf_1 _3751_ (.A(net103),
    .X(net333));
 sg13g2_buf_1 _3752_ (.A(net104),
    .X(net334));
 sg13g2_buf_1 _3753_ (.A(W6END[2]),
    .X(net335));
 sg13g2_buf_1 _3754_ (.A(W6END[3]),
    .X(net338));
 sg13g2_buf_1 _3755_ (.A(W6END[4]),
    .X(net339));
 sg13g2_buf_1 _3756_ (.A(W6END[5]),
    .X(net340));
 sg13g2_buf_1 _3757_ (.A(W6END[6]),
    .X(net341));
 sg13g2_buf_1 _3758_ (.A(W6END[7]),
    .X(net342));
 sg13g2_buf_1 _3759_ (.A(W6END[8]),
    .X(net343));
 sg13g2_buf_1 _3760_ (.A(W6END[9]),
    .X(net344));
 sg13g2_buf_1 _3761_ (.A(W6END[10]),
    .X(net345));
 sg13g2_buf_1 _3762_ (.A(W6END[11]),
    .X(net346));
 sg13g2_buf_1 _3763_ (.A(\Inst_RegFile_switch_matrix.W6BEG0 ),
    .X(net336));
 sg13g2_buf_2 rebuffer31 (.A(net531),
    .X(net529));
 sg13g2_buf_1 _3765_ (.A(WW4END[4]),
    .X(net347));
 sg13g2_buf_1 _3766_ (.A(WW4END[5]),
    .X(net354));
 sg13g2_buf_1 _3767_ (.A(WW4END[6]),
    .X(net355));
 sg13g2_buf_1 _3768_ (.A(WW4END[7]),
    .X(net356));
 sg13g2_buf_1 _3769_ (.A(WW4END[8]),
    .X(net357));
 sg13g2_buf_1 _3770_ (.A(WW4END[9]),
    .X(net358));
 sg13g2_buf_1 _3771_ (.A(WW4END[10]),
    .X(net359));
 sg13g2_buf_1 _3772_ (.A(WW4END[11]),
    .X(net360));
 sg13g2_buf_1 _3773_ (.A(WW4END[12]),
    .X(net361));
 sg13g2_buf_1 _3774_ (.A(WW4END[13]),
    .X(net362));
 sg13g2_buf_1 _3775_ (.A(WW4END[14]),
    .X(net348));
 sg13g2_buf_1 _3776_ (.A(WW4END[15]),
    .X(net349));
 sg13g2_buf_1 _3777_ (.A(\Inst_RegFile_switch_matrix.WW4BEG0 ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold235 (.A(\Inst_RegFile_32x4.mem[2][3] ),
    .X(net733));
 sg13g2_buf_1 _3779_ (.A(\Inst_RegFile_switch_matrix.WW4BEG2 ),
    .X(net352));
 sg13g2_buf_1 _3780_ (.A(\Inst_RegFile_switch_matrix.WW4BEG3 ),
    .X(net353));
 sg13g2_buf_16 fanout921 (.X(net921),
    .A(net922));
 sg13g2_buf_8 fanout922 (.A(A_ADR0),
    .X(net922));
 sg13g2_buf_1 fanout923 (.A(net925),
    .X(net923));
 sg13g2_buf_1 fanout924 (.A(net925),
    .X(net924));
 sg13g2_buf_1 fanout925 (.A(net927),
    .X(net925));
 sg13g2_buf_1 fanout926 (.A(net927),
    .X(net926));
 sg13g2_buf_1 fanout927 (.A(A_ADR0),
    .X(net927));
 sg13g2_buf_1 fanout928 (.A(net931),
    .X(net928));
 sg13g2_buf_1 fanout929 (.A(net930),
    .X(net929));
 sg13g2_buf_1 fanout930 (.A(net931),
    .X(net930));
 sg13g2_buf_1 fanout931 (.A(A_ADR0),
    .X(net931));
 sg13g2_buf_8 fanout932 (.A(net933),
    .X(net932));
 sg13g2_buf_8 fanout933 (.A(net936),
    .X(net933));
 sg13g2_buf_1 fanout934 (.A(net936),
    .X(net934));
 sg13g2_buf_1 fanout935 (.A(net936),
    .X(net935));
 sg13g2_buf_2 fanout936 (.A(_1087_),
    .X(net936));
 sg13g2_buf_1 fanout937 (.A(net938),
    .X(net937));
 sg13g2_buf_1 fanout938 (.A(net939),
    .X(net938));
 sg13g2_buf_1 fanout939 (.A(_1065_),
    .X(net939));
 sg13g2_buf_1 fanout940 (.A(net942),
    .X(net940));
 sg13g2_buf_1 fanout941 (.A(net942),
    .X(net941));
 sg13g2_buf_1 fanout942 (.A(_1065_),
    .X(net942));
 sg13g2_buf_8 fanout943 (.A(_0460_),
    .X(net943));
 sg13g2_buf_1 fanout944 (.A(net946),
    .X(net944));
 sg13g2_buf_1 fanout945 (.A(net946),
    .X(net945));
 sg13g2_buf_1 fanout946 (.A(_0368_),
    .X(net946));
 sg13g2_buf_1 fanout947 (.A(net948),
    .X(net947));
 sg13g2_buf_1 fanout948 (.A(_0368_),
    .X(net948));
 sg13g2_buf_1 fanout949 (.A(net951),
    .X(net949));
 sg13g2_buf_1 fanout950 (.A(net951),
    .X(net950));
 sg13g2_buf_1 fanout951 (.A(net954),
    .X(net951));
 sg13g2_buf_1 fanout952 (.A(net954),
    .X(net952));
 sg13g2_buf_1 fanout953 (.A(net954),
    .X(net953));
 sg13g2_buf_1 fanout954 (.A(_1067_),
    .X(net954));
 sg13g2_buf_1 fanout955 (.A(_0143_),
    .X(net955));
 sg13g2_buf_1 fanout956 (.A(_0143_),
    .X(net956));
 sg13g2_buf_2 rebuffer32 (.A(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .X(net530));
 sg13g2_buf_1 fanout958 (.A(net962),
    .X(net958));
 sg13g2_buf_1 fanout959 (.A(net962),
    .X(net959));
 sg13g2_buf_1 fanout960 (.A(net962),
    .X(net960));
 sg13g2_buf_1 fanout961 (.A(net962),
    .X(net961));
 sg13g2_buf_1 fanout962 (.A(_1069_),
    .X(net962));
 sg13g2_buf_8 fanout963 (.A(net504),
    .X(net963));
 sg13g2_dlygate4sd1_1 rebuffer13 (.A(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .X(net511));
 sg13g2_buf_16 fanout965 (.X(net965),
    .A(net513));
 sg13g2_buf_1 fanout966 (.A(net513),
    .X(net966));
 sg13g2_buf_1 fanout967 (.A(net513),
    .X(net967));
 sg13g2_dlygate4sd1_1 rebuffer5 (.A(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .X(net503));
 sg13g2_buf_8 fanout969 (.A(net520),
    .X(net969));
 sg13g2_buf_1 fanout970 (.A(net973),
    .X(net970));
 sg13g2_buf_1 fanout971 (.A(net972),
    .X(net971));
 sg13g2_buf_1 fanout972 (.A(net973),
    .X(net972));
 sg13g2_buf_8 fanout973 (.A(AD3),
    .X(net973));
 sg13g2_buf_16 fanout974 (.X(net974),
    .A(net975));
 sg13g2_buf_16 fanout975 (.X(net975),
    .A(AD3));
 sg13g2_buf_8 fanout976 (.A(_1167_),
    .X(net976));
 sg13g2_buf_1 fanout977 (.A(_1167_),
    .X(net977));
 sg13g2_buf_8 fanout978 (.A(net979),
    .X(net978));
 sg13g2_buf_16 fanout979 (.X(net979),
    .A(AD1));
 sg13g2_buf_1 fanout980 (.A(AD1),
    .X(net980));
 sg13g2_dlygate4sd1_1 rebuffer7 (.A(net504),
    .X(net505));
 sg13g2_buf_16 fanout982 (.X(net982),
    .A(net983));
 sg13g2_buf_8 fanout983 (.A(_0142_),
    .X(net983));
 sg13g2_buf_1 fanout984 (.A(net985),
    .X(net984));
 sg13g2_buf_8 fanout985 (.A(BD2),
    .X(net985));
 sg13g2_buf_1 fanout986 (.A(net987),
    .X(net986));
 sg13g2_buf_1 fanout987 (.A(net989),
    .X(net987));
 sg13g2_buf_1 fanout988 (.A(net989),
    .X(net988));
 sg13g2_buf_1 fanout989 (.A(BD2),
    .X(net989));
 sg13g2_buf_16 fanout990 (.X(net990),
    .A(net992));
 sg13g2_buf_1 fanout991 (.A(net992),
    .X(net991));
 sg13g2_buf_8 fanout992 (.A(B_ADR0),
    .X(net992));
 sg13g2_buf_1 fanout993 (.A(net996),
    .X(net993));
 sg13g2_buf_1 fanout994 (.A(net996),
    .X(net994));
 sg13g2_buf_1 fanout995 (.A(net996),
    .X(net995));
 sg13g2_buf_1 fanout996 (.A(net997),
    .X(net996));
 sg13g2_buf_1 fanout997 (.A(net998),
    .X(net997));
 sg13g2_buf_1 fanout998 (.A(B_ADR0),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_1165_),
    .X(net999));
 sg13g2_buf_2 rebuffer20 (.A(_0458_),
    .X(net518));
 sg13g2_buf_1 fanout1001 (.A(net1002),
    .X(net1001));
 sg13g2_buf_1 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(BD3),
    .X(net1003));
 sg13g2_buf_1 fanout1004 (.A(net1006),
    .X(net1004));
 sg13g2_buf_16 fanout1005 (.X(net1005),
    .A(net1006));
 sg13g2_buf_16 fanout1006 (.X(net1006),
    .A(net1007));
 sg13g2_buf_8 fanout1007 (.A(_0409_),
    .X(net1007));
 sg13g2_buf_1 fanout1008 (.A(net1009),
    .X(net1008));
 sg13g2_buf_1 fanout1009 (.A(_0409_),
    .X(net1009));
 sg13g2_buf_16 fanout1010 (.X(net1010),
    .A(_1164_));
 sg13g2_buf_16 fanout1011 (.X(net1011),
    .A(_1164_));
 sg13g2_buf_16 fanout1012 (.X(net1012),
    .A(net1014));
 sg13g2_buf_16 fanout1013 (.X(net1013),
    .A(net1014));
 sg13g2_buf_16 fanout1014 (.X(net1014),
    .A(BD1));
 sg13g2_buf_16 fanout1015 (.X(net1015),
    .A(BD1));
 sg13g2_buf_1 fanout1016 (.A(_1166_),
    .X(net1016));
 sg13g2_buf_1 fanout1017 (.A(net1018),
    .X(net1017));
 sg13g2_buf_16 fanout1018 (.X(net1018),
    .A(AD0));
 sg13g2_buf_1 fanout1019 (.A(net1020),
    .X(net1019));
 sg13g2_buf_1 fanout1020 (.A(AD0),
    .X(net1020));
 sg13g2_buf_8 rebuffer6 (.A(net525),
    .X(net504));
 sg13g2_buf_1 fanout1022 (.A(net1025),
    .X(net1022));
 sg13g2_buf_1 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_1 fanout1024 (.A(net1025),
    .X(net1024));
 sg13g2_buf_1 fanout1025 (.A(_1210_),
    .X(net1025));
 sg13g2_buf_1 fanout1026 (.A(net1028),
    .X(net1026));
 sg13g2_buf_1 fanout1027 (.A(net1028),
    .X(net1027));
 sg13g2_buf_1 fanout1028 (.A(_1210_),
    .X(net1028));
 sg13g2_buf_1 fanout1029 (.A(net1030),
    .X(net1029));
 sg13g2_buf_1 fanout1030 (.A(BD0),
    .X(net1030));
 sg13g2_buf_1 fanout1031 (.A(BD0),
    .X(net1031));
 sg13g2_buf_8 fanout1032 (.A(BD0),
    .X(net1032));
 sg13g2_buf_1 fanout1033 (.A(net1034),
    .X(net1033));
 sg13g2_buf_1 fanout1034 (.A(BD0),
    .X(net1034));
 sg13g2_buf_2 rebuffer18 (.A(net537),
    .X(net516));
 sg13g2_buf_1 fanout1036 (.A(_0367_),
    .X(net1036));
 sg13g2_buf_1 fanout1037 (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .X(net1037));
 sg13g2_buf_1 fanout1038 (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .X(net1038));
 sg13g2_buf_1 fanout1039 (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .X(net1039));
 sg13g2_buf_1 fanout1040 (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .X(net1040));
 sg13g2_buf_1 fanout1041 (.A(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .X(net1041));
 sg13g2_buf_1 fanout1042 (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .X(net1042));
 sg13g2_buf_1 fanout1043 (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .X(net1043));
 sg13g2_buf_1 fanout1044 (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .X(net1044));
 sg13g2_buf_1 fanout1045 (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .X(net1045));
 sg13g2_buf_1 fanout1046 (.A(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .X(net1046));
 sg13g2_buf_1 fanout1047 (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .X(net1047));
 sg13g2_buf_1 fanout1048 (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .X(net1048));
 sg13g2_buf_1 fanout1049 (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .X(net1049));
 sg13g2_buf_1 fanout1050 (.A(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .X(net1050));
 sg13g2_buf_1 fanout1051 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .X(net1051));
 sg13g2_buf_1 fanout1052 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .X(net1052));
 sg13g2_buf_1 fanout1053 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .X(net1053));
 sg13g2_buf_1 fanout1054 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .X(net1054));
 sg13g2_buf_1 fanout1055 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .X(net1055));
 sg13g2_buf_1 fanout1056 (.A(net1057),
    .X(net1056));
 sg13g2_buf_1 fanout1057 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .X(net1057));
 sg13g2_buf_1 fanout1058 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .X(net1058));
 sg13g2_buf_1 fanout1059 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .X(net1059));
 sg13g2_buf_1 fanout1060 (.A(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .X(net1060));
 sg13g2_buf_1 fanout1061 (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(net1061));
 sg13g2_buf_1 fanout1062 (.A(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .X(net1062));
 sg13g2_buf_1 fanout1063 (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(net1063));
 sg13g2_buf_1 fanout1064 (.A(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .X(net1064));
 sg13g2_buf_1 fanout1065 (.A(net105),
    .X(net1065));
 sg13g2_buf_1 fanout1066 (.A(net1067),
    .X(net1066));
 sg13g2_buf_1 fanout1067 (.A(W6END[0]),
    .X(net1067));
 sg13g2_buf_1 fanout1068 (.A(net1069),
    .X(net1068));
 sg13g2_buf_1 fanout1069 (.A(W1END[3]),
    .X(net1069));
 sg13g2_buf_1 fanout1070 (.A(net88),
    .X(net1070));
 sg13g2_buf_8 fanout1071 (.A(net87),
    .X(net1071));
 sg13g2_buf_1 fanout1072 (.A(net86),
    .X(net1072));
 sg13g2_buf_1 fanout1073 (.A(net33),
    .X(net1073));
 sg13g2_buf_1 fanout1074 (.A(net32),
    .X(net1074));
 sg13g2_buf_16 fanout1075 (.X(net1075),
    .A(net31));
 sg13g2_buf_1 fanout1076 (.A(net30),
    .X(net1076));
 sg13g2_buf_1 fanout1077 (.A(net1081),
    .X(net1077));
 sg13g2_buf_1 fanout1078 (.A(net1080),
    .X(net1078));
 sg13g2_buf_1 fanout1079 (.A(net1080),
    .X(net1079));
 sg13g2_buf_1 fanout1080 (.A(net1081),
    .X(net1080));
 sg13g2_buf_1 fanout1081 (.A(net29),
    .X(net1081));
 sg13g2_buf_1 fanout1082 (.A(net29),
    .X(net1082));
 sg13g2_buf_1 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_1 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_1 fanout1085 (.A(FrameStrobe[8]),
    .X(net1085));
 sg13g2_buf_1 fanout1086 (.A(FrameStrobe[8]),
    .X(net1086));
 sg13g2_buf_1 fanout1087 (.A(FrameStrobe[8]),
    .X(net1087));
 sg13g2_buf_1 fanout1088 (.A(net1092),
    .X(net1088));
 sg13g2_buf_1 fanout1089 (.A(net1092),
    .X(net1089));
 sg13g2_buf_1 fanout1090 (.A(net1092),
    .X(net1090));
 sg13g2_buf_1 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_1 fanout1092 (.A(FrameStrobe[7]),
    .X(net1092));
 sg13g2_buf_1 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_1 fanout1094 (.A(net1097),
    .X(net1094));
 sg13g2_buf_1 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_buf_1 fanout1096 (.A(net1097),
    .X(net1096));
 sg13g2_buf_1 fanout1097 (.A(FrameStrobe[6]),
    .X(net1097));
 sg13g2_buf_1 fanout1098 (.A(net1102),
    .X(net1098));
 sg13g2_buf_1 fanout1099 (.A(net1102),
    .X(net1099));
 sg13g2_buf_1 fanout1100 (.A(net1101),
    .X(net1100));
 sg13g2_buf_1 fanout1101 (.A(net1102),
    .X(net1101));
 sg13g2_buf_1 fanout1102 (.A(net28),
    .X(net1102));
 sg13g2_buf_1 fanout1103 (.A(net1108),
    .X(net1103));
 sg13g2_buf_1 fanout1104 (.A(net1108),
    .X(net1104));
 sg13g2_buf_1 fanout1105 (.A(net1107),
    .X(net1105));
 sg13g2_buf_1 fanout1106 (.A(net1107),
    .X(net1106));
 sg13g2_buf_1 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_1 fanout1108 (.A(FrameStrobe[4]),
    .X(net1108));
 sg13g2_buf_1 fanout1109 (.A(net1114),
    .X(net1109));
 sg13g2_buf_1 fanout1110 (.A(net1114),
    .X(net1110));
 sg13g2_buf_1 fanout1111 (.A(net1113),
    .X(net1111));
 sg13g2_buf_1 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_buf_1 fanout1113 (.A(net1114),
    .X(net1113));
 sg13g2_buf_1 fanout1114 (.A(FrameStrobe[3]),
    .X(net1114));
 sg13g2_buf_1 fanout1115 (.A(net1120),
    .X(net1115));
 sg13g2_buf_1 fanout1116 (.A(net1120),
    .X(net1116));
 sg13g2_buf_1 fanout1117 (.A(net1119),
    .X(net1117));
 sg13g2_buf_1 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_buf_1 fanout1119 (.A(net1120),
    .X(net1119));
 sg13g2_buf_1 fanout1120 (.A(FrameStrobe[2]),
    .X(net1120));
 sg13g2_buf_1 fanout1121 (.A(net1125),
    .X(net1121));
 sg13g2_buf_1 fanout1122 (.A(net1125),
    .X(net1122));
 sg13g2_buf_1 fanout1123 (.A(net1124),
    .X(net1123));
 sg13g2_buf_1 fanout1124 (.A(net1125),
    .X(net1124));
 sg13g2_buf_1 fanout1125 (.A(net1126),
    .X(net1125));
 sg13g2_buf_1 fanout1126 (.A(FrameStrobe[1]),
    .X(net1126));
 sg13g2_buf_1 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_buf_1 fanout1128 (.A(net1130),
    .X(net1128));
 sg13g2_buf_1 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_buf_1 fanout1130 (.A(net27),
    .X(net1130));
 sg13g2_buf_1 fanout1131 (.A(net1136),
    .X(net1131));
 sg13g2_buf_1 fanout1132 (.A(net1135),
    .X(net1132));
 sg13g2_buf_1 fanout1133 (.A(net1135),
    .X(net1133));
 sg13g2_buf_1 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_1 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_buf_1 fanout1136 (.A(FrameStrobe[11]),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(net1141),
    .X(net1137));
 sg13g2_buf_1 fanout1138 (.A(net1141),
    .X(net1138));
 sg13g2_buf_1 fanout1139 (.A(net1140),
    .X(net1139));
 sg13g2_buf_1 fanout1140 (.A(net1141),
    .X(net1140));
 sg13g2_buf_1 fanout1141 (.A(FrameStrobe[10]),
    .X(net1141));
 sg13g2_buf_1 fanout1142 (.A(net1143),
    .X(net1142));
 sg13g2_buf_1 fanout1143 (.A(net1147),
    .X(net1143));
 sg13g2_buf_1 fanout1144 (.A(net1146),
    .X(net1144));
 sg13g2_buf_1 fanout1145 (.A(net1146),
    .X(net1145));
 sg13g2_buf_1 fanout1146 (.A(net1147),
    .X(net1146));
 sg13g2_buf_1 fanout1147 (.A(FrameStrobe[0]),
    .X(net1147));
 sg13g2_buf_1 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_1 fanout1149 (.A(FrameData[9]),
    .X(net1149));
 sg13g2_buf_1 fanout1150 (.A(net1151),
    .X(net1150));
 sg13g2_buf_1 fanout1151 (.A(FrameData[8]),
    .X(net1151));
 sg13g2_buf_1 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_1 fanout1153 (.A(net26),
    .X(net1153));
 sg13g2_buf_1 fanout1154 (.A(net1155),
    .X(net1154));
 sg13g2_buf_1 fanout1155 (.A(net25),
    .X(net1155));
 sg13g2_buf_1 fanout1156 (.A(net1157),
    .X(net1156));
 sg13g2_buf_1 fanout1157 (.A(FrameData[5]),
    .X(net1157));
 sg13g2_buf_1 fanout1158 (.A(net1159),
    .X(net1158));
 sg13g2_buf_1 fanout1159 (.A(FrameData[4]),
    .X(net1159));
 sg13g2_buf_1 fanout1160 (.A(FrameData[3]),
    .X(net1160));
 sg13g2_buf_1 fanout1161 (.A(FrameData[3]),
    .X(net1161));
 sg13g2_buf_1 fanout1162 (.A(FrameData[31]),
    .X(net1162));
 sg13g2_buf_1 fanout1163 (.A(FrameData[31]),
    .X(net1163));
 sg13g2_buf_1 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_buf_1 fanout1165 (.A(FrameData[30]),
    .X(net1165));
 sg13g2_buf_1 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_buf_1 fanout1167 (.A(FrameData[2]),
    .X(net1167));
 sg13g2_buf_1 fanout1168 (.A(FrameData[29]),
    .X(net1168));
 sg13g2_buf_1 fanout1169 (.A(FrameData[29]),
    .X(net1169));
 sg13g2_buf_1 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_buf_1 fanout1171 (.A(FrameData[28]),
    .X(net1171));
 sg13g2_buf_1 fanout1172 (.A(FrameData[27]),
    .X(net1172));
 sg13g2_buf_1 fanout1173 (.A(FrameData[27]),
    .X(net1173));
 sg13g2_buf_1 fanout1174 (.A(net1175),
    .X(net1174));
 sg13g2_buf_1 fanout1175 (.A(FrameData[26]),
    .X(net1175));
 sg13g2_buf_1 fanout1176 (.A(FrameData[25]),
    .X(net1176));
 sg13g2_buf_1 fanout1177 (.A(FrameData[25]),
    .X(net1177));
 sg13g2_buf_1 fanout1178 (.A(FrameData[24]),
    .X(net1178));
 sg13g2_buf_1 fanout1179 (.A(FrameData[24]),
    .X(net1179));
 sg13g2_buf_1 fanout1180 (.A(net1181),
    .X(net1180));
 sg13g2_buf_1 fanout1181 (.A(FrameData[23]),
    .X(net1181));
 sg13g2_buf_1 fanout1182 (.A(FrameData[22]),
    .X(net1182));
 sg13g2_buf_1 fanout1183 (.A(FrameData[22]),
    .X(net1183));
 sg13g2_buf_1 fanout1184 (.A(FrameData[21]),
    .X(net1184));
 sg13g2_buf_1 fanout1185 (.A(FrameData[21]),
    .X(net1185));
 sg13g2_buf_1 fanout1186 (.A(FrameData[20]),
    .X(net1186));
 sg13g2_buf_1 fanout1187 (.A(FrameData[20]),
    .X(net1187));
 sg13g2_buf_1 fanout1188 (.A(FrameData[1]),
    .X(net1188));
 sg13g2_buf_1 fanout1189 (.A(FrameData[1]),
    .X(net1189));
 sg13g2_buf_1 fanout1190 (.A(net1191),
    .X(net1190));
 sg13g2_buf_1 fanout1191 (.A(FrameData[19]),
    .X(net1191));
 sg13g2_buf_1 fanout1192 (.A(net1193),
    .X(net1192));
 sg13g2_buf_1 fanout1193 (.A(FrameData[18]),
    .X(net1193));
 sg13g2_buf_1 fanout1194 (.A(net1195),
    .X(net1194));
 sg13g2_buf_1 fanout1195 (.A(FrameData[17]),
    .X(net1195));
 sg13g2_buf_1 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_1 fanout1197 (.A(FrameData[16]),
    .X(net1197));
 sg13g2_buf_1 fanout1198 (.A(net1200),
    .X(net1198));
 sg13g2_buf_1 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_1 fanout1200 (.A(FrameData[15]),
    .X(net1200));
 sg13g2_buf_1 fanout1201 (.A(net1202),
    .X(net1201));
 sg13g2_buf_1 fanout1202 (.A(FrameData[14]),
    .X(net1202));
 sg13g2_buf_1 fanout1203 (.A(net1205),
    .X(net1203));
 sg13g2_buf_1 fanout1204 (.A(net1205),
    .X(net1204));
 sg13g2_buf_1 fanout1205 (.A(FrameData[13]),
    .X(net1205));
 sg13g2_buf_1 fanout1206 (.A(FrameData[12]),
    .X(net1206));
 sg13g2_buf_1 fanout1207 (.A(FrameData[12]),
    .X(net1207));
 sg13g2_buf_1 fanout1208 (.A(net1209),
    .X(net1208));
 sg13g2_buf_1 fanout1209 (.A(FrameData[11]),
    .X(net1209));
 sg13g2_buf_1 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_1 fanout1211 (.A(FrameData[10]),
    .X(net1211));
 sg13g2_buf_1 fanout1212 (.A(FrameData[0]),
    .X(net1212));
 sg13g2_buf_1 fanout1213 (.A(FrameData[0]),
    .X(net1213));
 sg13g2_buf_1 fanout1214 (.A(E6END[1]),
    .X(net1214));
 sg13g2_buf_1 fanout1215 (.A(E6END[1]),
    .X(net1215));
 sg13g2_buf_1 fanout1216 (.A(E6END[0]),
    .X(net1216));
 sg13g2_buf_1 fanout1217 (.A(E6END[0]),
    .X(net1217));
 sg13g2_buf_1 fanout1218 (.A(net4),
    .X(net1218));
 sg13g2_buf_1 fanout1219 (.A(net3),
    .X(net1219));
 sg13g2_buf_16 fanout1220 (.X(net1220),
    .A(net2));
 sg13g2_buf_1 fanout1221 (.A(net1),
    .X(net1221));
 sg13g2_buf_1 input1 (.A(E1END[0]),
    .X(net1));
 sg13g2_buf_16 input2 (.X(net2),
    .A(E1END[1]));
 sg13g2_buf_1 input3 (.A(E1END[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(E1END[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(E2END[0]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(E2END[1]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(E2END[2]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(E2END[3]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(E2END[4]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(E2END[5]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(E2END[6]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(E2END[7]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(E2MID[0]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(E2MID[1]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(E2MID[2]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(E2MID[3]),
    .X(net16));
 sg13g2_buf_1 input17 (.A(E2MID[4]),
    .X(net17));
 sg13g2_buf_1 input18 (.A(E2MID[5]),
    .X(net18));
 sg13g2_buf_1 input19 (.A(E2MID[6]),
    .X(net19));
 sg13g2_buf_1 input20 (.A(E2MID[7]),
    .X(net20));
 sg13g2_buf_1 input21 (.A(EE4END[0]),
    .X(net21));
 sg13g2_buf_1 input22 (.A(EE4END[1]),
    .X(net22));
 sg13g2_buf_1 input23 (.A(EE4END[2]),
    .X(net23));
 sg13g2_buf_1 input24 (.A(EE4END[3]),
    .X(net24));
 sg13g2_buf_1 input25 (.A(FrameData[6]),
    .X(net25));
 sg13g2_buf_1 input26 (.A(FrameData[7]),
    .X(net26));
 sg13g2_buf_1 input27 (.A(FrameStrobe[12]),
    .X(net27));
 sg13g2_buf_1 input28 (.A(FrameStrobe[5]),
    .X(net28));
 sg13g2_buf_1 input29 (.A(FrameStrobe[9]),
    .X(net29));
 sg13g2_buf_1 input30 (.A(N1END[0]),
    .X(net30));
 sg13g2_buf_16 input31 (.X(net31),
    .A(N1END[1]));
 sg13g2_buf_1 input32 (.A(N1END[2]),
    .X(net32));
 sg13g2_buf_1 input33 (.A(N1END[3]),
    .X(net33));
 sg13g2_buf_1 input34 (.A(N2END[0]),
    .X(net34));
 sg13g2_buf_1 input35 (.A(N2END[1]),
    .X(net35));
 sg13g2_buf_1 input36 (.A(N2END[2]),
    .X(net36));
 sg13g2_buf_1 input37 (.A(N2END[3]),
    .X(net37));
 sg13g2_buf_1 input38 (.A(N2END[4]),
    .X(net38));
 sg13g2_buf_2 input39 (.A(N2END[5]),
    .X(net39));
 sg13g2_buf_1 input40 (.A(N2END[6]),
    .X(net40));
 sg13g2_buf_1 input41 (.A(N2END[7]),
    .X(net41));
 sg13g2_buf_1 input42 (.A(N2MID[0]),
    .X(net42));
 sg13g2_buf_1 input43 (.A(N2MID[1]),
    .X(net43));
 sg13g2_buf_1 input44 (.A(N2MID[2]),
    .X(net44));
 sg13g2_buf_1 input45 (.A(N2MID[3]),
    .X(net45));
 sg13g2_buf_1 input46 (.A(N2MID[4]),
    .X(net46));
 sg13g2_buf_1 input47 (.A(N2MID[5]),
    .X(net47));
 sg13g2_buf_1 input48 (.A(N2MID[6]),
    .X(net48));
 sg13g2_buf_1 input49 (.A(N2MID[7]),
    .X(net49));
 sg13g2_buf_1 input50 (.A(N4END[0]),
    .X(net50));
 sg13g2_buf_1 input51 (.A(N4END[1]),
    .X(net51));
 sg13g2_buf_1 input52 (.A(N4END[2]),
    .X(net52));
 sg13g2_buf_1 input53 (.A(N4END[3]),
    .X(net53));
 sg13g2_buf_1 input54 (.A(NN4END[0]),
    .X(net54));
 sg13g2_buf_1 input55 (.A(NN4END[1]),
    .X(net55));
 sg13g2_buf_1 input56 (.A(NN4END[2]),
    .X(net56));
 sg13g2_buf_8 input57 (.A(NN4END[3]),
    .X(net57));
 sg13g2_buf_1 input58 (.A(S1END[0]),
    .X(net58));
 sg13g2_buf_2 input59 (.A(S1END[1]),
    .X(net59));
 sg13g2_buf_1 input60 (.A(S1END[2]),
    .X(net60));
 sg13g2_buf_1 input61 (.A(S1END[3]),
    .X(net61));
 sg13g2_buf_1 input62 (.A(S2END[0]),
    .X(net62));
 sg13g2_buf_1 input63 (.A(S2END[1]),
    .X(net63));
 sg13g2_buf_1 input64 (.A(S2END[2]),
    .X(net64));
 sg13g2_buf_1 input65 (.A(S2END[3]),
    .X(net65));
 sg13g2_buf_1 input66 (.A(S2END[4]),
    .X(net66));
 sg13g2_buf_1 input67 (.A(S2END[5]),
    .X(net67));
 sg13g2_buf_1 input68 (.A(S2END[6]),
    .X(net68));
 sg13g2_buf_1 input69 (.A(S2END[7]),
    .X(net69));
 sg13g2_buf_1 input70 (.A(S2MID[0]),
    .X(net70));
 sg13g2_buf_1 input71 (.A(S2MID[1]),
    .X(net71));
 sg13g2_buf_1 input72 (.A(S2MID[2]),
    .X(net72));
 sg13g2_buf_1 input73 (.A(S2MID[3]),
    .X(net73));
 sg13g2_buf_1 input74 (.A(S2MID[4]),
    .X(net74));
 sg13g2_buf_1 input75 (.A(S2MID[5]),
    .X(net75));
 sg13g2_buf_1 input76 (.A(S2MID[6]),
    .X(net76));
 sg13g2_buf_1 input77 (.A(S2MID[7]),
    .X(net77));
 sg13g2_buf_1 input78 (.A(S4END[0]),
    .X(net78));
 sg13g2_buf_1 input79 (.A(S4END[1]),
    .X(net79));
 sg13g2_buf_1 input80 (.A(S4END[2]),
    .X(net80));
 sg13g2_buf_1 input81 (.A(S4END[3]),
    .X(net81));
 sg13g2_buf_1 input82 (.A(SS4END[0]),
    .X(net82));
 sg13g2_buf_1 input83 (.A(SS4END[1]),
    .X(net83));
 sg13g2_buf_1 input84 (.A(SS4END[2]),
    .X(net84));
 sg13g2_buf_1 input85 (.A(SS4END[3]),
    .X(net85));
 sg13g2_buf_1 input86 (.A(W1END[0]),
    .X(net86));
 sg13g2_buf_8 input87 (.A(W1END[1]),
    .X(net87));
 sg13g2_buf_1 input88 (.A(W1END[2]),
    .X(net88));
 sg13g2_buf_1 input89 (.A(W2END[0]),
    .X(net89));
 sg13g2_buf_1 input90 (.A(W2END[1]),
    .X(net90));
 sg13g2_buf_1 input91 (.A(W2END[2]),
    .X(net91));
 sg13g2_buf_1 input92 (.A(W2END[3]),
    .X(net92));
 sg13g2_buf_1 input93 (.A(W2END[4]),
    .X(net93));
 sg13g2_buf_1 input94 (.A(W2END[5]),
    .X(net94));
 sg13g2_buf_1 input95 (.A(W2END[6]),
    .X(net95));
 sg13g2_buf_1 input96 (.A(W2END[7]),
    .X(net96));
 sg13g2_buf_1 input97 (.A(W2MID[0]),
    .X(net97));
 sg13g2_buf_1 input98 (.A(W2MID[1]),
    .X(net98));
 sg13g2_buf_1 input99 (.A(W2MID[2]),
    .X(net99));
 sg13g2_buf_1 input100 (.A(W2MID[3]),
    .X(net100));
 sg13g2_buf_1 input101 (.A(W2MID[4]),
    .X(net101));
 sg13g2_buf_1 input102 (.A(W2MID[5]),
    .X(net102));
 sg13g2_buf_1 input103 (.A(W2MID[6]),
    .X(net103));
 sg13g2_buf_1 input104 (.A(W2MID[7]),
    .X(net104));
 sg13g2_buf_1 input105 (.A(W6END[1]),
    .X(net105));
 sg13g2_buf_1 input106 (.A(WW4END[0]),
    .X(net106));
 sg13g2_buf_1 input107 (.A(WW4END[1]),
    .X(net107));
 sg13g2_buf_1 input108 (.A(WW4END[2]),
    .X(net108));
 sg13g2_buf_1 input109 (.A(WW4END[3]),
    .X(net109));
 sg13g2_buf_1 output110 (.A(\Inst_RegFile_switch_matrix.E1BEG0 ),
    .X(E1BEG[0]));
 sg13g2_buf_1 output111 (.A(\Inst_RegFile_switch_matrix.E1BEG1 ),
    .X(E1BEG[1]));
 sg13g2_buf_1 output112 (.A(\Inst_RegFile_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sg13g2_buf_1 output113 (.A(\Inst_RegFile_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sg13g2_buf_1 output114 (.A(net114),
    .X(E2BEG[0]));
 sg13g2_buf_1 output115 (.A(net115),
    .X(E2BEG[1]));
 sg13g2_buf_1 output116 (.A(net116),
    .X(E2BEG[2]));
 sg13g2_buf_1 output117 (.A(net117),
    .X(E2BEG[3]));
 sg13g2_buf_1 output118 (.A(net118),
    .X(E2BEG[4]));
 sg13g2_buf_8 output119 (.A(net119),
    .X(E2BEG[5]));
 sg13g2_buf_1 output120 (.A(net120),
    .X(E2BEG[6]));
 sg13g2_buf_1 output121 (.A(net121),
    .X(E2BEG[7]));
 sg13g2_buf_1 output122 (.A(net122),
    .X(E2BEGb[0]));
 sg13g2_buf_1 output123 (.A(net123),
    .X(E2BEGb[1]));
 sg13g2_buf_1 output124 (.A(net124),
    .X(E2BEGb[2]));
 sg13g2_buf_1 output125 (.A(net125),
    .X(E2BEGb[3]));
 sg13g2_buf_1 output126 (.A(net126),
    .X(E2BEGb[4]));
 sg13g2_buf_1 output127 (.A(net127),
    .X(E2BEGb[5]));
 sg13g2_buf_1 output128 (.A(net128),
    .X(E2BEGb[6]));
 sg13g2_buf_1 output129 (.A(net129),
    .X(E2BEGb[7]));
 sg13g2_buf_1 output130 (.A(net130),
    .X(E6BEG[0]));
 sg13g2_buf_1 output131 (.A(\Inst_RegFile_switch_matrix.E6BEG0 ),
    .X(E6BEG[10]));
 sg13g2_buf_1 output132 (.A(\Inst_RegFile_switch_matrix.E6BEG1 ),
    .X(E6BEG[11]));
 sg13g2_buf_1 output133 (.A(net133),
    .X(E6BEG[1]));
 sg13g2_buf_1 output134 (.A(net134),
    .X(E6BEG[2]));
 sg13g2_buf_1 output135 (.A(net135),
    .X(E6BEG[3]));
 sg13g2_buf_1 output136 (.A(net136),
    .X(E6BEG[4]));
 sg13g2_buf_1 output137 (.A(net137),
    .X(E6BEG[5]));
 sg13g2_buf_1 output138 (.A(net138),
    .X(E6BEG[6]));
 sg13g2_buf_1 output139 (.A(net139),
    .X(E6BEG[7]));
 sg13g2_buf_1 output140 (.A(net140),
    .X(E6BEG[8]));
 sg13g2_buf_1 output141 (.A(net141),
    .X(E6BEG[9]));
 sg13g2_buf_1 output142 (.A(net142),
    .X(EE4BEG[0]));
 sg13g2_buf_1 output143 (.A(net143),
    .X(EE4BEG[10]));
 sg13g2_buf_1 output144 (.A(net144),
    .X(EE4BEG[11]));
 sg13g2_buf_1 output145 (.A(\Inst_RegFile_switch_matrix.EE4BEG0 ),
    .X(EE4BEG[12]));
 sg13g2_buf_1 output146 (.A(\Inst_RegFile_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[13]));
 sg13g2_buf_1 output147 (.A(net147),
    .X(EE4BEG[14]));
 sg13g2_buf_1 output148 (.A(net148),
    .X(EE4BEG[15]));
 sg13g2_buf_1 output149 (.A(net149),
    .X(EE4BEG[1]));
 sg13g2_buf_1 output150 (.A(net150),
    .X(EE4BEG[2]));
 sg13g2_buf_1 output151 (.A(net151),
    .X(EE4BEG[3]));
 sg13g2_buf_1 output152 (.A(net152),
    .X(EE4BEG[4]));
 sg13g2_buf_1 output153 (.A(net153),
    .X(EE4BEG[5]));
 sg13g2_buf_1 output154 (.A(net154),
    .X(EE4BEG[6]));
 sg13g2_buf_1 output155 (.A(net155),
    .X(EE4BEG[7]));
 sg13g2_buf_1 output156 (.A(net156),
    .X(EE4BEG[8]));
 sg13g2_buf_1 output157 (.A(net157),
    .X(EE4BEG[9]));
 sg13g2_buf_1 output158 (.A(net158),
    .X(FrameData_O[0]));
 sg13g2_buf_1 output159 (.A(net159),
    .X(FrameData_O[10]));
 sg13g2_buf_1 output160 (.A(net160),
    .X(FrameData_O[11]));
 sg13g2_buf_1 output161 (.A(net161),
    .X(FrameData_O[12]));
 sg13g2_buf_1 output162 (.A(net162),
    .X(FrameData_O[13]));
 sg13g2_buf_1 output163 (.A(net163),
    .X(FrameData_O[14]));
 sg13g2_buf_1 output164 (.A(net164),
    .X(FrameData_O[15]));
 sg13g2_buf_1 output165 (.A(net165),
    .X(FrameData_O[16]));
 sg13g2_buf_1 output166 (.A(net166),
    .X(FrameData_O[17]));
 sg13g2_buf_1 output167 (.A(net167),
    .X(FrameData_O[18]));
 sg13g2_buf_1 output168 (.A(net168),
    .X(FrameData_O[19]));
 sg13g2_buf_1 output169 (.A(net169),
    .X(FrameData_O[1]));
 sg13g2_buf_1 output170 (.A(net170),
    .X(FrameData_O[20]));
 sg13g2_buf_1 output171 (.A(net171),
    .X(FrameData_O[21]));
 sg13g2_buf_1 output172 (.A(net172),
    .X(FrameData_O[22]));
 sg13g2_buf_1 output173 (.A(net173),
    .X(FrameData_O[23]));
 sg13g2_buf_1 output174 (.A(net174),
    .X(FrameData_O[24]));
 sg13g2_buf_1 output175 (.A(net175),
    .X(FrameData_O[25]));
 sg13g2_buf_1 output176 (.A(net176),
    .X(FrameData_O[26]));
 sg13g2_buf_1 output177 (.A(net177),
    .X(FrameData_O[27]));
 sg13g2_buf_1 output178 (.A(net178),
    .X(FrameData_O[28]));
 sg13g2_buf_1 output179 (.A(net179),
    .X(FrameData_O[29]));
 sg13g2_buf_1 output180 (.A(net180),
    .X(FrameData_O[2]));
 sg13g2_buf_1 output181 (.A(net181),
    .X(FrameData_O[30]));
 sg13g2_buf_1 output182 (.A(net182),
    .X(FrameData_O[31]));
 sg13g2_buf_1 output183 (.A(net183),
    .X(FrameData_O[3]));
 sg13g2_buf_1 output184 (.A(net184),
    .X(FrameData_O[4]));
 sg13g2_buf_1 output185 (.A(net185),
    .X(FrameData_O[5]));
 sg13g2_buf_1 output186 (.A(net186),
    .X(FrameData_O[6]));
 sg13g2_buf_1 output187 (.A(net187),
    .X(FrameData_O[7]));
 sg13g2_buf_1 output188 (.A(net188),
    .X(FrameData_O[8]));
 sg13g2_buf_1 output189 (.A(net189),
    .X(FrameData_O[9]));
 sg13g2_buf_1 output190 (.A(net190),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 output191 (.A(net191),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 output192 (.A(net192),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 output193 (.A(net193),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 output194 (.A(net194),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 output195 (.A(net195),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 output196 (.A(net196),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 output197 (.A(net197),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 output198 (.A(net198),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 output199 (.A(net199),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 output200 (.A(net200),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 output201 (.A(net201),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 output202 (.A(net202),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 output203 (.A(net203),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 output204 (.A(net204),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 output205 (.A(net205),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 output206 (.A(net206),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 output207 (.A(net207),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 output208 (.A(net208),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 output209 (.A(net209),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 output210 (.A(net210),
    .X(N1BEG[0]));
 sg13g2_buf_1 output211 (.A(\Inst_RegFile_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]));
 sg13g2_buf_1 output212 (.A(\Inst_RegFile_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]));
 sg13g2_buf_1 output213 (.A(\Inst_RegFile_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]));
 sg13g2_buf_1 output214 (.A(net214),
    .X(N2BEG[0]));
 sg13g2_buf_1 output215 (.A(net215),
    .X(N2BEG[1]));
 sg13g2_buf_1 output216 (.A(net216),
    .X(N2BEG[2]));
 sg13g2_buf_1 output217 (.A(net217),
    .X(N2BEG[3]));
 sg13g2_buf_1 output218 (.A(net218),
    .X(N2BEG[4]));
 sg13g2_buf_1 output219 (.A(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .X(N2BEG[5]));
 sg13g2_buf_1 output220 (.A(net510),
    .X(N2BEG[6]));
 sg13g2_buf_1 output221 (.A(net221),
    .X(N2BEG[7]));
 sg13g2_buf_1 output222 (.A(net222),
    .X(N2BEGb[0]));
 sg13g2_buf_1 output223 (.A(net223),
    .X(N2BEGb[1]));
 sg13g2_buf_1 output224 (.A(net224),
    .X(N2BEGb[2]));
 sg13g2_buf_1 output225 (.A(net225),
    .X(N2BEGb[3]));
 sg13g2_buf_1 output226 (.A(net226),
    .X(N2BEGb[4]));
 sg13g2_buf_1 output227 (.A(net227),
    .X(N2BEGb[5]));
 sg13g2_buf_1 output228 (.A(net228),
    .X(N2BEGb[6]));
 sg13g2_buf_1 output229 (.A(net229),
    .X(N2BEGb[7]));
 sg13g2_buf_1 output230 (.A(net230),
    .X(N4BEG[0]));
 sg13g2_buf_1 output231 (.A(net231),
    .X(N4BEG[10]));
 sg13g2_buf_1 output232 (.A(net232),
    .X(N4BEG[11]));
 sg13g2_buf_1 output233 (.A(net233),
    .X(N4BEG[12]));
 sg13g2_buf_1 output234 (.A(net234),
    .X(N4BEG[13]));
 sg13g2_buf_1 output235 (.A(net235),
    .X(N4BEG[14]));
 sg13g2_buf_1 output236 (.A(net236),
    .X(N4BEG[15]));
 sg13g2_buf_1 output237 (.A(net237),
    .X(N4BEG[1]));
 sg13g2_buf_1 output238 (.A(net238),
    .X(N4BEG[2]));
 sg13g2_buf_1 output239 (.A(net239),
    .X(N4BEG[3]));
 sg13g2_buf_1 output240 (.A(net240),
    .X(N4BEG[4]));
 sg13g2_buf_1 output241 (.A(net241),
    .X(N4BEG[5]));
 sg13g2_buf_1 output242 (.A(net242),
    .X(N4BEG[6]));
 sg13g2_buf_1 output243 (.A(net243),
    .X(N4BEG[7]));
 sg13g2_buf_1 output244 (.A(net244),
    .X(N4BEG[8]));
 sg13g2_buf_1 output245 (.A(net245),
    .X(N4BEG[9]));
 sg13g2_buf_1 output246 (.A(net246),
    .X(NN4BEG[0]));
 sg13g2_buf_1 output247 (.A(net247),
    .X(NN4BEG[10]));
 sg13g2_buf_1 output248 (.A(net248),
    .X(NN4BEG[11]));
 sg13g2_buf_1 output249 (.A(\Inst_RegFile_switch_matrix.NN4BEG0 ),
    .X(NN4BEG[12]));
 sg13g2_buf_1 output250 (.A(\Inst_RegFile_switch_matrix.NN4BEG1 ),
    .X(NN4BEG[13]));
 sg13g2_buf_1 output251 (.A(net251),
    .X(NN4BEG[14]));
 sg13g2_buf_1 output252 (.A(net252),
    .X(NN4BEG[15]));
 sg13g2_buf_1 output253 (.A(net253),
    .X(NN4BEG[1]));
 sg13g2_buf_1 output254 (.A(net254),
    .X(NN4BEG[2]));
 sg13g2_buf_1 output255 (.A(net255),
    .X(NN4BEG[3]));
 sg13g2_buf_1 output256 (.A(net256),
    .X(NN4BEG[4]));
 sg13g2_buf_1 output257 (.A(net257),
    .X(NN4BEG[5]));
 sg13g2_buf_1 output258 (.A(net258),
    .X(NN4BEG[6]));
 sg13g2_buf_1 output259 (.A(net259),
    .X(NN4BEG[7]));
 sg13g2_buf_1 output260 (.A(net260),
    .X(NN4BEG[8]));
 sg13g2_buf_1 output261 (.A(net261),
    .X(NN4BEG[9]));
 sg13g2_buf_1 output262 (.A(\Inst_RegFile_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]));
 sg13g2_buf_1 output263 (.A(\Inst_RegFile_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sg13g2_buf_1 output264 (.A(\Inst_RegFile_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sg13g2_buf_1 output265 (.A(\Inst_RegFile_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sg13g2_buf_1 output266 (.A(net266),
    .X(S2BEG[0]));
 sg13g2_buf_1 output267 (.A(net267),
    .X(S2BEG[1]));
 sg13g2_buf_1 output268 (.A(net268),
    .X(S2BEG[2]));
 sg13g2_buf_1 output269 (.A(net269),
    .X(S2BEG[3]));
 sg13g2_buf_1 output270 (.A(net270),
    .X(S2BEG[4]));
 sg13g2_buf_1 output271 (.A(net271),
    .X(S2BEG[5]));
 sg13g2_buf_1 output272 (.A(net272),
    .X(S2BEG[6]));
 sg13g2_buf_1 output273 (.A(net273),
    .X(S2BEG[7]));
 sg13g2_buf_1 output274 (.A(net274),
    .X(S2BEGb[0]));
 sg13g2_buf_1 output275 (.A(net275),
    .X(S2BEGb[1]));
 sg13g2_buf_1 output276 (.A(net276),
    .X(S2BEGb[2]));
 sg13g2_buf_1 output277 (.A(net277),
    .X(S2BEGb[3]));
 sg13g2_buf_1 output278 (.A(net278),
    .X(S2BEGb[4]));
 sg13g2_buf_1 output279 (.A(net279),
    .X(S2BEGb[5]));
 sg13g2_buf_1 output280 (.A(net280),
    .X(S2BEGb[6]));
 sg13g2_buf_1 output281 (.A(net281),
    .X(S2BEGb[7]));
 sg13g2_buf_1 output282 (.A(net282),
    .X(S4BEG[0]));
 sg13g2_buf_1 output283 (.A(net283),
    .X(S4BEG[10]));
 sg13g2_buf_1 output284 (.A(net284),
    .X(S4BEG[11]));
 sg13g2_buf_1 output285 (.A(net285),
    .X(S4BEG[12]));
 sg13g2_buf_1 output286 (.A(net286),
    .X(S4BEG[13]));
 sg13g2_buf_1 output287 (.A(net287),
    .X(S4BEG[14]));
 sg13g2_buf_1 output288 (.A(net288),
    .X(S4BEG[15]));
 sg13g2_buf_1 output289 (.A(net289),
    .X(S4BEG[1]));
 sg13g2_buf_1 output290 (.A(net290),
    .X(S4BEG[2]));
 sg13g2_buf_1 output291 (.A(net291),
    .X(S4BEG[3]));
 sg13g2_buf_1 output292 (.A(net292),
    .X(S4BEG[4]));
 sg13g2_buf_1 output293 (.A(net293),
    .X(S4BEG[5]));
 sg13g2_buf_1 output294 (.A(net294),
    .X(S4BEG[6]));
 sg13g2_buf_1 output295 (.A(net295),
    .X(S4BEG[7]));
 sg13g2_buf_1 output296 (.A(net296),
    .X(S4BEG[8]));
 sg13g2_buf_1 output297 (.A(net297),
    .X(S4BEG[9]));
 sg13g2_buf_1 output298 (.A(net298),
    .X(SS4BEG[0]));
 sg13g2_buf_1 output299 (.A(net299),
    .X(SS4BEG[10]));
 sg13g2_buf_1 output300 (.A(net300),
    .X(SS4BEG[11]));
 sg13g2_buf_1 output301 (.A(\Inst_RegFile_switch_matrix.SS4BEG0 ),
    .X(SS4BEG[12]));
 sg13g2_buf_1 output302 (.A(\Inst_RegFile_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[13]));
 sg13g2_buf_1 output303 (.A(net303),
    .X(SS4BEG[14]));
 sg13g2_buf_1 output304 (.A(net304),
    .X(SS4BEG[15]));
 sg13g2_buf_1 output305 (.A(net305),
    .X(SS4BEG[1]));
 sg13g2_buf_1 output306 (.A(net306),
    .X(SS4BEG[2]));
 sg13g2_buf_1 output307 (.A(net307),
    .X(SS4BEG[3]));
 sg13g2_buf_1 output308 (.A(net308),
    .X(SS4BEG[4]));
 sg13g2_buf_1 output309 (.A(net309),
    .X(SS4BEG[5]));
 sg13g2_buf_1 output310 (.A(net310),
    .X(SS4BEG[6]));
 sg13g2_buf_1 output311 (.A(net311),
    .X(SS4BEG[7]));
 sg13g2_buf_1 output312 (.A(net312),
    .X(SS4BEG[8]));
 sg13g2_buf_1 output313 (.A(net313),
    .X(SS4BEG[9]));
 sg13g2_buf_1 output314 (.A(net314),
    .X(UserCLKo));
 sg13g2_buf_1 output315 (.A(\Inst_RegFile_switch_matrix.W1BEG0 ),
    .X(W1BEG[0]));
 sg13g2_buf_1 output316 (.A(\Inst_RegFile_switch_matrix.W1BEG1 ),
    .X(W1BEG[1]));
 sg13g2_buf_1 output317 (.A(\Inst_RegFile_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]));
 sg13g2_buf_1 output318 (.A(\Inst_RegFile_switch_matrix.W1BEG3 ),
    .X(W1BEG[3]));
 sg13g2_buf_1 output319 (.A(net319),
    .X(W2BEG[0]));
 sg13g2_buf_1 output320 (.A(net320),
    .X(W2BEG[1]));
 sg13g2_buf_1 output321 (.A(net321),
    .X(W2BEG[2]));
 sg13g2_buf_1 output322 (.A(net507),
    .X(W2BEG[3]));
 sg13g2_buf_1 output323 (.A(net323),
    .X(W2BEG[4]));
 sg13g2_buf_1 output324 (.A(net324),
    .X(W2BEG[5]));
 sg13g2_buf_1 output325 (.A(net325),
    .X(W2BEG[6]));
 sg13g2_buf_1 output326 (.A(net326),
    .X(W2BEG[7]));
 sg13g2_buf_1 output327 (.A(net327),
    .X(W2BEGb[0]));
 sg13g2_buf_1 output328 (.A(net328),
    .X(W2BEGb[1]));
 sg13g2_buf_1 output329 (.A(net329),
    .X(W2BEGb[2]));
 sg13g2_buf_1 output330 (.A(net330),
    .X(W2BEGb[3]));
 sg13g2_buf_1 output331 (.A(net331),
    .X(W2BEGb[4]));
 sg13g2_buf_1 output332 (.A(net332),
    .X(W2BEGb[5]));
 sg13g2_buf_1 output333 (.A(net333),
    .X(W2BEGb[6]));
 sg13g2_buf_1 output334 (.A(net334),
    .X(W2BEGb[7]));
 sg13g2_buf_1 output335 (.A(net335),
    .X(W6BEG[0]));
 sg13g2_buf_1 output336 (.A(net336),
    .X(W6BEG[10]));
 sg13g2_buf_1 output337 (.A(\Inst_RegFile_switch_matrix.W6BEG1 ),
    .X(W6BEG[11]));
 sg13g2_buf_1 output338 (.A(net338),
    .X(W6BEG[1]));
 sg13g2_buf_1 output339 (.A(net339),
    .X(W6BEG[2]));
 sg13g2_buf_1 output340 (.A(net340),
    .X(W6BEG[3]));
 sg13g2_buf_1 output341 (.A(net341),
    .X(W6BEG[4]));
 sg13g2_buf_1 output342 (.A(net342),
    .X(W6BEG[5]));
 sg13g2_buf_1 output343 (.A(net343),
    .X(W6BEG[6]));
 sg13g2_buf_1 output344 (.A(net344),
    .X(W6BEG[7]));
 sg13g2_buf_1 output345 (.A(net345),
    .X(W6BEG[8]));
 sg13g2_buf_1 output346 (.A(net346),
    .X(W6BEG[9]));
 sg13g2_buf_1 output347 (.A(net347),
    .X(WW4BEG[0]));
 sg13g2_buf_1 output348 (.A(net348),
    .X(WW4BEG[10]));
 sg13g2_buf_1 output349 (.A(net349),
    .X(WW4BEG[11]));
 sg13g2_buf_1 output350 (.A(net350),
    .X(WW4BEG[12]));
 sg13g2_buf_1 output351 (.A(\Inst_RegFile_switch_matrix.WW4BEG1 ),
    .X(WW4BEG[13]));
 sg13g2_buf_1 output352 (.A(net352),
    .X(WW4BEG[14]));
 sg13g2_buf_1 output353 (.A(net353),
    .X(WW4BEG[15]));
 sg13g2_buf_1 output354 (.A(net354),
    .X(WW4BEG[1]));
 sg13g2_buf_1 output355 (.A(net355),
    .X(WW4BEG[2]));
 sg13g2_buf_1 output356 (.A(net356),
    .X(WW4BEG[3]));
 sg13g2_buf_1 output357 (.A(net357),
    .X(WW4BEG[4]));
 sg13g2_buf_1 output358 (.A(net358),
    .X(WW4BEG[5]));
 sg13g2_buf_1 output359 (.A(net359),
    .X(WW4BEG[6]));
 sg13g2_buf_1 output360 (.A(net360),
    .X(WW4BEG[7]));
 sg13g2_buf_1 output361 (.A(net361),
    .X(WW4BEG[8]));
 sg13g2_buf_1 output362 (.A(net362),
    .X(WW4BEG[9]));
 sg13g2_tiehi _3381__363 (.L_HI(net363));
 sg13g2_dlygate4sd1_1 rebuffer2 (.A(_0388_),
    .X(net500));
 sg13g2_dlygate4sd1_1 rebuffer3 (.A(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .X(net501));
 sg13g2_dlygate4sd1_1 rebuffer4 (.A(_0137_),
    .X(net502));
 sg13g2_buf_2 rebuffer8 (.A(AD0),
    .X(net506));
 sg13g2_buf_2 rebuffer9 (.A(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .X(net507));
 sg13g2_dlygate4sd1_1 rebuffer10 (.A(net526),
    .X(net508));
 sg13g2_buf_2 rebuffer11 (.A(net527),
    .X(net509));
 sg13g2_buf_8 rebuffer12 (.A(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .X(net510));
 sg13g2_dlygate4sd1_1 rebuffer14 (.A(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .X(net512));
 sg13g2_buf_16 rebuffer15 (.X(net513),
    .A(net533));
 sg13g2_dlygate4sd1_1 rebuffer16 (.A(net513),
    .X(net514));
 sg13g2_buf_8 rebuffer17 (.A(AD1),
    .X(net515));
 sg13g2_dlygate4sd1_1 rebuffer19 (.A(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .X(net517));
 sg13g2_buf_2 rebuffer21 (.A(_0491_),
    .X(net519));
 sg13g2_buf_8 rebuffer22 (.A(_0186_),
    .X(net520));
 sg13g2_dlygate4sd1_1 rebuffer23 (.A(_0429_),
    .X(net521));
 sg13g2_dlygate4sd1_1 rebuffer24 (.A(_0429_),
    .X(net522));
 sg13g2_dlygate4sd1_1 rebuffer25 (.A(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .X(net523));
 sg13g2_dlygate4sd1_1 rebuffer26 (.A(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .X(net524));
 sg13g2_buf_8 rebuffer34 (.A(_0491_),
    .X(net532));
 sg13g2_buf_8 rebuffer35 (.A(AD2),
    .X(net533));
 sg13g2_dlygate4sd1_1 rebuffer39 (.A(net538),
    .X(net537));
 sg13g2_dlygate4sd1_1 rebuffer40 (.A(net539),
    .X(net538));
 sg13g2_dlygate4sd1_1 rebuffer41 (.A(net540),
    .X(net539));
 sg13g2_dlygate4sd1_1 rebuffer42 (.A(net541),
    .X(net540));
 sg13g2_dlygate4sd1_1 rebuffer43 (.A(net542),
    .X(net541));
 sg13g2_dlygate4sd1_1 rebuffer44 (.A(net543),
    .X(net542));
 sg13g2_dlygate4sd1_1 rebuffer45 (.A(net544),
    .X(net543));
 sg13g2_dlygate4sd1_1 rebuffer46 (.A(net545),
    .X(net544));
 sg13g2_dlygate4sd1_1 rebuffer47 (.A(net546),
    .X(net545));
 sg13g2_dlygate4sd1_1 rebuffer48 (.A(net547),
    .X(net546));
 sg13g2_dlygate4sd1_1 rebuffer49 (.A(net548),
    .X(net547));
 sg13g2_dlygate4sd1_1 rebuffer50 (.A(net549),
    .X(net548));
 sg13g2_dlygate4sd1_1 rebuffer51 (.A(net550),
    .X(net549));
 sg13g2_dlygate4sd1_1 rebuffer52 (.A(net551),
    .X(net550));
 sg13g2_buf_2 rebuffer53 (.A(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .X(net551));
 sg13g2_buf_2 rebuffer65 (.A(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .X(net563));
 sg13g2_dlygate4sd1_1 rebuffer219 (.A(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .X(net717));
 sg13g2_dlygate4sd1_1 rebuffer220 (.A(net965),
    .X(net718));
 sg13g2_dlygate4sd1_1 rebuffer221 (.A(net965),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold245 (.A(\Inst_RegFile_32x4.mem[10][3] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold246 (.A(\Inst_RegFile_32x4.mem[26][3] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold247 (.A(\Inst_RegFile_32x4.mem[2][2] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold248 (.A(\Inst_RegFile_32x4.mem[6][1] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold249 (.A(\Inst_RegFile_32x4.mem[8][1] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold250 (.A(\Inst_RegFile_32x4.mem[8][3] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold251 (.A(\Inst_RegFile_32x4.mem[0][3] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold252 (.A(\Inst_RegFile_32x4.mem[15][1] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold253 (.A(\Inst_RegFile_32x4.mem[13][1] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold254 (.A(\Inst_RegFile_32x4.mem[15][2] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold255 (.A(\Inst_RegFile_32x4.mem[13][2] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold256 (.A(\Inst_RegFile_32x4.mem[10][1] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold257 (.A(\Inst_RegFile_32x4.mem[26][1] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold258 (.A(\Inst_RegFile_32x4.mem[14][0] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold259 (.A(\Inst_RegFile_32x4.mem[26][0] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold260 (.A(\Inst_RegFile_32x4.mem[22][0] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold261 (.A(\Inst_RegFile_32x4.mem[10][0] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold262 (.A(\Inst_RegFile_32x4.mem[15][0] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold263 (.A(\Inst_RegFile_32x4.mem[20][2] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold264 (.A(\Inst_RegFile_32x4.mem[20][0] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold265 (.A(\Inst_RegFile_32x4.mem[20][1] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold266 (.A(\Inst_RegFile_32x4.mem[5][2] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold267 (.A(\Inst_RegFile_32x4.mem[1][1] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold268 (.A(\Inst_RegFile_32x4.mem[14][2] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold269 (.A(\Inst_RegFile_32x4.mem[24][1] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold270 (.A(\Inst_RegFile_32x4.mem[26][2] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold271 (.A(\Inst_RegFile_32x4.mem[28][1] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold272 (.A(\Inst_RegFile_32x4.mem[7][1] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold273 (.A(\Inst_RegFile_32x4.mem[12][1] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold274 (.A(\Inst_RegFile_32x4.mem[29][0] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold275 (.A(\Inst_RegFile_32x4.mem[1][3] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold276 (.A(\Inst_RegFile_32x4.mem[16][0] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold277 (.A(\Inst_RegFile_32x4.mem[30][0] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold278 (.A(\Inst_RegFile_32x4.mem[28][2] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold279 (.A(\Inst_RegFile_32x4.mem[5][0] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold280 (.A(\Inst_RegFile_32x4.mem[14][3] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold281 (.A(\Inst_RegFile_32x4.mem[18][0] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold282 (.A(\Inst_RegFile_32x4.mem[3][2] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold283 (.A(\Inst_RegFile_32x4.mem[19][0] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold284 (.A(\Inst_RegFile_32x4.mem[25][2] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold285 (.A(\Inst_RegFile_32x4.mem[19][3] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold286 (.A(\Inst_RegFile_32x4.mem[1][2] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold287 (.A(\Inst_RegFile_32x4.mem[17][2] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold288 (.A(\Inst_RegFile_32x4.mem[7][3] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold289 (.A(\Inst_RegFile_32x4.mem[30][3] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold290 (.A(\Inst_RegFile_32x4.mem[5][1] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold291 (.A(\Inst_RegFile_32x4.mem[28][3] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold292 (.A(\Inst_RegFile_32x4.mem[11][3] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold293 (.A(\Inst_RegFile_32x4.mem[3][3] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold294 (.A(\Inst_RegFile_32x4.mem[3][0] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold295 (.A(\Inst_RegFile_32x4.mem[22][1] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold296 (.A(\Inst_RegFile_32x4.mem[27][1] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold297 (.A(\Inst_RegFile_32x4.mem[22][3] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold298 (.A(\Inst_RegFile_32x4.mem[11][1] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold299 (.A(\Inst_RegFile_32x4.mem[5][3] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold300 (.A(\Inst_RegFile_32x4.mem[17][0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold301 (.A(\Inst_RegFile_32x4.mem[24][3] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold302 (.A(\Inst_RegFile_32x4.mem[29][1] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold303 (.A(\Inst_RegFile_32x4.mem[3][1] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold304 (.A(\Inst_RegFile_32x4.mem[21][2] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold305 (.A(\Inst_RegFile_32x4.mem[7][2] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold306 (.A(\Inst_RegFile_32x4.mem[11][0] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold307 (.A(\Inst_RegFile_32x4.mem[24][2] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold308 (.A(\Inst_RegFile_32x4.mem[14][1] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold309 (.A(\Inst_RegFile_32x4.mem[27][0] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold310 (.A(\Inst_RegFile_32x4.mem[29][2] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold311 (.A(\Inst_RegFile_32x4.mem[29][3] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold312 (.A(\Inst_RegFile_32x4.mem[25][1] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold313 (.A(\Inst_RegFile_32x4.mem[9][3] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold314 (.A(\Inst_RegFile_32x4.mem[28][0] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold315 (.A(\Inst_RegFile_32x4.mem[12][2] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold316 (.A(\Inst_RegFile_32x4.mem[21][3] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold317 (.A(\Inst_RegFile_32x4.mem[21][0] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold318 (.A(\Inst_RegFile_32x4.mem[12][3] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold319 (.A(\Inst_RegFile_32x4.mem[20][3] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold320 (.A(\Inst_RegFile_32x4.mem[16][3] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold321 (.A(\Inst_RegFile_32x4.mem[27][2] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold322 (.A(\Inst_RegFile_32x4.mem[30][1] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold323 (.A(\Inst_RegFile_32x4.mem[9][0] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold324 (.A(\Inst_RegFile_32x4.mem[17][3] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold325 (.A(\Inst_RegFile_32x4.mem[9][2] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold326 (.A(\Inst_RegFile_32x4.mem[31][0] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold327 (.A(\Inst_RegFile_32x4.mem[12][0] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold328 (.A(\Inst_RegFile_32x4.mem[19][1] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold329 (.A(\Inst_RegFile_32x4.mem[31][1] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold330 (.A(\Inst_RegFile_32x4.mem[23][3] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold331 (.A(\Inst_RegFile_32x4.mem[31][2] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold332 (.A(\Inst_RegFile_32x4.mem[25][3] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold333 (.A(\Inst_RegFile_32x4.mem[9][1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold334 (.A(\Inst_RegFile_32x4.mem[23][1] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold335 (.A(\Inst_RegFile_32x4.mem[11][2] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold336 (.A(\Inst_RegFile_32x4.mem[17][1] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold337 (.A(\Inst_RegFile_32x4.mem[7][0] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold338 (.A(\Inst_RegFile_32x4.mem[18][1] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold339 (.A(\Inst_RegFile_32x4.mem[18][3] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold340 (.A(\Inst_RegFile_32x4.mem[21][1] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold341 (.A(\Inst_RegFile_32x4.mem[19][2] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold342 (.A(\Inst_RegFile_32x4.mem[22][2] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold343 (.A(\Inst_RegFile_32x4.mem[23][0] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold344 (.A(\Inst_RegFile_32x4.mem[30][2] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold345 (.A(\Inst_RegFile_32x4.mem[1][0] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold346 (.A(\Inst_RegFile_32x4.mem[24][0] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold347 (.A(\Inst_RegFile_32x4.mem[16][1] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold348 (.A(\Inst_RegFile_32x4.mem[18][2] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold349 (.A(\Inst_RegFile_32x4.mem[23][2] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold350 (.A(\Inst_RegFile_32x4.mem[16][2] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold351 (.A(\Inst_RegFile_32x4.mem[27][3] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold352 (.A(\Inst_RegFile_32x4.mem[25][0] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold353 (.A(\Inst_RegFile_32x4.mem[31][3] ),
    .X(net851));
 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_2 ();
 sg13g2_fill_2 FILLER_0_44 ();
 sg13g2_fill_1 FILLER_0_46 ();
 sg13g2_fill_2 FILLER_0_88 ();
 sg13g2_fill_1 FILLER_0_90 ();
 sg13g2_fill_2 FILLER_0_111 ();
 sg13g2_fill_2 FILLER_0_285 ();
 sg13g2_fill_1 FILLER_0_287 ();
 sg13g2_fill_2 FILLER_0_375 ();
 sg13g2_fill_2 FILLER_0_518 ();
 sg13g2_fill_2 FILLER_0_528 ();
 sg13g2_fill_1 FILLER_0_530 ();
 sg13g2_fill_2 FILLER_1_16 ();
 sg13g2_fill_1 FILLER_1_18 ();
 sg13g2_fill_2 FILLER_1_63 ();
 sg13g2_fill_2 FILLER_1_69 ();
 sg13g2_fill_1 FILLER_1_71 ();
 sg13g2_fill_2 FILLER_1_80 ();
 sg13g2_fill_1 FILLER_1_82 ();
 sg13g2_fill_1 FILLER_1_95 ();
 sg13g2_fill_2 FILLER_1_120 ();
 sg13g2_fill_1 FILLER_1_126 ();
 sg13g2_fill_2 FILLER_1_143 ();
 sg13g2_fill_2 FILLER_1_219 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_fill_2 FILLER_1_402 ();
 sg13g2_fill_1 FILLER_1_404 ();
 sg13g2_fill_2 FILLER_1_524 ();
 sg13g2_fill_1 FILLER_1_526 ();
 sg13g2_fill_2 FILLER_2_40 ();
 sg13g2_fill_1 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_fill_2 FILLER_2_77 ();
 sg13g2_fill_1 FILLER_2_140 ();
 sg13g2_fill_2 FILLER_2_177 ();
 sg13g2_fill_1 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_217 ();
 sg13g2_fill_1 FILLER_2_265 ();
 sg13g2_fill_2 FILLER_2_271 ();
 sg13g2_fill_2 FILLER_2_338 ();
 sg13g2_fill_1 FILLER_2_376 ();
 sg13g2_fill_2 FILLER_2_403 ();
 sg13g2_fill_1 FILLER_2_425 ();
 sg13g2_fill_1 FILLER_2_513 ();
 sg13g2_fill_2 FILLER_3_36 ();
 sg13g2_decap_8 FILLER_3_58 ();
 sg13g2_decap_8 FILLER_3_65 ();
 sg13g2_decap_8 FILLER_3_72 ();
 sg13g2_fill_2 FILLER_3_79 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_104 ();
 sg13g2_fill_2 FILLER_3_123 ();
 sg13g2_fill_1 FILLER_3_125 ();
 sg13g2_fill_1 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_191 ();
 sg13g2_fill_1 FILLER_3_205 ();
 sg13g2_fill_2 FILLER_3_227 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_303 ();
 sg13g2_fill_2 FILLER_3_314 ();
 sg13g2_fill_1 FILLER_3_316 ();
 sg13g2_fill_2 FILLER_3_342 ();
 sg13g2_fill_1 FILLER_3_354 ();
 sg13g2_fill_2 FILLER_3_411 ();
 sg13g2_fill_1 FILLER_3_413 ();
 sg13g2_fill_2 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_505 ();
 sg13g2_fill_1 FILLER_3_507 ();
 sg13g2_fill_2 FILLER_3_512 ();
 sg13g2_fill_1 FILLER_3_518 ();
 sg13g2_fill_2 FILLER_4_8 ();
 sg13g2_fill_1 FILLER_4_10 ();
 sg13g2_fill_2 FILLER_4_31 ();
 sg13g2_fill_1 FILLER_4_38 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_4 FILLER_4_60 ();
 sg13g2_fill_2 FILLER_4_64 ();
 sg13g2_decap_8 FILLER_4_71 ();
 sg13g2_decap_4 FILLER_4_78 ();
 sg13g2_fill_2 FILLER_4_82 ();
 sg13g2_fill_2 FILLER_4_122 ();
 sg13g2_fill_1 FILLER_4_145 ();
 sg13g2_fill_2 FILLER_4_155 ();
 sg13g2_fill_1 FILLER_4_157 ();
 sg13g2_fill_1 FILLER_4_222 ();
 sg13g2_fill_2 FILLER_4_261 ();
 sg13g2_fill_2 FILLER_4_351 ();
 sg13g2_fill_1 FILLER_4_353 ();
 sg13g2_fill_1 FILLER_4_409 ();
 sg13g2_fill_1 FILLER_4_460 ();
 sg13g2_fill_2 FILLER_4_522 ();
 sg13g2_fill_1 FILLER_4_524 ();
 sg13g2_fill_2 FILLER_4_529 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_2 ();
 sg13g2_fill_1 FILLER_5_20 ();
 sg13g2_fill_1 FILLER_5_26 ();
 sg13g2_fill_1 FILLER_5_71 ();
 sg13g2_fill_2 FILLER_5_89 ();
 sg13g2_fill_1 FILLER_5_108 ();
 sg13g2_fill_2 FILLER_5_114 ();
 sg13g2_fill_1 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_1 FILLER_5_150 ();
 sg13g2_fill_2 FILLER_5_173 ();
 sg13g2_fill_2 FILLER_5_268 ();
 sg13g2_fill_2 FILLER_5_310 ();
 sg13g2_fill_2 FILLER_5_338 ();
 sg13g2_fill_1 FILLER_5_340 ();
 sg13g2_fill_2 FILLER_5_412 ();
 sg13g2_fill_1 FILLER_5_475 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_44 ();
 sg13g2_fill_1 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_91 ();
 sg13g2_fill_1 FILLER_6_112 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_274 ();
 sg13g2_fill_2 FILLER_6_319 ();
 sg13g2_fill_2 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_358 ();
 sg13g2_fill_2 FILLER_6_381 ();
 sg13g2_fill_1 FILLER_6_383 ();
 sg13g2_fill_2 FILLER_6_405 ();
 sg13g2_fill_1 FILLER_6_407 ();
 sg13g2_fill_2 FILLER_6_449 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_fill_2 FILLER_7_32 ();
 sg13g2_fill_2 FILLER_7_57 ();
 sg13g2_fill_2 FILLER_7_69 ();
 sg13g2_fill_1 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_210 ();
 sg13g2_fill_2 FILLER_7_257 ();
 sg13g2_fill_2 FILLER_7_303 ();
 sg13g2_fill_1 FILLER_7_358 ();
 sg13g2_fill_2 FILLER_7_460 ();
 sg13g2_fill_2 FILLER_7_501 ();
 sg13g2_fill_1 FILLER_7_503 ();
 sg13g2_fill_1 FILLER_7_530 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_50 ();
 sg13g2_fill_1 FILLER_8_52 ();
 sg13g2_fill_2 FILLER_8_99 ();
 sg13g2_fill_1 FILLER_8_101 ();
 sg13g2_fill_2 FILLER_8_156 ();
 sg13g2_fill_2 FILLER_8_188 ();
 sg13g2_fill_2 FILLER_8_207 ();
 sg13g2_fill_2 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_339 ();
 sg13g2_fill_2 FILLER_8_457 ();
 sg13g2_fill_1 FILLER_8_459 ();
 sg13g2_fill_2 FILLER_8_481 ();
 sg13g2_fill_1 FILLER_8_483 ();
 sg13g2_fill_2 FILLER_8_494 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_2 ();
 sg13g2_fill_2 FILLER_9_20 ();
 sg13g2_fill_1 FILLER_9_22 ();
 sg13g2_fill_2 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_132 ();
 sg13g2_fill_2 FILLER_9_164 ();
 sg13g2_fill_1 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_244 ();
 sg13g2_fill_2 FILLER_9_318 ();
 sg13g2_fill_1 FILLER_9_320 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_fill_2 FILLER_9_398 ();
 sg13g2_fill_1 FILLER_9_458 ();
 sg13g2_fill_1 FILLER_9_530 ();
 sg13g2_fill_2 FILLER_10_37 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_fill_2 FILLER_10_55 ();
 sg13g2_fill_1 FILLER_10_82 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_152 ();
 sg13g2_fill_1 FILLER_10_179 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_266 ();
 sg13g2_fill_1 FILLER_10_363 ();
 sg13g2_fill_1 FILLER_10_374 ();
 sg13g2_fill_1 FILLER_10_419 ();
 sg13g2_fill_2 FILLER_10_446 ();
 sg13g2_fill_1 FILLER_10_448 ();
 sg13g2_fill_1 FILLER_10_469 ();
 sg13g2_fill_2 FILLER_10_489 ();
 sg13g2_fill_1 FILLER_10_491 ();
 sg13g2_fill_2 FILLER_10_502 ();
 sg13g2_fill_1 FILLER_10_530 ();
 sg13g2_fill_2 FILLER_11_8 ();
 sg13g2_fill_1 FILLER_11_10 ();
 sg13g2_fill_1 FILLER_11_59 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_117 ();
 sg13g2_fill_2 FILLER_11_123 ();
 sg13g2_fill_1 FILLER_11_125 ();
 sg13g2_fill_2 FILLER_11_129 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_287 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_fill_1 FILLER_11_396 ();
 sg13g2_fill_1 FILLER_11_450 ();
 sg13g2_fill_2 FILLER_11_456 ();
 sg13g2_fill_1 FILLER_11_458 ();
 sg13g2_fill_1 FILLER_11_485 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_166 ();
 sg13g2_fill_2 FILLER_12_194 ();
 sg13g2_fill_2 FILLER_12_319 ();
 sg13g2_fill_1 FILLER_12_321 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_439 ();
 sg13g2_fill_1 FILLER_12_441 ();
 sg13g2_fill_2 FILLER_12_448 ();
 sg13g2_fill_1 FILLER_12_450 ();
 sg13g2_fill_2 FILLER_12_477 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_23 ();
 sg13g2_fill_2 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_133 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_decap_4 FILLER_13_153 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_fill_1 FILLER_13_285 ();
 sg13g2_fill_1 FILLER_13_332 ();
 sg13g2_fill_2 FILLER_13_402 ();
 sg13g2_fill_1 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_421 ();
 sg13g2_fill_2 FILLER_13_447 ();
 sg13g2_fill_1 FILLER_13_449 ();
 sg13g2_fill_1 FILLER_13_530 ();
 sg13g2_fill_1 FILLER_14_8 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_63 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_243 ();
 sg13g2_fill_2 FILLER_14_282 ();
 sg13g2_fill_1 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_301 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_fill_2 FILLER_14_395 ();
 sg13g2_fill_2 FILLER_14_480 ();
 sg13g2_fill_1 FILLER_14_482 ();
 sg13g2_fill_2 FILLER_14_498 ();
 sg13g2_fill_1 FILLER_14_509 ();
 sg13g2_fill_1 FILLER_14_530 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_49 ();
 sg13g2_fill_2 FILLER_15_74 ();
 sg13g2_fill_1 FILLER_15_76 ();
 sg13g2_fill_2 FILLER_15_111 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_fill_2 FILLER_15_158 ();
 sg13g2_fill_2 FILLER_15_181 ();
 sg13g2_fill_2 FILLER_15_208 ();
 sg13g2_fill_1 FILLER_15_210 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_1 FILLER_15_260 ();
 sg13g2_fill_1 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_323 ();
 sg13g2_fill_2 FILLER_15_360 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_15_438 ();
 sg13g2_fill_2 FILLER_15_449 ();
 sg13g2_fill_1 FILLER_15_487 ();
 sg13g2_fill_2 FILLER_15_528 ();
 sg13g2_fill_1 FILLER_15_530 ();
 sg13g2_fill_2 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_51 ();
 sg13g2_fill_2 FILLER_16_72 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_101 ();
 sg13g2_decap_4 FILLER_16_108 ();
 sg13g2_fill_2 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_131 ();
 sg13g2_decap_4 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_fill_2 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_258 ();
 sg13g2_fill_2 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_fill_2 FILLER_16_411 ();
 sg13g2_fill_1 FILLER_16_413 ();
 sg13g2_fill_1 FILLER_16_444 ();
 sg13g2_fill_2 FILLER_16_457 ();
 sg13g2_fill_1 FILLER_16_459 ();
 sg13g2_fill_2 FILLER_16_481 ();
 sg13g2_fill_1 FILLER_16_483 ();
 sg13g2_fill_2 FILLER_16_519 ();
 sg13g2_fill_1 FILLER_16_530 ();
 sg13g2_fill_2 FILLER_17_38 ();
 sg13g2_fill_2 FILLER_17_82 ();
 sg13g2_fill_2 FILLER_17_135 ();
 sg13g2_fill_1 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_8 FILLER_17_183 ();
 sg13g2_decap_4 FILLER_17_190 ();
 sg13g2_fill_1 FILLER_17_194 ();
 sg13g2_fill_2 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_267 ();
 sg13g2_fill_2 FILLER_17_314 ();
 sg13g2_fill_1 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_360 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_1 FILLER_17_463 ();
 sg13g2_fill_2 FILLER_17_474 ();
 sg13g2_fill_1 FILLER_17_530 ();
 sg13g2_fill_1 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_73 ();
 sg13g2_decap_4 FILLER_18_100 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_decap_4 FILLER_18_130 ();
 sg13g2_fill_1 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_fill_1 FILLER_18_305 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_441 ();
 sg13g2_fill_2 FILLER_18_471 ();
 sg13g2_fill_2 FILLER_18_492 ();
 sg13g2_fill_1 FILLER_18_494 ();
 sg13g2_fill_2 FILLER_19_8 ();
 sg13g2_fill_1 FILLER_19_47 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_fill_2 FILLER_19_107 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_decap_4 FILLER_19_127 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_257 ();
 sg13g2_fill_2 FILLER_19_283 ();
 sg13g2_fill_1 FILLER_19_285 ();
 sg13g2_fill_1 FILLER_19_307 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_fill_1 FILLER_19_337 ();
 sg13g2_fill_2 FILLER_19_352 ();
 sg13g2_fill_1 FILLER_19_354 ();
 sg13g2_fill_2 FILLER_19_379 ();
 sg13g2_fill_1 FILLER_19_381 ();
 sg13g2_fill_2 FILLER_19_419 ();
 sg13g2_fill_1 FILLER_19_421 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_37 ();
 sg13g2_fill_2 FILLER_20_111 ();
 sg13g2_fill_2 FILLER_20_159 ();
 sg13g2_fill_2 FILLER_20_224 ();
 sg13g2_fill_1 FILLER_20_226 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_264 ();
 sg13g2_fill_1 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_308 ();
 sg13g2_fill_1 FILLER_20_310 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_fill_1 FILLER_20_338 ();
 sg13g2_fill_2 FILLER_20_365 ();
 sg13g2_fill_1 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_1 FILLER_21_20 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_78 ();
 sg13g2_decap_8 FILLER_21_115 ();
 sg13g2_fill_2 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_2 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_186 ();
 sg13g2_fill_2 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_436 ();
 sg13g2_fill_1 FILLER_21_448 ();
 sg13g2_fill_1 FILLER_21_483 ();
 sg13g2_fill_2 FILLER_21_503 ();
 sg13g2_decap_4 FILLER_22_70 ();
 sg13g2_decap_4 FILLER_22_120 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_278 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_351 ();
 sg13g2_fill_1 FILLER_22_436 ();
 sg13g2_fill_2 FILLER_22_491 ();
 sg13g2_fill_2 FILLER_22_529 ();
 sg13g2_fill_2 FILLER_23_38 ();
 sg13g2_fill_1 FILLER_23_40 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_decap_8 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_decap_4 FILLER_23_216 ();
 sg13g2_fill_2 FILLER_23_220 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_fill_2 FILLER_23_405 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_2 FILLER_23_465 ();
 sg13g2_fill_1 FILLER_23_467 ();
 sg13g2_fill_2 FILLER_23_489 ();
 sg13g2_fill_2 FILLER_23_501 ();
 sg13g2_fill_2 FILLER_23_529 ();
 sg13g2_fill_2 FILLER_24_8 ();
 sg13g2_fill_1 FILLER_24_10 ();
 sg13g2_fill_2 FILLER_24_28 ();
 sg13g2_fill_1 FILLER_24_65 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_113 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_fill_2 FILLER_24_185 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_fill_2 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_fill_1 FILLER_24_432 ();
 sg13g2_fill_2 FILLER_24_454 ();
 sg13g2_fill_1 FILLER_24_498 ();
 sg13g2_fill_2 FILLER_24_529 ();
 sg13g2_fill_2 FILLER_25_8 ();
 sg13g2_fill_1 FILLER_25_10 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_34 ();
 sg13g2_decap_4 FILLER_25_78 ();
 sg13g2_fill_2 FILLER_25_82 ();
 sg13g2_decap_8 FILLER_25_135 ();
 sg13g2_decap_4 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_274 ();
 sg13g2_fill_1 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_340 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_2 FILLER_25_362 ();
 sg13g2_fill_2 FILLER_25_420 ();
 sg13g2_fill_2 FILLER_25_503 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_decap_4 FILLER_26_69 ();
 sg13g2_fill_2 FILLER_26_115 ();
 sg13g2_fill_1 FILLER_26_127 ();
 sg13g2_decap_8 FILLER_26_145 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_fill_2 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_fill_1 FILLER_26_363 ();
 sg13g2_fill_1 FILLER_26_451 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_2 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_fill_2 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_fill_2 FILLER_27_335 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_348 ();
 sg13g2_fill_2 FILLER_27_375 ();
 sg13g2_fill_1 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_fill_2 FILLER_27_435 ();
 sg13g2_fill_1 FILLER_27_437 ();
 sg13g2_fill_1 FILLER_27_495 ();
 sg13g2_decap_8 FILLER_28_36 ();
 sg13g2_fill_1 FILLER_28_43 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_fill_1 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_fill_2 FILLER_28_154 ();
 sg13g2_fill_1 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_decap_4 FILLER_28_296 ();
 sg13g2_fill_2 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_348 ();
 sg13g2_fill_1 FILLER_28_350 ();
 sg13g2_fill_2 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_377 ();
 sg13g2_fill_2 FILLER_28_443 ();
 sg13g2_fill_1 FILLER_28_445 ();
 sg13g2_fill_1 FILLER_28_464 ();
 sg13g2_fill_2 FILLER_28_474 ();
 sg13g2_fill_2 FILLER_28_529 ();
 sg13g2_fill_1 FILLER_29_38 ();
 sg13g2_decap_4 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_71 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_fill_1 FILLER_29_78 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_210 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_308 ();
 sg13g2_fill_2 FILLER_29_334 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_352 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_466 ();
 sg13g2_fill_1 FILLER_29_530 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_73 ();
 sg13g2_fill_2 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_fill_1 FILLER_30_112 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_fill_1 FILLER_30_123 ();
 sg13g2_fill_2 FILLER_30_158 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_decap_4 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_484 ();
 sg13g2_fill_1 FILLER_30_496 ();
 sg13g2_fill_2 FILLER_31_8 ();
 sg13g2_fill_2 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_90 ();
 sg13g2_decap_8 FILLER_31_139 ();
 sg13g2_decap_4 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_150 ();
 sg13g2_fill_2 FILLER_31_193 ();
 sg13g2_decap_4 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_31_377 ();
 sg13g2_fill_2 FILLER_31_445 ();
 sg13g2_fill_1 FILLER_31_447 ();
 sg13g2_fill_2 FILLER_31_490 ();
 sg13g2_fill_2 FILLER_31_511 ();
 sg13g2_fill_1 FILLER_31_530 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_2 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_41 ();
 sg13g2_decap_8 FILLER_32_48 ();
 sg13g2_decap_4 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_decap_4 FILLER_32_113 ();
 sg13g2_fill_1 FILLER_32_117 ();
 sg13g2_decap_4 FILLER_32_143 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_fill_1 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_330 ();
 sg13g2_fill_1 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_fill_1 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_476 ();
 sg13g2_fill_1 FILLER_32_487 ();
 sg13g2_fill_1 FILLER_32_503 ();
 sg13g2_fill_1 FILLER_32_530 ();
 sg13g2_fill_1 FILLER_33_55 ();
 sg13g2_decap_4 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_decap_4 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_137 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_274 ();
 sg13g2_decap_4 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_346 ();
 sg13g2_fill_1 FILLER_33_348 ();
 sg13g2_fill_1 FILLER_33_383 ();
 sg13g2_fill_1 FILLER_33_407 ();
 sg13g2_fill_2 FILLER_33_433 ();
 sg13g2_fill_2 FILLER_33_462 ();
 sg13g2_fill_1 FILLER_33_530 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_20 ();
 sg13g2_decap_8 FILLER_34_76 ();
 sg13g2_decap_8 FILLER_34_83 ();
 sg13g2_decap_8 FILLER_34_150 ();
 sg13g2_decap_4 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_184 ();
 sg13g2_fill_1 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_396 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_fill_1 FILLER_34_409 ();
 sg13g2_fill_1 FILLER_34_423 ();
 sg13g2_fill_1 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_34_444 ();
 sg13g2_fill_2 FILLER_34_453 ();
 sg13g2_fill_1 FILLER_34_455 ();
 sg13g2_fill_2 FILLER_34_473 ();
 sg13g2_fill_1 FILLER_34_475 ();
 sg13g2_fill_2 FILLER_34_528 ();
 sg13g2_fill_1 FILLER_34_530 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_47 ();
 sg13g2_fill_2 FILLER_35_54 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_decap_4 FILLER_35_81 ();
 sg13g2_fill_2 FILLER_35_106 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_212 ();
 sg13g2_fill_1 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_250 ();
 sg13g2_decap_8 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_277 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_291 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_fill_2 FILLER_35_356 ();
 sg13g2_fill_2 FILLER_35_391 ();
 sg13g2_fill_2 FILLER_35_413 ();
 sg13g2_fill_1 FILLER_35_469 ();
 sg13g2_fill_2 FILLER_35_484 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_decap_8 FILLER_36_45 ();
 sg13g2_fill_2 FILLER_36_52 ();
 sg13g2_fill_2 FILLER_36_71 ();
 sg13g2_fill_1 FILLER_36_73 ();
 sg13g2_fill_2 FILLER_36_113 ();
 sg13g2_fill_2 FILLER_36_133 ();
 sg13g2_decap_4 FILLER_36_164 ();
 sg13g2_fill_2 FILLER_36_168 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_231 ();
 sg13g2_fill_1 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_412 ();
 sg13g2_fill_1 FILLER_36_414 ();
 sg13g2_fill_1 FILLER_36_456 ();
 sg13g2_fill_2 FILLER_36_477 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_24 ();
 sg13g2_decap_8 FILLER_37_43 ();
 sg13g2_decap_4 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_54 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_96 ();
 sg13g2_fill_2 FILLER_37_111 ();
 sg13g2_fill_1 FILLER_37_125 ();
 sg13g2_decap_4 FILLER_37_173 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_fill_2 FILLER_37_233 ();
 sg13g2_fill_1 FILLER_37_235 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_fill_1 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_295 ();
 sg13g2_decap_8 FILLER_37_300 ();
 sg13g2_fill_2 FILLER_37_311 ();
 sg13g2_decap_4 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_344 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_423 ();
 sg13g2_fill_1 FILLER_37_425 ();
 sg13g2_fill_2 FILLER_37_463 ();
 sg13g2_fill_1 FILLER_37_465 ();
 sg13g2_fill_2 FILLER_37_492 ();
 sg13g2_fill_1 FILLER_37_494 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_decap_8 FILLER_38_41 ();
 sg13g2_decap_4 FILLER_38_48 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_decap_4 FILLER_38_278 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_decap_4 FILLER_38_339 ();
 sg13g2_fill_2 FILLER_38_458 ();
 sg13g2_fill_1 FILLER_38_514 ();
 sg13g2_fill_2 FILLER_38_529 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_fill_2 FILLER_39_23 ();
 sg13g2_decap_8 FILLER_39_46 ();
 sg13g2_fill_2 FILLER_39_53 ();
 sg13g2_fill_2 FILLER_39_82 ();
 sg13g2_fill_2 FILLER_39_105 ();
 sg13g2_fill_1 FILLER_39_107 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_4 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_234 ();
 sg13g2_decap_8 FILLER_39_298 ();
 sg13g2_decap_4 FILLER_39_305 ();
 sg13g2_fill_1 FILLER_39_309 ();
 sg13g2_fill_1 FILLER_39_359 ();
 sg13g2_fill_2 FILLER_39_426 ();
 sg13g2_fill_2 FILLER_39_456 ();
 sg13g2_fill_2 FILLER_39_475 ();
 sg13g2_fill_1 FILLER_39_477 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_7 ();
 sg13g2_decap_4 FILLER_40_25 ();
 sg13g2_decap_8 FILLER_40_39 ();
 sg13g2_fill_1 FILLER_40_67 ();
 sg13g2_fill_2 FILLER_40_115 ();
 sg13g2_fill_1 FILLER_40_117 ();
 sg13g2_fill_1 FILLER_40_183 ();
 sg13g2_decap_8 FILLER_40_194 ();
 sg13g2_fill_1 FILLER_40_201 ();
 sg13g2_fill_2 FILLER_40_223 ();
 sg13g2_decap_8 FILLER_40_242 ();
 sg13g2_decap_8 FILLER_40_249 ();
 sg13g2_decap_8 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_263 ();
 sg13g2_decap_8 FILLER_40_285 ();
 sg13g2_decap_4 FILLER_40_292 ();
 sg13g2_fill_2 FILLER_40_296 ();
 sg13g2_fill_1 FILLER_40_341 ();
 sg13g2_fill_2 FILLER_40_402 ();
 sg13g2_fill_1 FILLER_40_414 ();
 sg13g2_fill_2 FILLER_40_425 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_29 ();
 sg13g2_fill_1 FILLER_41_36 ();
 sg13g2_fill_2 FILLER_41_79 ();
 sg13g2_fill_1 FILLER_41_81 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_89 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_fill_2 FILLER_41_130 ();
 sg13g2_fill_1 FILLER_41_200 ();
 sg13g2_fill_1 FILLER_41_218 ();
 sg13g2_fill_2 FILLER_41_223 ();
 sg13g2_fill_1 FILLER_41_242 ();
 sg13g2_decap_8 FILLER_41_281 ();
 sg13g2_decap_4 FILLER_41_288 ();
 sg13g2_fill_2 FILLER_41_292 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_fill_2 FILLER_41_322 ();
 sg13g2_fill_2 FILLER_41_362 ();
 sg13g2_fill_1 FILLER_41_402 ();
 sg13g2_fill_1 FILLER_41_426 ();
 sg13g2_fill_1 FILLER_41_530 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_4 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_11 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_2 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_94 ();
 sg13g2_decap_8 FILLER_42_101 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_184 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_fill_1 FILLER_42_196 ();
 sg13g2_decap_4 FILLER_42_218 ();
 sg13g2_fill_2 FILLER_42_237 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_decap_4 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_306 ();
 sg13g2_fill_1 FILLER_42_324 ();
 sg13g2_fill_1 FILLER_42_353 ();
 sg13g2_fill_1 FILLER_42_380 ();
 sg13g2_fill_1 FILLER_42_393 ();
 sg13g2_fill_1 FILLER_42_437 ();
 sg13g2_fill_2 FILLER_42_489 ();
 sg13g2_decap_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_65 ();
 sg13g2_decap_8 FILLER_43_97 ();
 sg13g2_fill_2 FILLER_43_104 ();
 sg13g2_fill_1 FILLER_43_106 ();
 sg13g2_fill_2 FILLER_43_148 ();
 sg13g2_fill_1 FILLER_43_150 ();
 sg13g2_decap_4 FILLER_43_191 ();
 sg13g2_fill_1 FILLER_43_195 ();
 sg13g2_fill_2 FILLER_43_217 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_281 ();
 sg13g2_fill_1 FILLER_43_283 ();
 sg13g2_decap_4 FILLER_43_301 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_fill_1 FILLER_43_346 ();
 sg13g2_fill_2 FILLER_43_380 ();
 sg13g2_fill_1 FILLER_43_407 ();
 sg13g2_fill_2 FILLER_43_465 ();
 sg13g2_fill_1 FILLER_44_20 ();
 sg13g2_fill_1 FILLER_44_73 ();
 sg13g2_fill_2 FILLER_44_153 ();
 sg13g2_fill_2 FILLER_44_176 ();
 sg13g2_fill_1 FILLER_44_192 ();
 sg13g2_fill_2 FILLER_44_241 ();
 sg13g2_decap_4 FILLER_44_294 ();
 sg13g2_fill_1 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_324 ();
 sg13g2_fill_1 FILLER_44_326 ();
 sg13g2_fill_2 FILLER_44_354 ();
 sg13g2_fill_1 FILLER_44_356 ();
 sg13g2_fill_2 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_1 FILLER_44_423 ();
 sg13g2_fill_2 FILLER_44_448 ();
 sg13g2_fill_1 FILLER_44_450 ();
 sg13g2_fill_2 FILLER_44_483 ();
 sg13g2_fill_1 FILLER_44_485 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_4 ();
 sg13g2_fill_2 FILLER_45_63 ();
 sg13g2_fill_1 FILLER_45_65 ();
 sg13g2_fill_2 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_208 ();
 sg13g2_decap_4 FILLER_45_215 ();
 sg13g2_fill_2 FILLER_45_229 ();
 sg13g2_fill_1 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_259 ();
 sg13g2_fill_1 FILLER_45_261 ();
 sg13g2_fill_1 FILLER_45_297 ();
 sg13g2_decap_4 FILLER_45_332 ();
 sg13g2_fill_1 FILLER_45_336 ();
 sg13g2_fill_2 FILLER_45_362 ();
 sg13g2_fill_1 FILLER_45_364 ();
 sg13g2_fill_1 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_411 ();
 sg13g2_fill_2 FILLER_45_430 ();
 sg13g2_fill_1 FILLER_45_458 ();
 sg13g2_fill_2 FILLER_45_494 ();
 sg13g2_fill_1 FILLER_45_496 ();
 sg13g2_fill_1 FILLER_45_530 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_33 ();
 sg13g2_decap_4 FILLER_46_61 ();
 sg13g2_fill_2 FILLER_46_69 ();
 sg13g2_fill_1 FILLER_46_71 ();
 sg13g2_decap_4 FILLER_46_92 ();
 sg13g2_fill_2 FILLER_46_96 ();
 sg13g2_fill_2 FILLER_46_147 ();
 sg13g2_fill_1 FILLER_46_149 ();
 sg13g2_fill_2 FILLER_46_160 ();
 sg13g2_decap_8 FILLER_46_206 ();
 sg13g2_fill_1 FILLER_46_213 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_292 ();
 sg13g2_fill_1 FILLER_46_310 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_326 ();
 sg13g2_decap_4 FILLER_46_333 ();
 sg13g2_fill_2 FILLER_46_337 ();
 sg13g2_fill_2 FILLER_46_356 ();
 sg13g2_fill_1 FILLER_46_358 ();
 sg13g2_fill_1 FILLER_46_391 ();
 sg13g2_fill_2 FILLER_46_413 ();
 sg13g2_fill_2 FILLER_46_445 ();
 sg13g2_fill_1 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_47_8 ();
 sg13g2_decap_8 FILLER_47_15 ();
 sg13g2_decap_8 FILLER_47_22 ();
 sg13g2_fill_2 FILLER_47_29 ();
 sg13g2_fill_1 FILLER_47_31 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_fill_1 FILLER_47_49 ();
 sg13g2_decap_4 FILLER_47_89 ();
 sg13g2_fill_2 FILLER_47_93 ();
 sg13g2_fill_2 FILLER_47_117 ();
 sg13g2_fill_2 FILLER_47_124 ();
 sg13g2_fill_2 FILLER_47_156 ();
 sg13g2_fill_1 FILLER_47_158 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_220 ();
 sg13g2_decap_8 FILLER_47_289 ();
 sg13g2_decap_4 FILLER_47_300 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_decap_8 FILLER_47_326 ();
 sg13g2_fill_1 FILLER_47_333 ();
 sg13g2_decap_4 FILLER_47_338 ();
 sg13g2_fill_1 FILLER_47_342 ();
 sg13g2_fill_1 FILLER_47_351 ();
 sg13g2_fill_2 FILLER_47_360 ();
 sg13g2_fill_2 FILLER_47_384 ();
 sg13g2_fill_1 FILLER_47_386 ();
 sg13g2_fill_2 FILLER_47_529 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_4 FILLER_48_28 ();
 sg13g2_fill_2 FILLER_48_32 ();
 sg13g2_fill_1 FILLER_48_54 ();
 sg13g2_fill_1 FILLER_48_75 ();
 sg13g2_fill_2 FILLER_48_102 ();
 sg13g2_fill_2 FILLER_48_148 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_fill_1 FILLER_48_189 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_264 ();
 sg13g2_fill_1 FILLER_48_266 ();
 sg13g2_decap_4 FILLER_48_342 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_fill_2 FILLER_48_374 ();
 sg13g2_fill_1 FILLER_48_418 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_55 ();
 sg13g2_fill_1 FILLER_49_57 ();
 sg13g2_fill_1 FILLER_49_79 ();
 sg13g2_fill_1 FILLER_49_120 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_2 FILLER_49_202 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_fill_2 FILLER_49_279 ();
 sg13g2_fill_1 FILLER_49_281 ();
 sg13g2_decap_4 FILLER_49_320 ();
 sg13g2_decap_4 FILLER_49_389 ();
 sg13g2_fill_2 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_412 ();
 sg13g2_fill_1 FILLER_49_419 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_4 FILLER_50_28 ();
 sg13g2_fill_1 FILLER_50_36 ();
 sg13g2_fill_1 FILLER_50_58 ();
 sg13g2_fill_2 FILLER_50_275 ();
 sg13g2_fill_2 FILLER_50_287 ();
 sg13g2_fill_1 FILLER_50_289 ();
 sg13g2_decap_8 FILLER_50_311 ();
 sg13g2_decap_8 FILLER_50_318 ();
 sg13g2_decap_8 FILLER_50_325 ();
 sg13g2_fill_2 FILLER_50_332 ();
 sg13g2_fill_1 FILLER_50_334 ();
 sg13g2_fill_2 FILLER_50_360 ();
 sg13g2_fill_1 FILLER_50_380 ();
 sg13g2_decap_8 FILLER_50_415 ();
 sg13g2_fill_2 FILLER_50_422 ();
 sg13g2_fill_2 FILLER_50_434 ();
 sg13g2_fill_1 FILLER_50_436 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_18 ();
 sg13g2_fill_2 FILLER_51_23 ();
 sg13g2_fill_1 FILLER_51_25 ();
 sg13g2_fill_1 FILLER_51_48 ();
 sg13g2_fill_2 FILLER_51_54 ();
 sg13g2_fill_1 FILLER_51_56 ();
 sg13g2_fill_1 FILLER_51_62 ();
 sg13g2_fill_1 FILLER_51_124 ();
 sg13g2_fill_1 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_152 ();
 sg13g2_fill_1 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_fill_2 FILLER_51_302 ();
 sg13g2_fill_1 FILLER_51_304 ();
 sg13g2_decap_8 FILLER_51_313 ();
 sg13g2_fill_2 FILLER_51_320 ();
 sg13g2_fill_1 FILLER_51_322 ();
 sg13g2_fill_2 FILLER_51_327 ();
 sg13g2_fill_1 FILLER_51_351 ();
 sg13g2_decap_4 FILLER_51_384 ();
 sg13g2_fill_1 FILLER_51_388 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_4 FILLER_51_400 ();
 sg13g2_fill_1 FILLER_51_404 ();
 sg13g2_decap_8 FILLER_51_409 ();
 sg13g2_decap_8 FILLER_51_416 ();
 sg13g2_decap_8 FILLER_51_423 ();
 sg13g2_decap_4 FILLER_51_430 ();
 sg13g2_fill_2 FILLER_51_446 ();
 sg13g2_fill_1 FILLER_51_448 ();
 sg13g2_fill_1 FILLER_51_494 ();
 sg13g2_fill_2 FILLER_51_509 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_18 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_2 FILLER_52_63 ();
 sg13g2_fill_1 FILLER_52_65 ();
 sg13g2_fill_2 FILLER_52_128 ();
 sg13g2_fill_2 FILLER_52_156 ();
 sg13g2_fill_1 FILLER_52_158 ();
 sg13g2_fill_2 FILLER_52_232 ();
 sg13g2_fill_1 FILLER_52_248 ();
 sg13g2_fill_1 FILLER_52_253 ();
 sg13g2_fill_1 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_290 ();
 sg13g2_decap_4 FILLER_52_302 ();
 sg13g2_fill_1 FILLER_52_306 ();
 sg13g2_decap_4 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_419 ();
 sg13g2_decap_8 FILLER_52_426 ();
 sg13g2_decap_8 FILLER_52_433 ();
 sg13g2_decap_8 FILLER_52_440 ();
 sg13g2_decap_8 FILLER_52_447 ();
 sg13g2_decap_4 FILLER_52_454 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_fill_1 FILLER_52_469 ();
 sg13g2_fill_2 FILLER_52_487 ();
 sg13g2_fill_1 FILLER_52_489 ();
 sg13g2_fill_1 FILLER_52_498 ();
 sg13g2_fill_1 FILLER_52_503 ();
 sg13g2_fill_2 FILLER_52_520 ();
 sg13g2_fill_1 FILLER_52_522 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_21 ();
 sg13g2_fill_1 FILLER_53_87 ();
 sg13g2_fill_2 FILLER_53_118 ();
 sg13g2_fill_2 FILLER_53_130 ();
 sg13g2_fill_1 FILLER_53_132 ();
 sg13g2_fill_1 FILLER_53_199 ();
 sg13g2_fill_2 FILLER_53_235 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_1 FILLER_53_362 ();
 sg13g2_decap_8 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_53_409 ();
 sg13g2_decap_8 FILLER_53_416 ();
 sg13g2_fill_2 FILLER_53_423 ();
 sg13g2_decap_8 FILLER_53_429 ();
 sg13g2_decap_4 FILLER_53_436 ();
 sg13g2_fill_2 FILLER_53_440 ();
 sg13g2_decap_8 FILLER_53_450 ();
 sg13g2_decap_8 FILLER_53_457 ();
 sg13g2_decap_8 FILLER_53_464 ();
 sg13g2_decap_4 FILLER_53_471 ();
 sg13g2_fill_1 FILLER_53_475 ();
 sg13g2_fill_2 FILLER_53_484 ();
 sg13g2_fill_1 FILLER_53_490 ();
 sg13g2_fill_2 FILLER_53_499 ();
 sg13g2_fill_2 FILLER_53_509 ();
 sg13g2_fill_1 FILLER_53_511 ();
 sg13g2_fill_2 FILLER_53_516 ();
 sg13g2_fill_1 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_fill_2 FILLER_54_28 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_109 ();
 sg13g2_fill_2 FILLER_54_125 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_1 FILLER_54_146 ();
 sg13g2_fill_2 FILLER_54_240 ();
 sg13g2_fill_2 FILLER_54_284 ();
 sg13g2_fill_1 FILLER_54_356 ();
 sg13g2_decap_8 FILLER_54_395 ();
 sg13g2_decap_8 FILLER_54_402 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_decap_4 FILLER_54_434 ();
 sg13g2_decap_8 FILLER_54_446 ();
 sg13g2_decap_8 FILLER_54_453 ();
 sg13g2_decap_8 FILLER_54_460 ();
 sg13g2_decap_8 FILLER_54_467 ();
 sg13g2_decap_4 FILLER_54_474 ();
 sg13g2_fill_2 FILLER_54_478 ();
 sg13g2_fill_2 FILLER_54_496 ();
 sg13g2_fill_1 FILLER_54_498 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_4 FILLER_55_28 ();
 sg13g2_fill_2 FILLER_55_32 ();
 sg13g2_fill_2 FILLER_55_55 ();
 sg13g2_fill_1 FILLER_55_57 ();
 sg13g2_fill_2 FILLER_55_80 ();
 sg13g2_fill_1 FILLER_55_102 ();
 sg13g2_fill_1 FILLER_55_108 ();
 sg13g2_fill_1 FILLER_55_195 ();
 sg13g2_fill_2 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_263 ();
 sg13g2_fill_2 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_381 ();
 sg13g2_decap_8 FILLER_55_388 ();
 sg13g2_decap_8 FILLER_55_395 ();
 sg13g2_fill_2 FILLER_55_402 ();
 sg13g2_decap_8 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_55_415 ();
 sg13g2_decap_8 FILLER_55_422 ();
 sg13g2_fill_2 FILLER_55_429 ();
 sg13g2_decap_4 FILLER_55_439 ();
 sg13g2_decap_8 FILLER_55_451 ();
 sg13g2_decap_8 FILLER_55_458 ();
 sg13g2_decap_8 FILLER_55_465 ();
 sg13g2_decap_8 FILLER_55_472 ();
 sg13g2_fill_2 FILLER_55_479 ();
 sg13g2_fill_1 FILLER_55_481 ();
 sg13g2_fill_1 FILLER_55_498 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_90 ();
 sg13g2_fill_2 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_101 ();
 sg13g2_fill_2 FILLER_56_127 ();
 sg13g2_fill_1 FILLER_56_129 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_198 ();
 sg13g2_fill_2 FILLER_56_226 ();
 sg13g2_fill_1 FILLER_56_293 ();
 sg13g2_fill_1 FILLER_56_346 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_decap_8 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_388 ();
 sg13g2_decap_8 FILLER_56_395 ();
 sg13g2_decap_8 FILLER_56_402 ();
 sg13g2_decap_4 FILLER_56_409 ();
 sg13g2_fill_2 FILLER_56_413 ();
 sg13g2_fill_2 FILLER_56_419 ();
 sg13g2_fill_1 FILLER_56_421 ();
 sg13g2_fill_1 FILLER_56_426 ();
 sg13g2_decap_8 FILLER_56_435 ();
 sg13g2_decap_8 FILLER_56_442 ();
 sg13g2_decap_8 FILLER_56_449 ();
 sg13g2_decap_8 FILLER_56_456 ();
 sg13g2_decap_8 FILLER_56_463 ();
 sg13g2_decap_8 FILLER_56_470 ();
 sg13g2_fill_1 FILLER_56_477 ();
 sg13g2_fill_1 FILLER_56_506 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_4 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_18 ();
 sg13g2_fill_1 FILLER_57_23 ();
 sg13g2_fill_2 FILLER_57_44 ();
 sg13g2_fill_2 FILLER_57_75 ();
 sg13g2_fill_2 FILLER_57_108 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_188 ();
 sg13g2_fill_2 FILLER_57_193 ();
 sg13g2_fill_2 FILLER_57_246 ();
 sg13g2_decap_4 FILLER_57_314 ();
 sg13g2_fill_1 FILLER_57_343 ();
 sg13g2_decap_8 FILLER_57_366 ();
 sg13g2_decap_8 FILLER_57_373 ();
 sg13g2_decap_8 FILLER_57_380 ();
 sg13g2_decap_8 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_decap_8 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_57_415 ();
 sg13g2_decap_8 FILLER_57_422 ();
 sg13g2_decap_8 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_57_436 ();
 sg13g2_decap_8 FILLER_57_443 ();
 sg13g2_decap_8 FILLER_57_450 ();
 sg13g2_decap_8 FILLER_57_457 ();
 sg13g2_decap_8 FILLER_57_464 ();
 sg13g2_fill_2 FILLER_57_471 ();
 sg13g2_fill_1 FILLER_57_501 ();
 sg13g2_fill_1 FILLER_57_510 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_132 ();
 sg13g2_fill_1 FILLER_58_212 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_fill_1 FILLER_58_324 ();
 sg13g2_decap_8 FILLER_58_367 ();
 sg13g2_decap_8 FILLER_58_374 ();
 sg13g2_decap_8 FILLER_58_381 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_4 FILLER_58_395 ();
 sg13g2_fill_2 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_405 ();
 sg13g2_fill_2 FILLER_58_412 ();
 sg13g2_decap_8 FILLER_58_418 ();
 sg13g2_fill_1 FILLER_58_425 ();
 sg13g2_decap_8 FILLER_58_438 ();
 sg13g2_decap_4 FILLER_58_445 ();
 sg13g2_decap_8 FILLER_58_453 ();
 sg13g2_fill_1 FILLER_58_460 ();
 sg13g2_fill_2 FILLER_58_489 ();
 sg13g2_fill_1 FILLER_58_491 ();
 sg13g2_fill_1 FILLER_58_496 ();
 sg13g2_fill_2 FILLER_58_513 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_2 ();
 sg13g2_fill_2 FILLER_59_100 ();
 sg13g2_fill_1 FILLER_59_102 ();
 sg13g2_fill_2 FILLER_59_129 ();
 sg13g2_fill_2 FILLER_59_156 ();
 sg13g2_fill_1 FILLER_59_175 ();
 sg13g2_fill_2 FILLER_59_206 ();
 sg13g2_fill_1 FILLER_59_208 ();
 sg13g2_fill_2 FILLER_59_239 ();
 sg13g2_fill_1 FILLER_59_253 ();
 sg13g2_fill_2 FILLER_59_275 ();
 sg13g2_fill_1 FILLER_59_289 ();
 sg13g2_fill_2 FILLER_59_338 ();
 sg13g2_fill_2 FILLER_59_353 ();
 sg13g2_fill_1 FILLER_59_355 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_fill_2 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_decap_4 FILLER_59_427 ();
 sg13g2_fill_2 FILLER_59_431 ();
 sg13g2_fill_1 FILLER_59_505 ();
 sg13g2_fill_2 FILLER_59_510 ();
 sg13g2_fill_1 FILLER_59_512 ();
 sg13g2_fill_2 FILLER_59_517 ();
endmodule
