magic
tech sky130A
magscale 1 2
timestamp 1740383996
<< viali >>
rect 2513 8585 2547 8619
rect 2973 8585 3007 8619
rect 4629 8585 4663 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6469 8585 6503 8619
rect 7021 8585 7055 8619
rect 9045 8585 9079 8619
rect 9597 8585 9631 8619
rect 10701 8585 10735 8619
rect 11897 8585 11931 8619
rect 12633 8585 12667 8619
rect 14197 8585 14231 8619
rect 15117 8585 15151 8619
rect 15669 8585 15703 8619
rect 16221 8585 16255 8619
rect 16865 8585 16899 8619
rect 17049 8585 17083 8619
rect 18521 8585 18555 8619
rect 19625 8585 19659 8619
rect 21925 8585 21959 8619
rect 22385 8585 22419 8619
rect 23673 8585 23707 8619
rect 24041 8585 24075 8619
rect 24501 8585 24535 8619
rect 26157 8585 26191 8619
rect 30021 8585 30055 8619
rect 30573 8585 30607 8619
rect 32229 8585 32263 8619
rect 32781 8585 32815 8619
rect 33885 8585 33919 8619
rect 34989 8585 35023 8619
rect 36093 8585 36127 8619
rect 36645 8585 36679 8619
rect 37013 8585 37047 8619
rect 37381 8585 37415 8619
rect 38393 8585 38427 8619
rect 39405 8585 39439 8619
rect 3341 8517 3375 8551
rect 3893 8517 3927 8551
rect 4261 8517 4295 8551
rect 4445 8517 4479 8551
rect 5549 8517 5583 8551
rect 8401 8517 8435 8551
rect 8585 8517 8619 8551
rect 11253 8517 11287 8551
rect 1409 8449 1443 8483
rect 2329 8449 2363 8483
rect 3157 8449 3191 8483
rect 4813 8449 4847 8483
rect 5089 8449 5123 8483
rect 6653 8449 6687 8483
rect 6837 8449 6871 8483
rect 7481 8449 7515 8483
rect 9229 8449 9263 8483
rect 9781 8449 9815 8483
rect 10885 8449 10919 8483
rect 11069 8449 11103 8483
rect 11713 8449 11747 8483
rect 12817 8449 12851 8483
rect 13185 8449 13219 8483
rect 14381 8449 14415 8483
rect 15301 8449 15335 8483
rect 15485 8449 15519 8483
rect 16405 8449 16439 8483
rect 16681 8449 16715 8483
rect 17233 8449 17267 8483
rect 17601 8449 17635 8483
rect 18705 8449 18739 8483
rect 19441 8449 19475 8483
rect 20269 8449 20303 8483
rect 20545 8449 20579 8483
rect 21373 8449 21407 8483
rect 22109 8449 22143 8483
rect 22201 8449 22235 8483
rect 22753 8449 22787 8483
rect 23857 8449 23891 8483
rect 24225 8449 24259 8483
rect 24685 8449 24719 8483
rect 25053 8449 25087 8483
rect 26341 8449 26375 8483
rect 27445 8449 27479 8483
rect 28549 8449 28583 8483
rect 29837 8449 29871 8483
rect 30205 8449 30239 8483
rect 30757 8449 30791 8483
rect 31217 8449 31251 8483
rect 32413 8449 32447 8483
rect 32965 8449 32999 8483
rect 34069 8449 34103 8483
rect 35173 8449 35207 8483
rect 36277 8449 36311 8483
rect 36737 8449 36771 8483
rect 36829 8449 36863 8483
rect 37565 8449 37599 8483
rect 37841 8449 37875 8483
rect 38209 8449 38243 8483
rect 38761 8449 38795 8483
rect 38853 8449 38887 8483
rect 39221 8449 39255 8483
rect 1685 8381 1719 8415
rect 3525 8381 3559 8415
rect 7205 8381 7239 8415
rect 12909 8381 12943 8415
rect 17325 8381 17359 8415
rect 22477 8381 22511 8415
rect 24777 8381 24811 8415
rect 27169 8381 27203 8415
rect 28273 8381 28307 8415
rect 30941 8381 30975 8415
rect 8217 8313 8251 8347
rect 21557 8313 21591 8347
rect 29653 8313 29687 8347
rect 31953 8313 31987 8347
rect 38025 8313 38059 8347
rect 39037 8313 39071 8347
rect 3985 8245 4019 8279
rect 13921 8245 13955 8279
rect 18337 8245 18371 8279
rect 21281 8245 21315 8279
rect 23489 8245 23523 8279
rect 25789 8245 25823 8279
rect 28181 8245 28215 8279
rect 29285 8245 29319 8279
rect 38577 8245 38611 8279
rect 2697 8041 2731 8075
rect 4813 8041 4847 8075
rect 14289 8041 14323 8075
rect 16865 8041 16899 8075
rect 19625 8041 19659 8075
rect 22569 8041 22603 8075
rect 27261 8041 27295 8075
rect 33333 8041 33367 8075
rect 36277 8041 36311 8075
rect 36829 8041 36863 8075
rect 37657 8041 37691 8075
rect 38301 8041 38335 8075
rect 3617 7973 3651 8007
rect 6009 7973 6043 8007
rect 8769 7973 8803 8007
rect 10333 7973 10367 8007
rect 10701 7973 10735 8007
rect 11805 7973 11839 8007
rect 12541 7973 12575 8007
rect 21373 7973 21407 8007
rect 25513 7973 25547 8007
rect 28181 7973 28215 8007
rect 33241 7973 33275 8007
rect 37105 7973 37139 8007
rect 37933 7973 37967 8007
rect 3157 7905 3191 7939
rect 6377 7905 6411 7939
rect 7297 7905 7331 7939
rect 9965 7905 9999 7939
rect 12081 7905 12115 7939
rect 12817 7905 12851 7939
rect 15209 7905 15243 7939
rect 15669 7905 15703 7939
rect 15945 7905 15979 7939
rect 20913 7905 20947 7939
rect 21766 7905 21800 7939
rect 25053 7905 25087 7939
rect 25906 7905 25940 7939
rect 27537 7905 27571 7939
rect 31309 7905 31343 7939
rect 31769 7905 31803 7939
rect 32162 7905 32196 7939
rect 32321 7905 32355 7939
rect 38669 7905 38703 7939
rect 1869 7837 1903 7871
rect 2237 7837 2271 7871
rect 2605 7837 2639 7871
rect 2973 7837 3007 7871
rect 3801 7837 3835 7871
rect 4077 7837 4111 7871
rect 4997 7837 5031 7871
rect 5273 7837 5307 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 9689 7837 9723 7871
rect 10793 7837 10827 7871
rect 11069 7837 11103 7871
rect 11897 7837 11931 7871
rect 12955 7837 12989 7871
rect 13093 7837 13127 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 15025 7837 15059 7871
rect 16083 7837 16117 7871
rect 16221 7837 16255 7871
rect 17049 7837 17083 7871
rect 17325 7837 17359 7871
rect 17601 7837 17635 7871
rect 19441 7837 19475 7871
rect 20729 7837 20763 7871
rect 21649 7837 21683 7871
rect 21925 7837 21959 7871
rect 23397 7837 23431 7871
rect 23673 7837 23707 7871
rect 24041 7837 24075 7871
rect 24593 7837 24627 7871
rect 24869 7837 24903 7871
rect 25789 7837 25823 7871
rect 26065 7837 26099 7871
rect 26709 7837 26743 7871
rect 26801 7837 26835 7871
rect 27445 7837 27479 7871
rect 27721 7837 27755 7871
rect 28457 7837 28491 7871
rect 28574 7837 28608 7871
rect 28733 7837 28767 7871
rect 29377 7837 29411 7871
rect 29561 7837 29595 7871
rect 29929 7837 29963 7871
rect 31125 7837 31159 7871
rect 32045 7837 32079 7871
rect 32965 7837 32999 7871
rect 33057 7837 33091 7871
rect 33517 7837 33551 7871
rect 35449 7837 35483 7871
rect 35725 7837 35759 7871
rect 36461 7837 36495 7871
rect 37013 7837 37047 7871
rect 37289 7837 37323 7871
rect 37473 7837 37507 7871
rect 37749 7837 37783 7871
rect 38117 7837 38151 7871
rect 38761 7837 38795 7871
rect 38853 7837 38887 7871
rect 39221 7837 39255 7871
rect 1501 7769 1535 7803
rect 2053 7769 2087 7803
rect 2421 7769 2455 7803
rect 3433 7769 3467 7803
rect 6193 7769 6227 7803
rect 8585 7769 8619 7803
rect 10149 7769 10183 7803
rect 10517 7769 10551 7803
rect 17233 7769 17267 7803
rect 38577 7769 38611 7803
rect 1593 7701 1627 7735
rect 2697 7701 2731 7735
rect 7205 7701 7239 7735
rect 8309 7701 8343 7735
rect 8953 7701 8987 7735
rect 14565 7701 14599 7735
rect 18337 7701 18371 7735
rect 22661 7701 22695 7735
rect 24225 7701 24259 7735
rect 24777 7701 24811 7735
rect 26985 7701 27019 7735
rect 29745 7701 29779 7735
rect 30113 7701 30147 7735
rect 34713 7701 34747 7735
rect 38485 7701 38519 7735
rect 39037 7701 39071 7735
rect 39405 7701 39439 7735
rect 2513 7497 2547 7531
rect 9965 7497 9999 7531
rect 12541 7497 12575 7531
rect 15761 7497 15795 7531
rect 19809 7497 19843 7531
rect 21281 7497 21315 7531
rect 23397 7497 23431 7531
rect 26341 7497 26375 7531
rect 28181 7497 28215 7531
rect 30113 7497 30147 7531
rect 33977 7497 34011 7531
rect 37657 7497 37691 7531
rect 38669 7497 38703 7531
rect 5825 7429 5859 7463
rect 1685 7361 1719 7395
rect 2329 7361 2363 7395
rect 2605 7361 2639 7395
rect 2881 7361 2915 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 4997 7361 5031 7395
rect 5641 7361 5675 7395
rect 7205 7361 7239 7395
rect 8493 7361 8527 7395
rect 8769 7361 8803 7395
rect 9413 7361 9447 7395
rect 9505 7361 9539 7395
rect 9873 7361 9907 7395
rect 10609 7361 10643 7395
rect 11529 7361 11563 7395
rect 11805 7361 11839 7395
rect 13093 7361 13127 7395
rect 14841 7361 14875 7395
rect 15117 7361 15151 7395
rect 15853 7361 15887 7395
rect 17141 7361 17175 7395
rect 17969 7361 18003 7395
rect 18153 7361 18187 7395
rect 18889 7361 18923 7395
rect 19165 7361 19199 7395
rect 20545 7361 20579 7395
rect 22569 7361 22603 7395
rect 25053 7361 25087 7395
rect 25605 7361 25639 7395
rect 27169 7361 27203 7395
rect 27445 7361 27479 7395
rect 28273 7361 28307 7395
rect 28457 7361 28491 7395
rect 29469 7361 29503 7395
rect 30665 7361 30699 7395
rect 31217 7361 31251 7395
rect 32137 7361 32171 7395
rect 33057 7361 33091 7395
rect 34897 7361 34931 7395
rect 35173 7361 35207 7395
rect 35449 7361 35483 7395
rect 37841 7361 37875 7395
rect 38117 7361 38151 7395
rect 38485 7361 38519 7395
rect 39037 7361 39071 7395
rect 39221 7361 39255 7395
rect 1409 7293 1443 7327
rect 7481 7293 7515 7327
rect 7573 7293 7607 7327
rect 7757 7293 7791 7327
rect 8217 7293 8251 7327
rect 8631 7293 8665 7327
rect 10333 7293 10367 7327
rect 12817 7293 12851 7327
rect 13921 7293 13955 7327
rect 14105 7293 14139 7327
rect 14565 7293 14599 7327
rect 14958 7293 14992 7327
rect 16865 7293 16899 7327
rect 18613 7293 18647 7327
rect 19027 7293 19061 7327
rect 20269 7293 20303 7327
rect 22293 7293 22327 7327
rect 24041 7293 24075 7327
rect 24179 7293 24213 7327
rect 24317 7293 24351 7327
rect 25237 7293 25271 7327
rect 25325 7293 25359 7327
rect 29193 7293 29227 7327
rect 29310 7293 29344 7327
rect 30941 7293 30975 7327
rect 32321 7293 32355 7327
rect 33174 7293 33208 7327
rect 33333 7293 33367 7327
rect 4813 7225 4847 7259
rect 23305 7225 23339 7259
rect 24593 7225 24627 7259
rect 28917 7225 28951 7259
rect 31953 7225 31987 7259
rect 32781 7225 32815 7259
rect 35265 7225 35299 7259
rect 3617 7157 3651 7191
rect 4721 7157 4755 7191
rect 6469 7157 6503 7191
rect 9689 7157 9723 7191
rect 11345 7157 11379 7191
rect 13829 7157 13863 7191
rect 16037 7157 16071 7191
rect 17877 7157 17911 7191
rect 30849 7157 30883 7191
rect 34161 7157 34195 7191
rect 38301 7157 38335 7191
rect 39405 7157 39439 7191
rect 3617 6953 3651 6987
rect 13093 6953 13127 6987
rect 13829 6953 13863 6987
rect 15393 6953 15427 6987
rect 20085 6953 20119 6987
rect 28457 6953 28491 6987
rect 31401 6953 31435 6987
rect 38209 6953 38243 6987
rect 4445 6885 4479 6919
rect 15485 6885 15519 6919
rect 25237 6885 25271 6919
rect 1777 6817 1811 6851
rect 3157 6817 3191 6851
rect 4997 6817 5031 6851
rect 5733 6817 5767 6851
rect 6377 6817 6411 6851
rect 6536 6817 6570 6851
rect 6653 6817 6687 6851
rect 6929 6817 6963 6851
rect 7573 6817 7607 6851
rect 7757 6817 7791 6851
rect 9229 6817 9263 6851
rect 14381 6817 14415 6851
rect 17141 6817 17175 6851
rect 17233 6817 17267 6851
rect 21097 6817 21131 6851
rect 27445 6817 27479 6851
rect 29561 6817 29595 6851
rect 30205 6817 30239 6851
rect 30481 6817 30515 6851
rect 30598 6817 30632 6851
rect 1501 6749 1535 6783
rect 2053 6749 2087 6783
rect 3433 6749 3467 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 4721 6749 4755 6783
rect 4859 6749 4893 6783
rect 7389 6749 7423 6783
rect 8033 6749 8067 6783
rect 8953 6751 8987 6785
rect 9505 6749 9539 6783
rect 10517 6749 10551 6783
rect 10885 6749 10919 6783
rect 10977 6749 11011 6783
rect 11253 6749 11287 6783
rect 12265 6749 12299 6783
rect 12357 6749 12391 6783
rect 12633 6749 12667 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 13645 6749 13679 6783
rect 14105 6749 14139 6783
rect 14657 6749 14691 6783
rect 16221 6749 16255 6783
rect 16497 6749 16531 6783
rect 16957 6749 16991 6783
rect 17509 6749 17543 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 20269 6749 20303 6783
rect 20453 6749 20487 6783
rect 20637 6749 20671 6783
rect 21373 6749 21407 6783
rect 21490 6749 21524 6783
rect 21649 6749 21683 6783
rect 22293 6749 22327 6783
rect 22385 6749 22419 6783
rect 23489 6749 23523 6783
rect 23765 6749 23799 6783
rect 24869 6749 24903 6783
rect 25973 6749 26007 6783
rect 26249 6749 26283 6783
rect 26341 6749 26375 6783
rect 26617 6749 26651 6783
rect 27721 6749 27755 6783
rect 29745 6749 29779 6783
rect 30757 6749 30791 6783
rect 31953 6749 31987 6783
rect 32229 6749 32263 6783
rect 33057 6749 33091 6783
rect 33333 6749 33367 6783
rect 34437 6749 34471 6783
rect 34713 6749 34747 6783
rect 34989 6749 35023 6783
rect 36001 6749 36035 6783
rect 37933 6749 37967 6783
rect 38393 6765 38427 6799
rect 38669 6749 38703 6783
rect 38853 6749 38887 6783
rect 39221 6749 39255 6783
rect 1685 6681 1719 6715
rect 2973 6681 3007 6715
rect 9045 6681 9079 6715
rect 10609 6681 10643 6715
rect 10701 6681 10735 6715
rect 2789 6613 2823 6647
rect 5641 6613 5675 6647
rect 8769 6613 8803 6647
rect 10241 6613 10275 6647
rect 10333 6613 10367 6647
rect 11989 6613 12023 6647
rect 12173 6613 12207 6647
rect 12541 6613 12575 6647
rect 12817 6613 12851 6647
rect 13553 6613 13587 6647
rect 14289 6613 14323 6647
rect 18245 6613 18279 6647
rect 19257 6613 19291 6647
rect 19809 6613 19843 6647
rect 22569 6613 22603 6647
rect 22753 6613 22787 6647
rect 25053 6613 25087 6647
rect 27353 6613 27387 6647
rect 32965 6613 32999 6647
rect 34069 6613 34103 6647
rect 34253 6613 34287 6647
rect 35725 6613 35759 6647
rect 35817 6613 35851 6647
rect 38117 6613 38151 6647
rect 38485 6613 38519 6647
rect 39037 6613 39071 6647
rect 39405 6613 39439 6647
rect 10425 6409 10459 6443
rect 12357 6409 12391 6443
rect 16865 6409 16899 6443
rect 21097 6409 21131 6443
rect 34345 6409 34379 6443
rect 35541 6409 35575 6443
rect 36001 6409 36035 6443
rect 38301 6409 38335 6443
rect 39405 6409 39439 6443
rect 10885 6341 10919 6375
rect 1409 6273 1443 6307
rect 1685 6273 1719 6307
rect 2329 6273 2363 6307
rect 2881 6273 2915 6307
rect 4629 6273 4663 6307
rect 4767 6273 4801 6307
rect 5641 6273 5675 6307
rect 5917 6273 5951 6307
rect 6745 6273 6779 6307
rect 6837 6273 6871 6307
rect 7113 6273 7147 6307
rect 7665 6273 7699 6307
rect 8677 6273 8711 6307
rect 9551 6273 9585 6307
rect 10793 6273 10827 6307
rect 11646 6273 11680 6307
rect 11897 6273 11931 6307
rect 12173 6273 12207 6307
rect 12725 6273 12759 6307
rect 13829 6273 13863 6307
rect 14841 6273 14875 6307
rect 15577 6273 15611 6307
rect 16497 6273 16531 6307
rect 16681 6273 16715 6307
rect 16957 6273 16991 6307
rect 17233 6273 17267 6307
rect 18337 6273 18371 6307
rect 19349 6273 19383 6307
rect 20361 6273 20395 6307
rect 22201 6273 22235 6307
rect 23305 6273 23339 6307
rect 24869 6273 24903 6307
rect 25145 6273 25179 6307
rect 25973 6273 26007 6307
rect 26617 6273 26651 6307
rect 27721 6273 27755 6307
rect 27997 6273 28031 6307
rect 28089 6273 28123 6307
rect 28365 6273 28399 6307
rect 30251 6273 30285 6307
rect 30389 6273 30423 6307
rect 31033 6273 31067 6307
rect 31309 6273 31343 6307
rect 31769 6273 31803 6307
rect 32321 6273 32355 6307
rect 32505 6273 32539 6307
rect 33425 6273 33459 6307
rect 35173 6273 35207 6307
rect 35909 6273 35943 6307
rect 38485 6273 38519 6307
rect 38761 6273 38795 6307
rect 38853 6273 38887 6307
rect 39221 6273 39255 6307
rect 2605 6205 2639 6239
rect 3709 6205 3743 6239
rect 3893 6205 3927 6239
rect 4905 6205 4939 6239
rect 5549 6205 5583 6239
rect 7389 6205 7423 6239
rect 8493 6205 8527 6239
rect 9137 6205 9171 6239
rect 9413 6205 9447 6239
rect 9689 6205 9723 6239
rect 10977 6205 11011 6239
rect 12449 6205 12483 6239
rect 13553 6205 13587 6239
rect 14657 6205 14691 6239
rect 15694 6205 15728 6239
rect 15853 6205 15887 6239
rect 18153 6205 18187 6239
rect 18797 6205 18831 6239
rect 19073 6205 19107 6239
rect 19190 6205 19224 6239
rect 20085 6205 20119 6239
rect 21925 6205 21959 6239
rect 23029 6205 23063 6239
rect 26249 6205 26283 6239
rect 29193 6205 29227 6239
rect 29377 6205 29411 6239
rect 30113 6205 30147 6239
rect 32689 6205 32723 6239
rect 33149 6205 33183 6239
rect 33542 6205 33576 6239
rect 33701 6205 33735 6239
rect 35449 6205 35483 6239
rect 36093 6205 36127 6239
rect 2513 6137 2547 6171
rect 3617 6137 3651 6171
rect 4353 6137 4387 6171
rect 5825 6137 5859 6171
rect 7021 6137 7055 6171
rect 12081 6137 12115 6171
rect 15301 6137 15335 6171
rect 19993 6137 20027 6171
rect 24133 6137 24167 6171
rect 25237 6137 25271 6171
rect 29101 6137 29135 6171
rect 29837 6137 29871 6171
rect 38577 6137 38611 6171
rect 6101 6069 6135 6103
rect 6561 6069 6595 6103
rect 7297 6069 7331 6103
rect 8401 6069 8435 6103
rect 10333 6069 10367 6103
rect 11575 6069 11609 6103
rect 13461 6069 13495 6103
rect 14565 6069 14599 6103
rect 17969 6069 18003 6103
rect 22937 6069 22971 6103
rect 24041 6069 24075 6103
rect 26801 6069 26835 6103
rect 26985 6069 27019 6103
rect 31125 6069 31159 6103
rect 31953 6069 31987 6103
rect 34437 6069 34471 6103
rect 39037 6069 39071 6103
rect 3433 5865 3467 5899
rect 4813 5865 4847 5899
rect 5181 5865 5215 5899
rect 6377 5865 6411 5899
rect 8769 5865 8803 5899
rect 11437 5865 11471 5899
rect 15945 5865 15979 5899
rect 19073 5865 19107 5899
rect 21097 5865 21131 5899
rect 28917 5865 28951 5899
rect 30573 5865 30607 5899
rect 38393 5865 38427 5899
rect 39405 5865 39439 5899
rect 1685 5797 1719 5831
rect 2053 5797 2087 5831
rect 2789 5797 2823 5831
rect 3157 5797 3191 5831
rect 6285 5797 6319 5831
rect 9505 5797 9539 5831
rect 12173 5797 12207 5831
rect 13645 5797 13679 5831
rect 13737 5797 13771 5831
rect 17141 5797 17175 5831
rect 17877 5797 17911 5831
rect 21189 5797 21223 5831
rect 23029 5797 23063 5831
rect 26617 5797 26651 5831
rect 27813 5797 27847 5831
rect 31677 5797 31711 5831
rect 32321 5797 32355 5831
rect 36737 5797 36771 5831
rect 39037 5797 39071 5831
rect 3801 5729 3835 5763
rect 7021 5729 7055 5763
rect 7180 5729 7214 5763
rect 7573 5729 7607 5763
rect 8033 5729 8067 5763
rect 9045 5729 9079 5763
rect 9137 5729 9171 5763
rect 10241 5729 10275 5763
rect 10517 5729 10551 5763
rect 10655 5729 10689 5763
rect 12725 5729 12759 5763
rect 14289 5729 14323 5763
rect 14749 5729 14783 5763
rect 15025 5729 15059 5763
rect 15163 5729 15197 5763
rect 18429 5729 18463 5763
rect 20085 5729 20119 5763
rect 22569 5729 22603 5763
rect 23305 5729 23339 5763
rect 23579 5729 23613 5763
rect 25881 5729 25915 5763
rect 25973 5729 26007 5763
rect 26157 5729 26191 5763
rect 26893 5729 26927 5763
rect 27031 5729 27065 5763
rect 27169 5729 27203 5763
rect 27905 5729 27939 5763
rect 29285 5729 29319 5763
rect 29561 5729 29595 5763
rect 1869 5661 1903 5695
rect 2605 5661 2639 5695
rect 4077 5661 4111 5695
rect 4997 5661 5031 5695
rect 5273 5661 5307 5695
rect 5549 5661 5583 5695
rect 7297 5661 7331 5695
rect 8217 5661 8251 5695
rect 8309 5661 8343 5695
rect 8585 5661 8619 5695
rect 9321 5661 9355 5695
rect 9597 5661 9631 5695
rect 9781 5661 9815 5695
rect 10793 5661 10827 5695
rect 11529 5661 11563 5695
rect 11713 5661 11747 5695
rect 12449 5661 12483 5695
rect 12566 5661 12600 5695
rect 13461 5661 13495 5695
rect 13921 5661 13955 5695
rect 14105 5661 14139 5695
rect 15301 5661 15335 5695
rect 16129 5661 16163 5695
rect 16405 5661 16439 5695
rect 17233 5661 17267 5695
rect 17417 5661 17451 5695
rect 18153 5661 18187 5695
rect 18270 5661 18304 5695
rect 19257 5661 19291 5695
rect 19809 5661 19843 5695
rect 20361 5661 20395 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 22385 5661 22419 5695
rect 23443 5661 23477 5695
rect 24225 5661 24259 5695
rect 24409 5661 24443 5695
rect 24961 5661 24995 5695
rect 25605 5661 25639 5695
rect 28181 5661 28215 5695
rect 29837 5661 29871 5695
rect 30665 5661 30699 5695
rect 30941 5661 30975 5695
rect 32137 5661 32171 5695
rect 32597 5661 32631 5695
rect 34713 5661 34747 5695
rect 36553 5661 36587 5695
rect 38577 5661 38611 5695
rect 38853 5661 38887 5695
rect 39221 5661 39255 5695
rect 1501 5593 1535 5627
rect 2237 5593 2271 5627
rect 2421 5593 2455 5627
rect 2973 5593 3007 5627
rect 3341 5593 3375 5627
rect 13369 5593 13403 5627
rect 29101 5593 29135 5627
rect 34529 5593 34563 5627
rect 8493 5525 8527 5559
rect 19441 5525 19475 5559
rect 19993 5525 20027 5559
rect 21649 5525 21683 5559
rect 24593 5525 24627 5559
rect 24777 5525 24811 5559
rect 29193 5525 29227 5559
rect 32413 5525 32447 5559
rect 33241 5525 33275 5559
rect 36001 5525 36035 5559
rect 1961 5321 1995 5355
rect 3433 5321 3467 5355
rect 4353 5321 4387 5355
rect 6193 5321 6227 5355
rect 9229 5321 9263 5355
rect 12265 5321 12299 5355
rect 12541 5321 12575 5355
rect 12633 5321 12667 5355
rect 13093 5321 13127 5355
rect 15117 5321 15151 5355
rect 19717 5321 19751 5355
rect 29929 5321 29963 5355
rect 32321 5321 32355 5355
rect 34621 5321 34655 5355
rect 36185 5321 36219 5355
rect 39405 5321 39439 5355
rect 1501 5253 1535 5287
rect 1685 5253 1719 5287
rect 1869 5253 1903 5287
rect 2237 5253 2271 5287
rect 4169 5253 4203 5287
rect 33824 5253 33858 5287
rect 35909 5253 35943 5287
rect 2697 5185 2731 5219
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 3525 5185 3559 5219
rect 3801 5185 3835 5219
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 4537 5185 4571 5219
rect 4696 5185 4730 5219
rect 4972 5185 5006 5219
rect 5457 5185 5491 5219
rect 6653 5185 6687 5219
rect 6837 5185 6871 5219
rect 7113 5185 7147 5219
rect 7389 5185 7423 5219
rect 8426 5185 8460 5219
rect 8585 5185 8619 5219
rect 10241 5185 10275 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12081 5185 12115 5219
rect 12357 5185 12391 5219
rect 12817 5185 12851 5219
rect 12909 5185 12943 5219
rect 13185 5185 13219 5219
rect 13737 5185 13771 5219
rect 14565 5185 14599 5219
rect 14841 5185 14875 5219
rect 15853 5185 15887 5219
rect 16313 5185 16347 5219
rect 16773 5185 16807 5219
rect 17049 5185 17083 5219
rect 17877 5185 17911 5219
rect 18797 5185 18831 5219
rect 18914 5185 18948 5219
rect 19809 5185 19843 5219
rect 19993 5185 20027 5219
rect 20729 5185 20763 5219
rect 21649 5185 21683 5219
rect 22017 5185 22051 5219
rect 22477 5185 22511 5219
rect 23029 5185 23063 5219
rect 24593 5185 24627 5219
rect 25329 5185 25363 5219
rect 26157 5185 26191 5219
rect 26801 5185 26835 5219
rect 27353 5185 27387 5219
rect 27537 5185 27571 5219
rect 27813 5185 27847 5219
rect 28089 5215 28123 5249
rect 29193 5185 29227 5219
rect 30573 5185 30607 5219
rect 31033 5185 31067 5219
rect 31125 5185 31159 5219
rect 31493 5185 31527 5219
rect 32137 5185 32171 5219
rect 32413 5185 32447 5219
rect 34069 5185 34103 5219
rect 36001 5185 36035 5219
rect 38853 5185 38887 5219
rect 39221 5185 39255 5219
rect 5181 5117 5215 5151
rect 6377 5117 6411 5151
rect 7573 5117 7607 5151
rect 8309 5117 8343 5151
rect 9321 5117 9355 5151
rect 9505 5117 9539 5151
rect 10379 5117 10413 5151
rect 10517 5117 10551 5151
rect 13461 5117 13495 5151
rect 16129 5117 16163 5151
rect 18061 5117 18095 5151
rect 19073 5117 19107 5151
rect 20846 5117 20880 5151
rect 21005 5117 21039 5151
rect 22753 5117 22787 5151
rect 25053 5117 25087 5151
rect 28917 5117 28951 5151
rect 2421 5049 2455 5083
rect 3709 5049 3743 5083
rect 4767 5049 4801 5083
rect 6561 5049 6595 5083
rect 7021 5049 7055 5083
rect 8033 5049 8067 5083
rect 9965 5049 9999 5083
rect 11989 5049 12023 5083
rect 14473 5049 14507 5083
rect 17785 5049 17819 5083
rect 18521 5049 18555 5083
rect 20453 5049 20487 5083
rect 31677 5049 31711 5083
rect 2881 4981 2915 5015
rect 3157 4981 3191 5015
rect 3985 4981 4019 5015
rect 4353 4981 4387 5015
rect 5043 4981 5077 5015
rect 6469 4981 6503 5015
rect 7297 4981 7331 5015
rect 11161 4981 11195 5015
rect 11621 4981 11655 5015
rect 13369 4981 13403 5015
rect 14749 4981 14783 5015
rect 15025 4981 15059 5015
rect 16497 4981 16531 5015
rect 21833 4981 21867 5015
rect 22293 4981 22327 5015
rect 23765 4981 23799 5015
rect 24777 4981 24811 5015
rect 26065 4981 26099 5015
rect 26341 4981 26375 5015
rect 26617 4981 26651 5015
rect 27169 4981 27203 5015
rect 27721 4981 27755 5015
rect 28825 4981 28859 5015
rect 30389 4981 30423 5015
rect 30941 4981 30975 5015
rect 31309 4981 31343 5015
rect 32597 4981 32631 5015
rect 32689 4981 32723 5015
rect 39037 4981 39071 5015
rect 1961 4777 1995 4811
rect 2513 4777 2547 4811
rect 2881 4777 2915 4811
rect 8953 4777 8987 4811
rect 9137 4777 9171 4811
rect 9597 4777 9631 4811
rect 13093 4777 13127 4811
rect 13737 4777 13771 4811
rect 15945 4777 15979 4811
rect 16221 4777 16255 4811
rect 19257 4777 19291 4811
rect 27445 4777 27479 4811
rect 33241 4777 33275 4811
rect 33333 4777 33367 4811
rect 36001 4777 36035 4811
rect 36829 4777 36863 4811
rect 39405 4777 39439 4811
rect 21649 4709 21683 4743
rect 23765 4709 23799 4743
rect 26249 4709 26283 4743
rect 30021 4709 30055 4743
rect 32045 4709 32079 4743
rect 4445 4641 4479 4675
rect 4583 4641 4617 4675
rect 4997 4641 5031 4675
rect 5457 4641 5491 4675
rect 7113 4641 7147 4675
rect 7573 4641 7607 4675
rect 7966 4641 8000 4675
rect 10793 4641 10827 4675
rect 12081 4641 12115 4675
rect 14749 4641 14783 4675
rect 15025 4641 15059 4675
rect 15301 4641 15335 4675
rect 17141 4641 17175 4675
rect 17417 4641 17451 4675
rect 18061 4641 18095 4675
rect 21097 4641 21131 4675
rect 22661 4641 22695 4675
rect 25789 4641 25823 4675
rect 26525 4641 26559 4675
rect 27905 4641 27939 4675
rect 31401 4641 31435 4675
rect 31585 4641 31619 4675
rect 32321 4641 32355 4675
rect 32438 4641 32472 4675
rect 34345 4641 34379 4675
rect 1501 4573 1535 4607
rect 1869 4573 1903 4607
rect 2789 4573 2823 4607
rect 3065 4573 3099 4607
rect 3433 4573 3467 4607
rect 3801 4573 3835 4607
rect 4721 4573 4755 4607
rect 5641 4573 5675 4607
rect 5733 4573 5767 4607
rect 6009 4573 6043 4607
rect 6929 4573 6963 4607
rect 7849 4573 7883 4607
rect 8125 4573 8159 4607
rect 9137 4573 9171 4607
rect 9505 4573 9539 4607
rect 9781 4573 9815 4607
rect 9965 4573 9999 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 11069 4573 11103 4607
rect 11207 4573 11241 4607
rect 11345 4573 11379 4607
rect 12357 4573 12391 4607
rect 13921 4573 13955 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 15142 4573 15176 4607
rect 16865 4573 16899 4607
rect 17024 4573 17058 4607
rect 17877 4573 17911 4607
rect 18153 4573 18187 4607
rect 18705 4573 18739 4607
rect 18797 4573 18831 4607
rect 19993 4573 20027 4607
rect 20269 4573 20303 4607
rect 20729 4573 20763 4607
rect 21281 4573 21315 4607
rect 22385 4573 22419 4607
rect 22753 4573 22787 4607
rect 23029 4573 23063 4607
rect 23857 4573 23891 4607
rect 24409 4573 24443 4607
rect 24777 4573 24811 4607
rect 25145 4573 25179 4607
rect 25605 4573 25639 4607
rect 26642 4573 26676 4607
rect 26801 4573 26835 4607
rect 27813 4573 27847 4607
rect 28181 4573 28215 4607
rect 30757 4573 30791 4607
rect 31033 4573 31067 4607
rect 32597 4573 32631 4607
rect 34069 4573 34103 4607
rect 37013 4573 37047 4607
rect 38853 4573 38887 4607
rect 39221 4573 39255 4607
rect 1685 4505 1719 4539
rect 2237 4505 2271 4539
rect 2421 4505 2455 4539
rect 13369 4505 13403 4539
rect 20913 4505 20947 4539
rect 29193 4505 29227 4539
rect 34713 4505 34747 4539
rect 2513 4437 2547 4471
rect 3249 4437 3283 4471
rect 3617 4437 3651 4471
rect 6745 4437 6779 4471
rect 8769 4437 8803 4471
rect 11989 4437 12023 4471
rect 13461 4437 13495 4471
rect 18337 4437 18371 4471
rect 18521 4437 18555 4471
rect 18981 4437 19015 4471
rect 20545 4437 20579 4471
rect 21465 4437 21499 4471
rect 24041 4437 24075 4471
rect 24593 4437 24627 4471
rect 24961 4437 24995 4471
rect 25329 4437 25363 4471
rect 27629 4437 27663 4471
rect 28917 4437 28951 4471
rect 29101 4437 29135 4471
rect 39037 4437 39071 4471
rect 1961 4233 1995 4267
rect 3525 4233 3559 4267
rect 7297 4233 7331 4267
rect 11805 4233 11839 4267
rect 14473 4233 14507 4267
rect 22201 4233 22235 4267
rect 22569 4233 22603 4267
rect 30297 4233 30331 4267
rect 1501 4165 1535 4199
rect 1869 4165 1903 4199
rect 6009 4165 6043 4199
rect 9137 4165 9171 4199
rect 13093 4165 13127 4199
rect 20545 4165 20579 4199
rect 21649 4165 21683 4199
rect 36093 4165 36127 4199
rect 1685 4097 1719 4131
rect 2145 4097 2179 4131
rect 2697 4097 2731 4131
rect 4328 4097 4362 4131
rect 5365 4097 5399 4131
rect 5641 4097 5675 4131
rect 6469 4097 6503 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 8217 4097 8251 4131
rect 10333 4097 10367 4131
rect 10471 4097 10505 4131
rect 11253 4097 11287 4131
rect 11897 4097 11931 4131
rect 12357 4097 12391 4131
rect 12633 4097 12667 4131
rect 12909 4097 12943 4131
rect 13737 4097 13771 4131
rect 15018 4097 15052 4131
rect 15209 4097 15243 4131
rect 15761 4097 15795 4131
rect 17141 4097 17175 4131
rect 17509 4097 17543 4131
rect 17877 4097 17911 4131
rect 18889 4097 18923 4131
rect 19625 4097 19659 4131
rect 21465 4097 21499 4131
rect 21833 4097 21867 4131
rect 23029 4097 23063 4131
rect 24225 4097 24259 4131
rect 24869 4097 24903 4131
rect 25053 4097 25087 4131
rect 25329 4097 25363 4131
rect 26157 4097 26191 4131
rect 26525 4097 26559 4131
rect 27261 4097 27295 4131
rect 28273 4097 28307 4131
rect 29561 4097 29595 4131
rect 30205 4097 30239 4131
rect 31033 4097 31067 4131
rect 31309 4097 31343 4131
rect 31401 4097 31435 4131
rect 32137 4097 32171 4131
rect 32505 4097 32539 4131
rect 34078 4097 34112 4131
rect 34621 4097 34655 4131
rect 34989 4097 35023 4131
rect 36185 4097 36219 4131
rect 36829 4097 36863 4131
rect 38853 4097 38887 4131
rect 39221 4097 39255 4131
rect 2421 4029 2455 4063
rect 4169 4029 4203 4063
rect 4445 4029 4479 4063
rect 5181 4029 5215 4063
rect 7389 4029 7423 4063
rect 7481 4029 7515 4063
rect 7941 4029 7975 4063
rect 9413 4029 9447 4063
rect 9597 4029 9631 4063
rect 10057 4029 10091 4063
rect 10609 4029 10643 4063
rect 11713 4029 11747 4063
rect 13461 4029 13495 4063
rect 15393 4029 15427 4063
rect 15485 4029 15519 4063
rect 17601 4029 17635 4063
rect 18705 4029 18739 4063
rect 19742 4029 19776 4063
rect 19901 4029 19935 4063
rect 21189 4029 21223 4063
rect 22661 4029 22695 4063
rect 22845 4029 22879 4063
rect 23213 4029 23247 4063
rect 23673 4029 23707 4063
rect 23949 4029 23983 4063
rect 24066 4029 24100 4063
rect 26985 4029 27019 4063
rect 28365 4029 28399 4063
rect 28549 4029 28583 4063
rect 29009 4029 29043 4063
rect 29285 4029 29319 4063
rect 29423 4029 29457 4063
rect 34345 4029 34379 4063
rect 34713 4029 34747 4063
rect 35909 4029 35943 4063
rect 4721 3961 4755 3995
rect 6193 3961 6227 3995
rect 6561 3961 6595 3995
rect 6929 3961 6963 3995
rect 9321 3961 9355 3995
rect 12449 3961 12483 3995
rect 16957 3961 16991 3995
rect 18613 3961 18647 3995
rect 19349 3961 19383 3995
rect 26065 3961 26099 3995
rect 27997 3961 28031 3995
rect 32965 3961 32999 3995
rect 35725 3961 35759 3995
rect 36553 3961 36587 3995
rect 39405 3961 39439 3995
rect 2329 3893 2363 3927
rect 3433 3893 3467 3927
rect 6009 3893 6043 3927
rect 6469 3893 6503 3927
rect 8953 3893 8987 3927
rect 12265 3893 12299 3927
rect 12817 3893 12851 3927
rect 13277 3893 13311 3927
rect 14841 3893 14875 3927
rect 16497 3893 16531 3927
rect 17325 3893 17359 3927
rect 22017 3893 22051 3927
rect 26341 3893 26375 3927
rect 26709 3893 26743 3927
rect 28089 3893 28123 3927
rect 31585 3893 31619 3927
rect 32321 3893 32355 3927
rect 32689 3893 32723 3927
rect 34437 3893 34471 3927
rect 36645 3893 36679 3927
rect 39037 3893 39071 3927
rect 1593 3689 1627 3723
rect 3617 3689 3651 3723
rect 4629 3689 4663 3723
rect 6837 3689 6871 3723
rect 7665 3689 7699 3723
rect 7849 3689 7883 3723
rect 8585 3689 8619 3723
rect 11713 3689 11747 3723
rect 18981 3689 19015 3723
rect 21833 3689 21867 3723
rect 24501 3689 24535 3723
rect 27629 3689 27663 3723
rect 32873 3689 32907 3723
rect 36461 3689 36495 3723
rect 38485 3689 38519 3723
rect 39405 3689 39439 3723
rect 2053 3621 2087 3655
rect 6101 3621 6135 3655
rect 10517 3621 10551 3655
rect 12357 3621 12391 3655
rect 13093 3621 13127 3655
rect 15945 3621 15979 3655
rect 17233 3621 17267 3655
rect 19901 3621 19935 3655
rect 30941 3621 30975 3655
rect 33149 3621 33183 3655
rect 39037 3621 39071 3655
rect 2605 3553 2639 3587
rect 5089 3553 5123 3587
rect 6193 3553 6227 3587
rect 6285 3553 6319 3587
rect 6653 3553 6687 3587
rect 7205 3553 7239 3587
rect 7941 3553 7975 3587
rect 9229 3553 9263 3587
rect 10793 3553 10827 3587
rect 11069 3553 11103 3587
rect 13645 3553 13679 3587
rect 14749 3553 14783 3587
rect 15025 3553 15059 3587
rect 15163 3553 15197 3587
rect 16681 3553 16715 3587
rect 16840 3553 16874 3587
rect 17693 3553 17727 3587
rect 19441 3553 19475 3587
rect 20294 3553 20328 3587
rect 20453 3553 20487 3587
rect 25513 3553 25547 3587
rect 26433 3553 26467 3587
rect 26709 3553 26743 3587
rect 26826 3553 26860 3587
rect 27721 3553 27755 3587
rect 29929 3553 29963 3587
rect 31033 3553 31067 3587
rect 31677 3553 31711 3587
rect 32229 3553 32263 3587
rect 34345 3553 34379 3587
rect 1501 3485 1535 3519
rect 1869 3485 1903 3519
rect 2881 3485 2915 3519
rect 3893 3485 3927 3519
rect 4261 3485 4295 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 4813 3485 4847 3519
rect 5365 3485 5399 3519
rect 6561 3485 6595 3519
rect 6929 3485 6963 3519
rect 7021 3485 7055 3519
rect 7297 3485 7331 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 9321 3485 9355 3519
rect 9873 3485 9907 3519
rect 10057 3485 10091 3519
rect 10910 3485 10944 3519
rect 11805 3485 11839 3519
rect 11989 3485 12023 3519
rect 12081 3485 12115 3519
rect 12173 3485 12207 3519
rect 12909 3485 12943 3519
rect 13369 3485 13403 3519
rect 14105 3485 14139 3519
rect 14289 3485 14323 3519
rect 15301 3485 15335 3519
rect 16957 3485 16991 3519
rect 17877 3485 17911 3519
rect 17969 3485 18003 3519
rect 18245 3485 18279 3519
rect 19257 3485 19291 3519
rect 20177 3485 20211 3519
rect 21465 3485 21499 3519
rect 22569 3485 22603 3519
rect 22845 3485 22879 3519
rect 23857 3485 23891 3519
rect 24133 3485 24167 3519
rect 25237 3485 25271 3519
rect 25789 3485 25823 3519
rect 25973 3485 26007 3519
rect 26985 3485 27019 3519
rect 27997 3485 28031 3519
rect 28825 3485 28859 3519
rect 29193 3485 29227 3519
rect 29561 3485 29595 3519
rect 30205 3485 30239 3519
rect 31217 3485 31251 3519
rect 31953 3485 31987 3519
rect 32070 3485 32104 3519
rect 32965 3485 32999 3519
rect 34069 3485 34103 3519
rect 34713 3485 34747 3519
rect 35173 3485 35207 3519
rect 38669 3485 38703 3519
rect 38853 3485 38887 3519
rect 39221 3485 39255 3519
rect 2237 3417 2271 3451
rect 2421 3417 2455 3451
rect 7205 3417 7239 3451
rect 8033 3417 8067 3451
rect 12541 3417 12575 3451
rect 13829 3417 13863 3451
rect 21097 3417 21131 3451
rect 23029 3417 23063 3451
rect 3985 3349 4019 3383
rect 4445 3349 4479 3383
rect 4997 3349 5031 3383
rect 6469 3349 6503 3383
rect 7665 3349 7699 3383
rect 8217 3349 8251 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 9781 3349 9815 3383
rect 12633 3349 12667 3383
rect 13553 3349 13587 3383
rect 16037 3349 16071 3383
rect 21649 3349 21683 3383
rect 23121 3349 23155 3383
rect 28733 3349 28767 3383
rect 29009 3349 29043 3383
rect 29377 3349 29411 3383
rect 29745 3349 29779 3383
rect 33333 3349 33367 3383
rect 34897 3349 34931 3383
rect 1961 3145 1995 3179
rect 3249 3145 3283 3179
rect 4353 3145 4387 3179
rect 11345 3145 11379 3179
rect 13829 3145 13863 3179
rect 14105 3145 14139 3179
rect 16497 3145 16531 3179
rect 28825 3145 28859 3179
rect 31861 3145 31895 3179
rect 33701 3145 33735 3179
rect 33793 3145 33827 3179
rect 36093 3145 36127 3179
rect 36553 3145 36587 3179
rect 37749 3145 37783 3179
rect 38025 3145 38059 3179
rect 39405 3145 39439 3179
rect 1501 3077 1535 3111
rect 24685 3077 24719 3111
rect 38669 3077 38703 3111
rect 1869 3009 1903 3043
rect 2513 3009 2547 3043
rect 3617 3009 3651 3043
rect 4537 3009 4571 3043
rect 4997 3009 5031 3043
rect 5181 3009 5215 3043
rect 5457 3009 5491 3043
rect 6377 3009 6411 3043
rect 6653 3009 6687 3043
rect 7481 3009 7515 3043
rect 8033 3009 8067 3043
rect 8953 3009 8987 3043
rect 9505 3009 9539 3043
rect 10333 3009 10367 3043
rect 10609 3009 10643 3043
rect 12541 3009 12575 3043
rect 13093 3009 13127 3043
rect 13921 3009 13955 3043
rect 14473 3009 14507 3043
rect 15117 3009 15151 3043
rect 15761 3009 15795 3043
rect 16773 3009 16807 3043
rect 17141 3009 17175 3043
rect 17509 3009 17543 3043
rect 19349 3009 19383 3043
rect 19625 3009 19659 3043
rect 20361 3009 20395 3043
rect 21373 3009 21407 3043
rect 22109 3009 22143 3043
rect 23029 3009 23063 3043
rect 23765 3009 23799 3043
rect 24041 3009 24075 3043
rect 25513 3009 25547 3043
rect 25881 3009 25915 3043
rect 26525 3009 26559 3043
rect 26617 3009 26651 3043
rect 26985 3009 27019 3043
rect 27169 3009 27203 3043
rect 28181 3009 28215 3043
rect 29101 3009 29135 3043
rect 29954 3009 29988 3043
rect 31125 3009 31159 3043
rect 32413 3009 32447 3043
rect 33241 3009 33275 3043
rect 34253 3009 34287 3043
rect 34621 3009 34655 3043
rect 34989 3009 35023 3043
rect 35357 3009 35391 3043
rect 35725 3009 35759 3043
rect 36277 3009 36311 3043
rect 36369 3009 36403 3043
rect 37933 3009 37967 3043
rect 38209 3009 38243 3043
rect 38301 3009 38335 3043
rect 38761 3009 38795 3043
rect 38853 3009 38887 3043
rect 39221 3009 39255 3043
rect 2237 2941 2271 2975
rect 3341 2941 3375 2975
rect 7757 2941 7791 2975
rect 9229 2941 9263 2975
rect 11621 2941 11655 2975
rect 11897 2941 11931 2975
rect 12817 2941 12851 2975
rect 15393 2941 15427 2975
rect 15485 2941 15519 2975
rect 18153 2941 18187 2975
rect 18312 2941 18346 2975
rect 18429 2941 18463 2975
rect 19165 2941 19199 2975
rect 19441 2941 19475 2975
rect 20478 2941 20512 2975
rect 20637 2941 20671 2975
rect 21833 2941 21867 2975
rect 22845 2941 22879 2975
rect 23489 2941 23523 2975
rect 23903 2941 23937 2975
rect 25789 2941 25823 2975
rect 27629 2941 27663 2975
rect 27905 2941 27939 2975
rect 28043 2941 28077 2975
rect 28917 2941 28951 2975
rect 29837 2941 29871 2975
rect 30113 2941 30147 2975
rect 30849 2941 30883 2975
rect 32137 2941 32171 2975
rect 33517 2941 33551 2975
rect 1685 2873 1719 2907
rect 4721 2873 4755 2907
rect 6193 2873 6227 2907
rect 10241 2873 10275 2907
rect 12725 2873 12759 2907
rect 18705 2873 18739 2907
rect 20085 2873 20119 2907
rect 21557 2873 21591 2907
rect 24777 2873 24811 2907
rect 29561 2873 29595 2907
rect 33149 2873 33183 2907
rect 34437 2873 34471 2907
rect 38485 2873 38519 2907
rect 4905 2805 4939 2839
rect 7573 2805 7607 2839
rect 8769 2805 8803 2839
rect 9045 2805 9079 2839
rect 14289 2805 14323 2839
rect 16957 2805 16991 2839
rect 17325 2805 17359 2839
rect 21281 2805 21315 2839
rect 26065 2805 26099 2839
rect 26341 2805 26375 2839
rect 26801 2805 26835 2839
rect 30757 2805 30791 2839
rect 34161 2805 34195 2839
rect 34805 2805 34839 2839
rect 35173 2805 35207 2839
rect 35541 2805 35575 2839
rect 35909 2805 35943 2839
rect 39037 2805 39071 2839
rect 1593 2601 1627 2635
rect 3525 2601 3559 2635
rect 4629 2601 4663 2635
rect 7481 2601 7515 2635
rect 11805 2601 11839 2635
rect 13737 2601 13771 2635
rect 17233 2601 17267 2635
rect 17785 2601 17819 2635
rect 20269 2601 20303 2635
rect 21373 2601 21407 2635
rect 39405 2601 39439 2635
rect 7297 2533 7331 2567
rect 11989 2533 12023 2567
rect 13369 2533 13403 2567
rect 16497 2533 16531 2567
rect 16957 2533 16991 2567
rect 22845 2533 22879 2567
rect 23949 2533 23983 2567
rect 26249 2533 26283 2567
rect 26985 2533 27019 2567
rect 29377 2533 29411 2567
rect 30573 2533 30607 2567
rect 31861 2533 31895 2567
rect 32321 2533 32355 2567
rect 34529 2533 34563 2567
rect 36001 2533 36035 2567
rect 38301 2533 38335 2567
rect 2789 2465 2823 2499
rect 3157 2465 3191 2499
rect 6193 2465 6227 2499
rect 7573 2465 7607 2499
rect 8217 2465 8251 2499
rect 11897 2465 11931 2499
rect 12357 2465 12391 2499
rect 15485 2465 15519 2499
rect 19257 2465 19291 2499
rect 20361 2465 20395 2499
rect 22937 2465 22971 2499
rect 30849 2465 30883 2499
rect 1501 2397 1535 2431
rect 2237 2397 2271 2431
rect 2973 2397 3007 2431
rect 4537 2397 4571 2431
rect 5917 2397 5951 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 7849 2397 7883 2431
rect 7941 2397 7975 2431
rect 9413 2397 9447 2431
rect 9689 2397 9723 2431
rect 11069 2397 11103 2431
rect 11345 2397 11379 2431
rect 11529 2397 11563 2431
rect 12081 2397 12115 2431
rect 12633 2397 12667 2431
rect 13553 2397 13587 2431
rect 13921 2397 13955 2431
rect 14105 2397 14139 2431
rect 14381 2397 14415 2431
rect 14657 2397 14691 2431
rect 15761 2397 15795 2431
rect 17049 2397 17083 2431
rect 19073 2397 19107 2431
rect 19533 2397 19567 2431
rect 20637 2397 20671 2431
rect 21465 2397 21499 2431
rect 21833 2397 21867 2431
rect 22109 2397 22143 2431
rect 23213 2397 23247 2431
rect 24041 2397 24075 2431
rect 24685 2397 24719 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 25513 2397 25547 2431
rect 26341 2397 26375 2431
rect 27721 2397 27755 2431
rect 27997 2397 28031 2431
rect 28089 2397 28123 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 29561 2397 29595 2431
rect 29837 2397 29871 2431
rect 31125 2397 31159 2431
rect 32137 2397 32171 2431
rect 32505 2397 32539 2431
rect 33149 2397 33183 2431
rect 33241 2397 33275 2431
rect 33885 2397 33919 2431
rect 33977 2397 34011 2431
rect 34345 2397 34379 2431
rect 34713 2397 34747 2431
rect 35081 2397 35115 2431
rect 35449 2397 35483 2431
rect 35817 2397 35851 2431
rect 36369 2397 36403 2431
rect 37749 2397 37783 2431
rect 38117 2397 38151 2431
rect 38485 2397 38519 2431
rect 38853 2397 38887 2431
rect 39221 2397 39255 2431
rect 1869 2329 1903 2363
rect 2421 2329 2455 2363
rect 2605 2329 2639 2363
rect 3433 2329 3467 2363
rect 3985 2329 4019 2363
rect 4169 2329 4203 2363
rect 4905 2329 4939 2363
rect 9137 2329 9171 2363
rect 16773 2329 16807 2363
rect 1961 2261 1995 2295
rect 4997 2261 5031 2295
rect 5181 2261 5215 2295
rect 9229 2261 9263 2295
rect 11621 2261 11655 2295
rect 12265 2261 12299 2295
rect 14289 2261 14323 2295
rect 15393 2261 15427 2295
rect 21649 2261 21683 2295
rect 24225 2261 24259 2295
rect 24501 2261 24535 2295
rect 24961 2261 24995 2295
rect 26525 2261 26559 2295
rect 28273 2261 28307 2295
rect 32689 2261 32723 2295
rect 32965 2261 32999 2295
rect 33425 2261 33459 2295
rect 33793 2261 33827 2295
rect 34161 2261 34195 2295
rect 34897 2261 34931 2295
rect 35265 2261 35299 2295
rect 35633 2261 35667 2295
rect 36185 2261 36219 2295
rect 37933 2261 37967 2295
rect 38669 2261 38703 2295
rect 39037 2261 39071 2295
<< metal1 >>
rect 5626 10820 5632 10872
rect 5684 10860 5690 10872
rect 16390 10860 16396 10872
rect 5684 10832 16396 10860
rect 5684 10820 5690 10832
rect 16390 10820 16396 10832
rect 16448 10820 16454 10872
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 18322 10792 18328 10804
rect 2924 10764 18328 10792
rect 2924 10752 2930 10764
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 7650 10684 7656 10736
rect 7708 10724 7714 10736
rect 19426 10724 19432 10736
rect 7708 10696 19432 10724
rect 7708 10684 7714 10696
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 13354 10656 13360 10668
rect 12676 10628 13360 10656
rect 12676 10616 12682 10628
rect 13354 10616 13360 10628
rect 13412 10656 13418 10668
rect 28534 10656 28540 10668
rect 13412 10628 28540 10656
rect 13412 10616 13418 10628
rect 28534 10616 28540 10628
rect 28592 10616 28598 10668
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 23934 10588 23940 10600
rect 14424 10560 23940 10588
rect 14424 10548 14430 10560
rect 23934 10548 23940 10560
rect 23992 10548 23998 10600
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 17678 10520 17684 10532
rect 9824 10492 17684 10520
rect 9824 10480 9830 10492
rect 17678 10480 17684 10492
rect 17736 10480 17742 10532
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 17828 10492 31754 10520
rect 17828 10480 17834 10492
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 17034 10452 17040 10464
rect 6236 10424 17040 10452
rect 6236 10412 6242 10424
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 22738 10452 22744 10464
rect 17276 10424 22744 10452
rect 17276 10412 17282 10424
rect 22738 10412 22744 10424
rect 22796 10412 22802 10464
rect 31726 10452 31754 10492
rect 33778 10452 33784 10464
rect 31726 10424 33784 10452
rect 33778 10412 33784 10424
rect 33836 10412 33842 10464
rect 9306 10344 9312 10396
rect 9364 10384 9370 10396
rect 32398 10384 32404 10396
rect 9364 10356 32404 10384
rect 9364 10344 9370 10356
rect 32398 10344 32404 10356
rect 32456 10344 32462 10396
rect 28902 10316 28908 10328
rect 2746 10288 28908 10316
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 2746 10248 2774 10288
rect 28902 10276 28908 10288
rect 28960 10276 28966 10328
rect 31202 10248 31208 10260
rect 1636 10220 2774 10248
rect 7576 10220 31208 10248
rect 1636 10208 1642 10220
rect 2590 10072 2596 10124
rect 2648 10112 2654 10124
rect 7576 10112 7604 10220
rect 31202 10208 31208 10220
rect 31260 10208 31266 10260
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 17218 10180 17224 10192
rect 9640 10152 17224 10180
rect 9640 10140 9646 10152
rect 17218 10140 17224 10152
rect 17276 10140 17282 10192
rect 17954 10140 17960 10192
rect 18012 10180 18018 10192
rect 26694 10180 26700 10192
rect 18012 10152 26700 10180
rect 18012 10140 18018 10152
rect 26694 10140 26700 10152
rect 26752 10140 26758 10192
rect 35618 10180 35624 10192
rect 26804 10152 35624 10180
rect 2648 10084 7604 10112
rect 2648 10072 2654 10084
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 21910 10112 21916 10124
rect 12308 10084 21916 10112
rect 12308 10072 12314 10084
rect 21910 10072 21916 10084
rect 21968 10072 21974 10124
rect 26804 10112 26832 10152
rect 35618 10140 35624 10152
rect 35676 10140 35682 10192
rect 22296 10084 26832 10112
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 22296 10044 22324 10084
rect 27062 10072 27068 10124
rect 27120 10112 27126 10124
rect 36078 10112 36084 10124
rect 27120 10084 36084 10112
rect 27120 10072 27126 10084
rect 36078 10072 36084 10084
rect 36136 10072 36142 10124
rect 16540 10016 22324 10044
rect 16540 10004 16546 10016
rect 26970 10004 26976 10056
rect 27028 10044 27034 10056
rect 34054 10044 34060 10056
rect 27028 10016 34060 10044
rect 27028 10004 27034 10016
rect 34054 10004 34060 10016
rect 34112 10004 34118 10056
rect 1302 9936 1308 9988
rect 1360 9976 1366 9988
rect 21358 9976 21364 9988
rect 1360 9948 21364 9976
rect 1360 9936 1366 9948
rect 21358 9936 21364 9948
rect 21416 9936 21422 9988
rect 22462 9936 22468 9988
rect 22520 9976 22526 9988
rect 34238 9976 34244 9988
rect 22520 9948 34244 9976
rect 22520 9936 22526 9948
rect 34238 9936 34244 9948
rect 34296 9936 34302 9988
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 12342 9908 12348 9920
rect 2556 9880 12348 9908
rect 2556 9868 2562 9880
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 21910 9868 21916 9920
rect 21968 9908 21974 9920
rect 34422 9908 34428 9920
rect 21968 9880 34428 9908
rect 21968 9868 21974 9880
rect 34422 9868 34428 9880
rect 34480 9868 34486 9920
rect 2314 9800 2320 9852
rect 2372 9840 2378 9852
rect 9674 9840 9680 9852
rect 2372 9812 9680 9840
rect 2372 9800 2378 9812
rect 9674 9800 9680 9812
rect 9732 9800 9738 9852
rect 16574 9800 16580 9852
rect 16632 9840 16638 9852
rect 16632 9812 21588 9840
rect 16632 9800 16638 9812
rect 7374 9732 7380 9784
rect 7432 9772 7438 9784
rect 7432 9744 15332 9772
rect 7432 9732 7438 9744
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 15304 9704 15332 9744
rect 15378 9732 15384 9784
rect 15436 9772 15442 9784
rect 20714 9772 20720 9784
rect 15436 9744 20720 9772
rect 15436 9732 15442 9744
rect 20714 9732 20720 9744
rect 20772 9732 20778 9784
rect 15470 9704 15476 9716
rect 3844 9676 9720 9704
rect 15304 9676 15476 9704
rect 3844 9664 3850 9676
rect 9692 9636 9720 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 20438 9664 20444 9716
rect 20496 9704 20502 9716
rect 21450 9704 21456 9716
rect 20496 9676 21456 9704
rect 20496 9664 20502 9676
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 21560 9704 21588 9812
rect 22094 9800 22100 9852
rect 22152 9840 22158 9852
rect 35986 9840 35992 9852
rect 22152 9812 35992 9840
rect 22152 9800 22158 9812
rect 35986 9800 35992 9812
rect 36044 9800 36050 9852
rect 22646 9732 22652 9784
rect 22704 9772 22710 9784
rect 23658 9772 23664 9784
rect 22704 9744 23664 9772
rect 22704 9732 22710 9744
rect 23658 9732 23664 9744
rect 23716 9732 23722 9784
rect 24670 9732 24676 9784
rect 24728 9772 24734 9784
rect 24728 9744 31754 9772
rect 24728 9732 24734 9744
rect 26970 9704 26976 9716
rect 21560 9676 26976 9704
rect 26970 9664 26976 9676
rect 27028 9664 27034 9716
rect 28166 9664 28172 9716
rect 28224 9704 28230 9716
rect 29638 9704 29644 9716
rect 28224 9676 29644 9704
rect 28224 9664 28230 9676
rect 29638 9664 29644 9676
rect 29696 9664 29702 9716
rect 31726 9704 31754 9744
rect 33410 9704 33416 9716
rect 31726 9676 33416 9704
rect 33410 9664 33416 9676
rect 33468 9664 33474 9716
rect 16482 9636 16488 9648
rect 9692 9608 16488 9636
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 22830 9596 22836 9648
rect 22888 9636 22894 9648
rect 22888 9608 31754 9636
rect 22888 9596 22894 9608
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6328 9540 13216 9568
rect 6328 9528 6334 9540
rect 8662 9460 8668 9512
rect 8720 9500 8726 9512
rect 8720 9472 9674 9500
rect 8720 9460 8726 9472
rect 9646 9432 9674 9472
rect 13078 9432 13084 9444
rect 9646 9404 13084 9432
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 12066 9364 12072 9376
rect 3752 9336 12072 9364
rect 3752 9324 3758 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 2774 9256 2780 9308
rect 2832 9256 2838 9308
rect 4246 9256 4252 9308
rect 4304 9296 4310 9308
rect 9490 9296 9496 9308
rect 4304 9268 9496 9296
rect 4304 9256 4310 9268
rect 9490 9256 9496 9268
rect 9548 9256 9554 9308
rect 13188 9296 13216 9540
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 23566 9568 23572 9580
rect 15068 9540 23572 9568
rect 15068 9528 15074 9540
rect 23566 9528 23572 9540
rect 23624 9528 23630 9580
rect 13280 9500 13308 9528
rect 31478 9500 31484 9512
rect 13280 9472 31484 9500
rect 31478 9460 31484 9472
rect 31536 9460 31542 9512
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 20622 9432 20628 9444
rect 13320 9404 20628 9432
rect 13320 9392 13326 9404
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 30006 9432 30012 9444
rect 22244 9404 30012 9432
rect 22244 9392 22250 9404
rect 30006 9392 30012 9404
rect 30064 9392 30070 9444
rect 31726 9432 31754 9608
rect 35250 9432 35256 9444
rect 31726 9404 35256 9432
rect 35250 9392 35256 9404
rect 35308 9392 35314 9444
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 25682 9364 25688 9376
rect 16908 9336 25688 9364
rect 16908 9324 16914 9336
rect 25682 9324 25688 9336
rect 25740 9324 25746 9376
rect 25774 9324 25780 9376
rect 25832 9364 25838 9376
rect 36630 9364 36636 9376
rect 25832 9336 36636 9364
rect 25832 9324 25838 9336
rect 36630 9324 36636 9336
rect 36688 9324 36694 9376
rect 26694 9296 26700 9308
rect 13188 9268 26700 9296
rect 26694 9256 26700 9268
rect 26752 9256 26758 9308
rect 37182 9256 37188 9308
rect 37240 9296 37246 9308
rect 38562 9296 38568 9308
rect 37240 9268 38568 9296
rect 37240 9256 37246 9268
rect 38562 9256 38568 9268
rect 38620 9256 38626 9308
rect 2792 9092 2820 9256
rect 6638 9188 6644 9240
rect 6696 9228 6702 9240
rect 10870 9228 10876 9240
rect 6696 9200 10876 9228
rect 6696 9188 6702 9200
rect 10870 9188 10876 9200
rect 10928 9188 10934 9240
rect 12526 9188 12532 9240
rect 12584 9228 12590 9240
rect 15010 9228 15016 9240
rect 12584 9200 15016 9228
rect 12584 9188 12590 9200
rect 15010 9188 15016 9200
rect 15068 9188 15074 9240
rect 15102 9188 15108 9240
rect 15160 9228 15166 9240
rect 17954 9228 17960 9240
rect 15160 9200 17960 9228
rect 15160 9188 15166 9200
rect 17954 9188 17960 9200
rect 18012 9188 18018 9240
rect 19518 9188 19524 9240
rect 19576 9228 19582 9240
rect 24118 9228 24124 9240
rect 19576 9200 24124 9228
rect 19576 9188 19582 9200
rect 24118 9188 24124 9200
rect 24176 9188 24182 9240
rect 24210 9188 24216 9240
rect 24268 9228 24274 9240
rect 36814 9228 36820 9240
rect 24268 9200 36820 9228
rect 24268 9188 24274 9200
rect 36814 9188 36820 9200
rect 36872 9188 36878 9240
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 20530 9160 20536 9172
rect 8536 9132 20536 9160
rect 8536 9120 8542 9132
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 20622 9120 20628 9172
rect 20680 9160 20686 9172
rect 22186 9160 22192 9172
rect 20680 9132 22192 9160
rect 20680 9120 20686 9132
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 26786 9160 26792 9172
rect 22336 9132 26792 9160
rect 22336 9120 22342 9132
rect 26786 9120 26792 9132
rect 26844 9120 26850 9172
rect 31386 9160 31392 9172
rect 26896 9132 31392 9160
rect 2866 9092 2872 9104
rect 2792 9064 2872 9092
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 5626 9092 5632 9104
rect 4580 9064 5632 9092
rect 4580 9052 4586 9064
rect 5626 9052 5632 9064
rect 5684 9052 5690 9104
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 26896 9092 26924 9132
rect 31386 9120 31392 9132
rect 31444 9120 31450 9172
rect 8628 9064 26924 9092
rect 8628 9052 8634 9064
rect 4062 8984 4068 9036
rect 4120 9024 4126 9036
rect 10226 9024 10232 9036
rect 4120 8996 10232 9024
rect 4120 8984 4126 8996
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 14826 9024 14832 9036
rect 12728 8996 14832 9024
rect 2406 8916 2412 8968
rect 2464 8956 2470 8968
rect 12526 8956 12532 8968
rect 2464 8928 12532 8956
rect 2464 8916 2470 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 1912 8860 2774 8888
rect 1912 8848 1918 8860
rect 2746 8820 2774 8860
rect 5258 8848 5264 8900
rect 5316 8888 5322 8900
rect 12728 8888 12756 8996
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 15654 8984 15660 9036
rect 15712 9024 15718 9036
rect 15712 8996 23796 9024
rect 15712 8984 15718 8996
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 22002 8956 22008 8968
rect 14516 8928 22008 8956
rect 14516 8916 14522 8928
rect 22002 8916 22008 8928
rect 22060 8916 22066 8968
rect 23768 8956 23796 8996
rect 23842 8984 23848 9036
rect 23900 9024 23906 9036
rect 35802 9024 35808 9036
rect 23900 8996 35808 9024
rect 23900 8984 23906 8996
rect 35802 8984 35808 8996
rect 35860 8984 35866 9036
rect 24394 8956 24400 8968
rect 23768 8928 24400 8956
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 26326 8916 26332 8968
rect 26384 8956 26390 8968
rect 37366 8956 37372 8968
rect 26384 8928 37372 8956
rect 26384 8916 26390 8928
rect 37366 8916 37372 8928
rect 37424 8916 37430 8968
rect 5316 8860 12756 8888
rect 5316 8848 5322 8860
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 19702 8888 19708 8900
rect 12860 8860 19708 8888
rect 12860 8848 12866 8860
rect 19702 8848 19708 8860
rect 19760 8848 19766 8900
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 24578 8888 24584 8900
rect 20772 8860 24584 8888
rect 20772 8848 20778 8860
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 25866 8848 25872 8900
rect 25924 8888 25930 8900
rect 32858 8888 32864 8900
rect 25924 8860 32864 8888
rect 25924 8848 25930 8860
rect 32858 8848 32864 8860
rect 32916 8848 32922 8900
rect 33594 8848 33600 8900
rect 33652 8888 33658 8900
rect 36354 8888 36360 8900
rect 33652 8860 36360 8888
rect 33652 8848 33658 8860
rect 36354 8848 36360 8860
rect 36412 8848 36418 8900
rect 37734 8888 37740 8900
rect 36832 8860 37740 8888
rect 7466 8820 7472 8832
rect 2746 8792 7472 8820
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 16482 8820 16488 8832
rect 8444 8792 16488 8820
rect 8444 8780 8450 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 19610 8780 19616 8832
rect 19668 8820 19674 8832
rect 22278 8820 22284 8832
rect 19668 8792 22284 8820
rect 19668 8780 19674 8792
rect 22278 8780 22284 8792
rect 22336 8780 22342 8832
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 28350 8820 28356 8832
rect 22428 8792 28356 8820
rect 22428 8780 22434 8792
rect 28350 8780 28356 8792
rect 28408 8780 28414 8832
rect 28902 8780 28908 8832
rect 28960 8820 28966 8832
rect 30282 8820 30288 8832
rect 28960 8792 30288 8820
rect 28960 8780 28966 8792
rect 30282 8780 30288 8792
rect 30340 8780 30346 8832
rect 30742 8780 30748 8832
rect 30800 8820 30806 8832
rect 36832 8820 36860 8860
rect 37734 8848 37740 8860
rect 37792 8848 37798 8900
rect 30800 8792 36860 8820
rect 30800 8780 30806 8792
rect 36906 8780 36912 8832
rect 36964 8820 36970 8832
rect 38470 8820 38476 8832
rect 36964 8792 38476 8820
rect 36964 8780 36970 8792
rect 38470 8780 38476 8792
rect 38528 8780 38534 8832
rect 1104 8730 39836 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 9010 8730
rect 9062 8678 9074 8730
rect 9126 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 15010 8730
rect 15062 8678 15074 8730
rect 15126 8678 15138 8730
rect 15190 8678 15202 8730
rect 15254 8678 15266 8730
rect 15318 8678 21010 8730
rect 21062 8678 21074 8730
rect 21126 8678 21138 8730
rect 21190 8678 21202 8730
rect 21254 8678 21266 8730
rect 21318 8678 27010 8730
rect 27062 8678 27074 8730
rect 27126 8678 27138 8730
rect 27190 8678 27202 8730
rect 27254 8678 27266 8730
rect 27318 8678 33010 8730
rect 33062 8678 33074 8730
rect 33126 8678 33138 8730
rect 33190 8678 33202 8730
rect 33254 8678 33266 8730
rect 33318 8678 39010 8730
rect 39062 8678 39074 8730
rect 39126 8678 39138 8730
rect 39190 8678 39202 8730
rect 39254 8678 39266 8730
rect 39318 8678 39836 8730
rect 1104 8656 39836 8678
rect 2498 8576 2504 8628
rect 2556 8576 2562 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2924 8588 2973 8616
rect 2924 8576 2930 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 3694 8616 3700 8628
rect 2961 8579 3019 8585
rect 3252 8588 3700 8616
rect 1670 8508 1676 8560
rect 1728 8508 1734 8560
rect 3252 8548 3280 8588
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 4212 8588 4629 8616
rect 4212 8576 4218 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 4617 8579 4675 8585
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5994 8616 6000 8628
rect 5675 8588 6000 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6144 8588 6469 8616
rect 6144 8576 6150 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 7009 8619 7067 8625
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 7190 8616 7196 8628
rect 7055 8588 7196 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7524 8588 8156 8616
rect 7524 8576 7530 8588
rect 2746 8520 3280 8548
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1688 8480 1716 8508
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1688 8452 2329 8480
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2746 8412 2774 8520
rect 3326 8508 3332 8560
rect 3384 8508 3390 8560
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 4246 8508 4252 8560
rect 4304 8508 4310 8560
rect 4430 8508 4436 8560
rect 4488 8508 4494 8560
rect 5442 8548 5448 8560
rect 4724 8520 5448 8548
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 4062 8480 4068 8492
rect 3191 8452 4068 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 1719 8384 2774 8412
rect 3513 8415 3571 8421
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 4724 8412 4752 8520
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5534 8508 5540 8560
rect 5592 8508 5598 8560
rect 8128 8548 8156 8588
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8352 8588 9045 8616
rect 8352 8576 8358 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9033 8579 9091 8585
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9456 8588 9597 8616
rect 9456 8576 9462 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10560 8588 10701 8616
rect 10560 8576 10566 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11664 8588 11897 8616
rect 11664 8576 11670 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 12710 8616 12716 8628
rect 12667 8588 12716 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 13872 8588 14197 8616
rect 13872 8576 13878 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 15105 8619 15163 8625
rect 15105 8616 15117 8619
rect 14976 8588 15117 8616
rect 14976 8576 14982 8588
rect 15105 8585 15117 8588
rect 15151 8585 15163 8619
rect 15105 8579 15163 8585
rect 15654 8576 15660 8628
rect 15712 8576 15718 8628
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 16080 8588 16221 8616
rect 16080 8576 16086 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 16209 8579 16267 8585
rect 16850 8576 16856 8628
rect 16908 8576 16914 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17126 8616 17132 8628
rect 17083 8588 17132 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18509 8619 18567 8625
rect 18509 8616 18521 8619
rect 18288 8588 18521 8616
rect 18288 8576 18294 8588
rect 18509 8585 18521 8588
rect 18555 8585 18567 8619
rect 18509 8579 18567 8585
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 19392 8588 19625 8616
rect 19392 8576 19398 8588
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19613 8579 19671 8585
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 19760 8588 21404 8616
rect 19760 8576 19766 8588
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 5644 8520 7788 8548
rect 8128 8520 8401 8548
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 5040 8452 5089 8480
rect 5040 8440 5046 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 5644 8480 5672 8520
rect 5316 8452 5672 8480
rect 5316 8440 5322 8452
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 7466 8440 7472 8492
rect 7524 8440 7530 8492
rect 5718 8412 5724 8424
rect 3559 8384 4752 8412
rect 4816 8384 5724 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 4816 8344 4844 8384
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 7190 8372 7196 8424
rect 7248 8372 7254 8424
rect 7760 8412 7788 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 8389 8511 8447 8517
rect 8404 8480 8432 8511
rect 8570 8508 8576 8560
rect 8628 8508 8634 8560
rect 9674 8548 9680 8560
rect 9048 8520 9680 8548
rect 9048 8480 9076 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 11146 8548 11152 8560
rect 10888 8520 11152 8548
rect 8404 8452 9076 8480
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8480 9275 8483
rect 9582 8480 9588 8492
rect 9263 8452 9588 8480
rect 9263 8449 9275 8452
rect 9217 8443 9275 8449
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9766 8440 9772 8492
rect 9824 8440 9830 8492
rect 10888 8489 10916 8520
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 11238 8508 11244 8560
rect 11296 8508 11302 8560
rect 14642 8548 14648 8560
rect 12820 8520 14648 8548
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 12820 8489 12848 8520
rect 14642 8508 14648 8520
rect 14700 8508 14706 8560
rect 20898 8548 20904 8560
rect 14752 8520 17908 8548
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 11716 8412 11744 8443
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 7760 8384 11744 8412
rect 12894 8372 12900 8424
rect 12952 8372 12958 8424
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14752 8412 14780 8520
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 15378 8480 15384 8492
rect 15335 8452 15384 8480
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8480 15531 8483
rect 15746 8480 15752 8492
rect 15519 8452 15752 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16574 8480 16580 8492
rect 16439 8452 16580 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 17552 8452 17601 8480
rect 17552 8440 17558 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 14332 8384 14780 8412
rect 14332 8372 14338 8384
rect 17310 8372 17316 8424
rect 17368 8372 17374 8424
rect 17880 8412 17908 8520
rect 18708 8520 20904 8548
rect 18708 8489 18736 8520
rect 20898 8508 20904 8520
rect 20956 8508 20962 8560
rect 18693 8483 18751 8489
rect 18693 8449 18705 8483
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 20438 8480 20444 8492
rect 20303 8452 20444 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 19444 8412 19472 8443
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20530 8440 20536 8492
rect 20588 8440 20594 8492
rect 21376 8489 21404 8588
rect 21542 8576 21548 8628
rect 21600 8616 21606 8628
rect 21913 8619 21971 8625
rect 21913 8616 21925 8619
rect 21600 8588 21925 8616
rect 21600 8576 21606 8588
rect 21913 8585 21925 8588
rect 21959 8585 21971 8619
rect 21913 8579 21971 8585
rect 22370 8576 22376 8628
rect 22428 8576 22434 8628
rect 23658 8576 23664 8628
rect 23716 8576 23722 8628
rect 23750 8576 23756 8628
rect 23808 8616 23814 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 23808 8588 24041 8616
rect 23808 8576 23814 8588
rect 24029 8585 24041 8588
rect 24075 8585 24087 8619
rect 24029 8579 24087 8585
rect 24489 8619 24547 8625
rect 24489 8585 24501 8619
rect 24535 8616 24547 8619
rect 24762 8616 24768 8628
rect 24535 8588 24768 8616
rect 24535 8585 24547 8588
rect 24489 8579 24547 8585
rect 24762 8576 24768 8588
rect 24820 8576 24826 8628
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 26145 8619 26203 8625
rect 26145 8616 26157 8619
rect 26016 8588 26157 8616
rect 26016 8576 26022 8588
rect 26145 8585 26157 8588
rect 26191 8585 26203 8619
rect 26145 8579 26203 8585
rect 29270 8576 29276 8628
rect 29328 8616 29334 8628
rect 30009 8619 30067 8625
rect 30009 8616 30021 8619
rect 29328 8588 30021 8616
rect 29328 8576 29334 8588
rect 30009 8585 30021 8588
rect 30055 8585 30067 8619
rect 30009 8579 30067 8585
rect 30374 8576 30380 8628
rect 30432 8616 30438 8628
rect 30561 8619 30619 8625
rect 30561 8616 30573 8619
rect 30432 8588 30573 8616
rect 30432 8576 30438 8588
rect 30561 8585 30573 8588
rect 30607 8585 30619 8619
rect 31662 8616 31668 8628
rect 30561 8579 30619 8585
rect 30760 8588 31668 8616
rect 30760 8548 30788 8588
rect 31662 8576 31668 8588
rect 31720 8576 31726 8628
rect 31754 8576 31760 8628
rect 31812 8616 31818 8628
rect 32217 8619 32275 8625
rect 32217 8616 32229 8619
rect 31812 8588 32229 8616
rect 31812 8576 31818 8588
rect 32217 8585 32229 8588
rect 32263 8585 32275 8619
rect 32217 8579 32275 8585
rect 32582 8576 32588 8628
rect 32640 8616 32646 8628
rect 32769 8619 32827 8625
rect 32769 8616 32781 8619
rect 32640 8588 32781 8616
rect 32640 8576 32646 8588
rect 32769 8585 32781 8588
rect 32815 8585 32827 8619
rect 32769 8579 32827 8585
rect 33686 8576 33692 8628
rect 33744 8616 33750 8628
rect 33873 8619 33931 8625
rect 33873 8616 33885 8619
rect 33744 8588 33885 8616
rect 33744 8576 33750 8588
rect 33873 8585 33885 8588
rect 33919 8585 33931 8619
rect 33873 8579 33931 8585
rect 34790 8576 34796 8628
rect 34848 8616 34854 8628
rect 34977 8619 35035 8625
rect 34977 8616 34989 8619
rect 34848 8588 34989 8616
rect 34848 8576 34854 8588
rect 34977 8585 34989 8588
rect 35023 8585 35035 8619
rect 34977 8579 35035 8585
rect 35894 8576 35900 8628
rect 35952 8616 35958 8628
rect 36081 8619 36139 8625
rect 36081 8616 36093 8619
rect 35952 8588 36093 8616
rect 35952 8576 35958 8588
rect 36081 8585 36093 8588
rect 36127 8585 36139 8619
rect 36081 8579 36139 8585
rect 36630 8576 36636 8628
rect 36688 8576 36694 8628
rect 37001 8619 37059 8625
rect 37001 8585 37013 8619
rect 37047 8585 37059 8619
rect 37001 8579 37059 8585
rect 36170 8548 36176 8560
rect 21468 8520 22784 8548
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 17880 8384 19472 8412
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 21468 8412 21496 8520
rect 22094 8440 22100 8492
rect 22152 8440 22158 8492
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8480 22247 8483
rect 22370 8480 22376 8492
rect 22235 8452 22376 8480
rect 22235 8449 22247 8452
rect 22189 8443 22247 8449
rect 22370 8440 22376 8452
rect 22428 8440 22434 8492
rect 22756 8489 22784 8520
rect 24688 8520 29776 8548
rect 22741 8483 22799 8489
rect 22741 8449 22753 8483
rect 22787 8449 22799 8483
rect 22741 8443 22799 8449
rect 23842 8440 23848 8492
rect 23900 8440 23906 8492
rect 24210 8440 24216 8492
rect 24268 8440 24274 8492
rect 24688 8489 24716 8520
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 24946 8440 24952 8492
rect 25004 8480 25010 8492
rect 25041 8483 25099 8489
rect 25041 8480 25053 8483
rect 25004 8452 25053 8480
rect 25004 8440 25010 8452
rect 25041 8449 25053 8452
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 26326 8440 26332 8492
rect 26384 8440 26390 8492
rect 27430 8440 27436 8492
rect 27488 8480 27494 8492
rect 28537 8483 28595 8489
rect 28537 8480 28549 8483
rect 27488 8452 28549 8480
rect 27488 8440 27494 8452
rect 28537 8449 28549 8452
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 21048 8384 21496 8412
rect 22204 8384 22477 8412
rect 21048 8372 21054 8384
rect 22204 8356 22232 8384
rect 22465 8381 22477 8384
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 24765 8415 24823 8421
rect 24765 8381 24777 8415
rect 24811 8381 24823 8415
rect 24765 8375 24823 8381
rect 3988 8316 4844 8344
rect 8205 8347 8263 8353
rect 3988 8285 4016 8316
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 8754 8344 8760 8356
rect 8251 8316 8760 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 9674 8304 9680 8356
rect 9732 8344 9738 8356
rect 9732 8316 11560 8344
rect 9732 8304 9738 8316
rect 3973 8279 4031 8285
rect 3973 8245 3985 8279
rect 4019 8245 4031 8279
rect 3973 8239 4031 8245
rect 4798 8236 4804 8288
rect 4856 8276 4862 8288
rect 8294 8276 8300 8288
rect 4856 8248 8300 8276
rect 4856 8236 4862 8248
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 11422 8276 11428 8288
rect 8444 8248 11428 8276
rect 8444 8236 8450 8248
rect 11422 8236 11428 8248
rect 11480 8236 11486 8288
rect 11532 8276 11560 8316
rect 13556 8316 16252 8344
rect 13556 8276 13584 8316
rect 11532 8248 13584 8276
rect 13909 8279 13967 8285
rect 13909 8245 13921 8279
rect 13955 8276 13967 8279
rect 14550 8276 14556 8288
rect 13955 8248 14556 8276
rect 13955 8245 13967 8248
rect 13909 8239 13967 8245
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 16224 8276 16252 8316
rect 18230 8304 18236 8356
rect 18288 8344 18294 8356
rect 18288 8316 19334 8344
rect 18288 8304 18294 8316
rect 18046 8276 18052 8288
rect 16224 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18325 8279 18383 8285
rect 18325 8245 18337 8279
rect 18371 8276 18383 8279
rect 19150 8276 19156 8288
rect 18371 8248 19156 8276
rect 18371 8245 18383 8248
rect 18325 8239 18383 8245
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 19306 8276 19334 8316
rect 21192 8316 21404 8344
rect 21192 8276 21220 8316
rect 19306 8248 21220 8276
rect 21266 8236 21272 8288
rect 21324 8236 21330 8288
rect 21376 8276 21404 8316
rect 21450 8304 21456 8356
rect 21508 8344 21514 8356
rect 21545 8347 21603 8353
rect 21545 8344 21557 8347
rect 21508 8316 21557 8344
rect 21508 8304 21514 8316
rect 21545 8313 21557 8316
rect 21591 8313 21603 8347
rect 21545 8307 21603 8313
rect 22186 8304 22192 8356
rect 22244 8304 22250 8356
rect 23106 8276 23112 8288
rect 21376 8248 23112 8276
rect 23106 8236 23112 8248
rect 23164 8236 23170 8288
rect 23474 8236 23480 8288
rect 23532 8236 23538 8288
rect 24780 8276 24808 8375
rect 26878 8372 26884 8424
rect 26936 8412 26942 8424
rect 27157 8415 27215 8421
rect 27157 8412 27169 8415
rect 26936 8384 27169 8412
rect 26936 8372 26942 8384
rect 27157 8381 27169 8384
rect 27203 8381 27215 8415
rect 28261 8415 28319 8421
rect 28261 8412 28273 8415
rect 27157 8375 27215 8381
rect 27816 8384 28273 8412
rect 26326 8344 26332 8356
rect 25424 8316 26332 8344
rect 24854 8276 24860 8288
rect 24780 8248 24860 8276
rect 24854 8236 24860 8248
rect 24912 8276 24918 8288
rect 25424 8276 25452 8316
rect 26326 8304 26332 8316
rect 26384 8304 26390 8356
rect 24912 8248 25452 8276
rect 24912 8236 24918 8248
rect 25498 8236 25504 8288
rect 25556 8276 25562 8288
rect 25777 8279 25835 8285
rect 25777 8276 25789 8279
rect 25556 8248 25789 8276
rect 25556 8236 25562 8248
rect 25777 8245 25789 8248
rect 25823 8245 25835 8279
rect 26344 8276 26372 8304
rect 27816 8276 27844 8384
rect 28261 8381 28273 8384
rect 28307 8381 28319 8415
rect 28261 8375 28319 8381
rect 29638 8304 29644 8356
rect 29696 8304 29702 8356
rect 26344 8248 27844 8276
rect 25777 8239 25835 8245
rect 28166 8236 28172 8288
rect 28224 8236 28230 8288
rect 29273 8279 29331 8285
rect 29273 8245 29285 8279
rect 29319 8276 29331 8279
rect 29454 8276 29460 8288
rect 29319 8248 29460 8276
rect 29319 8245 29331 8248
rect 29273 8239 29331 8245
rect 29454 8236 29460 8248
rect 29512 8236 29518 8288
rect 29748 8276 29776 8520
rect 30208 8520 30788 8548
rect 30852 8520 36176 8548
rect 30208 8489 30236 8520
rect 29825 8483 29883 8489
rect 29825 8449 29837 8483
rect 29871 8449 29883 8483
rect 29825 8443 29883 8449
rect 30193 8483 30251 8489
rect 30193 8449 30205 8483
rect 30239 8449 30251 8483
rect 30193 8443 30251 8449
rect 29840 8412 29868 8443
rect 30742 8440 30748 8492
rect 30800 8440 30806 8492
rect 30852 8412 30880 8520
rect 36170 8508 36176 8520
rect 36228 8508 36234 8560
rect 37016 8548 37044 8579
rect 37274 8576 37280 8628
rect 37332 8616 37338 8628
rect 37369 8619 37427 8625
rect 37369 8616 37381 8619
rect 37332 8588 37381 8616
rect 37332 8576 37338 8588
rect 37369 8585 37381 8588
rect 37415 8585 37427 8619
rect 37369 8579 37427 8585
rect 38102 8576 38108 8628
rect 38160 8616 38166 8628
rect 38381 8619 38439 8625
rect 38381 8616 38393 8619
rect 38160 8588 38393 8616
rect 38160 8576 38166 8588
rect 38381 8585 38393 8588
rect 38427 8585 38439 8619
rect 38381 8579 38439 8585
rect 39390 8576 39396 8628
rect 39448 8576 39454 8628
rect 38654 8548 38660 8560
rect 37016 8520 38660 8548
rect 38654 8508 38660 8520
rect 38712 8508 38718 8560
rect 31202 8440 31208 8492
rect 31260 8440 31266 8492
rect 32401 8483 32459 8489
rect 32401 8449 32413 8483
rect 32447 8480 32459 8483
rect 32674 8480 32680 8492
rect 32447 8452 32680 8480
rect 32447 8449 32459 8452
rect 32401 8443 32459 8449
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8480 33011 8483
rect 33594 8480 33600 8492
rect 32999 8452 33600 8480
rect 32999 8449 33011 8452
rect 32953 8443 33011 8449
rect 33594 8440 33600 8452
rect 33652 8440 33658 8492
rect 33870 8440 33876 8492
rect 33928 8480 33934 8492
rect 34057 8483 34115 8489
rect 34057 8480 34069 8483
rect 33928 8452 34069 8480
rect 33928 8440 33934 8452
rect 34057 8449 34069 8452
rect 34103 8449 34115 8483
rect 34057 8443 34115 8449
rect 35158 8440 35164 8492
rect 35216 8440 35222 8492
rect 36265 8483 36323 8489
rect 36265 8449 36277 8483
rect 36311 8480 36323 8483
rect 36630 8480 36636 8492
rect 36311 8452 36636 8480
rect 36311 8449 36323 8452
rect 36265 8443 36323 8449
rect 36630 8440 36636 8452
rect 36688 8440 36694 8492
rect 36725 8483 36783 8489
rect 36725 8449 36737 8483
rect 36771 8480 36783 8483
rect 36817 8483 36875 8489
rect 36817 8480 36829 8483
rect 36771 8452 36829 8480
rect 36771 8449 36783 8452
rect 36725 8443 36783 8449
rect 36817 8449 36829 8452
rect 36863 8449 36875 8483
rect 36817 8443 36875 8449
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37826 8440 37832 8492
rect 37884 8440 37890 8492
rect 38197 8483 38255 8489
rect 38197 8449 38209 8483
rect 38243 8449 38255 8483
rect 38197 8443 38255 8449
rect 29840 8384 30880 8412
rect 30929 8415 30987 8421
rect 30929 8381 30941 8415
rect 30975 8381 30987 8415
rect 30929 8375 30987 8381
rect 30742 8304 30748 8356
rect 30800 8344 30806 8356
rect 30944 8344 30972 8375
rect 31662 8372 31668 8424
rect 31720 8412 31726 8424
rect 37090 8412 37096 8424
rect 31720 8384 37096 8412
rect 31720 8372 31726 8384
rect 37090 8372 37096 8384
rect 37148 8372 37154 8424
rect 37642 8372 37648 8424
rect 37700 8412 37706 8424
rect 38212 8412 38240 8443
rect 38470 8440 38476 8492
rect 38528 8480 38534 8492
rect 38749 8483 38807 8489
rect 38749 8480 38761 8483
rect 38528 8452 38761 8480
rect 38528 8440 38534 8452
rect 38749 8449 38761 8452
rect 38795 8449 38807 8483
rect 38749 8443 38807 8449
rect 38838 8440 38844 8492
rect 38896 8440 38902 8492
rect 38930 8440 38936 8492
rect 38988 8480 38994 8492
rect 39209 8483 39267 8489
rect 39209 8480 39221 8483
rect 38988 8452 39221 8480
rect 38988 8440 38994 8452
rect 39209 8449 39221 8452
rect 39255 8449 39267 8483
rect 39209 8443 39267 8449
rect 37700 8384 38240 8412
rect 37700 8372 37706 8384
rect 30800 8316 30972 8344
rect 31941 8347 31999 8353
rect 30800 8304 30806 8316
rect 31941 8313 31953 8347
rect 31987 8344 31999 8347
rect 32306 8344 32312 8356
rect 31987 8316 32312 8344
rect 31987 8313 31999 8316
rect 31941 8307 31999 8313
rect 32306 8304 32312 8316
rect 32364 8304 32370 8356
rect 38013 8347 38071 8353
rect 32416 8316 37964 8344
rect 32416 8276 32444 8316
rect 29748 8248 32444 8276
rect 34422 8236 34428 8288
rect 34480 8276 34486 8288
rect 37826 8276 37832 8288
rect 34480 8248 37832 8276
rect 34480 8236 34486 8248
rect 37826 8236 37832 8248
rect 37884 8236 37890 8288
rect 37936 8276 37964 8316
rect 38013 8313 38025 8347
rect 38059 8344 38071 8347
rect 38470 8344 38476 8356
rect 38059 8316 38476 8344
rect 38059 8313 38071 8316
rect 38013 8307 38071 8313
rect 38470 8304 38476 8316
rect 38528 8304 38534 8356
rect 39022 8304 39028 8356
rect 39080 8304 39086 8356
rect 38565 8279 38623 8285
rect 38565 8276 38577 8279
rect 37936 8248 38577 8276
rect 38565 8245 38577 8248
rect 38611 8245 38623 8279
rect 38565 8239 38623 8245
rect 1104 8186 39836 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 13950 8186
rect 14002 8134 14014 8186
rect 14066 8134 14078 8186
rect 14130 8134 14142 8186
rect 14194 8134 14206 8186
rect 14258 8134 19950 8186
rect 20002 8134 20014 8186
rect 20066 8134 20078 8186
rect 20130 8134 20142 8186
rect 20194 8134 20206 8186
rect 20258 8134 25950 8186
rect 26002 8134 26014 8186
rect 26066 8134 26078 8186
rect 26130 8134 26142 8186
rect 26194 8134 26206 8186
rect 26258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 37950 8186
rect 38002 8134 38014 8186
rect 38066 8134 38078 8186
rect 38130 8134 38142 8186
rect 38194 8134 38206 8186
rect 38258 8134 39836 8186
rect 1104 8112 39836 8134
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 4522 8072 4528 8084
rect 2731 8044 4528 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 4801 8075 4859 8081
rect 4801 8041 4813 8075
rect 4847 8072 4859 8075
rect 5258 8072 5264 8084
rect 4847 8044 5264 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 10778 8072 10784 8084
rect 5408 8044 10784 8072
rect 5408 8032 5414 8044
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 14277 8075 14335 8081
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14458 8072 14464 8084
rect 14323 8044 14464 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 14752 8044 16620 8072
rect 1394 7964 1400 8016
rect 1452 8004 1458 8016
rect 1452 7976 2636 8004
rect 1452 7964 1458 7976
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1452 7840 1869 7868
rect 1452 7828 1458 7840
rect 1857 7837 1869 7840
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2608 7877 2636 7976
rect 3602 7964 3608 8016
rect 3660 7964 3666 8016
rect 5997 8007 6055 8013
rect 5997 7973 6009 8007
rect 6043 8004 6055 8007
rect 6914 8004 6920 8016
rect 6043 7976 6920 8004
rect 6043 7973 6055 7976
rect 5997 7967 6055 7973
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 8570 8004 8576 8016
rect 8312 7976 8576 8004
rect 3145 7939 3203 7945
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3694 7936 3700 7948
rect 3191 7908 3700 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3694 7896 3700 7908
rect 3752 7896 3758 7948
rect 6362 7896 6368 7948
rect 6420 7896 6426 7948
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7248 7908 7297 7936
rect 7248 7896 7254 7908
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 8312 7936 8340 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 8757 8007 8815 8013
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 8846 8004 8852 8016
rect 8803 7976 8852 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 10318 7964 10324 8016
rect 10376 7964 10382 8016
rect 10686 7964 10692 8016
rect 10744 7964 10750 8016
rect 11793 8007 11851 8013
rect 11793 7973 11805 8007
rect 11839 8004 11851 8007
rect 12529 8007 12587 8013
rect 12529 8004 12541 8007
rect 11839 7976 12541 8004
rect 11839 7973 11851 7976
rect 11793 7967 11851 7973
rect 12529 7973 12541 7976
rect 12575 7973 12587 8007
rect 12529 7967 12587 7973
rect 13538 7964 13544 8016
rect 13596 8004 13602 8016
rect 14752 8004 14780 8044
rect 13596 7976 14780 8004
rect 13596 7964 13602 7976
rect 14826 7964 14832 8016
rect 14884 8004 14890 8016
rect 16592 8004 16620 8044
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 16853 8075 16911 8081
rect 16853 8072 16865 8075
rect 16724 8044 16865 8072
rect 16724 8032 16730 8044
rect 16853 8041 16865 8044
rect 16899 8041 16911 8075
rect 16853 8035 16911 8041
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17000 8044 19334 8072
rect 17000 8032 17006 8044
rect 19306 8004 19334 8044
rect 19610 8032 19616 8084
rect 19668 8032 19674 8084
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20990 8072 20996 8084
rect 20220 8044 20996 8072
rect 20220 8032 20226 8044
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 21634 8072 21640 8084
rect 21100 8044 21640 8072
rect 21100 8004 21128 8044
rect 21634 8032 21640 8044
rect 21692 8072 21698 8084
rect 21692 8044 22324 8072
rect 21692 8032 21698 8044
rect 14884 7976 15792 8004
rect 16592 7976 17080 8004
rect 19306 7976 21128 8004
rect 14884 7964 14890 7976
rect 9953 7939 10011 7945
rect 7285 7899 7343 7905
rect 7852 7908 8340 7936
rect 8404 7908 9168 7936
rect 7852 7880 7880 7908
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2832 7840 2973 7868
rect 2832 7828 2838 7840
rect 2961 7837 2973 7840
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3568 7840 3801 7868
rect 3568 7828 3574 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3789 7831 3847 7837
rect 3896 7840 4077 7868
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 2038 7760 2044 7812
rect 2096 7760 2102 7812
rect 2409 7803 2467 7809
rect 2409 7769 2421 7803
rect 2455 7800 2467 7803
rect 2455 7772 2820 7800
rect 2455 7769 2467 7772
rect 2409 7763 2467 7769
rect 2792 7744 2820 7772
rect 2866 7760 2872 7812
rect 2924 7800 2930 7812
rect 3421 7803 3479 7809
rect 3421 7800 3433 7803
rect 2924 7772 3433 7800
rect 2924 7760 2930 7772
rect 3421 7769 3433 7772
rect 3467 7800 3479 7803
rect 3896 7800 3924 7840
rect 4065 7837 4077 7840
rect 4111 7868 4123 7871
rect 4614 7868 4620 7880
rect 4111 7840 4620 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 4338 7800 4344 7812
rect 3467 7772 3924 7800
rect 4080 7772 4344 7800
rect 3467 7769 3479 7772
rect 3421 7763 3479 7769
rect 1026 7692 1032 7744
rect 1084 7732 1090 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1084 7704 1593 7732
rect 1084 7692 1090 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 1581 7695 1639 7701
rect 2590 7692 2596 7744
rect 2648 7732 2654 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2648 7704 2697 7732
rect 2648 7692 2654 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 4080 7732 4108 7772
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 4890 7760 4896 7812
rect 4948 7800 4954 7812
rect 5000 7800 5028 7831
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5316 7840 5580 7868
rect 5316 7828 5322 7840
rect 5350 7800 5356 7812
rect 4948 7772 5356 7800
rect 4948 7760 4954 7772
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5552 7800 5580 7840
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 5776 7840 7021 7868
rect 5776 7828 5782 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7834 7868 7840 7880
rect 7607 7840 7840 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 6181 7803 6239 7809
rect 6181 7800 6193 7803
rect 5552 7772 6193 7800
rect 6181 7769 6193 7772
rect 6227 7800 6239 7803
rect 6270 7800 6276 7812
rect 6227 7772 6276 7800
rect 6227 7769 6239 7772
rect 6181 7763 6239 7769
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 8404 7800 8432 7908
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 9140 7868 9168 7908
rect 9953 7905 9965 7939
rect 9999 7936 10011 7939
rect 10410 7936 10416 7948
rect 9999 7908 10416 7936
rect 9999 7905 10011 7908
rect 9953 7899 10011 7905
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11756 7908 12081 7936
rect 11756 7896 11762 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 12434 7936 12440 7948
rect 12069 7899 12127 7905
rect 12268 7908 12440 7936
rect 9582 7868 9588 7880
rect 8536 7840 9076 7868
rect 9140 7840 9588 7868
rect 8536 7828 8542 7840
rect 6380 7772 8432 7800
rect 2832 7704 4108 7732
rect 2832 7692 2838 7704
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 6380 7732 6408 7772
rect 8570 7760 8576 7812
rect 8628 7760 8634 7812
rect 4212 7704 6408 7732
rect 4212 7692 4218 7704
rect 7190 7692 7196 7744
rect 7248 7692 7254 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 8260 7704 8309 7732
rect 8260 7692 8266 7704
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8297 7695 8355 7701
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8904 7704 8953 7732
rect 8904 7692 8910 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 9048 7732 9076 7840
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9674 7828 9680 7880
rect 9732 7828 9738 7880
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 9824 7840 10548 7868
rect 9824 7828 9830 7840
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 10134 7800 10140 7812
rect 9548 7772 10140 7800
rect 9548 7760 9554 7772
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 10520 7809 10548 7840
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11330 7868 11336 7880
rect 11103 7840 11336 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 10505 7803 10563 7809
rect 10505 7769 10517 7803
rect 10551 7800 10563 7803
rect 11072 7800 11100 7831
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12268 7868 12296 7908
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12805 7939 12863 7945
rect 12805 7936 12817 7939
rect 12676 7908 12817 7936
rect 12676 7896 12682 7908
rect 12805 7905 12817 7908
rect 12851 7905 12863 7939
rect 12805 7899 12863 7905
rect 13630 7896 13636 7948
rect 13688 7936 13694 7948
rect 15197 7939 15255 7945
rect 15197 7936 15209 7939
rect 13688 7908 15209 7936
rect 13688 7896 13694 7908
rect 15197 7905 15209 7908
rect 15243 7936 15255 7939
rect 15562 7936 15568 7948
rect 15243 7908 15568 7936
rect 15243 7905 15255 7908
rect 15197 7899 15255 7905
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 15654 7896 15660 7948
rect 15712 7896 15718 7948
rect 15764 7936 15792 7976
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15764 7908 15945 7936
rect 15933 7905 15945 7908
rect 15979 7936 15991 7939
rect 16942 7936 16948 7948
rect 15979 7908 16948 7936
rect 15979 7905 15991 7908
rect 15933 7899 15991 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 12986 7877 12992 7880
rect 11940 7840 12296 7868
rect 12943 7871 12992 7877
rect 11940 7828 11946 7840
rect 12943 7837 12955 7871
rect 12989 7837 12992 7871
rect 12943 7831 12992 7837
rect 12986 7828 12992 7831
rect 13044 7828 13050 7880
rect 13078 7828 13084 7880
rect 13136 7828 13142 7880
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13771 7840 14105 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14366 7828 14372 7880
rect 14424 7828 14430 7880
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14918 7868 14924 7880
rect 14516 7840 14924 7868
rect 14516 7828 14522 7840
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 16114 7877 16120 7880
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 16071 7871 16120 7877
rect 16071 7837 16083 7871
rect 16117 7837 16120 7871
rect 16071 7831 16120 7837
rect 15028 7800 15056 7831
rect 16114 7828 16120 7831
rect 16172 7828 16178 7880
rect 16206 7828 16212 7880
rect 16264 7828 16270 7880
rect 17052 7877 17080 7976
rect 21266 7964 21272 8016
rect 21324 8004 21330 8016
rect 21361 8007 21419 8013
rect 21361 8004 21373 8007
rect 21324 7976 21373 8004
rect 21324 7964 21330 7976
rect 21361 7973 21373 7976
rect 21407 7973 21419 8007
rect 22296 8004 22324 8044
rect 22370 8032 22376 8084
rect 22428 8072 22434 8084
rect 22557 8075 22615 8081
rect 22557 8072 22569 8075
rect 22428 8044 22569 8072
rect 22428 8032 22434 8044
rect 22557 8041 22569 8044
rect 22603 8041 22615 8075
rect 24302 8072 24308 8084
rect 22557 8035 22615 8041
rect 22664 8044 24308 8072
rect 22664 8004 22692 8044
rect 24302 8032 24308 8044
rect 24360 8032 24366 8084
rect 25038 8032 25044 8084
rect 25096 8072 25102 8084
rect 26142 8072 26148 8084
rect 25096 8044 26148 8072
rect 25096 8032 25102 8044
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 27249 8075 27307 8081
rect 27249 8041 27261 8075
rect 27295 8072 27307 8075
rect 27338 8072 27344 8084
rect 27295 8044 27344 8072
rect 27295 8041 27307 8044
rect 27249 8035 27307 8041
rect 27338 8032 27344 8044
rect 27396 8032 27402 8084
rect 30742 8072 30748 8084
rect 27448 8044 30748 8072
rect 22296 7976 22692 8004
rect 21361 7967 21419 7973
rect 24118 7964 24124 8016
rect 24176 8004 24182 8016
rect 24176 7976 25176 8004
rect 24176 7964 24182 7976
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 18012 7908 20913 7936
rect 18012 7896 18018 7908
rect 20901 7905 20913 7908
rect 20947 7936 20959 7939
rect 20990 7936 20996 7948
rect 20947 7908 20996 7936
rect 20947 7905 20959 7908
rect 20901 7899 20959 7905
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 21754 7939 21812 7945
rect 21754 7936 21766 7939
rect 21100 7908 21766 7936
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 10551 7772 11100 7800
rect 13556 7772 15056 7800
rect 10551 7769 10563 7772
rect 10505 7763 10563 7769
rect 11974 7732 11980 7744
rect 9048 7704 11980 7732
rect 8941 7695 8999 7701
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 13556 7732 13584 7772
rect 12584 7704 13584 7732
rect 14553 7735 14611 7741
rect 12584 7692 12590 7704
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 16298 7732 16304 7744
rect 14599 7704 16304 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 17052 7732 17080 7831
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 19794 7868 19800 7880
rect 19475 7840 19800 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 20714 7828 20720 7880
rect 20772 7828 20778 7880
rect 21100 7868 21128 7908
rect 21754 7905 21766 7908
rect 21800 7905 21812 7939
rect 24946 7936 24952 7948
rect 21754 7899 21812 7905
rect 24596 7908 24952 7936
rect 20824 7840 21128 7868
rect 17221 7803 17279 7809
rect 17221 7769 17233 7803
rect 17267 7800 17279 7803
rect 17328 7800 17356 7828
rect 17862 7800 17868 7812
rect 17267 7772 17868 7800
rect 17267 7769 17279 7772
rect 17221 7763 17279 7769
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 18248 7772 19334 7800
rect 18248 7732 18276 7772
rect 17052 7704 18276 7732
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18598 7732 18604 7744
rect 18371 7704 18604 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 19306 7732 19334 7772
rect 20254 7760 20260 7812
rect 20312 7800 20318 7812
rect 20824 7800 20852 7840
rect 21634 7828 21640 7880
rect 21692 7828 21698 7880
rect 21910 7828 21916 7880
rect 21968 7828 21974 7880
rect 23382 7828 23388 7880
rect 23440 7828 23446 7880
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7868 23719 7871
rect 23750 7868 23756 7880
rect 23707 7840 23756 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 23750 7828 23756 7840
rect 23808 7828 23814 7880
rect 24026 7828 24032 7880
rect 24084 7828 24090 7880
rect 24486 7828 24492 7880
rect 24544 7868 24550 7880
rect 24596 7877 24624 7908
rect 24946 7896 24952 7908
rect 25004 7896 25010 7948
rect 25038 7896 25044 7948
rect 25096 7896 25102 7948
rect 25148 7936 25176 7976
rect 25498 7964 25504 8016
rect 25556 7964 25562 8016
rect 26878 7964 26884 8016
rect 26936 8004 26942 8016
rect 27448 8004 27476 8044
rect 30742 8032 30748 8044
rect 30800 8072 30806 8084
rect 31570 8072 31576 8084
rect 30800 8044 31576 8072
rect 30800 8032 30806 8044
rect 31570 8032 31576 8044
rect 31628 8032 31634 8084
rect 32122 8032 32128 8084
rect 32180 8072 32186 8084
rect 33321 8075 33379 8081
rect 33321 8072 33333 8075
rect 32180 8044 33333 8072
rect 32180 8032 32186 8044
rect 33321 8041 33333 8044
rect 33367 8041 33379 8075
rect 33321 8035 33379 8041
rect 33962 8032 33968 8084
rect 34020 8072 34026 8084
rect 34422 8072 34428 8084
rect 34020 8044 34428 8072
rect 34020 8032 34026 8044
rect 34422 8032 34428 8044
rect 34480 8032 34486 8084
rect 36170 8032 36176 8084
rect 36228 8072 36234 8084
rect 36265 8075 36323 8081
rect 36265 8072 36277 8075
rect 36228 8044 36277 8072
rect 36228 8032 36234 8044
rect 36265 8041 36277 8044
rect 36311 8041 36323 8075
rect 36265 8035 36323 8041
rect 36814 8032 36820 8084
rect 36872 8032 36878 8084
rect 37642 8032 37648 8084
rect 37700 8032 37706 8084
rect 38286 8032 38292 8084
rect 38344 8032 38350 8084
rect 26936 7976 27476 8004
rect 26936 7964 26942 7976
rect 28166 7964 28172 8016
rect 28224 7964 28230 8016
rect 33229 8007 33287 8013
rect 31036 7976 31892 8004
rect 25406 7936 25412 7948
rect 25148 7908 25412 7936
rect 25406 7896 25412 7908
rect 25464 7936 25470 7948
rect 25894 7939 25952 7945
rect 25894 7936 25906 7939
rect 25464 7908 25906 7936
rect 25464 7896 25470 7908
rect 25894 7905 25906 7908
rect 25940 7905 25952 7939
rect 25894 7899 25952 7905
rect 27338 7896 27344 7948
rect 27396 7936 27402 7948
rect 27525 7939 27583 7945
rect 27525 7936 27537 7939
rect 27396 7908 27537 7936
rect 27396 7896 27402 7908
rect 27525 7905 27537 7908
rect 27571 7905 27583 7939
rect 27525 7899 27583 7905
rect 29086 7896 29092 7948
rect 29144 7936 29150 7948
rect 30282 7936 30288 7948
rect 29144 7908 30288 7936
rect 29144 7896 29150 7908
rect 30282 7896 30288 7908
rect 30340 7936 30346 7948
rect 31036 7936 31064 7976
rect 30340 7908 31064 7936
rect 30340 7896 30346 7908
rect 31294 7896 31300 7948
rect 31352 7896 31358 7948
rect 31754 7896 31760 7948
rect 31812 7896 31818 7948
rect 31864 7936 31892 7976
rect 33229 7973 33241 8007
rect 33275 8004 33287 8007
rect 34146 8004 34152 8016
rect 33275 7976 34152 8004
rect 33275 7973 33287 7976
rect 33229 7967 33287 7973
rect 34146 7964 34152 7976
rect 34204 7964 34210 8016
rect 35802 7964 35808 8016
rect 35860 8004 35866 8016
rect 37093 8007 37151 8013
rect 37093 8004 37105 8007
rect 35860 7976 37105 8004
rect 35860 7964 35866 7976
rect 37093 7973 37105 7976
rect 37139 7973 37151 8007
rect 37093 7967 37151 7973
rect 37921 8007 37979 8013
rect 37921 7973 37933 8007
rect 37967 8004 37979 8007
rect 38378 8004 38384 8016
rect 37967 7976 38384 8004
rect 37967 7973 37979 7976
rect 37921 7967 37979 7973
rect 38378 7964 38384 7976
rect 38436 7964 38442 8016
rect 32150 7939 32208 7945
rect 32150 7936 32162 7939
rect 31864 7908 32162 7936
rect 32150 7905 32162 7908
rect 32196 7905 32208 7939
rect 32150 7899 32208 7905
rect 32306 7896 32312 7948
rect 32364 7896 32370 7948
rect 35820 7908 37780 7936
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24544 7840 24593 7868
rect 24544 7828 24550 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24857 7871 24915 7877
rect 24857 7837 24869 7871
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 20312 7772 20852 7800
rect 20312 7760 20318 7772
rect 23106 7760 23112 7812
rect 23164 7800 23170 7812
rect 24872 7800 24900 7831
rect 25774 7828 25780 7880
rect 25832 7828 25838 7880
rect 26050 7828 26056 7880
rect 26108 7828 26114 7880
rect 26697 7871 26755 7877
rect 26697 7837 26709 7871
rect 26743 7868 26755 7871
rect 26789 7871 26847 7877
rect 26789 7868 26801 7871
rect 26743 7840 26801 7868
rect 26743 7837 26755 7840
rect 26697 7831 26755 7837
rect 26789 7837 26801 7840
rect 26835 7837 26847 7871
rect 26789 7831 26847 7837
rect 27430 7828 27436 7880
rect 27488 7828 27494 7880
rect 27709 7871 27767 7877
rect 27709 7837 27721 7871
rect 27755 7868 27767 7871
rect 27890 7868 27896 7880
rect 27755 7840 27896 7868
rect 27755 7837 27767 7840
rect 27709 7831 27767 7837
rect 27724 7800 27752 7831
rect 27890 7828 27896 7840
rect 27948 7828 27954 7880
rect 28442 7828 28448 7880
rect 28500 7828 28506 7880
rect 28534 7828 28540 7880
rect 28592 7877 28598 7880
rect 28592 7871 28620 7877
rect 28608 7837 28620 7871
rect 28592 7831 28620 7837
rect 28592 7828 28598 7831
rect 28718 7828 28724 7880
rect 28776 7828 28782 7880
rect 29365 7871 29423 7877
rect 29365 7837 29377 7871
rect 29411 7868 29423 7871
rect 29549 7871 29607 7877
rect 29549 7868 29561 7871
rect 29411 7840 29561 7868
rect 29411 7837 29423 7840
rect 29365 7831 29423 7837
rect 29549 7837 29561 7840
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 29917 7871 29975 7877
rect 29917 7837 29929 7871
rect 29963 7868 29975 7871
rect 30098 7868 30104 7880
rect 29963 7840 30104 7868
rect 29963 7837 29975 7840
rect 29917 7831 29975 7837
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 31110 7828 31116 7880
rect 31168 7828 31174 7880
rect 32030 7828 32036 7880
rect 32088 7828 32094 7880
rect 32953 7871 33011 7877
rect 32953 7837 32965 7871
rect 32999 7868 33011 7871
rect 33045 7871 33103 7877
rect 33045 7868 33057 7871
rect 32999 7840 33057 7868
rect 32999 7837 33011 7840
rect 32953 7831 33011 7837
rect 33045 7837 33057 7840
rect 33091 7837 33103 7871
rect 33045 7831 33103 7837
rect 33505 7871 33563 7877
rect 33505 7837 33517 7871
rect 33551 7868 33563 7871
rect 33962 7868 33968 7880
rect 33551 7840 33968 7868
rect 33551 7837 33563 7840
rect 33505 7831 33563 7837
rect 33962 7828 33968 7840
rect 34020 7828 34026 7880
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 35437 7871 35495 7877
rect 35437 7868 35449 7871
rect 34848 7840 35449 7868
rect 34848 7828 34854 7840
rect 35437 7837 35449 7840
rect 35483 7837 35495 7871
rect 35437 7831 35495 7837
rect 35710 7828 35716 7880
rect 35768 7828 35774 7880
rect 35820 7800 35848 7908
rect 36262 7828 36268 7880
rect 36320 7868 36326 7880
rect 36449 7871 36507 7877
rect 36449 7868 36461 7871
rect 36320 7840 36461 7868
rect 36320 7828 36326 7840
rect 36449 7837 36461 7840
rect 36495 7837 36507 7871
rect 36449 7831 36507 7837
rect 37001 7871 37059 7877
rect 37001 7837 37013 7871
rect 37047 7837 37059 7871
rect 37001 7831 37059 7837
rect 37277 7871 37335 7877
rect 37277 7837 37289 7871
rect 37323 7837 37335 7871
rect 37277 7831 37335 7837
rect 23164 7772 24900 7800
rect 26528 7772 27752 7800
rect 32784 7772 35848 7800
rect 23164 7760 23170 7772
rect 22186 7732 22192 7744
rect 19306 7704 22192 7732
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22646 7692 22652 7744
rect 22704 7692 22710 7744
rect 23290 7692 23296 7744
rect 23348 7732 23354 7744
rect 24118 7732 24124 7744
rect 23348 7704 24124 7732
rect 23348 7692 23354 7704
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 24210 7692 24216 7744
rect 24268 7692 24274 7744
rect 24765 7735 24823 7741
rect 24765 7701 24777 7735
rect 24811 7732 24823 7735
rect 25590 7732 25596 7744
rect 24811 7704 25596 7732
rect 24811 7701 24823 7704
rect 24765 7695 24823 7701
rect 25590 7692 25596 7704
rect 25648 7692 25654 7744
rect 25958 7692 25964 7744
rect 26016 7732 26022 7744
rect 26528 7732 26556 7772
rect 32784 7744 32812 7772
rect 26016 7704 26556 7732
rect 26016 7692 26022 7704
rect 26602 7692 26608 7744
rect 26660 7732 26666 7744
rect 26973 7735 27031 7741
rect 26973 7732 26985 7735
rect 26660 7704 26985 7732
rect 26660 7692 26666 7704
rect 26973 7701 26985 7704
rect 27019 7701 27031 7735
rect 26973 7695 27031 7701
rect 29733 7735 29791 7741
rect 29733 7701 29745 7735
rect 29779 7732 29791 7735
rect 29914 7732 29920 7744
rect 29779 7704 29920 7732
rect 29779 7701 29791 7704
rect 29733 7695 29791 7701
rect 29914 7692 29920 7704
rect 29972 7692 29978 7744
rect 30101 7735 30159 7741
rect 30101 7701 30113 7735
rect 30147 7732 30159 7735
rect 31754 7732 31760 7744
rect 30147 7704 31760 7732
rect 30147 7701 30159 7704
rect 30101 7695 30159 7701
rect 31754 7692 31760 7704
rect 31812 7692 31818 7744
rect 32766 7692 32772 7744
rect 32824 7692 32830 7744
rect 33502 7692 33508 7744
rect 33560 7732 33566 7744
rect 34701 7735 34759 7741
rect 34701 7732 34713 7735
rect 33560 7704 34713 7732
rect 33560 7692 33566 7704
rect 34701 7701 34713 7704
rect 34747 7701 34759 7735
rect 34701 7695 34759 7701
rect 34882 7692 34888 7744
rect 34940 7732 34946 7744
rect 37016 7732 37044 7831
rect 37292 7800 37320 7831
rect 37458 7828 37464 7880
rect 37516 7828 37522 7880
rect 37752 7877 37780 7908
rect 37826 7896 37832 7948
rect 37884 7936 37890 7948
rect 37884 7908 38148 7936
rect 37884 7896 37890 7908
rect 38120 7877 38148 7908
rect 38654 7896 38660 7948
rect 38712 7896 38718 7948
rect 37737 7871 37795 7877
rect 37737 7837 37749 7871
rect 37783 7837 37795 7871
rect 37737 7831 37795 7837
rect 38105 7871 38163 7877
rect 38105 7837 38117 7871
rect 38151 7837 38163 7871
rect 38105 7831 38163 7837
rect 38749 7871 38807 7877
rect 38749 7837 38761 7871
rect 38795 7868 38807 7871
rect 38841 7871 38899 7877
rect 38841 7868 38853 7871
rect 38795 7840 38853 7868
rect 38795 7837 38807 7840
rect 38749 7831 38807 7837
rect 38841 7837 38853 7840
rect 38887 7837 38899 7871
rect 38841 7831 38899 7837
rect 39209 7871 39267 7877
rect 39209 7837 39221 7871
rect 39255 7837 39267 7871
rect 39209 7831 39267 7837
rect 37826 7800 37832 7812
rect 37292 7772 37832 7800
rect 37826 7760 37832 7772
rect 37884 7760 37890 7812
rect 38565 7803 38623 7809
rect 38565 7769 38577 7803
rect 38611 7800 38623 7803
rect 39224 7800 39252 7831
rect 38611 7772 39252 7800
rect 38611 7769 38623 7772
rect 38565 7763 38623 7769
rect 34940 7704 37044 7732
rect 34940 7692 34946 7704
rect 37274 7692 37280 7744
rect 37332 7732 37338 7744
rect 38473 7735 38531 7741
rect 38473 7732 38485 7735
rect 37332 7704 38485 7732
rect 37332 7692 37338 7704
rect 38473 7701 38485 7704
rect 38519 7701 38531 7735
rect 38473 7695 38531 7701
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 39025 7735 39083 7741
rect 39025 7732 39037 7735
rect 38988 7704 39037 7732
rect 38988 7692 38994 7704
rect 39025 7701 39037 7704
rect 39071 7701 39083 7735
rect 39025 7695 39083 7701
rect 39390 7692 39396 7744
rect 39448 7692 39454 7744
rect 1104 7642 39836 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 9010 7642
rect 9062 7590 9074 7642
rect 9126 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 15010 7642
rect 15062 7590 15074 7642
rect 15126 7590 15138 7642
rect 15190 7590 15202 7642
rect 15254 7590 15266 7642
rect 15318 7590 21010 7642
rect 21062 7590 21074 7642
rect 21126 7590 21138 7642
rect 21190 7590 21202 7642
rect 21254 7590 21266 7642
rect 21318 7590 27010 7642
rect 27062 7590 27074 7642
rect 27126 7590 27138 7642
rect 27190 7590 27202 7642
rect 27254 7590 27266 7642
rect 27318 7590 33010 7642
rect 33062 7590 33074 7642
rect 33126 7590 33138 7642
rect 33190 7590 33202 7642
rect 33254 7590 33266 7642
rect 33318 7590 39010 7642
rect 39062 7590 39074 7642
rect 39126 7590 39138 7642
rect 39190 7590 39202 7642
rect 39254 7590 39266 7642
rect 39318 7590 39836 7642
rect 1104 7568 39836 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 9766 7528 9772 7540
rect 2547 7500 9772 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 9950 7488 9956 7540
rect 10008 7488 10014 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11790 7528 11796 7540
rect 11112 7500 11796 7528
rect 11112 7488 11118 7500
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 11974 7488 11980 7540
rect 12032 7528 12038 7540
rect 12529 7531 12587 7537
rect 12032 7500 12480 7528
rect 12032 7488 12038 7500
rect 750 7420 756 7472
rect 808 7460 814 7472
rect 4890 7460 4896 7472
rect 808 7432 2360 7460
rect 808 7420 814 7432
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 2332 7401 2360 7432
rect 2608 7432 4896 7460
rect 2608 7401 2636 7432
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1578 7324 1584 7336
rect 1443 7296 1584 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 2608 7324 2636 7355
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3712 7401 3740 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 5810 7420 5816 7472
rect 5868 7420 5874 7472
rect 7374 7420 7380 7472
rect 7432 7420 7438 7472
rect 12342 7460 12348 7472
rect 9324 7432 12348 7460
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 4246 7392 4252 7404
rect 4019 7364 4252 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 4246 7352 4252 7364
rect 4304 7392 4310 7404
rect 4614 7392 4620 7404
rect 4304 7364 4620 7392
rect 4304 7352 4310 7364
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 5736 7364 7205 7392
rect 1820 7296 2636 7324
rect 1820 7284 1826 7296
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 5736 7324 5764 7364
rect 7193 7361 7205 7364
rect 7239 7392 7251 7395
rect 7392 7392 7420 7420
rect 7239 7364 7420 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 8478 7352 8484 7404
rect 8536 7352 8542 7404
rect 8754 7352 8760 7404
rect 8812 7352 8818 7404
rect 4396 7296 5764 7324
rect 4396 7284 4402 7296
rect 7466 7284 7472 7336
rect 7524 7284 7530 7336
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 7742 7284 7748 7336
rect 7800 7284 7806 7336
rect 8202 7284 8208 7336
rect 8260 7284 8266 7336
rect 8619 7327 8677 7333
rect 8619 7293 8631 7327
rect 8665 7324 8677 7327
rect 9324 7324 9352 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 12452 7460 12480 7500
rect 12529 7497 12541 7531
rect 12575 7528 12587 7531
rect 13078 7528 13084 7540
rect 12575 7500 13084 7528
rect 12575 7497 12587 7500
rect 12529 7491 12587 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 14458 7528 14464 7540
rect 14108 7500 14464 7528
rect 14108 7460 14136 7500
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14792 7500 15700 7528
rect 14792 7488 14798 7500
rect 12452 7432 14136 7460
rect 15672 7460 15700 7500
rect 15746 7488 15752 7540
rect 15804 7488 15810 7540
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 17954 7528 17960 7540
rect 16080 7500 17960 7528
rect 16080 7488 16086 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18104 7500 19748 7528
rect 18104 7488 18110 7500
rect 17586 7460 17592 7472
rect 15672 7432 16252 7460
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7392 9459 7395
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9447 7364 9505 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9493 7361 9505 7364
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10042 7392 10048 7404
rect 9907 7364 10048 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10152 7364 10609 7392
rect 8665 7296 9352 7324
rect 8665 7293 8677 7296
rect 8619 7287 8677 7293
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4801 7259 4859 7265
rect 4801 7256 4813 7259
rect 4580 7228 4813 7256
rect 4580 7216 4586 7228
rect 4801 7225 4813 7228
rect 4847 7225 4859 7259
rect 4801 7219 4859 7225
rect 1118 7148 1124 7200
rect 1176 7188 1182 7200
rect 2958 7188 2964 7200
rect 1176 7160 2964 7188
rect 1176 7148 1182 7160
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 4338 7188 4344 7200
rect 3651 7160 4344 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4488 7160 4721 7188
rect 4488 7148 4494 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 5132 7160 6469 7188
rect 5132 7148 5138 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 6457 7151 6515 7157
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 9140 7188 9168 7296
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 10152 7324 10180 7364
rect 10597 7361 10609 7364
rect 10643 7392 10655 7395
rect 10643 7364 10916 7392
rect 10643 7361 10655 7364
rect 10597 7355 10655 7361
rect 9640 7296 10180 7324
rect 10321 7327 10379 7333
rect 9640 7284 9646 7296
rect 10321 7293 10333 7327
rect 10367 7293 10379 7327
rect 10888 7324 10916 7364
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 12452 7392 12572 7396
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 11848 7368 13093 7392
rect 11848 7364 12480 7368
rect 12544 7364 13093 7368
rect 11848 7352 11854 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 15841 7395 15899 7401
rect 15841 7361 15853 7395
rect 15887 7392 15899 7395
rect 16114 7392 16120 7404
rect 15887 7364 16120 7392
rect 15887 7361 15899 7364
rect 15841 7355 15899 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16224 7392 16252 7432
rect 17328 7432 17592 7460
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 16224 7364 17141 7392
rect 17129 7361 17141 7364
rect 17175 7392 17187 7395
rect 17218 7392 17224 7404
rect 17175 7364 17224 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17218 7352 17224 7364
rect 17276 7396 17282 7404
rect 17328 7396 17356 7432
rect 17586 7420 17592 7432
rect 17644 7420 17650 7472
rect 19720 7460 19748 7500
rect 19794 7488 19800 7540
rect 19852 7488 19858 7540
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 21269 7531 21327 7537
rect 19944 7500 21220 7528
rect 19944 7488 19950 7500
rect 20162 7460 20168 7472
rect 19720 7432 20168 7460
rect 20162 7420 20168 7432
rect 20220 7460 20226 7472
rect 21192 7460 21220 7500
rect 21269 7497 21281 7531
rect 21315 7528 21327 7531
rect 21910 7528 21916 7540
rect 21315 7500 21916 7528
rect 21315 7497 21327 7500
rect 21269 7491 21327 7497
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 23385 7531 23443 7537
rect 23385 7497 23397 7531
rect 23431 7528 23443 7531
rect 24026 7528 24032 7540
rect 23431 7500 24032 7528
rect 23431 7497 23443 7500
rect 23385 7491 23443 7497
rect 24026 7488 24032 7500
rect 24084 7488 24090 7540
rect 24118 7488 24124 7540
rect 24176 7528 24182 7540
rect 24176 7500 25084 7528
rect 24176 7488 24182 7500
rect 23290 7460 23296 7472
rect 20220 7432 20576 7460
rect 21192 7432 23296 7460
rect 20220 7420 20226 7432
rect 17276 7368 17356 7396
rect 17276 7352 17282 7368
rect 17402 7352 17408 7404
rect 17460 7392 17466 7404
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17460 7364 17969 7392
rect 17460 7352 17466 7364
rect 17957 7361 17969 7364
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 11054 7324 11060 7336
rect 10888 7296 11060 7324
rect 10321 7287 10379 7293
rect 6604 7160 9168 7188
rect 6604 7148 6610 7160
rect 9674 7148 9680 7200
rect 9732 7148 9738 7200
rect 10336 7188 10364 7287
rect 11054 7284 11060 7296
rect 11112 7284 11118 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7324 14151 7327
rect 14458 7324 14464 7336
rect 14139 7296 14464 7324
rect 14139 7293 14151 7296
rect 14093 7287 14151 7293
rect 10410 7188 10416 7200
rect 10336 7160 10416 7188
rect 10410 7148 10416 7160
rect 10468 7188 10474 7200
rect 10962 7188 10968 7200
rect 10468 7160 10968 7188
rect 10468 7148 10474 7160
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11330 7148 11336 7200
rect 11388 7148 11394 7200
rect 12820 7188 12848 7287
rect 13924 7256 13952 7287
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14550 7284 14556 7336
rect 14608 7284 14614 7336
rect 14918 7284 14924 7336
rect 14976 7333 14982 7336
rect 14976 7327 15004 7333
rect 14992 7324 15004 7327
rect 15286 7324 15292 7336
rect 14992 7296 15292 7324
rect 14992 7293 15004 7296
rect 14976 7287 15004 7293
rect 14976 7284 14982 7287
rect 15286 7284 15292 7296
rect 15344 7324 15350 7336
rect 16022 7324 16028 7336
rect 15344 7296 16028 7324
rect 15344 7284 15350 7296
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16850 7284 16856 7336
rect 16908 7284 16914 7336
rect 17972 7324 18000 7355
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 18874 7352 18880 7404
rect 18932 7352 18938 7404
rect 19150 7352 19156 7404
rect 19208 7352 19214 7404
rect 20438 7392 20444 7404
rect 20272 7364 20444 7392
rect 18230 7324 18236 7336
rect 17972 7296 18236 7324
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 18598 7284 18604 7336
rect 18656 7284 18662 7336
rect 19058 7333 19064 7336
rect 19015 7327 19064 7333
rect 19015 7293 19027 7327
rect 19061 7293 19064 7327
rect 19015 7287 19064 7293
rect 19058 7284 19064 7287
rect 19116 7284 19122 7336
rect 20162 7284 20168 7336
rect 20220 7324 20226 7336
rect 20272 7333 20300 7364
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 20548 7401 20576 7432
rect 23290 7420 23296 7432
rect 23348 7420 23354 7472
rect 25056 7460 25084 7500
rect 25130 7488 25136 7540
rect 25188 7528 25194 7540
rect 25958 7528 25964 7540
rect 25188 7500 25964 7528
rect 25188 7488 25194 7500
rect 25958 7488 25964 7500
rect 26016 7488 26022 7540
rect 26050 7488 26056 7540
rect 26108 7528 26114 7540
rect 26329 7531 26387 7537
rect 26329 7528 26341 7531
rect 26108 7500 26341 7528
rect 26108 7488 26114 7500
rect 26329 7497 26341 7500
rect 26375 7497 26387 7531
rect 26329 7491 26387 7497
rect 26786 7488 26792 7540
rect 26844 7528 26850 7540
rect 28074 7528 28080 7540
rect 26844 7500 28080 7528
rect 26844 7488 26850 7500
rect 28074 7488 28080 7500
rect 28132 7488 28138 7540
rect 28169 7531 28227 7537
rect 28169 7497 28181 7531
rect 28215 7528 28227 7531
rect 28718 7528 28724 7540
rect 28215 7500 28724 7528
rect 28215 7497 28227 7500
rect 28169 7491 28227 7497
rect 28718 7488 28724 7500
rect 28776 7488 28782 7540
rect 28810 7488 28816 7540
rect 28868 7528 28874 7540
rect 28868 7500 30052 7528
rect 28868 7488 28874 7500
rect 30024 7460 30052 7500
rect 30098 7488 30104 7540
rect 30156 7488 30162 7540
rect 33042 7528 33048 7540
rect 30208 7500 33048 7528
rect 30208 7460 30236 7500
rect 33042 7488 33048 7500
rect 33100 7488 33106 7540
rect 33410 7488 33416 7540
rect 33468 7528 33474 7540
rect 33468 7500 33824 7528
rect 33468 7488 33474 7500
rect 25056 7432 28488 7460
rect 30024 7432 30236 7460
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7361 20591 7395
rect 20533 7355 20591 7361
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 25056 7401 25084 7432
rect 22557 7395 22615 7401
rect 22557 7392 22569 7395
rect 20680 7364 22569 7392
rect 20680 7352 20686 7364
rect 22557 7361 22569 7364
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 25130 7352 25136 7404
rect 25188 7392 25194 7404
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 25188 7364 25605 7392
rect 25188 7352 25194 7364
rect 25593 7361 25605 7364
rect 25639 7361 25651 7395
rect 25593 7355 25651 7361
rect 25866 7352 25872 7404
rect 25924 7392 25930 7404
rect 26878 7392 26884 7404
rect 25924 7364 26884 7392
rect 25924 7352 25930 7364
rect 26878 7352 26884 7364
rect 26936 7392 26942 7404
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 26936 7364 27169 7392
rect 26936 7352 26942 7364
rect 27157 7361 27169 7364
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27430 7352 27436 7404
rect 27488 7392 27494 7404
rect 27706 7392 27712 7404
rect 27488 7364 27712 7392
rect 27488 7352 27494 7364
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 27890 7352 27896 7404
rect 27948 7392 27954 7404
rect 28258 7392 28264 7404
rect 27948 7364 28264 7392
rect 27948 7352 27954 7364
rect 28258 7352 28264 7364
rect 28316 7352 28322 7404
rect 28460 7401 28488 7432
rect 30374 7420 30380 7472
rect 30432 7460 30438 7472
rect 30432 7432 30788 7460
rect 30432 7420 30438 7432
rect 28445 7395 28503 7401
rect 28445 7361 28457 7395
rect 28491 7392 28503 7395
rect 28626 7392 28632 7404
rect 28491 7364 28632 7392
rect 28491 7361 28503 7364
rect 28445 7355 28503 7361
rect 28626 7352 28632 7364
rect 28684 7352 28690 7404
rect 29454 7352 29460 7404
rect 29512 7352 29518 7404
rect 30650 7352 30656 7404
rect 30708 7352 30714 7404
rect 30760 7392 30788 7432
rect 31018 7420 31024 7472
rect 31076 7420 31082 7472
rect 31110 7420 31116 7472
rect 31168 7460 31174 7472
rect 33796 7460 33824 7500
rect 33962 7488 33968 7540
rect 34020 7488 34026 7540
rect 34238 7488 34244 7540
rect 34296 7528 34302 7540
rect 37274 7528 37280 7540
rect 34296 7500 37280 7528
rect 34296 7488 34302 7500
rect 37274 7488 37280 7500
rect 37332 7488 37338 7540
rect 37366 7488 37372 7540
rect 37424 7528 37430 7540
rect 37645 7531 37703 7537
rect 37645 7528 37657 7531
rect 37424 7500 37657 7528
rect 37424 7488 37430 7500
rect 37645 7497 37657 7500
rect 37691 7497 37703 7531
rect 37645 7491 37703 7497
rect 38657 7531 38715 7537
rect 38657 7497 38669 7531
rect 38703 7528 38715 7531
rect 38746 7528 38752 7540
rect 38703 7500 38752 7528
rect 38703 7497 38715 7500
rect 38657 7491 38715 7497
rect 38746 7488 38752 7500
rect 38804 7488 38810 7540
rect 31168 7432 32352 7460
rect 33796 7432 34008 7460
rect 31168 7420 31174 7432
rect 31036 7392 31064 7420
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30760 7364 31217 7392
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 31294 7352 31300 7404
rect 31352 7392 31358 7404
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31352 7364 32137 7392
rect 31352 7352 31358 7364
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32324 7392 32352 7432
rect 33980 7404 34008 7432
rect 34330 7420 34336 7472
rect 34388 7460 34394 7472
rect 34388 7432 38148 7460
rect 34388 7420 34394 7432
rect 32324 7364 32536 7392
rect 32125 7355 32183 7361
rect 20257 7327 20315 7333
rect 20257 7324 20269 7327
rect 20220 7296 20269 7324
rect 20220 7284 20226 7296
rect 20257 7293 20269 7296
rect 20303 7293 20315 7327
rect 20257 7287 20315 7293
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 21542 7324 21548 7336
rect 21324 7296 21548 7324
rect 21324 7284 21330 7296
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 22186 7284 22192 7336
rect 22244 7324 22250 7336
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 22244 7296 22293 7324
rect 22244 7284 22250 7296
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 23474 7284 23480 7336
rect 23532 7324 23538 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23532 7296 24041 7324
rect 23532 7284 23538 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 24118 7284 24124 7336
rect 24176 7333 24182 7336
rect 24176 7327 24225 7333
rect 24176 7293 24179 7327
rect 24213 7293 24225 7327
rect 24176 7287 24225 7293
rect 24176 7284 24182 7287
rect 24302 7284 24308 7336
rect 24360 7324 24366 7336
rect 24360 7296 24716 7324
rect 24360 7284 24366 7296
rect 14642 7256 14648 7268
rect 13924 7228 14648 7256
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 16758 7256 16764 7268
rect 15988 7228 16764 7256
rect 15988 7216 15994 7228
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 17788 7228 18736 7256
rect 12894 7188 12900 7200
rect 12820 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7188 12958 7200
rect 13170 7188 13176 7200
rect 12952 7160 13176 7188
rect 12952 7148 12958 7160
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 15102 7188 15108 7200
rect 13863 7160 15108 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 16022 7148 16028 7200
rect 16080 7148 16086 7200
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 17788 7188 17816 7228
rect 16448 7160 17816 7188
rect 17865 7191 17923 7197
rect 16448 7148 16454 7160
rect 17865 7157 17877 7191
rect 17911 7188 17923 7191
rect 18506 7188 18512 7200
rect 17911 7160 18512 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 18708 7188 18736 7228
rect 21174 7216 21180 7268
rect 21232 7256 21238 7268
rect 22094 7256 22100 7268
rect 21232 7228 22100 7256
rect 21232 7216 21238 7228
rect 22094 7216 22100 7228
rect 22152 7216 22158 7268
rect 23293 7259 23351 7265
rect 23293 7225 23305 7259
rect 23339 7256 23351 7259
rect 24581 7259 24639 7265
rect 23339 7228 23704 7256
rect 23339 7225 23351 7228
rect 23293 7219 23351 7225
rect 21266 7188 21272 7200
rect 18708 7160 21272 7188
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 23676 7188 23704 7228
rect 24581 7225 24593 7259
rect 24627 7225 24639 7259
rect 24581 7219 24639 7225
rect 24596 7188 24624 7219
rect 23676 7160 24624 7188
rect 24688 7188 24716 7296
rect 24946 7284 24952 7336
rect 25004 7324 25010 7336
rect 25225 7327 25283 7333
rect 25225 7324 25237 7327
rect 25004 7296 25237 7324
rect 25004 7284 25010 7296
rect 25225 7293 25237 7296
rect 25271 7293 25283 7327
rect 25225 7287 25283 7293
rect 25313 7327 25371 7333
rect 25313 7293 25325 7327
rect 25359 7293 25371 7327
rect 29178 7324 29184 7336
rect 25313 7287 25371 7293
rect 27816 7296 29184 7324
rect 24854 7216 24860 7268
rect 24912 7256 24918 7268
rect 25328 7256 25356 7287
rect 24912 7228 25356 7256
rect 24912 7216 24918 7228
rect 26326 7216 26332 7268
rect 26384 7256 26390 7268
rect 27154 7256 27160 7268
rect 26384 7228 27160 7256
rect 26384 7216 26390 7228
rect 27154 7216 27160 7228
rect 27212 7216 27218 7268
rect 27816 7188 27844 7296
rect 29178 7284 29184 7296
rect 29236 7284 29242 7336
rect 29270 7284 29276 7336
rect 29328 7333 29334 7336
rect 29328 7327 29356 7333
rect 29344 7293 29356 7327
rect 29328 7287 29356 7293
rect 30929 7327 30987 7333
rect 30929 7293 30941 7327
rect 30975 7293 30987 7327
rect 30929 7287 30987 7293
rect 32309 7327 32367 7333
rect 32309 7293 32321 7327
rect 32355 7324 32367 7327
rect 32398 7324 32404 7336
rect 32355 7296 32404 7324
rect 32355 7293 32367 7296
rect 32309 7287 32367 7293
rect 29328 7284 29334 7287
rect 28902 7216 28908 7268
rect 28960 7216 28966 7268
rect 30742 7216 30748 7268
rect 30800 7256 30806 7268
rect 30944 7256 30972 7287
rect 32398 7284 32404 7296
rect 32456 7284 32462 7336
rect 32508 7324 32536 7364
rect 33042 7352 33048 7404
rect 33100 7352 33106 7404
rect 33962 7352 33968 7404
rect 34020 7352 34026 7404
rect 34606 7352 34612 7404
rect 34664 7392 34670 7404
rect 34885 7395 34943 7401
rect 34885 7392 34897 7395
rect 34664 7364 34897 7392
rect 34664 7352 34670 7364
rect 34885 7361 34897 7364
rect 34931 7361 34943 7395
rect 34885 7355 34943 7361
rect 34974 7352 34980 7404
rect 35032 7392 35038 7404
rect 35161 7395 35219 7401
rect 35161 7392 35173 7395
rect 35032 7364 35173 7392
rect 35032 7352 35038 7364
rect 35161 7361 35173 7364
rect 35207 7361 35219 7395
rect 35161 7355 35219 7361
rect 33162 7327 33220 7333
rect 33162 7324 33174 7327
rect 32508 7296 33174 7324
rect 33162 7293 33174 7296
rect 33208 7293 33220 7327
rect 33162 7287 33220 7293
rect 33321 7327 33379 7333
rect 33321 7293 33333 7327
rect 33367 7324 33379 7327
rect 33502 7324 33508 7336
rect 33367 7296 33508 7324
rect 33367 7293 33379 7296
rect 33321 7287 33379 7293
rect 33502 7284 33508 7296
rect 33560 7284 33566 7336
rect 35176 7324 35204 7355
rect 35434 7352 35440 7404
rect 35492 7352 35498 7404
rect 36538 7352 36544 7404
rect 36596 7392 36602 7404
rect 38120 7401 38148 7432
rect 37829 7395 37887 7401
rect 37829 7392 37841 7395
rect 36596 7364 37841 7392
rect 36596 7352 36602 7364
rect 37829 7361 37841 7364
rect 37875 7361 37887 7395
rect 37829 7355 37887 7361
rect 38105 7395 38163 7401
rect 38105 7361 38117 7395
rect 38151 7361 38163 7395
rect 38105 7355 38163 7361
rect 38470 7352 38476 7404
rect 38528 7352 38534 7404
rect 38654 7352 38660 7404
rect 38712 7392 38718 7404
rect 39025 7395 39083 7401
rect 39025 7392 39037 7395
rect 38712 7364 39037 7392
rect 38712 7352 38718 7364
rect 39025 7361 39037 7364
rect 39071 7392 39083 7395
rect 39209 7395 39267 7401
rect 39209 7392 39221 7395
rect 39071 7364 39221 7392
rect 39071 7361 39083 7364
rect 39025 7355 39083 7361
rect 39209 7361 39221 7364
rect 39255 7361 39267 7395
rect 39209 7355 39267 7361
rect 35710 7324 35716 7336
rect 35176 7296 35716 7324
rect 35710 7284 35716 7296
rect 35768 7284 35774 7336
rect 30800 7228 30972 7256
rect 30800 7216 30806 7228
rect 31846 7216 31852 7268
rect 31904 7256 31910 7268
rect 31941 7259 31999 7265
rect 31941 7256 31953 7259
rect 31904 7228 31953 7256
rect 31904 7216 31910 7228
rect 31941 7225 31953 7228
rect 31987 7225 31999 7259
rect 31941 7219 31999 7225
rect 32030 7216 32036 7268
rect 32088 7256 32094 7268
rect 32490 7256 32496 7268
rect 32088 7228 32496 7256
rect 32088 7216 32094 7228
rect 32490 7216 32496 7228
rect 32548 7216 32554 7268
rect 32769 7259 32827 7265
rect 32769 7225 32781 7259
rect 32815 7225 32827 7259
rect 32769 7219 32827 7225
rect 24688 7160 27844 7188
rect 28626 7148 28632 7200
rect 28684 7188 28690 7200
rect 30558 7188 30564 7200
rect 28684 7160 30564 7188
rect 28684 7148 28690 7160
rect 30558 7148 30564 7160
rect 30616 7148 30622 7200
rect 30837 7191 30895 7197
rect 30837 7157 30849 7191
rect 30883 7188 30895 7191
rect 31570 7188 31576 7200
rect 30883 7160 31576 7188
rect 30883 7157 30895 7160
rect 30837 7151 30895 7157
rect 31570 7148 31576 7160
rect 31628 7148 31634 7200
rect 32784 7188 32812 7219
rect 35250 7216 35256 7268
rect 35308 7216 35314 7268
rect 35342 7216 35348 7268
rect 35400 7256 35406 7268
rect 36722 7256 36728 7268
rect 35400 7228 36728 7256
rect 35400 7216 35406 7228
rect 36722 7216 36728 7228
rect 36780 7216 36786 7268
rect 40034 7256 40040 7268
rect 38626 7228 40040 7256
rect 34149 7191 34207 7197
rect 34149 7188 34161 7191
rect 32784 7160 34161 7188
rect 34149 7157 34161 7160
rect 34195 7157 34207 7191
rect 34149 7151 34207 7157
rect 38289 7191 38347 7197
rect 38289 7157 38301 7191
rect 38335 7188 38347 7191
rect 38626 7188 38654 7228
rect 40034 7216 40040 7228
rect 40092 7216 40098 7268
rect 38335 7160 38654 7188
rect 38335 7157 38347 7160
rect 38289 7151 38347 7157
rect 39390 7148 39396 7200
rect 39448 7148 39454 7200
rect 1104 7098 39836 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 13950 7098
rect 14002 7046 14014 7098
rect 14066 7046 14078 7098
rect 14130 7046 14142 7098
rect 14194 7046 14206 7098
rect 14258 7046 19950 7098
rect 20002 7046 20014 7098
rect 20066 7046 20078 7098
rect 20130 7046 20142 7098
rect 20194 7046 20206 7098
rect 20258 7046 25950 7098
rect 26002 7046 26014 7098
rect 26066 7046 26078 7098
rect 26130 7046 26142 7098
rect 26194 7046 26206 7098
rect 26258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 37950 7098
rect 38002 7046 38014 7098
rect 38066 7046 38078 7098
rect 38130 7046 38142 7098
rect 38194 7046 38206 7098
rect 38258 7046 39836 7098
rect 1104 7024 39836 7046
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 2406 6984 2412 6996
rect 2096 6956 2412 6984
rect 2096 6944 2102 6956
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 3605 6987 3663 6993
rect 3605 6984 3617 6987
rect 2740 6956 3617 6984
rect 2740 6944 2746 6956
rect 3605 6953 3617 6956
rect 3651 6953 3663 6987
rect 3605 6947 3663 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 11054 6984 11060 6996
rect 4304 6956 11060 6984
rect 4304 6944 4310 6956
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 13078 6944 13084 6996
rect 13136 6944 13142 6996
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13817 6987 13875 6993
rect 13817 6984 13829 6987
rect 13228 6956 13829 6984
rect 13228 6944 13234 6956
rect 13817 6953 13829 6956
rect 13863 6984 13875 6987
rect 15010 6984 15016 6996
rect 13863 6956 15016 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 15381 6987 15439 6993
rect 15381 6953 15393 6987
rect 15427 6984 15439 6987
rect 15654 6984 15660 6996
rect 15427 6956 15660 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16206 6984 16212 6996
rect 15856 6956 16212 6984
rect 1486 6876 1492 6928
rect 1544 6876 1550 6928
rect 4430 6876 4436 6928
rect 4488 6876 4494 6928
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 7432 6888 7788 6916
rect 7432 6876 7438 6888
rect 1504 6789 1532 6876
rect 1762 6808 1768 6860
rect 1820 6808 1826 6860
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3510 6848 3516 6860
rect 3191 6820 3516 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4396 6820 4997 6848
rect 4396 6808 4402 6820
rect 4985 6817 4997 6820
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5718 6808 5724 6860
rect 5776 6808 5782 6860
rect 6362 6808 6368 6860
rect 6420 6808 6426 6860
rect 6546 6857 6552 6860
rect 6524 6851 6552 6857
rect 6524 6817 6536 6851
rect 6524 6811 6552 6817
rect 6546 6808 6552 6811
rect 6604 6808 6610 6860
rect 6638 6808 6644 6860
rect 6696 6808 6702 6860
rect 6914 6808 6920 6860
rect 6972 6808 6978 6860
rect 7558 6808 7564 6860
rect 7616 6808 7622 6860
rect 7760 6857 7788 6888
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 12768 6888 14136 6916
rect 12768 6876 12774 6888
rect 7745 6851 7803 6857
rect 7745 6817 7757 6851
rect 7791 6817 7803 6851
rect 9217 6851 9275 6857
rect 9217 6848 9229 6851
rect 7745 6811 7803 6817
rect 8312 6820 9229 6848
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2314 6780 2320 6792
rect 2087 6752 2320 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3694 6780 3700 6792
rect 3467 6752 3700 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1854 6712 1860 6724
rect 1719 6684 1860 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 2961 6715 3019 6721
rect 2961 6681 2973 6715
rect 3007 6712 3019 6715
rect 3234 6712 3240 6724
rect 3007 6684 3240 6712
rect 3007 6681 3019 6684
rect 2961 6675 3019 6681
rect 3234 6672 3240 6684
rect 3292 6672 3298 6724
rect 3804 6712 3832 6743
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 4890 6789 4896 6792
rect 4847 6783 4896 6789
rect 4847 6749 4859 6783
rect 4893 6749 4896 6783
rect 4847 6743 4896 6749
rect 4890 6740 4896 6743
rect 4948 6740 4954 6792
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 3712 6684 3832 6712
rect 3712 6656 3740 6684
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2740 6616 2789 6644
rect 2740 6604 2746 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 3694 6604 3700 6656
rect 3752 6604 3758 6656
rect 5626 6604 5632 6656
rect 5684 6604 5690 6656
rect 6546 6604 6552 6656
rect 6604 6644 6610 6656
rect 7392 6644 7420 6743
rect 7760 6712 7788 6811
rect 8018 6740 8024 6792
rect 8076 6740 8082 6792
rect 8312 6780 8340 6820
rect 9217 6817 9229 6820
rect 9263 6817 9275 6851
rect 14108 6848 14136 6888
rect 14182 6876 14188 6928
rect 14240 6916 14246 6928
rect 15473 6919 15531 6925
rect 14240 6888 14412 6916
rect 14240 6876 14246 6888
rect 14384 6857 14412 6888
rect 15473 6885 15485 6919
rect 15519 6916 15531 6919
rect 15856 6916 15884 6956
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 16574 6944 16580 6996
rect 16632 6984 16638 6996
rect 19978 6984 19984 6996
rect 16632 6956 19984 6984
rect 16632 6944 16638 6956
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 20070 6944 20076 6996
rect 20128 6944 20134 6996
rect 20162 6944 20168 6996
rect 20220 6984 20226 6996
rect 24118 6984 24124 6996
rect 20220 6956 24124 6984
rect 20220 6944 20226 6956
rect 24118 6944 24124 6956
rect 24176 6984 24182 6996
rect 28445 6987 28503 6993
rect 24176 6956 28120 6984
rect 24176 6944 24182 6956
rect 15519 6888 15884 6916
rect 15519 6885 15531 6888
rect 15473 6879 15531 6885
rect 17954 6876 17960 6928
rect 18012 6916 18018 6928
rect 20530 6916 20536 6928
rect 18012 6888 20536 6916
rect 18012 6876 18018 6888
rect 20530 6876 20536 6888
rect 20588 6876 20594 6928
rect 20732 6888 21220 6916
rect 14369 6851 14427 6857
rect 9217 6811 9275 6817
rect 10428 6820 10916 6848
rect 8128 6752 8340 6780
rect 8128 6712 8156 6752
rect 8846 6740 8852 6792
rect 8904 6782 8910 6792
rect 8941 6785 8999 6791
rect 8941 6782 8953 6785
rect 8904 6754 8953 6782
rect 8904 6740 8910 6754
rect 8941 6751 8953 6754
rect 8987 6751 8999 6785
rect 8941 6745 8999 6751
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 7760 6684 8156 6712
rect 9033 6715 9091 6721
rect 9033 6681 9045 6715
rect 9079 6712 9091 6715
rect 10428 6712 10456 6820
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 10888 6789 10916 6820
rect 11532 6820 12756 6848
rect 14108 6820 14228 6848
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 10962 6740 10968 6792
rect 11020 6740 11026 6792
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 9079 6684 10456 6712
rect 9079 6681 9091 6684
rect 9033 6675 9091 6681
rect 10594 6672 10600 6724
rect 10652 6672 10658 6724
rect 10686 6672 10692 6724
rect 10744 6672 10750 6724
rect 10778 6672 10784 6724
rect 10836 6712 10842 6724
rect 11532 6712 11560 6820
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11664 6752 12265 6780
rect 11664 6740 11670 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 12342 6740 12348 6792
rect 12400 6740 12406 6792
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12728 6780 12756 6820
rect 12986 6780 12992 6792
rect 12728 6752 12992 6780
rect 12621 6743 12679 6749
rect 10836 6684 11560 6712
rect 12636 6712 12664 6743
rect 12986 6740 12992 6752
rect 13044 6740 13050 6792
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13446 6780 13452 6792
rect 13403 6752 13452 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 13630 6740 13636 6792
rect 13688 6740 13694 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13872 6752 14105 6780
rect 13872 6740 13878 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14200 6780 14228 6820
rect 14369 6817 14381 6851
rect 14415 6817 14427 6851
rect 14369 6811 14427 6817
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16850 6848 16856 6860
rect 16632 6820 16856 6848
rect 16632 6808 16638 6820
rect 16850 6808 16856 6820
rect 16908 6848 16914 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 16908 6820 17141 6848
rect 16908 6808 16914 6820
rect 17129 6817 17141 6820
rect 17175 6848 17187 6851
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 17175 6820 17233 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 20732 6848 20760 6888
rect 17920 6820 20760 6848
rect 17920 6808 17926 6820
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 20864 6820 21097 6848
rect 20864 6808 20870 6820
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 21192 6848 21220 6888
rect 24578 6876 24584 6928
rect 24636 6916 24642 6928
rect 25225 6919 25283 6925
rect 25225 6916 25237 6919
rect 24636 6888 25237 6916
rect 24636 6876 24642 6888
rect 25225 6885 25237 6888
rect 25271 6885 25283 6919
rect 25225 6879 25283 6885
rect 26326 6876 26332 6928
rect 26384 6876 26390 6928
rect 28092 6916 28120 6956
rect 28445 6953 28457 6987
rect 28491 6984 28503 6987
rect 28902 6984 28908 6996
rect 28491 6956 28908 6984
rect 28491 6953 28503 6956
rect 28445 6947 28503 6953
rect 28902 6944 28908 6956
rect 28960 6944 28966 6996
rect 30650 6944 30656 6996
rect 30708 6984 30714 6996
rect 31389 6987 31447 6993
rect 31389 6984 31401 6987
rect 30708 6956 31401 6984
rect 30708 6944 30714 6956
rect 31389 6953 31401 6956
rect 31435 6953 31447 6987
rect 34606 6984 34612 6996
rect 31389 6947 31447 6953
rect 31726 6956 34612 6984
rect 29270 6916 29276 6928
rect 28092 6888 29276 6916
rect 29270 6876 29276 6888
rect 29328 6916 29334 6928
rect 29328 6888 30328 6916
rect 29328 6876 29334 6888
rect 21818 6848 21824 6860
rect 21192 6820 21824 6848
rect 21085 6811 21143 6817
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 14200 6752 14657 6780
rect 14093 6743 14151 6749
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 15562 6780 15568 6792
rect 14976 6752 15568 6780
rect 14976 6740 14982 6752
rect 15562 6740 15568 6752
rect 15620 6740 15626 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6780 16543 6783
rect 16758 6780 16764 6792
rect 16531 6752 16764 6780
rect 16531 6749 16543 6752
rect 16485 6743 16543 6749
rect 12636 6684 13676 6712
rect 10836 6672 10842 6684
rect 6604 6616 7420 6644
rect 8757 6647 8815 6653
rect 6604 6604 6610 6616
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9858 6644 9864 6656
rect 8803 6616 9864 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 10008 6616 10241 6644
rect 10008 6604 10014 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10229 6607 10287 6613
rect 10318 6604 10324 6656
rect 10376 6604 10382 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11514 6644 11520 6656
rect 11020 6616 11520 6644
rect 11020 6604 11026 6616
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 11977 6647 12035 6653
rect 11977 6644 11989 6647
rect 11940 6616 11989 6644
rect 11940 6604 11946 6616
rect 11977 6613 11989 6616
rect 12023 6613 12035 6647
rect 11977 6607 12035 6613
rect 12158 6604 12164 6656
rect 12216 6604 12222 6656
rect 12526 6604 12532 6656
rect 12584 6604 12590 6656
rect 12802 6604 12808 6656
rect 12860 6604 12866 6656
rect 13538 6604 13544 6656
rect 13596 6604 13602 6656
rect 13648 6644 13676 6684
rect 13722 6672 13728 6724
rect 13780 6712 13786 6724
rect 16224 6712 16252 6743
rect 16758 6740 16764 6752
rect 16816 6780 16822 6792
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16816 6752 16957 6780
rect 16816 6740 16822 6752
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 17494 6740 17500 6792
rect 17552 6740 17558 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19116 6752 19441 6780
rect 19116 6740 19122 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19576 6752 19625 6780
rect 19576 6740 19582 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 20346 6780 20352 6792
rect 20303 6752 20352 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 20346 6740 20352 6752
rect 20404 6740 20410 6792
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6780 20499 6783
rect 20530 6780 20536 6792
rect 20487 6752 20536 6780
rect 20487 6749 20499 6752
rect 20441 6743 20499 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20625 6783 20683 6789
rect 20625 6749 20637 6783
rect 20671 6749 20683 6783
rect 20625 6743 20683 6749
rect 13780 6684 16252 6712
rect 13780 6672 13786 6684
rect 16298 6672 16304 6724
rect 16356 6712 16362 6724
rect 17512 6712 17540 6740
rect 19334 6712 19340 6724
rect 16356 6684 17540 6712
rect 18248 6684 19340 6712
rect 16356 6672 16362 6684
rect 14182 6644 14188 6656
rect 13648 6616 14188 6644
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 14277 6647 14335 6653
rect 14277 6613 14289 6647
rect 14323 6644 14335 6647
rect 14826 6644 14832 6656
rect 14323 6616 14832 6644
rect 14323 6613 14335 6616
rect 14277 6607 14335 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 16942 6644 16948 6656
rect 15068 6616 16948 6644
rect 15068 6604 15074 6616
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 18248 6653 18276 6684
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 20162 6672 20168 6724
rect 20220 6712 20226 6724
rect 20640 6712 20668 6743
rect 21358 6740 21364 6792
rect 21416 6740 21422 6792
rect 21450 6740 21456 6792
rect 21508 6789 21514 6792
rect 21508 6783 21536 6789
rect 21524 6749 21536 6783
rect 21508 6743 21536 6749
rect 21508 6740 21514 6743
rect 21634 6740 21640 6792
rect 21692 6740 21698 6792
rect 22281 6783 22339 6789
rect 22281 6749 22293 6783
rect 22327 6780 22339 6783
rect 22373 6783 22431 6789
rect 22373 6780 22385 6783
rect 22327 6752 22385 6780
rect 22327 6749 22339 6752
rect 22281 6743 22339 6749
rect 22373 6749 22385 6752
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 23106 6712 23112 6724
rect 20220 6684 20668 6712
rect 22480 6684 23112 6712
rect 20220 6672 20226 6684
rect 18233 6647 18291 6653
rect 18233 6613 18245 6647
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 19242 6604 19248 6656
rect 19300 6604 19306 6656
rect 19797 6647 19855 6653
rect 19797 6613 19809 6647
rect 19843 6644 19855 6647
rect 22480 6644 22508 6684
rect 23106 6672 23112 6684
rect 23164 6672 23170 6724
rect 23492 6712 23520 6743
rect 23750 6740 23756 6792
rect 23808 6780 23814 6792
rect 24762 6780 24768 6792
rect 23808 6752 24768 6780
rect 23808 6740 23814 6752
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 24854 6740 24860 6792
rect 24912 6780 24918 6792
rect 25130 6780 25136 6792
rect 24912 6752 25136 6780
rect 24912 6740 24918 6752
rect 25130 6740 25136 6752
rect 25188 6740 25194 6792
rect 25866 6780 25872 6792
rect 25332 6752 25872 6780
rect 24026 6712 24032 6724
rect 23492 6684 24032 6712
rect 24026 6672 24032 6684
rect 24084 6712 24090 6724
rect 24486 6712 24492 6724
rect 24084 6684 24492 6712
rect 24084 6672 24090 6684
rect 24486 6672 24492 6684
rect 24544 6672 24550 6724
rect 25332 6712 25360 6752
rect 25866 6740 25872 6752
rect 25924 6740 25930 6792
rect 25958 6740 25964 6792
rect 26016 6740 26022 6792
rect 26234 6740 26240 6792
rect 26292 6740 26298 6792
rect 26344 6789 26372 6876
rect 27154 6808 27160 6860
rect 27212 6848 27218 6860
rect 27433 6851 27491 6857
rect 27433 6848 27445 6851
rect 27212 6820 27445 6848
rect 27212 6808 27218 6820
rect 27433 6817 27445 6820
rect 27479 6817 27491 6851
rect 27433 6811 27491 6817
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6749 26387 6783
rect 26329 6743 26387 6749
rect 26510 6740 26516 6792
rect 26568 6780 26574 6792
rect 26605 6783 26663 6789
rect 26605 6780 26617 6783
rect 26568 6752 26617 6780
rect 26568 6740 26574 6752
rect 26605 6749 26617 6752
rect 26651 6749 26663 6783
rect 26605 6743 26663 6749
rect 26694 6740 26700 6792
rect 26752 6780 26758 6792
rect 27338 6780 27344 6792
rect 26752 6752 27344 6780
rect 26752 6740 26758 6752
rect 27338 6740 27344 6752
rect 27396 6740 27402 6792
rect 27448 6780 27476 6811
rect 28258 6808 28264 6860
rect 28316 6848 28322 6860
rect 29549 6851 29607 6857
rect 29549 6848 29561 6851
rect 28316 6820 29561 6848
rect 28316 6808 28322 6820
rect 29549 6817 29561 6820
rect 29595 6817 29607 6851
rect 29549 6811 29607 6817
rect 30190 6808 30196 6860
rect 30248 6808 30254 6860
rect 30300 6848 30328 6888
rect 31202 6876 31208 6928
rect 31260 6916 31266 6928
rect 31726 6916 31754 6956
rect 34606 6944 34612 6956
rect 34664 6944 34670 6996
rect 37734 6944 37740 6996
rect 37792 6984 37798 6996
rect 38197 6987 38255 6993
rect 38197 6984 38209 6987
rect 37792 6956 38209 6984
rect 37792 6944 37798 6956
rect 38197 6953 38209 6956
rect 38243 6953 38255 6987
rect 38197 6947 38255 6953
rect 31260 6888 31754 6916
rect 31260 6876 31266 6888
rect 30469 6851 30527 6857
rect 30469 6848 30481 6851
rect 30300 6820 30481 6848
rect 30469 6817 30481 6820
rect 30515 6817 30527 6851
rect 30469 6811 30527 6817
rect 30558 6808 30564 6860
rect 30616 6857 30622 6860
rect 30616 6851 30644 6857
rect 30632 6817 30644 6851
rect 30616 6811 30644 6817
rect 30616 6808 30622 6811
rect 38304 6805 38424 6814
rect 38562 6808 38568 6860
rect 38620 6848 38626 6860
rect 38620 6820 39252 6848
rect 38620 6808 38626 6820
rect 38304 6799 38439 6805
rect 38304 6796 38393 6799
rect 27614 6780 27620 6792
rect 27448 6752 27620 6780
rect 27614 6740 27620 6752
rect 27672 6740 27678 6792
rect 27706 6740 27712 6792
rect 27764 6740 27770 6792
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 24964 6684 25360 6712
rect 19843 6616 22508 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 22554 6604 22560 6656
rect 22612 6604 22618 6656
rect 22738 6604 22744 6656
rect 22796 6604 22802 6656
rect 23014 6604 23020 6656
rect 23072 6644 23078 6656
rect 24964 6644 24992 6684
rect 25406 6672 25412 6724
rect 25464 6712 25470 6724
rect 29748 6712 29776 6743
rect 30742 6740 30748 6792
rect 30800 6740 30806 6792
rect 31662 6740 31668 6792
rect 31720 6780 31726 6792
rect 31941 6783 31999 6789
rect 31941 6780 31953 6783
rect 31720 6752 31953 6780
rect 31720 6740 31726 6752
rect 31941 6749 31953 6752
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 25464 6684 29776 6712
rect 31956 6712 31984 6743
rect 32214 6740 32220 6792
rect 32272 6740 32278 6792
rect 33045 6783 33103 6789
rect 33045 6780 33057 6783
rect 32324 6752 33057 6780
rect 32324 6712 32352 6752
rect 33045 6749 33057 6752
rect 33091 6749 33103 6783
rect 33045 6743 33103 6749
rect 33321 6783 33379 6789
rect 33321 6749 33333 6783
rect 33367 6780 33379 6783
rect 33410 6780 33416 6792
rect 33367 6752 33416 6780
rect 33367 6749 33379 6752
rect 33321 6743 33379 6749
rect 33410 6740 33416 6752
rect 33468 6740 33474 6792
rect 34054 6740 34060 6792
rect 34112 6780 34118 6792
rect 34238 6780 34244 6792
rect 34112 6752 34244 6780
rect 34112 6740 34118 6752
rect 34238 6740 34244 6752
rect 34296 6740 34302 6792
rect 34425 6783 34483 6789
rect 34425 6749 34437 6783
rect 34471 6780 34483 6783
rect 34606 6780 34612 6792
rect 34471 6752 34612 6780
rect 34471 6749 34483 6752
rect 34425 6743 34483 6749
rect 34606 6740 34612 6752
rect 34664 6740 34670 6792
rect 34701 6783 34759 6789
rect 34701 6749 34713 6783
rect 34747 6749 34759 6783
rect 34977 6783 35035 6789
rect 34977 6780 34989 6783
rect 34701 6743 34759 6749
rect 34808 6752 34989 6780
rect 31956 6684 32352 6712
rect 25464 6672 25470 6684
rect 23072 6616 24992 6644
rect 25041 6647 25099 6653
rect 23072 6604 23078 6616
rect 25041 6613 25053 6647
rect 25087 6644 25099 6647
rect 25866 6644 25872 6656
rect 25087 6616 25872 6644
rect 25087 6613 25099 6616
rect 25041 6607 25099 6613
rect 25866 6604 25872 6616
rect 25924 6604 25930 6656
rect 27338 6604 27344 6656
rect 27396 6604 27402 6656
rect 27430 6604 27436 6656
rect 27488 6644 27494 6656
rect 28258 6644 28264 6656
rect 27488 6616 28264 6644
rect 27488 6604 27494 6616
rect 28258 6604 28264 6616
rect 28316 6604 28322 6656
rect 29748 6644 29776 6684
rect 32858 6672 32864 6724
rect 32916 6712 32922 6724
rect 32916 6684 34284 6712
rect 32916 6672 32922 6684
rect 32582 6644 32588 6656
rect 29748 6616 32588 6644
rect 32582 6604 32588 6616
rect 32640 6604 32646 6656
rect 32766 6604 32772 6656
rect 32824 6644 32830 6656
rect 32953 6647 33011 6653
rect 32953 6644 32965 6647
rect 32824 6616 32965 6644
rect 32824 6604 32830 6616
rect 32953 6613 32965 6616
rect 32999 6613 33011 6647
rect 32953 6607 33011 6613
rect 33686 6604 33692 6656
rect 33744 6644 33750 6656
rect 34256 6653 34284 6684
rect 34057 6647 34115 6653
rect 34057 6644 34069 6647
rect 33744 6616 34069 6644
rect 33744 6604 33750 6616
rect 34057 6613 34069 6616
rect 34103 6613 34115 6647
rect 34057 6607 34115 6613
rect 34241 6647 34299 6653
rect 34241 6613 34253 6647
rect 34287 6613 34299 6647
rect 34716 6644 34744 6743
rect 34808 6724 34836 6752
rect 34977 6749 34989 6752
rect 35023 6749 35035 6783
rect 34977 6743 35035 6749
rect 35066 6740 35072 6792
rect 35124 6780 35130 6792
rect 35989 6783 36047 6789
rect 35989 6780 36001 6783
rect 35124 6752 36001 6780
rect 35124 6740 35130 6752
rect 35989 6749 36001 6752
rect 36035 6749 36047 6783
rect 35989 6743 36047 6749
rect 37734 6740 37740 6792
rect 37792 6780 37798 6792
rect 37921 6783 37979 6789
rect 37921 6780 37933 6783
rect 37792 6752 37933 6780
rect 37792 6740 37798 6752
rect 37921 6749 37933 6752
rect 37967 6749 37979 6783
rect 37921 6743 37979 6749
rect 38120 6786 38393 6796
rect 38120 6768 38332 6786
rect 34790 6672 34796 6724
rect 34848 6672 34854 6724
rect 35526 6672 35532 6724
rect 35584 6712 35590 6724
rect 38120 6712 38148 6768
rect 38381 6765 38393 6786
rect 38427 6765 38439 6799
rect 38381 6759 38439 6765
rect 38470 6740 38476 6792
rect 38528 6776 38534 6792
rect 39224 6789 39252 6820
rect 38657 6783 38715 6789
rect 38657 6780 38669 6783
rect 38580 6776 38669 6780
rect 38528 6752 38669 6776
rect 38528 6748 38608 6752
rect 38657 6749 38669 6752
rect 38703 6749 38715 6783
rect 38528 6740 38534 6748
rect 38657 6743 38715 6749
rect 38841 6783 38899 6789
rect 38841 6749 38853 6783
rect 38887 6749 38899 6783
rect 38841 6743 38899 6749
rect 39209 6783 39267 6789
rect 39209 6749 39221 6783
rect 39255 6749 39267 6783
rect 39209 6743 39267 6749
rect 38746 6712 38752 6724
rect 35584 6684 38148 6712
rect 38212 6684 38752 6712
rect 35584 6672 35590 6684
rect 35342 6644 35348 6656
rect 34716 6616 35348 6644
rect 34241 6607 34299 6613
rect 35342 6604 35348 6616
rect 35400 6604 35406 6656
rect 35710 6604 35716 6656
rect 35768 6604 35774 6656
rect 35802 6604 35808 6656
rect 35860 6604 35866 6656
rect 38105 6647 38163 6653
rect 38105 6613 38117 6647
rect 38151 6644 38163 6647
rect 38212 6644 38240 6684
rect 38746 6672 38752 6684
rect 38804 6672 38810 6724
rect 38151 6616 38240 6644
rect 38151 6613 38163 6616
rect 38105 6607 38163 6613
rect 38378 6604 38384 6656
rect 38436 6644 38442 6656
rect 38473 6647 38531 6653
rect 38473 6644 38485 6647
rect 38436 6616 38485 6644
rect 38436 6604 38442 6616
rect 38473 6613 38485 6616
rect 38519 6613 38531 6647
rect 38473 6607 38531 6613
rect 38562 6604 38568 6656
rect 38620 6644 38626 6656
rect 38856 6644 38884 6743
rect 39574 6712 39580 6724
rect 39040 6684 39580 6712
rect 39040 6653 39068 6684
rect 39574 6672 39580 6684
rect 39632 6672 39638 6724
rect 38620 6616 38884 6644
rect 39025 6647 39083 6653
rect 38620 6604 38626 6616
rect 39025 6613 39037 6647
rect 39071 6613 39083 6647
rect 39025 6607 39083 6613
rect 39390 6604 39396 6656
rect 39448 6604 39454 6656
rect 1104 6554 39836 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 9010 6554
rect 9062 6502 9074 6554
rect 9126 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 15010 6554
rect 15062 6502 15074 6554
rect 15126 6502 15138 6554
rect 15190 6502 15202 6554
rect 15254 6502 15266 6554
rect 15318 6502 21010 6554
rect 21062 6502 21074 6554
rect 21126 6502 21138 6554
rect 21190 6502 21202 6554
rect 21254 6502 21266 6554
rect 21318 6502 27010 6554
rect 27062 6502 27074 6554
rect 27126 6502 27138 6554
rect 27190 6502 27202 6554
rect 27254 6502 27266 6554
rect 27318 6502 33010 6554
rect 33062 6502 33074 6554
rect 33126 6502 33138 6554
rect 33190 6502 33202 6554
rect 33254 6502 33266 6554
rect 33318 6502 39010 6554
rect 39062 6502 39074 6554
rect 39126 6502 39138 6554
rect 39190 6502 39202 6554
rect 39254 6502 39266 6554
rect 39318 6502 39836 6554
rect 1104 6480 39836 6502
rect 7190 6440 7196 6452
rect 1688 6412 7196 6440
rect 1394 6264 1400 6316
rect 1452 6264 1458 6316
rect 1688 6313 1716 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 9950 6440 9956 6452
rect 9180 6412 9956 6440
rect 9180 6400 9186 6412
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 10686 6440 10692 6452
rect 10459 6412 10692 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 11480 6412 11836 6440
rect 11480 6400 11486 6412
rect 2792 6344 3924 6372
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6273 2375 6307
rect 2792 6304 2820 6344
rect 2317 6267 2375 6273
rect 2516 6276 2820 6304
rect 1210 6196 1216 6248
rect 1268 6236 1274 6248
rect 2332 6236 2360 6267
rect 1268 6208 2360 6236
rect 1268 6196 1274 6208
rect 2516 6177 2544 6276
rect 2866 6264 2872 6316
rect 2924 6264 2930 6316
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 3896 6304 3924 6344
rect 6086 6332 6092 6384
rect 6144 6372 6150 6384
rect 10873 6375 10931 6381
rect 6144 6344 7997 6372
rect 6144 6332 6150 6344
rect 4062 6304 4068 6316
rect 3896 6276 4068 6304
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4798 6313 4804 6316
rect 4755 6307 4804 6313
rect 4755 6273 4767 6307
rect 4801 6273 4804 6307
rect 4755 6267 4804 6273
rect 4798 6264 4804 6267
rect 4856 6264 4862 6316
rect 5626 6264 5632 6316
rect 5684 6264 5690 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6205 2651 6239
rect 3620 6236 3648 6264
rect 2593 6199 2651 6205
rect 3252 6208 3648 6236
rect 2501 6171 2559 6177
rect 2501 6137 2513 6171
rect 2547 6137 2559 6171
rect 2608 6168 2636 6199
rect 2608 6140 2728 6168
rect 2501 6131 2559 6137
rect 2700 6100 2728 6140
rect 3252 6100 3280 6208
rect 3694 6196 3700 6248
rect 3752 6196 3758 6248
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 4430 6236 4436 6248
rect 3927 6208 4436 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4890 6196 4896 6248
rect 4948 6196 4954 6248
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 5920 6236 5948 6267
rect 6730 6264 6736 6316
rect 6788 6264 6794 6316
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 5583 6208 5948 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6840 6236 6868 6267
rect 7098 6264 7104 6316
rect 7156 6264 7162 6316
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7650 6304 7656 6316
rect 7248 6276 7656 6304
rect 7248 6264 7254 6276
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 6696 6208 6868 6236
rect 6696 6196 6702 6208
rect 7374 6196 7380 6248
rect 7432 6196 7438 6248
rect 7969 6236 7997 6344
rect 10873 6341 10885 6375
rect 10919 6372 10931 6375
rect 10962 6372 10968 6384
rect 10919 6344 10968 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9582 6313 9588 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8628 6276 8677 6304
rect 8628 6264 8634 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 9539 6307 9588 6313
rect 9539 6273 9551 6307
rect 9585 6273 9588 6307
rect 9539 6267 9588 6273
rect 9582 6264 9588 6267
rect 9640 6264 9646 6316
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10594 6304 10600 6316
rect 10376 6276 10600 6304
rect 10376 6264 10382 6276
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11422 6304 11428 6316
rect 10827 6276 11428 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 11634 6307 11692 6313
rect 11634 6304 11646 6307
rect 11532 6276 11646 6304
rect 8481 6239 8539 6245
rect 7969 6208 8432 6236
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6168 3663 6171
rect 4341 6171 4399 6177
rect 4341 6168 4353 6171
rect 3651 6140 4353 6168
rect 3651 6137 3663 6140
rect 3605 6131 3663 6137
rect 4341 6137 4353 6140
rect 4387 6137 4399 6171
rect 4341 6131 4399 6137
rect 5813 6171 5871 6177
rect 5813 6137 5825 6171
rect 5859 6168 5871 6171
rect 6362 6168 6368 6180
rect 5859 6140 6368 6168
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 7009 6171 7067 6177
rect 7009 6137 7021 6171
rect 7055 6168 7067 6171
rect 8404 6168 8432 6208
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8754 6236 8760 6248
rect 8527 6208 8760 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 9232 6208 9413 6236
rect 8938 6168 8944 6180
rect 7055 6140 7512 6168
rect 8404 6140 8944 6168
rect 7055 6137 7067 6140
rect 7009 6131 7067 6137
rect 2700 6072 3280 6100
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 3970 6100 3976 6112
rect 3568 6072 3976 6100
rect 3568 6060 3574 6072
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 6089 6103 6147 6109
rect 6089 6069 6101 6103
rect 6135 6100 6147 6103
rect 6178 6100 6184 6112
rect 6135 6072 6184 6100
rect 6135 6069 6147 6072
rect 6089 6063 6147 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6546 6060 6552 6112
rect 6604 6060 6610 6112
rect 7282 6060 7288 6112
rect 7340 6060 7346 6112
rect 7484 6100 7512 6140
rect 8938 6128 8944 6140
rect 8996 6168 9002 6180
rect 9232 6168 9260 6208
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 9674 6196 9680 6248
rect 9732 6196 9738 6248
rect 9858 6196 9864 6248
rect 9916 6236 9922 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 9916 6208 10977 6236
rect 9916 6196 9922 6208
rect 10965 6205 10977 6208
rect 11011 6236 11023 6239
rect 11532 6236 11560 6276
rect 11634 6273 11646 6276
rect 11680 6273 11692 6307
rect 11634 6267 11692 6273
rect 11011 6208 11560 6236
rect 11808 6236 11836 6412
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 12308 6412 12357 6440
rect 12308 6400 12314 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12492 6412 13952 6440
rect 12492 6400 12498 6412
rect 13722 6372 13728 6384
rect 12176 6344 13728 6372
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 11974 6304 11980 6316
rect 11931 6276 11980 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 12176 6313 12204 6344
rect 13722 6332 13728 6344
rect 13780 6372 13786 6384
rect 13780 6344 13860 6372
rect 13780 6332 13786 6344
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 12124 6276 12173 6304
rect 12124 6264 12130 6276
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 13832 6313 13860 6344
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13924 6304 13952 6412
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 15930 6440 15936 6452
rect 14424 6412 15936 6440
rect 14424 6400 14430 6412
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16114 6400 16120 6452
rect 16172 6440 16178 6452
rect 16172 6412 16804 6440
rect 16172 6400 16178 6412
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 13924 6276 14841 6304
rect 13817 6267 13875 6273
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15562 6264 15568 6316
rect 15620 6264 15626 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16531 6276 16681 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16776 6304 16804 6412
rect 16850 6400 16856 6452
rect 16908 6400 16914 6452
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 20990 6440 20996 6452
rect 17000 6412 20996 6440
rect 17000 6400 17006 6412
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 21085 6443 21143 6449
rect 21085 6409 21097 6443
rect 21131 6440 21143 6443
rect 21634 6440 21640 6452
rect 21131 6412 21640 6440
rect 21131 6409 21143 6412
rect 21085 6403 21143 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 23014 6440 23020 6452
rect 21968 6412 23020 6440
rect 21968 6400 21974 6412
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 24854 6400 24860 6452
rect 24912 6400 24918 6452
rect 25958 6400 25964 6452
rect 26016 6440 26022 6452
rect 33410 6440 33416 6452
rect 26016 6412 33416 6440
rect 26016 6400 26022 6412
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 21450 6372 21456 6384
rect 20036 6344 21456 6372
rect 20036 6332 20042 6344
rect 21450 6332 21456 6344
rect 21508 6332 21514 6384
rect 21560 6344 24256 6372
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16776 6276 16957 6304
rect 16669 6267 16727 6273
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17218 6264 17224 6316
rect 17276 6264 17282 6316
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18322 6304 18328 6316
rect 18104 6276 18328 6304
rect 18104 6264 18110 6276
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 19334 6264 19340 6316
rect 19392 6264 19398 6316
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 19904 6276 20361 6304
rect 19904 6248 19932 6276
rect 20349 6273 20361 6276
rect 20395 6304 20407 6307
rect 20395 6276 20668 6304
rect 20395 6273 20407 6276
rect 20349 6267 20407 6273
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11808 6208 12449 6236
rect 11011 6205 11023 6208
rect 10965 6199 11023 6205
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 8996 6140 9260 6168
rect 8996 6128 9002 6140
rect 10686 6128 10692 6180
rect 10744 6168 10750 6180
rect 11054 6168 11060 6180
rect 10744 6140 11060 6168
rect 10744 6128 10750 6140
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 12069 6171 12127 6177
rect 12069 6137 12081 6171
rect 12115 6168 12127 6171
rect 12250 6168 12256 6180
rect 12115 6140 12256 6168
rect 12115 6137 12127 6140
rect 12069 6131 12127 6137
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 12452 6168 12480 6199
rect 13538 6196 13544 6248
rect 13596 6196 13602 6248
rect 14182 6196 14188 6248
rect 14240 6196 14246 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14424 6208 14657 6236
rect 14424 6196 14430 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 14645 6199 14703 6205
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 15194 6236 15200 6248
rect 14792 6208 15200 6236
rect 14792 6196 14798 6208
rect 15194 6196 15200 6208
rect 15252 6236 15258 6248
rect 15682 6239 15740 6245
rect 15682 6236 15694 6239
rect 15252 6208 15694 6236
rect 15252 6196 15258 6208
rect 15682 6205 15694 6208
rect 15728 6205 15740 6239
rect 15682 6199 15740 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16390 6236 16396 6248
rect 15887 6208 16396 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 18138 6196 18144 6248
rect 18196 6196 18202 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 18564 6208 18797 6236
rect 18564 6196 18570 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18932 6208 19073 6236
rect 18932 6196 18938 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 19150 6196 19156 6248
rect 19208 6245 19214 6248
rect 19208 6239 19236 6245
rect 19224 6205 19236 6239
rect 19208 6199 19236 6205
rect 19208 6196 19214 6199
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 19576 6208 19748 6236
rect 19576 6196 19582 6208
rect 14200 6168 14228 6196
rect 12452 6140 12572 6168
rect 14200 6140 14872 6168
rect 7834 6100 7840 6112
rect 7484 6072 7840 6100
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6100 8447 6103
rect 9582 6100 9588 6112
rect 8435 6072 9588 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10321 6103 10379 6109
rect 10321 6100 10333 6103
rect 10100 6072 10333 6100
rect 10100 6060 10106 6072
rect 10321 6069 10333 6072
rect 10367 6069 10379 6103
rect 10321 6063 10379 6069
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 11563 6103 11621 6109
rect 11563 6100 11575 6103
rect 10560 6072 11575 6100
rect 10560 6060 10566 6072
rect 11563 6069 11575 6072
rect 11609 6069 11621 6103
rect 12544 6100 12572 6140
rect 13170 6100 13176 6112
rect 12544 6072 13176 6100
rect 11563 6063 11621 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13449 6103 13507 6109
rect 13449 6069 13461 6103
rect 13495 6100 13507 6103
rect 14458 6100 14464 6112
rect 13495 6072 14464 6100
rect 13495 6069 13507 6072
rect 13449 6063 13507 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14734 6100 14740 6112
rect 14599 6072 14740 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 14844 6100 14872 6140
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 15289 6171 15347 6177
rect 15289 6168 15301 6171
rect 14976 6140 15301 6168
rect 14976 6128 14982 6140
rect 15289 6137 15301 6140
rect 15335 6137 15347 6171
rect 19720 6168 19748 6208
rect 19886 6196 19892 6248
rect 19944 6196 19950 6248
rect 20070 6196 20076 6248
rect 20128 6196 20134 6248
rect 20640 6236 20668 6276
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 21560 6304 21588 6344
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 20772 6276 21588 6304
rect 21652 6276 22201 6304
rect 20772 6264 20778 6276
rect 21652 6236 21680 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 23293 6307 23351 6313
rect 23293 6304 23305 6307
rect 22189 6267 22247 6273
rect 22572 6276 23305 6304
rect 20640 6208 21680 6236
rect 21910 6196 21916 6248
rect 21968 6196 21974 6248
rect 19981 6171 20039 6177
rect 19981 6168 19993 6171
rect 19720 6140 19993 6168
rect 15289 6131 15347 6137
rect 19981 6137 19993 6140
rect 20027 6137 20039 6171
rect 19981 6131 20039 6137
rect 16574 6100 16580 6112
rect 14844 6072 16580 6100
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 17957 6103 18015 6109
rect 17957 6100 17969 6103
rect 17920 6072 17969 6100
rect 17920 6060 17926 6072
rect 17957 6069 17969 6072
rect 18003 6069 18015 6103
rect 17957 6063 18015 6069
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 19150 6100 19156 6112
rect 18196 6072 19156 6100
rect 18196 6060 18202 6072
rect 19150 6060 19156 6072
rect 19208 6100 19214 6112
rect 20714 6100 20720 6112
rect 19208 6072 20720 6100
rect 19208 6060 19214 6072
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 21358 6060 21364 6112
rect 21416 6100 21422 6112
rect 22572 6100 22600 6276
rect 23293 6273 23305 6276
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 23014 6196 23020 6248
rect 23072 6196 23078 6248
rect 24118 6128 24124 6180
rect 24176 6128 24182 6180
rect 21416 6072 22600 6100
rect 21416 6060 21422 6072
rect 22922 6060 22928 6112
rect 22980 6060 22986 6112
rect 23658 6060 23664 6112
rect 23716 6100 23722 6112
rect 24029 6103 24087 6109
rect 24029 6100 24041 6103
rect 23716 6072 24041 6100
rect 23716 6060 23722 6072
rect 24029 6069 24041 6072
rect 24075 6069 24087 6103
rect 24228 6100 24256 6344
rect 24302 6264 24308 6316
rect 24360 6304 24366 6316
rect 24872 6313 24900 6400
rect 26510 6372 26516 6384
rect 26436 6344 26516 6372
rect 24857 6307 24915 6313
rect 24857 6304 24869 6307
rect 24360 6276 24869 6304
rect 24360 6264 24366 6276
rect 24857 6273 24869 6276
rect 24903 6273 24915 6307
rect 24857 6267 24915 6273
rect 24946 6264 24952 6316
rect 25004 6304 25010 6316
rect 25133 6307 25191 6313
rect 25133 6304 25145 6307
rect 25004 6276 25145 6304
rect 25004 6264 25010 6276
rect 25133 6273 25145 6276
rect 25179 6273 25191 6307
rect 25133 6267 25191 6273
rect 25498 6264 25504 6316
rect 25556 6304 25562 6316
rect 25961 6307 26019 6313
rect 25961 6304 25973 6307
rect 25556 6276 25973 6304
rect 25556 6264 25562 6276
rect 25961 6273 25973 6276
rect 26007 6304 26019 6307
rect 26436 6304 26464 6344
rect 26510 6332 26516 6344
rect 26568 6332 26574 6384
rect 26694 6332 26700 6384
rect 26752 6372 26758 6384
rect 27430 6372 27436 6384
rect 26752 6344 27436 6372
rect 26752 6332 26758 6344
rect 27430 6332 27436 6344
rect 27488 6332 27494 6384
rect 27724 6313 27752 6412
rect 28534 6372 28540 6384
rect 28000 6344 28540 6372
rect 26605 6307 26663 6313
rect 26605 6304 26617 6307
rect 26007 6276 26617 6304
rect 26007 6273 26019 6276
rect 25961 6267 26019 6273
rect 26605 6273 26617 6276
rect 26651 6273 26663 6307
rect 26605 6267 26663 6273
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6273 27767 6307
rect 27709 6267 27767 6273
rect 27798 6264 27804 6316
rect 27856 6304 27862 6316
rect 28000 6313 28028 6344
rect 28534 6332 28540 6344
rect 28592 6332 28598 6384
rect 27985 6307 28043 6313
rect 27985 6304 27997 6307
rect 27856 6276 27997 6304
rect 27856 6264 27862 6276
rect 27985 6273 27997 6276
rect 28031 6273 28043 6307
rect 27985 6267 28043 6273
rect 28074 6264 28080 6316
rect 28132 6264 28138 6316
rect 28258 6264 28264 6316
rect 28316 6304 28322 6316
rect 28353 6307 28411 6313
rect 28353 6304 28365 6307
rect 28316 6276 28365 6304
rect 28316 6264 28322 6276
rect 28353 6273 28365 6276
rect 28399 6273 28411 6307
rect 28353 6267 28411 6273
rect 28442 6264 28448 6316
rect 28500 6304 28506 6316
rect 30282 6313 30288 6316
rect 30239 6307 30288 6313
rect 28500 6276 29592 6304
rect 28500 6264 28506 6276
rect 26237 6239 26295 6245
rect 26237 6205 26249 6239
rect 26283 6236 26295 6239
rect 26418 6236 26424 6248
rect 26283 6208 26424 6236
rect 26283 6205 26295 6208
rect 26237 6199 26295 6205
rect 26418 6196 26424 6208
rect 26476 6196 26482 6248
rect 26510 6196 26516 6248
rect 26568 6236 26574 6248
rect 26568 6208 27292 6236
rect 26568 6196 26574 6208
rect 25225 6171 25283 6177
rect 25225 6137 25237 6171
rect 25271 6168 25283 6171
rect 25406 6168 25412 6180
rect 25271 6140 25412 6168
rect 25271 6137 25283 6140
rect 25225 6131 25283 6137
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 27154 6168 27160 6180
rect 26160 6140 27160 6168
rect 25590 6100 25596 6112
rect 24228 6072 25596 6100
rect 24029 6063 24087 6069
rect 25590 6060 25596 6072
rect 25648 6100 25654 6112
rect 26160 6100 26188 6140
rect 27154 6128 27160 6140
rect 27212 6128 27218 6180
rect 25648 6072 26188 6100
rect 26789 6103 26847 6109
rect 25648 6060 25654 6072
rect 26789 6069 26801 6103
rect 26835 6100 26847 6103
rect 26878 6100 26884 6112
rect 26835 6072 26884 6100
rect 26835 6069 26847 6072
rect 26789 6063 26847 6069
rect 26878 6060 26884 6072
rect 26936 6060 26942 6112
rect 26970 6060 26976 6112
rect 27028 6060 27034 6112
rect 27264 6100 27292 6208
rect 29178 6196 29184 6248
rect 29236 6196 29242 6248
rect 29270 6196 29276 6248
rect 29328 6236 29334 6248
rect 29365 6239 29423 6245
rect 29365 6236 29377 6239
rect 29328 6208 29377 6236
rect 29328 6196 29334 6208
rect 29365 6205 29377 6208
rect 29411 6205 29423 6239
rect 29564 6236 29592 6276
rect 30239 6273 30251 6307
rect 30285 6273 30288 6307
rect 30239 6267 30288 6273
rect 30282 6264 30288 6267
rect 30340 6264 30346 6316
rect 30374 6264 30380 6316
rect 30432 6264 30438 6316
rect 31772 6313 31800 6412
rect 33410 6400 33416 6412
rect 33468 6400 33474 6452
rect 34333 6443 34391 6449
rect 34333 6409 34345 6443
rect 34379 6440 34391 6443
rect 35066 6440 35072 6452
rect 34379 6412 35072 6440
rect 34379 6409 34391 6412
rect 34333 6403 34391 6409
rect 35066 6400 35072 6412
rect 35124 6400 35130 6452
rect 35434 6400 35440 6452
rect 35492 6440 35498 6452
rect 35529 6443 35587 6449
rect 35529 6440 35541 6443
rect 35492 6412 35541 6440
rect 35492 6400 35498 6412
rect 35529 6409 35541 6412
rect 35575 6409 35587 6443
rect 35529 6403 35587 6409
rect 35894 6400 35900 6452
rect 35952 6440 35958 6452
rect 35989 6443 36047 6449
rect 35989 6440 36001 6443
rect 35952 6412 36001 6440
rect 35952 6400 35958 6412
rect 35989 6409 36001 6412
rect 36035 6409 36047 6443
rect 35989 6403 36047 6409
rect 37550 6400 37556 6452
rect 37608 6440 37614 6452
rect 38289 6443 38347 6449
rect 38289 6440 38301 6443
rect 37608 6412 38301 6440
rect 37608 6400 37614 6412
rect 38289 6409 38301 6412
rect 38335 6409 38347 6443
rect 38289 6403 38347 6409
rect 39393 6443 39451 6449
rect 39393 6409 39405 6443
rect 39439 6440 39451 6443
rect 39482 6440 39488 6452
rect 39439 6412 39488 6440
rect 39439 6409 39451 6412
rect 39393 6403 39451 6409
rect 39482 6400 39488 6412
rect 39540 6400 39546 6452
rect 35710 6332 35716 6384
rect 35768 6372 35774 6384
rect 35768 6344 36124 6372
rect 35768 6332 35774 6344
rect 31021 6307 31079 6313
rect 31021 6273 31033 6307
rect 31067 6304 31079 6307
rect 31297 6307 31355 6313
rect 31297 6304 31309 6307
rect 31067 6276 31309 6304
rect 31067 6273 31079 6276
rect 31021 6267 31079 6273
rect 31297 6273 31309 6276
rect 31343 6273 31355 6307
rect 31297 6267 31355 6273
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6273 31815 6307
rect 31757 6267 31815 6273
rect 32306 6264 32312 6316
rect 32364 6304 32370 6316
rect 32493 6307 32551 6313
rect 32493 6304 32505 6307
rect 32364 6276 32505 6304
rect 32364 6264 32370 6276
rect 32493 6273 32505 6276
rect 32539 6273 32551 6307
rect 32493 6267 32551 6273
rect 33410 6264 33416 6316
rect 33468 6264 33474 6316
rect 34514 6264 34520 6316
rect 34572 6304 34578 6316
rect 35161 6307 35219 6313
rect 35161 6304 35173 6307
rect 34572 6276 35173 6304
rect 34572 6264 34578 6276
rect 35161 6273 35173 6276
rect 35207 6273 35219 6307
rect 35161 6267 35219 6273
rect 35897 6307 35955 6313
rect 35897 6273 35909 6307
rect 35943 6273 35955 6307
rect 35897 6267 35955 6273
rect 30101 6239 30159 6245
rect 30101 6236 30113 6239
rect 29564 6208 30113 6236
rect 29365 6199 29423 6205
rect 30101 6205 30113 6208
rect 30147 6236 30159 6239
rect 32398 6236 32404 6248
rect 30147 6208 32404 6236
rect 30147 6205 30159 6208
rect 30101 6199 30159 6205
rect 32398 6196 32404 6208
rect 32456 6196 32462 6248
rect 32677 6239 32735 6245
rect 32677 6236 32689 6239
rect 32508 6208 32689 6236
rect 29089 6171 29147 6177
rect 29089 6137 29101 6171
rect 29135 6168 29147 6171
rect 29825 6171 29883 6177
rect 29825 6168 29837 6171
rect 29135 6140 29837 6168
rect 29135 6137 29147 6140
rect 29089 6131 29147 6137
rect 29825 6137 29837 6140
rect 29871 6137 29883 6171
rect 29825 6131 29883 6137
rect 30834 6128 30840 6180
rect 30892 6168 30898 6180
rect 32508 6168 32536 6208
rect 32677 6205 32689 6208
rect 32723 6205 32735 6239
rect 32677 6199 32735 6205
rect 32766 6196 32772 6248
rect 32824 6236 32830 6248
rect 33137 6239 33195 6245
rect 33137 6236 33149 6239
rect 32824 6208 33149 6236
rect 32824 6196 32830 6208
rect 33137 6205 33149 6208
rect 33183 6205 33195 6239
rect 33530 6239 33588 6245
rect 33530 6236 33542 6239
rect 33137 6199 33195 6205
rect 33244 6208 33542 6236
rect 30892 6140 32536 6168
rect 30892 6128 30898 6140
rect 28994 6100 29000 6112
rect 27264 6072 29000 6100
rect 28994 6060 29000 6072
rect 29052 6060 29058 6112
rect 31110 6060 31116 6112
rect 31168 6060 31174 6112
rect 31941 6103 31999 6109
rect 31941 6069 31953 6103
rect 31987 6100 31999 6103
rect 32306 6100 32312 6112
rect 31987 6072 32312 6100
rect 31987 6069 31999 6072
rect 31941 6063 31999 6069
rect 32306 6060 32312 6072
rect 32364 6060 32370 6112
rect 32508 6100 32536 6140
rect 32582 6128 32588 6180
rect 32640 6168 32646 6180
rect 33244 6168 33272 6208
rect 33530 6205 33542 6208
rect 33576 6205 33588 6239
rect 33530 6199 33588 6205
rect 33686 6196 33692 6248
rect 33744 6196 33750 6248
rect 35434 6196 35440 6248
rect 35492 6196 35498 6248
rect 32640 6140 33272 6168
rect 34072 6140 34560 6168
rect 32640 6128 32646 6140
rect 34072 6100 34100 6140
rect 32508 6072 34100 6100
rect 34238 6060 34244 6112
rect 34296 6100 34302 6112
rect 34425 6103 34483 6109
rect 34425 6100 34437 6103
rect 34296 6072 34437 6100
rect 34296 6060 34302 6072
rect 34425 6069 34437 6072
rect 34471 6069 34483 6103
rect 34532 6100 34560 6140
rect 35912 6100 35940 6267
rect 36096 6245 36124 6344
rect 37366 6264 37372 6316
rect 37424 6304 37430 6316
rect 38473 6307 38531 6313
rect 38473 6304 38485 6307
rect 37424 6276 38485 6304
rect 37424 6264 37430 6276
rect 38473 6273 38485 6276
rect 38519 6273 38531 6307
rect 38473 6267 38531 6273
rect 38746 6264 38752 6316
rect 38804 6264 38810 6316
rect 38841 6307 38899 6313
rect 38841 6273 38853 6307
rect 38887 6273 38899 6307
rect 38841 6267 38899 6273
rect 36081 6239 36139 6245
rect 36081 6205 36093 6239
rect 36127 6205 36139 6239
rect 36081 6199 36139 6205
rect 36170 6196 36176 6248
rect 36228 6236 36234 6248
rect 38856 6236 38884 6267
rect 39206 6264 39212 6316
rect 39264 6264 39270 6316
rect 36228 6208 38884 6236
rect 36228 6196 36234 6208
rect 37090 6128 37096 6180
rect 37148 6168 37154 6180
rect 38565 6171 38623 6177
rect 38565 6168 38577 6171
rect 37148 6140 38577 6168
rect 37148 6128 37154 6140
rect 38565 6137 38577 6140
rect 38611 6137 38623 6171
rect 38565 6131 38623 6137
rect 34532 6072 35940 6100
rect 34425 6063 34483 6069
rect 39022 6060 39028 6112
rect 39080 6060 39086 6112
rect 1104 6010 39836 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 13950 6010
rect 14002 5958 14014 6010
rect 14066 5958 14078 6010
rect 14130 5958 14142 6010
rect 14194 5958 14206 6010
rect 14258 5958 19950 6010
rect 20002 5958 20014 6010
rect 20066 5958 20078 6010
rect 20130 5958 20142 6010
rect 20194 5958 20206 6010
rect 20258 5958 25950 6010
rect 26002 5958 26014 6010
rect 26066 5958 26078 6010
rect 26130 5958 26142 6010
rect 26194 5958 26206 6010
rect 26258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 37950 6010
rect 38002 5958 38014 6010
rect 38066 5958 38078 6010
rect 38130 5958 38142 6010
rect 38194 5958 38206 6010
rect 38258 5958 39836 6010
rect 1104 5936 39836 5958
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 4062 5896 4068 5908
rect 3467 5868 4068 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 4890 5896 4896 5908
rect 4847 5868 4896 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 4890 5856 4896 5868
rect 4948 5856 4954 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 6086 5896 6092 5908
rect 5215 5868 6092 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 7098 5896 7104 5908
rect 6411 5868 7104 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 8202 5896 8208 5908
rect 7248 5868 8208 5896
rect 7248 5856 7254 5868
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8720 5868 8769 5896
rect 8720 5856 8726 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 10502 5896 10508 5908
rect 8757 5859 8815 5865
rect 9048 5868 10508 5896
rect 1673 5831 1731 5837
rect 1673 5797 1685 5831
rect 1719 5828 1731 5831
rect 1762 5828 1768 5840
rect 1719 5800 1768 5828
rect 1719 5797 1731 5800
rect 1673 5791 1731 5797
rect 1762 5788 1768 5800
rect 1820 5788 1826 5840
rect 2041 5831 2099 5837
rect 2041 5797 2053 5831
rect 2087 5828 2099 5831
rect 2498 5828 2504 5840
rect 2087 5800 2504 5828
rect 2087 5797 2099 5800
rect 2041 5791 2099 5797
rect 2498 5788 2504 5800
rect 2556 5788 2562 5840
rect 2774 5788 2780 5840
rect 2832 5788 2838 5840
rect 3142 5788 3148 5840
rect 3200 5788 3206 5840
rect 6273 5831 6331 5837
rect 6273 5797 6285 5831
rect 6319 5797 6331 5831
rect 6273 5791 6331 5797
rect 2958 5720 2964 5772
rect 3016 5760 3022 5772
rect 3016 5732 3556 5760
rect 3016 5720 3022 5732
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1857 5695 1915 5701
rect 1857 5692 1869 5695
rect 1452 5664 1869 5692
rect 1452 5652 1458 5664
rect 1857 5661 1869 5664
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3528 5692 3556 5732
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 3660 5732 3801 5760
rect 3660 5720 3666 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 3789 5723 3847 5729
rect 5902 5720 5908 5772
rect 5960 5720 5966 5772
rect 6288 5760 6316 5791
rect 8570 5788 8576 5840
rect 8628 5788 8634 5840
rect 7009 5763 7067 5769
rect 7009 5760 7021 5763
rect 6288 5732 7021 5760
rect 7009 5729 7021 5732
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 7168 5763 7226 5769
rect 7168 5729 7180 5763
rect 7214 5760 7226 5763
rect 7466 5760 7472 5772
rect 7214 5732 7472 5760
rect 7214 5729 7226 5732
rect 7168 5723 7226 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 7558 5720 7564 5772
rect 7616 5720 7622 5772
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8588 5760 8616 5788
rect 9048 5769 9076 5868
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 11422 5856 11428 5908
rect 11480 5856 11486 5908
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 15933 5899 15991 5905
rect 11848 5868 14320 5896
rect 11848 5856 11854 5868
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 10134 5828 10140 5840
rect 9539 5800 10140 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 11238 5788 11244 5840
rect 11296 5788 11302 5840
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 12161 5831 12219 5837
rect 12161 5828 12173 5831
rect 11388 5800 12173 5828
rect 11388 5788 11394 5800
rect 12161 5797 12173 5800
rect 12207 5797 12219 5831
rect 13633 5831 13691 5837
rect 13633 5828 13645 5831
rect 12161 5791 12219 5797
rect 13096 5800 13645 5828
rect 8067 5732 8616 5760
rect 9033 5763 9091 5769
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 9033 5729 9045 5763
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 9398 5760 9404 5772
rect 9171 5732 9404 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 9674 5760 9680 5772
rect 9508 5732 9680 5760
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 2639 5664 3464 5692
rect 3528 5664 4077 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 1670 5624 1676 5636
rect 1535 5596 1676 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 1670 5584 1676 5596
rect 1728 5584 1734 5636
rect 2222 5584 2228 5636
rect 2280 5584 2286 5636
rect 2409 5627 2467 5633
rect 2409 5593 2421 5627
rect 2455 5624 2467 5627
rect 2682 5624 2688 5636
rect 2455 5596 2688 5624
rect 2455 5593 2467 5596
rect 2409 5587 2467 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 2958 5624 2964 5636
rect 2792 5596 2964 5624
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 2792 5556 2820 5596
rect 2958 5584 2964 5596
rect 3016 5584 3022 5636
rect 3329 5627 3387 5633
rect 3329 5593 3341 5627
rect 3375 5593 3387 5627
rect 3436 5624 3464 5664
rect 4065 5661 4077 5664
rect 4111 5692 4123 5695
rect 4111 5664 4936 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4908 5624 4936 5664
rect 4982 5652 4988 5704
rect 5040 5652 5046 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5692 5595 5695
rect 5626 5692 5632 5704
rect 5583 5664 5632 5692
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 5626 5652 5632 5664
rect 5684 5692 5690 5704
rect 5920 5692 5948 5720
rect 9508 5704 9536 5732
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10229 5763 10287 5769
rect 10229 5760 10241 5763
rect 10008 5732 10241 5760
rect 10008 5720 10014 5732
rect 10229 5729 10241 5732
rect 10275 5729 10287 5763
rect 10229 5723 10287 5729
rect 10502 5720 10508 5772
rect 10560 5720 10566 5772
rect 10643 5763 10701 5769
rect 10643 5729 10655 5763
rect 10689 5760 10701 5763
rect 11256 5760 11284 5788
rect 13096 5772 13124 5800
rect 13633 5797 13645 5800
rect 13679 5797 13691 5831
rect 13633 5791 13691 5797
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 11790 5760 11796 5772
rect 10689 5732 11796 5760
rect 10689 5729 10701 5732
rect 10643 5723 10701 5729
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 11940 5732 12725 5760
rect 11940 5720 11946 5732
rect 12713 5729 12725 5732
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 13078 5720 13084 5772
rect 13136 5720 13142 5772
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 13740 5760 13768 5791
rect 14292 5769 14320 5868
rect 14384 5868 15884 5896
rect 14277 5763 14335 5769
rect 13412 5732 13768 5760
rect 13832 5732 14228 5760
rect 13412 5720 13418 5732
rect 5684 5664 5948 5692
rect 5684 5652 5690 5664
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8478 5692 8484 5704
rect 8343 5664 8484 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9309 5695 9367 5701
rect 9309 5692 9321 5695
rect 8904 5664 9321 5692
rect 8904 5652 8910 5664
rect 9309 5661 9321 5664
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 5902 5624 5908 5636
rect 3436 5596 4108 5624
rect 4908 5596 5908 5624
rect 3329 5587 3387 5593
rect 2648 5528 2820 5556
rect 2648 5516 2654 5528
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3344 5556 3372 5587
rect 4080 5568 4108 5596
rect 5902 5584 5908 5596
rect 5960 5584 5966 5636
rect 8220 5624 8248 5652
rect 8220 5596 8800 5624
rect 2924 5528 3372 5556
rect 2924 5516 2930 5528
rect 4062 5516 4068 5568
rect 4120 5516 4126 5568
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 5534 5556 5540 5568
rect 5132 5528 5540 5556
rect 5132 5516 5138 5528
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7282 5556 7288 5568
rect 6604 5528 7288 5556
rect 6604 5516 6610 5528
rect 7282 5516 7288 5528
rect 7340 5556 7346 5568
rect 8386 5556 8392 5568
rect 7340 5528 8392 5556
rect 7340 5516 7346 5528
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 8662 5556 8668 5568
rect 8527 5528 8668 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 8772 5556 8800 5596
rect 9490 5556 9496 5568
rect 8772 5528 9496 5556
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 9600 5556 9628 5655
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 11716 5624 11744 5655
rect 12434 5652 12440 5704
rect 12492 5652 12498 5704
rect 12526 5652 12532 5704
rect 12584 5701 12590 5704
rect 12584 5695 12612 5701
rect 12600 5661 12612 5695
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 12584 5655 12612 5661
rect 13372 5664 13461 5692
rect 12584 5652 12590 5655
rect 13372 5633 13400 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 11388 5596 11744 5624
rect 13357 5627 13415 5633
rect 11388 5584 11394 5596
rect 13357 5593 13369 5627
rect 13403 5593 13415 5627
rect 13357 5587 13415 5593
rect 10134 5556 10140 5568
rect 9600 5528 10140 5556
rect 10134 5516 10140 5528
rect 10192 5556 10198 5568
rect 11348 5556 11376 5584
rect 10192 5528 11376 5556
rect 10192 5516 10198 5528
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 13832 5556 13860 5732
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14200 5692 14228 5732
rect 14277 5729 14289 5763
rect 14323 5729 14335 5763
rect 14277 5723 14335 5729
rect 14384 5692 14412 5868
rect 14458 5788 14464 5840
rect 14516 5828 14522 5840
rect 14826 5828 14832 5840
rect 14516 5800 14832 5828
rect 14516 5788 14522 5800
rect 14826 5788 14832 5800
rect 14884 5788 14890 5840
rect 14734 5720 14740 5772
rect 14792 5720 14798 5772
rect 15010 5720 15016 5772
rect 15068 5720 15074 5772
rect 15194 5769 15200 5772
rect 15151 5763 15200 5769
rect 15151 5729 15163 5763
rect 15197 5729 15200 5763
rect 15151 5723 15200 5729
rect 15194 5720 15200 5723
rect 15252 5720 15258 5772
rect 14200 5664 14412 5692
rect 14093 5655 14151 5661
rect 12492 5528 13860 5556
rect 13924 5556 13952 5655
rect 14108 5624 14136 5655
rect 15286 5652 15292 5704
rect 15344 5652 15350 5704
rect 14274 5624 14280 5636
rect 14108 5596 14280 5624
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 15856 5624 15884 5868
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 16206 5896 16212 5908
rect 15979 5868 16212 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 16758 5856 16764 5908
rect 16816 5896 16822 5908
rect 16816 5868 18828 5896
rect 16816 5856 16822 5868
rect 17129 5831 17187 5837
rect 17129 5797 17141 5831
rect 17175 5797 17187 5831
rect 17129 5791 17187 5797
rect 17144 5760 17172 5791
rect 17862 5788 17868 5840
rect 17920 5788 17926 5840
rect 18417 5763 18475 5769
rect 18417 5760 18429 5763
rect 17144 5732 18429 5760
rect 18417 5729 18429 5732
rect 18463 5729 18475 5763
rect 18800 5760 18828 5868
rect 19058 5856 19064 5908
rect 19116 5856 19122 5908
rect 19334 5856 19340 5908
rect 19392 5896 19398 5908
rect 20530 5896 20536 5908
rect 19392 5868 20536 5896
rect 19392 5856 19398 5868
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 21085 5899 21143 5905
rect 21085 5896 21097 5899
rect 20864 5868 21097 5896
rect 20864 5856 20870 5868
rect 21085 5865 21097 5868
rect 21131 5865 21143 5899
rect 26970 5896 26976 5908
rect 21085 5859 21143 5865
rect 22296 5868 25937 5896
rect 20898 5788 20904 5840
rect 20956 5828 20962 5840
rect 21177 5831 21235 5837
rect 21177 5828 21189 5831
rect 20956 5800 21189 5828
rect 20956 5788 20962 5800
rect 21177 5797 21189 5800
rect 21223 5797 21235 5831
rect 22186 5828 22192 5840
rect 21177 5791 21235 5797
rect 21284 5800 22192 5828
rect 19702 5760 19708 5772
rect 18800 5732 19708 5760
rect 18417 5723 18475 5729
rect 19702 5720 19708 5732
rect 19760 5760 19766 5772
rect 20073 5763 20131 5769
rect 20073 5760 20085 5763
rect 19760 5732 20085 5760
rect 19760 5720 19766 5732
rect 20073 5729 20085 5732
rect 20119 5729 20131 5763
rect 20073 5723 20131 5729
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 21284 5760 21312 5800
rect 22186 5788 22192 5800
rect 22244 5788 22250 5840
rect 21048 5732 21312 5760
rect 21048 5720 21054 5732
rect 16114 5652 16120 5704
rect 16172 5652 16178 5704
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 16356 5664 16405 5692
rect 16356 5652 16362 5664
rect 16393 5661 16405 5664
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 17218 5652 17224 5704
rect 17276 5652 17282 5704
rect 17402 5652 17408 5704
rect 17460 5652 17466 5704
rect 18138 5652 18144 5704
rect 18196 5652 18202 5704
rect 18230 5652 18236 5704
rect 18288 5701 18294 5704
rect 18288 5695 18316 5701
rect 18304 5661 18316 5695
rect 18288 5655 18316 5661
rect 18288 5652 18294 5655
rect 19242 5652 19248 5704
rect 19300 5652 19306 5704
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 20349 5695 20407 5701
rect 20349 5661 20361 5695
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 17420 5624 17448 5652
rect 19610 5624 19616 5636
rect 15856 5596 17448 5624
rect 18892 5596 19616 5624
rect 14734 5556 14740 5568
rect 13924 5528 14740 5556
rect 12492 5516 12498 5528
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 14826 5516 14832 5568
rect 14884 5556 14890 5568
rect 15286 5556 15292 5568
rect 14884 5528 15292 5556
rect 14884 5516 14890 5528
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 18892 5556 18920 5596
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 19812 5624 19840 5655
rect 20070 5624 20076 5636
rect 19812 5596 20076 5624
rect 20070 5584 20076 5596
rect 20128 5584 20134 5636
rect 20364 5624 20392 5655
rect 20438 5652 20444 5704
rect 20496 5692 20502 5704
rect 20496 5664 21312 5692
rect 20496 5652 20502 5664
rect 21174 5624 21180 5636
rect 20364 5596 21180 5624
rect 21174 5584 21180 5596
rect 21232 5584 21238 5636
rect 21284 5624 21312 5664
rect 21358 5652 21364 5704
rect 21416 5652 21422 5704
rect 21450 5652 21456 5704
rect 21508 5652 21514 5704
rect 21542 5652 21548 5704
rect 21600 5692 21606 5704
rect 22296 5692 22324 5868
rect 22370 5788 22376 5840
rect 22428 5828 22434 5840
rect 22428 5800 22600 5828
rect 22428 5788 22434 5800
rect 22572 5769 22600 5800
rect 22922 5788 22928 5840
rect 22980 5828 22986 5840
rect 23017 5831 23075 5837
rect 23017 5828 23029 5831
rect 22980 5800 23029 5828
rect 22980 5788 22986 5800
rect 23017 5797 23029 5800
rect 23063 5797 23075 5831
rect 25909 5828 25937 5868
rect 26620 5868 26976 5896
rect 26510 5828 26516 5840
rect 25909 5800 26004 5828
rect 23017 5791 23075 5797
rect 22557 5763 22615 5769
rect 22557 5729 22569 5763
rect 22603 5729 22615 5763
rect 22557 5723 22615 5729
rect 23290 5720 23296 5772
rect 23348 5720 23354 5772
rect 23566 5760 23572 5772
rect 23527 5732 23572 5760
rect 23566 5720 23572 5732
rect 23624 5720 23630 5772
rect 25976 5769 26004 5800
rect 26160 5800 26516 5828
rect 26160 5772 26188 5800
rect 26510 5788 26516 5800
rect 26568 5788 26574 5840
rect 26620 5837 26648 5868
rect 26970 5856 26976 5868
rect 27028 5856 27034 5908
rect 27154 5856 27160 5908
rect 27212 5896 27218 5908
rect 28905 5899 28963 5905
rect 27212 5868 28580 5896
rect 27212 5856 27218 5868
rect 26605 5831 26663 5837
rect 26605 5797 26617 5831
rect 26651 5797 26663 5831
rect 26605 5791 26663 5797
rect 27614 5788 27620 5840
rect 27672 5828 27678 5840
rect 27801 5831 27859 5837
rect 27801 5828 27813 5831
rect 27672 5800 27813 5828
rect 27672 5788 27678 5800
rect 27801 5797 27813 5800
rect 27847 5797 27859 5831
rect 28552 5828 28580 5868
rect 28905 5865 28917 5899
rect 28951 5896 28963 5899
rect 30374 5896 30380 5908
rect 28951 5868 30380 5896
rect 28951 5865 28963 5868
rect 28905 5859 28963 5865
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 30561 5899 30619 5905
rect 30561 5865 30573 5899
rect 30607 5896 30619 5899
rect 30742 5896 30748 5908
rect 30607 5868 30748 5896
rect 30607 5865 30619 5868
rect 30561 5859 30619 5865
rect 30742 5856 30748 5868
rect 30800 5856 30806 5908
rect 34698 5856 34704 5908
rect 34756 5896 34762 5908
rect 35066 5896 35072 5908
rect 34756 5868 35072 5896
rect 34756 5856 34762 5868
rect 35066 5856 35072 5868
rect 35124 5856 35130 5908
rect 35158 5856 35164 5908
rect 35216 5896 35222 5908
rect 38381 5899 38439 5905
rect 38381 5896 38393 5899
rect 35216 5868 38393 5896
rect 35216 5856 35222 5868
rect 38381 5865 38393 5868
rect 38427 5865 38439 5899
rect 38381 5859 38439 5865
rect 39390 5856 39396 5908
rect 39448 5856 39454 5908
rect 29454 5828 29460 5840
rect 28552 5800 29460 5828
rect 27801 5791 27859 5797
rect 29454 5788 29460 5800
rect 29512 5788 29518 5840
rect 31665 5831 31723 5837
rect 31665 5797 31677 5831
rect 31711 5797 31723 5831
rect 31665 5791 31723 5797
rect 32309 5831 32367 5837
rect 32309 5797 32321 5831
rect 32355 5828 32367 5831
rect 32858 5828 32864 5840
rect 32355 5800 32864 5828
rect 32355 5797 32367 5800
rect 32309 5791 32367 5797
rect 25869 5763 25927 5769
rect 25869 5760 25881 5763
rect 25056 5732 25881 5760
rect 25056 5704 25084 5732
rect 25869 5729 25881 5732
rect 25915 5729 25927 5763
rect 25869 5723 25927 5729
rect 25961 5763 26019 5769
rect 25961 5729 25973 5763
rect 26007 5729 26019 5763
rect 25961 5723 26019 5729
rect 26142 5720 26148 5772
rect 26200 5720 26206 5772
rect 26694 5760 26700 5772
rect 26252 5732 26700 5760
rect 23474 5701 23480 5704
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 21600 5664 22385 5692
rect 21600 5652 21606 5664
rect 22373 5661 22385 5664
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 23431 5695 23480 5701
rect 23431 5661 23443 5695
rect 23477 5661 23480 5695
rect 23431 5655 23480 5661
rect 23446 5654 23480 5655
rect 23474 5652 23480 5654
rect 23532 5652 23538 5704
rect 24213 5695 24271 5701
rect 24213 5661 24225 5695
rect 24259 5692 24271 5695
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 24259 5664 24409 5692
rect 24259 5661 24271 5664
rect 24213 5655 24271 5661
rect 24397 5661 24409 5664
rect 24443 5661 24455 5695
rect 24397 5655 24455 5661
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5688 25007 5695
rect 25038 5688 25044 5704
rect 24995 5661 25044 5688
rect 24949 5660 25044 5661
rect 24949 5655 25007 5660
rect 25038 5652 25044 5660
rect 25096 5652 25102 5704
rect 25590 5652 25596 5704
rect 25648 5652 25654 5704
rect 26252 5692 26280 5732
rect 26694 5720 26700 5732
rect 26752 5760 26758 5772
rect 27062 5769 27068 5772
rect 26881 5763 26939 5769
rect 26881 5760 26893 5763
rect 26752 5732 26893 5760
rect 26752 5720 26758 5732
rect 26881 5729 26893 5732
rect 26927 5729 26939 5763
rect 26881 5723 26939 5729
rect 27019 5763 27068 5769
rect 27019 5729 27031 5763
rect 27065 5729 27068 5763
rect 27019 5723 27068 5729
rect 27062 5720 27068 5723
rect 27120 5720 27126 5772
rect 27157 5763 27215 5769
rect 27157 5729 27169 5763
rect 27203 5760 27215 5763
rect 27338 5760 27344 5772
rect 27203 5732 27344 5760
rect 27203 5729 27215 5732
rect 27157 5723 27215 5729
rect 27338 5720 27344 5732
rect 27396 5720 27402 5772
rect 27890 5720 27896 5772
rect 27948 5720 27954 5772
rect 29273 5763 29331 5769
rect 29273 5729 29285 5763
rect 29319 5760 29331 5763
rect 29549 5763 29607 5769
rect 29549 5760 29561 5763
rect 29319 5732 29561 5760
rect 29319 5729 29331 5732
rect 29273 5723 29331 5729
rect 29549 5729 29561 5732
rect 29595 5729 29607 5763
rect 31680 5760 31708 5791
rect 32858 5788 32864 5800
rect 32916 5788 32922 5840
rect 33870 5788 33876 5840
rect 33928 5828 33934 5840
rect 35710 5828 35716 5840
rect 33928 5800 35716 5828
rect 33928 5788 33934 5800
rect 35710 5788 35716 5800
rect 35768 5788 35774 5840
rect 36725 5831 36783 5837
rect 36725 5797 36737 5831
rect 36771 5828 36783 5831
rect 38930 5828 38936 5840
rect 36771 5800 38936 5828
rect 36771 5797 36783 5800
rect 36725 5791 36783 5797
rect 38930 5788 38936 5800
rect 38988 5788 38994 5840
rect 39025 5831 39083 5837
rect 39025 5797 39037 5831
rect 39071 5828 39083 5831
rect 39942 5828 39948 5840
rect 39071 5800 39948 5828
rect 39071 5797 39083 5800
rect 39025 5791 39083 5797
rect 39942 5788 39948 5800
rect 40000 5788 40006 5840
rect 32490 5760 32496 5772
rect 31680 5732 32496 5760
rect 29549 5723 29607 5729
rect 32490 5720 32496 5732
rect 32548 5720 32554 5772
rect 32674 5720 32680 5772
rect 32732 5760 32738 5772
rect 38470 5760 38476 5772
rect 32732 5732 38476 5760
rect 32732 5720 32738 5732
rect 38470 5720 38476 5732
rect 38528 5720 38534 5772
rect 25909 5664 26280 5692
rect 22278 5624 22284 5636
rect 21284 5596 22284 5624
rect 22278 5584 22284 5596
rect 22336 5584 22342 5636
rect 25130 5624 25136 5636
rect 24044 5596 25136 5624
rect 15620 5528 18920 5556
rect 15620 5516 15626 5528
rect 18966 5516 18972 5568
rect 19024 5556 19030 5568
rect 19429 5559 19487 5565
rect 19429 5556 19441 5559
rect 19024 5528 19441 5556
rect 19024 5516 19030 5528
rect 19429 5525 19441 5528
rect 19475 5525 19487 5559
rect 19429 5519 19487 5525
rect 19981 5559 20039 5565
rect 19981 5525 19993 5559
rect 20027 5556 20039 5559
rect 20898 5556 20904 5568
rect 20027 5528 20904 5556
rect 20027 5525 20039 5528
rect 19981 5519 20039 5525
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 21637 5559 21695 5565
rect 21637 5525 21649 5559
rect 21683 5556 21695 5559
rect 24044 5556 24072 5596
rect 25130 5584 25136 5596
rect 25188 5584 25194 5636
rect 25222 5584 25228 5636
rect 25280 5624 25286 5636
rect 25909 5624 25937 5664
rect 28074 5652 28080 5704
rect 28132 5692 28138 5704
rect 28169 5695 28227 5701
rect 28169 5692 28181 5695
rect 28132 5664 28181 5692
rect 28132 5652 28138 5664
rect 28169 5661 28181 5664
rect 28215 5661 28227 5695
rect 28169 5655 28227 5661
rect 29012 5664 29316 5692
rect 29012 5624 29040 5664
rect 25280 5596 25937 5624
rect 27632 5596 29040 5624
rect 25280 5584 25286 5596
rect 21683 5528 24072 5556
rect 21683 5525 21695 5528
rect 21637 5519 21695 5525
rect 24578 5516 24584 5568
rect 24636 5516 24642 5568
rect 24670 5516 24676 5568
rect 24728 5556 24734 5568
rect 24765 5559 24823 5565
rect 24765 5556 24777 5559
rect 24728 5528 24777 5556
rect 24728 5516 24734 5528
rect 24765 5525 24777 5528
rect 24811 5556 24823 5559
rect 26418 5556 26424 5568
rect 24811 5528 26424 5556
rect 24811 5525 24823 5528
rect 24765 5519 24823 5525
rect 26418 5516 26424 5528
rect 26476 5516 26482 5568
rect 26786 5516 26792 5568
rect 26844 5556 26850 5568
rect 27632 5556 27660 5596
rect 29086 5584 29092 5636
rect 29144 5584 29150 5636
rect 29288 5624 29316 5664
rect 29822 5652 29828 5704
rect 29880 5652 29886 5704
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 30653 5695 30711 5701
rect 30653 5692 30665 5695
rect 30524 5664 30665 5692
rect 30524 5652 30530 5664
rect 30653 5661 30665 5664
rect 30699 5661 30711 5695
rect 30653 5655 30711 5661
rect 30834 5652 30840 5704
rect 30892 5692 30898 5704
rect 30929 5695 30987 5701
rect 30929 5692 30941 5695
rect 30892 5664 30941 5692
rect 30892 5652 30898 5664
rect 30929 5661 30941 5664
rect 30975 5661 30987 5695
rect 30929 5655 30987 5661
rect 31018 5652 31024 5704
rect 31076 5692 31082 5704
rect 32125 5695 32183 5701
rect 32125 5692 32137 5695
rect 31076 5664 32137 5692
rect 31076 5652 31082 5664
rect 32125 5661 32137 5664
rect 32171 5661 32183 5695
rect 32125 5655 32183 5661
rect 32214 5652 32220 5704
rect 32272 5692 32278 5704
rect 32585 5695 32643 5701
rect 32272 5664 32536 5692
rect 32272 5652 32278 5664
rect 32508 5624 32536 5664
rect 32585 5661 32597 5695
rect 32631 5692 32643 5695
rect 32766 5692 32772 5704
rect 32631 5664 32772 5692
rect 32631 5661 32643 5664
rect 32585 5655 32643 5661
rect 32766 5652 32772 5664
rect 32824 5652 32830 5704
rect 33410 5652 33416 5704
rect 33468 5692 33474 5704
rect 34701 5695 34759 5701
rect 34701 5692 34713 5695
rect 33468 5664 34713 5692
rect 33468 5652 33474 5664
rect 34701 5661 34713 5664
rect 34747 5661 34759 5695
rect 34701 5655 34759 5661
rect 35066 5652 35072 5704
rect 35124 5692 35130 5704
rect 36541 5695 36599 5701
rect 36541 5692 36553 5695
rect 35124 5664 36553 5692
rect 35124 5652 35130 5664
rect 36541 5661 36553 5664
rect 36587 5661 36599 5695
rect 36541 5655 36599 5661
rect 37550 5652 37556 5704
rect 37608 5692 37614 5704
rect 38565 5695 38623 5701
rect 38565 5692 38577 5695
rect 37608 5664 38577 5692
rect 37608 5652 37614 5664
rect 38565 5661 38577 5664
rect 38611 5661 38623 5695
rect 38565 5655 38623 5661
rect 38841 5695 38899 5701
rect 38841 5661 38853 5695
rect 38887 5661 38899 5695
rect 38841 5655 38899 5661
rect 39209 5695 39267 5701
rect 39209 5661 39221 5695
rect 39255 5661 39267 5695
rect 39209 5655 39267 5661
rect 29288 5596 32260 5624
rect 32508 5596 34468 5624
rect 26844 5528 27660 5556
rect 26844 5516 26850 5528
rect 27706 5516 27712 5568
rect 27764 5556 27770 5568
rect 28442 5556 28448 5568
rect 27764 5528 28448 5556
rect 27764 5516 27770 5528
rect 28442 5516 28448 5528
rect 28500 5516 28506 5568
rect 28534 5516 28540 5568
rect 28592 5556 28598 5568
rect 28902 5556 28908 5568
rect 28592 5528 28908 5556
rect 28592 5516 28598 5528
rect 28902 5516 28908 5528
rect 28960 5556 28966 5568
rect 29181 5559 29239 5565
rect 29181 5556 29193 5559
rect 28960 5528 29193 5556
rect 28960 5516 28966 5528
rect 29181 5525 29193 5528
rect 29227 5525 29239 5559
rect 29181 5519 29239 5525
rect 29454 5516 29460 5568
rect 29512 5556 29518 5568
rect 32122 5556 32128 5568
rect 29512 5528 32128 5556
rect 29512 5516 29518 5528
rect 32122 5516 32128 5528
rect 32180 5516 32186 5568
rect 32232 5556 32260 5596
rect 32401 5559 32459 5565
rect 32401 5556 32413 5559
rect 32232 5528 32413 5556
rect 32401 5525 32413 5528
rect 32447 5525 32459 5559
rect 32401 5519 32459 5525
rect 33229 5559 33287 5565
rect 33229 5525 33241 5559
rect 33275 5556 33287 5559
rect 34054 5556 34060 5568
rect 33275 5528 34060 5556
rect 33275 5525 33287 5528
rect 33229 5519 33287 5525
rect 34054 5516 34060 5528
rect 34112 5516 34118 5568
rect 34440 5556 34468 5596
rect 34514 5584 34520 5636
rect 34572 5584 34578 5636
rect 36078 5584 36084 5636
rect 36136 5624 36142 5636
rect 38856 5624 38884 5655
rect 36136 5596 38884 5624
rect 36136 5584 36142 5596
rect 34974 5556 34980 5568
rect 34440 5528 34980 5556
rect 34974 5516 34980 5528
rect 35032 5516 35038 5568
rect 35894 5516 35900 5568
rect 35952 5556 35958 5568
rect 35989 5559 36047 5565
rect 35989 5556 36001 5559
rect 35952 5528 36001 5556
rect 35952 5516 35958 5528
rect 35989 5525 36001 5528
rect 36035 5525 36047 5559
rect 35989 5519 36047 5525
rect 36446 5516 36452 5568
rect 36504 5556 36510 5568
rect 39224 5556 39252 5655
rect 36504 5528 39252 5556
rect 36504 5516 36510 5528
rect 1104 5466 39836 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 9010 5466
rect 9062 5414 9074 5466
rect 9126 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 15010 5466
rect 15062 5414 15074 5466
rect 15126 5414 15138 5466
rect 15190 5414 15202 5466
rect 15254 5414 15266 5466
rect 15318 5414 21010 5466
rect 21062 5414 21074 5466
rect 21126 5414 21138 5466
rect 21190 5414 21202 5466
rect 21254 5414 21266 5466
rect 21318 5414 27010 5466
rect 27062 5414 27074 5466
rect 27126 5414 27138 5466
rect 27190 5414 27202 5466
rect 27254 5414 27266 5466
rect 27318 5414 33010 5466
rect 33062 5414 33074 5466
rect 33126 5414 33138 5466
rect 33190 5414 33202 5466
rect 33254 5414 33266 5466
rect 33318 5414 39010 5466
rect 39062 5414 39074 5466
rect 39126 5414 39138 5466
rect 39190 5414 39202 5466
rect 39254 5414 39266 5466
rect 39318 5414 39836 5466
rect 1104 5392 39836 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1946 5352 1952 5364
rect 1452 5324 1952 5352
rect 1452 5312 1458 5324
rect 1946 5312 1952 5324
rect 2004 5312 2010 5364
rect 3418 5312 3424 5364
rect 3476 5312 3482 5364
rect 3878 5312 3884 5364
rect 3936 5352 3942 5364
rect 4341 5355 4399 5361
rect 4341 5352 4353 5355
rect 3936 5324 4353 5352
rect 3936 5312 3942 5324
rect 4341 5321 4353 5324
rect 4387 5321 4399 5355
rect 4341 5315 4399 5321
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 6086 5352 6092 5364
rect 4856 5324 6092 5352
rect 4856 5312 4862 5324
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 7558 5352 7564 5364
rect 6227 5324 7564 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 7558 5312 7564 5324
rect 7616 5312 7622 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 9217 5355 9275 5361
rect 7800 5324 9168 5352
rect 7800 5312 7806 5324
rect 1486 5244 1492 5296
rect 1544 5244 1550 5296
rect 1670 5244 1676 5296
rect 1728 5244 1734 5296
rect 1854 5244 1860 5296
rect 1912 5244 1918 5296
rect 2225 5287 2283 5293
rect 2225 5284 2237 5287
rect 1964 5256 2237 5284
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 1964 5216 1992 5256
rect 2225 5253 2237 5256
rect 2271 5284 2283 5287
rect 2314 5284 2320 5296
rect 2271 5256 2320 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 1636 5188 1992 5216
rect 1636 5176 1642 5188
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 2648 5188 2697 5216
rect 2648 5176 2654 5188
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 2924 5188 2973 5216
rect 2924 5176 2930 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3234 5176 3240 5228
rect 3292 5176 3298 5228
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 3602 5176 3608 5228
rect 3660 5216 3666 5228
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3660 5188 3801 5216
rect 3660 5176 3666 5188
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3896 5216 3924 5312
rect 4157 5287 4215 5293
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 5074 5284 5080 5296
rect 4203 5256 4384 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 4356 5228 4384 5256
rect 4975 5256 5080 5284
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3896 5188 4077 5216
rect 3789 5179 3847 5185
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 2424 5148 2452 5176
rect 1912 5120 2452 5148
rect 4264 5148 4292 5179
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 4522 5176 4528 5228
rect 4580 5176 4586 5228
rect 4684 5219 4742 5225
rect 4684 5185 4696 5219
rect 4730 5216 4742 5219
rect 4798 5216 4804 5228
rect 4730 5188 4804 5216
rect 4730 5185 4742 5188
rect 4684 5179 4742 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4975 5225 5003 5256
rect 5074 5244 5080 5256
rect 5132 5244 5138 5296
rect 5994 5284 6000 5296
rect 5460 5256 6000 5284
rect 5460 5228 5488 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 6914 5284 6920 5296
rect 6196 5256 6920 5284
rect 6196 5228 6224 5256
rect 6914 5244 6920 5256
rect 6972 5284 6978 5296
rect 6972 5256 7420 5284
rect 6972 5244 6978 5256
rect 4960 5219 5018 5225
rect 4960 5185 4972 5219
rect 5006 5185 5018 5219
rect 4960 5179 5018 5185
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6604 5188 6653 5216
rect 6604 5176 6610 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6788 5188 6837 5216
rect 6788 5176 6794 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7190 5216 7196 5228
rect 7147 5188 7196 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7392 5225 7420 5256
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 8386 5176 8392 5228
rect 8444 5225 8450 5228
rect 8444 5219 8472 5225
rect 8460 5185 8472 5219
rect 8444 5179 8472 5185
rect 8573 5219 8631 5225
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 9140 5216 9168 5324
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9398 5352 9404 5364
rect 9263 5324 9404 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 11514 5352 11520 5364
rect 9508 5324 11520 5352
rect 9306 5244 9312 5296
rect 9364 5284 9370 5296
rect 9508 5284 9536 5324
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 11756 5324 12112 5352
rect 11756 5312 11762 5324
rect 9364 5256 9536 5284
rect 9364 5244 9370 5256
rect 9140 5188 9674 5216
rect 8573 5179 8631 5185
rect 8444 5176 8450 5179
rect 5074 5148 5080 5160
rect 4264 5120 5080 5148
rect 1912 5108 1918 5120
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5166 5108 5172 5160
rect 5224 5108 5230 5160
rect 5736 5148 5764 5176
rect 5736 5120 6040 5148
rect 2406 5040 2412 5092
rect 2464 5040 2470 5092
rect 3697 5083 3755 5089
rect 3697 5080 3709 5083
rect 2746 5052 3709 5080
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2746 5012 2774 5052
rect 3697 5049 3709 5052
rect 3743 5049 3755 5083
rect 4154 5080 4160 5092
rect 3697 5043 3755 5049
rect 3896 5052 4160 5080
rect 2372 4984 2774 5012
rect 2869 5015 2927 5021
rect 2372 4972 2378 4984
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 2958 5012 2964 5024
rect 2915 4984 2964 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 3896 5012 3924 5052
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 4755 5083 4813 5089
rect 4264 5052 4660 5080
rect 3191 4984 3924 5012
rect 3973 5015 4031 5021
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 3973 4981 3985 5015
rect 4019 5012 4031 5015
rect 4264 5012 4292 5052
rect 4019 4984 4292 5012
rect 4019 4981 4031 4984
rect 3973 4975 4031 4981
rect 4338 4972 4344 5024
rect 4396 4972 4402 5024
rect 4632 5012 4660 5052
rect 4755 5049 4767 5083
rect 4801 5080 4813 5083
rect 6012 5080 6040 5120
rect 6086 5108 6092 5160
rect 6144 5148 6150 5160
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 6144 5120 6377 5148
rect 6144 5108 6150 5120
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7524 5120 7573 5148
rect 7524 5108 7530 5120
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 7742 5108 7748 5160
rect 7800 5108 7806 5160
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8110 5148 8116 5160
rect 7984 5120 8116 5148
rect 7984 5108 7990 5120
rect 8110 5108 8116 5120
rect 8168 5148 8174 5160
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 8168 5120 8309 5148
rect 8168 5108 8174 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8588 5148 8616 5179
rect 8938 5148 8944 5160
rect 8588 5120 8944 5148
rect 8297 5111 8355 5117
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 9122 5108 9128 5160
rect 9180 5148 9186 5160
rect 9306 5148 9312 5160
rect 9180 5120 9312 5148
rect 9180 5108 9186 5120
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 9490 5108 9496 5160
rect 9548 5108 9554 5160
rect 9646 5148 9674 5188
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 11882 5216 11888 5228
rect 11839 5188 11888 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 10410 5157 10416 5160
rect 10367 5151 10416 5157
rect 10367 5148 10379 5151
rect 9646 5120 10379 5148
rect 10367 5117 10379 5120
rect 10413 5117 10416 5151
rect 10367 5111 10416 5117
rect 10410 5108 10416 5111
rect 10468 5108 10474 5160
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 10686 5148 10692 5160
rect 10551 5120 10692 5148
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 10686 5108 10692 5120
rect 10744 5148 10750 5160
rect 11716 5148 11744 5179
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 12084 5225 12112 5324
rect 12250 5312 12256 5364
rect 12308 5312 12314 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12529 5355 12587 5361
rect 12529 5352 12541 5355
rect 12492 5324 12541 5352
rect 12492 5312 12498 5324
rect 12529 5321 12541 5324
rect 12575 5321 12587 5355
rect 12529 5315 12587 5321
rect 12618 5312 12624 5364
rect 12676 5312 12682 5364
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 13081 5355 13139 5361
rect 13081 5321 13093 5355
rect 13127 5352 13139 5355
rect 13127 5324 14872 5352
rect 13127 5321 13139 5324
rect 13081 5315 13139 5321
rect 12820 5284 12848 5312
rect 14844 5284 14872 5324
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 14976 5324 15117 5352
rect 14976 5312 14982 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 19705 5355 19763 5361
rect 15252 5324 19564 5352
rect 15252 5312 15258 5324
rect 19536 5284 19564 5324
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 21450 5352 21456 5364
rect 19751 5324 21456 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 23750 5352 23756 5364
rect 22704 5324 23756 5352
rect 22704 5312 22710 5324
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 24118 5312 24124 5364
rect 24176 5352 24182 5364
rect 25222 5352 25228 5364
rect 24176 5324 25228 5352
rect 24176 5312 24182 5324
rect 25222 5312 25228 5324
rect 25280 5312 25286 5364
rect 25314 5312 25320 5364
rect 25372 5352 25378 5364
rect 26510 5352 26516 5364
rect 25372 5324 26516 5352
rect 25372 5312 25378 5324
rect 26510 5312 26516 5324
rect 26568 5312 26574 5364
rect 26602 5312 26608 5364
rect 26660 5352 26666 5364
rect 27430 5352 27436 5364
rect 26660 5324 27436 5352
rect 26660 5312 26666 5324
rect 27430 5312 27436 5324
rect 27488 5312 27494 5364
rect 27890 5352 27896 5364
rect 27816 5324 27896 5352
rect 12820 5256 13584 5284
rect 14844 5256 17908 5284
rect 19536 5256 20024 5284
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12069 5179 12127 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 12710 5216 12716 5228
rect 12391 5188 12716 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 12802 5176 12808 5228
rect 12860 5176 12866 5228
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5216 12955 5219
rect 13078 5216 13084 5228
rect 12943 5188 13084 5216
rect 12943 5185 12955 5188
rect 12897 5179 12955 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5185 13231 5219
rect 13556 5216 13584 5256
rect 13725 5219 13783 5225
rect 13725 5216 13737 5219
rect 13556 5188 13737 5216
rect 13173 5179 13231 5185
rect 13725 5185 13737 5188
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 12618 5148 12624 5160
rect 10744 5120 10916 5148
rect 11716 5120 12624 5148
rect 10744 5108 10750 5120
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 4801 5052 5304 5080
rect 6012 5052 6561 5080
rect 4801 5049 4813 5052
rect 4755 5043 4813 5049
rect 4890 5012 4896 5024
rect 4632 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5031 5015 5089 5021
rect 5031 4981 5043 5015
rect 5077 5012 5089 5015
rect 5166 5012 5172 5024
rect 5077 4984 5172 5012
rect 5077 4981 5089 4984
rect 5031 4975 5089 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5276 5012 5304 5052
rect 6549 5049 6561 5052
rect 6595 5049 6607 5083
rect 6549 5043 6607 5049
rect 7006 5040 7012 5092
rect 7064 5040 7070 5092
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7760 5080 7788 5108
rect 7156 5052 7788 5080
rect 8021 5083 8079 5089
rect 7156 5040 7162 5052
rect 8021 5049 8033 5083
rect 8067 5049 8079 5083
rect 9950 5080 9956 5092
rect 8021 5043 8079 5049
rect 8956 5052 9956 5080
rect 5442 5012 5448 5024
rect 5276 4984 5448 5012
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6457 5015 6515 5021
rect 6457 5012 6469 5015
rect 6328 4984 6469 5012
rect 6328 4972 6334 4984
rect 6457 4981 6469 4984
rect 6503 4981 6515 5015
rect 6457 4975 6515 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7650 5012 7656 5024
rect 7331 4984 7656 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 8036 5012 8064 5043
rect 8956 5012 8984 5052
rect 9950 5040 9956 5052
rect 10008 5040 10014 5092
rect 8036 4984 8984 5012
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9582 5012 9588 5024
rect 9088 4984 9588 5012
rect 9088 4972 9094 4984
rect 9582 4972 9588 4984
rect 9640 5012 9646 5024
rect 10888 5012 10916 5120
rect 12618 5108 12624 5120
rect 12676 5148 12682 5160
rect 12986 5148 12992 5160
rect 12676 5120 12992 5148
rect 12676 5108 12682 5120
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13188 5148 13216 5179
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 14826 5176 14832 5228
rect 14884 5176 14890 5228
rect 15746 5176 15752 5228
rect 15804 5214 15810 5228
rect 15841 5219 15899 5225
rect 15841 5214 15853 5219
rect 15804 5186 15853 5214
rect 15804 5176 15810 5186
rect 15841 5185 15853 5186
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 16206 5176 16212 5228
rect 16264 5216 16270 5228
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 16264 5188 16313 5216
rect 16264 5176 16270 5188
rect 16301 5185 16313 5188
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16758 5176 16764 5228
rect 16816 5176 16822 5228
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17880 5225 17908 5256
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 17000 5188 17049 5216
rect 17000 5176 17006 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 18230 5216 18236 5228
rect 17911 5188 18236 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 18782 5176 18788 5228
rect 18840 5176 18846 5228
rect 18874 5176 18880 5228
rect 18932 5225 18938 5228
rect 18932 5219 18960 5225
rect 18948 5185 18960 5219
rect 18932 5179 18960 5185
rect 19797 5219 19855 5225
rect 19797 5185 19809 5219
rect 19843 5216 19855 5219
rect 19886 5216 19892 5228
rect 19843 5188 19892 5216
rect 19843 5185 19855 5188
rect 19797 5179 19855 5185
rect 18932 5176 18938 5179
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 19996 5225 20024 5256
rect 22664 5256 26924 5284
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 20714 5176 20720 5228
rect 20772 5176 20778 5228
rect 21637 5219 21695 5225
rect 21637 5185 21649 5219
rect 21683 5216 21695 5219
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21683 5188 22017 5216
rect 21683 5185 21695 5188
rect 21637 5179 21695 5185
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22462 5176 22468 5228
rect 22520 5176 22526 5228
rect 13354 5148 13360 5160
rect 13188 5120 13360 5148
rect 13354 5108 13360 5120
rect 13412 5148 13418 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 13412 5120 13461 5148
rect 13412 5108 13418 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 16117 5151 16175 5157
rect 14424 5120 15424 5148
rect 14424 5108 14430 5120
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 11977 5083 12035 5089
rect 11112 5052 11928 5080
rect 11112 5040 11118 5052
rect 9640 4984 10916 5012
rect 9640 4972 9646 4984
rect 10962 4972 10968 5024
rect 11020 5012 11026 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 11020 4984 11161 5012
rect 11020 4972 11026 4984
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11149 4975 11207 4981
rect 11609 5015 11667 5021
rect 11609 4981 11621 5015
rect 11655 5012 11667 5015
rect 11790 5012 11796 5024
rect 11655 4984 11796 5012
rect 11655 4981 11667 4984
rect 11609 4975 11667 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 11900 5012 11928 5052
rect 11977 5049 11989 5083
rect 12023 5080 12035 5083
rect 13262 5080 13268 5092
rect 12023 5052 13268 5080
rect 12023 5049 12035 5052
rect 11977 5043 12035 5049
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 14461 5083 14519 5089
rect 14461 5049 14473 5083
rect 14507 5080 14519 5083
rect 15286 5080 15292 5092
rect 14507 5052 15292 5080
rect 14507 5049 14519 5052
rect 14461 5043 14519 5049
rect 15286 5040 15292 5052
rect 15344 5040 15350 5092
rect 12526 5012 12532 5024
rect 11900 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 14090 5012 14096 5024
rect 13403 4984 14096 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14737 5015 14795 5021
rect 14737 4981 14749 5015
rect 14783 5012 14795 5015
rect 14918 5012 14924 5024
rect 14783 4984 14924 5012
rect 14783 4981 14795 4984
rect 14737 4975 14795 4981
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15013 5015 15071 5021
rect 15013 4981 15025 5015
rect 15059 5012 15071 5015
rect 15102 5012 15108 5024
rect 15059 4984 15108 5012
rect 15059 4981 15071 4984
rect 15013 4975 15071 4981
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 15396 5012 15424 5120
rect 16117 5117 16129 5151
rect 16163 5148 16175 5151
rect 16390 5148 16396 5160
rect 16163 5120 16396 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 18046 5108 18052 5160
rect 18104 5108 18110 5160
rect 18414 5108 18420 5160
rect 18472 5148 18478 5160
rect 18892 5148 18920 5176
rect 18472 5120 18920 5148
rect 19061 5151 19119 5157
rect 18472 5108 18478 5120
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 19242 5148 19248 5160
rect 19107 5120 19248 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 20834 5151 20892 5157
rect 20834 5148 20846 5151
rect 19996 5120 20846 5148
rect 17773 5083 17831 5089
rect 16040 5052 16620 5080
rect 16040 5012 16068 5052
rect 15396 4984 16068 5012
rect 16298 4972 16304 5024
rect 16356 5012 16362 5024
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 16356 4984 16497 5012
rect 16356 4972 16362 4984
rect 16485 4981 16497 4984
rect 16531 4981 16543 5015
rect 16592 5012 16620 5052
rect 17773 5049 17785 5083
rect 17819 5080 17831 5083
rect 18509 5083 18567 5089
rect 18509 5080 18521 5083
rect 17819 5052 18521 5080
rect 17819 5049 17831 5052
rect 17773 5043 17831 5049
rect 18509 5049 18521 5052
rect 18555 5049 18567 5083
rect 18509 5043 18567 5049
rect 17862 5012 17868 5024
rect 16592 4984 17868 5012
rect 16485 4975 16543 4981
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 18230 4972 18236 5024
rect 18288 5012 18294 5024
rect 19996 5012 20024 5120
rect 20834 5117 20846 5120
rect 20880 5117 20892 5151
rect 20834 5111 20892 5117
rect 20993 5151 21051 5157
rect 20993 5117 21005 5151
rect 21039 5148 21051 5151
rect 22664 5148 22692 5256
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 23017 5219 23075 5225
rect 23017 5216 23029 5219
rect 22980 5188 23029 5216
rect 22980 5176 22986 5188
rect 23017 5185 23029 5188
rect 23063 5216 23075 5219
rect 24302 5216 24308 5228
rect 23063 5188 24308 5216
rect 23063 5185 23075 5188
rect 23017 5179 23075 5185
rect 24302 5176 24308 5188
rect 24360 5176 24366 5228
rect 24581 5219 24639 5225
rect 24581 5185 24593 5219
rect 24627 5216 24639 5219
rect 24854 5216 24860 5228
rect 24627 5188 24860 5216
rect 24627 5185 24639 5188
rect 24581 5179 24639 5185
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 25317 5219 25375 5225
rect 25317 5216 25329 5219
rect 24964 5188 25329 5216
rect 21039 5120 22692 5148
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 22738 5108 22744 5160
rect 22796 5108 22802 5160
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 24026 5148 24032 5160
rect 23440 5120 24032 5148
rect 23440 5108 23446 5120
rect 24026 5108 24032 5120
rect 24084 5148 24090 5160
rect 24964 5148 24992 5188
rect 25317 5185 25329 5188
rect 25363 5185 25375 5219
rect 25317 5179 25375 5185
rect 25406 5176 25412 5228
rect 25464 5216 25470 5228
rect 26145 5219 26203 5225
rect 26145 5216 26157 5219
rect 25464 5188 26157 5216
rect 25464 5176 25470 5188
rect 26145 5185 26157 5188
rect 26191 5185 26203 5219
rect 26145 5179 26203 5185
rect 26786 5176 26792 5228
rect 26844 5176 26850 5228
rect 24084 5120 24992 5148
rect 24084 5108 24090 5120
rect 25038 5108 25044 5160
rect 25096 5108 25102 5160
rect 26896 5148 26924 5256
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5216 27399 5219
rect 27430 5216 27436 5228
rect 27387 5188 27436 5216
rect 27387 5185 27399 5188
rect 27341 5179 27399 5185
rect 27430 5176 27436 5188
rect 27488 5176 27494 5228
rect 27525 5219 27583 5225
rect 27525 5185 27537 5219
rect 27571 5216 27583 5219
rect 27614 5216 27620 5228
rect 27571 5188 27620 5216
rect 27571 5185 27583 5188
rect 27525 5179 27583 5185
rect 27614 5176 27620 5188
rect 27672 5176 27678 5228
rect 27816 5225 27844 5324
rect 27890 5312 27896 5324
rect 27948 5352 27954 5364
rect 29086 5352 29092 5364
rect 27948 5324 29092 5352
rect 27948 5312 27954 5324
rect 29086 5312 29092 5324
rect 29144 5352 29150 5364
rect 29638 5352 29644 5364
rect 29144 5324 29644 5352
rect 29144 5312 29150 5324
rect 29638 5312 29644 5324
rect 29696 5312 29702 5364
rect 29917 5355 29975 5361
rect 29917 5321 29929 5355
rect 29963 5352 29975 5355
rect 30190 5352 30196 5364
rect 29963 5324 30196 5352
rect 29963 5321 29975 5324
rect 29917 5315 29975 5321
rect 30190 5312 30196 5324
rect 30248 5312 30254 5364
rect 32309 5355 32367 5361
rect 30760 5324 32168 5352
rect 28074 5244 28080 5296
rect 28132 5244 28138 5296
rect 28166 5244 28172 5296
rect 28224 5284 28230 5296
rect 28224 5256 30512 5284
rect 28224 5244 28230 5256
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5185 27859 5219
rect 28077 5215 28089 5244
rect 28123 5215 28135 5244
rect 28077 5209 28135 5215
rect 27801 5179 27859 5185
rect 27706 5148 27712 5160
rect 26896 5120 27712 5148
rect 27706 5108 27712 5120
rect 27764 5108 27770 5160
rect 20438 5040 20444 5092
rect 20496 5040 20502 5092
rect 21542 5040 21548 5092
rect 21600 5080 21606 5092
rect 22646 5080 22652 5092
rect 21600 5052 22652 5080
rect 21600 5040 21606 5052
rect 22646 5040 22652 5052
rect 22704 5040 22710 5092
rect 27816 5080 27844 5179
rect 28442 5176 28448 5228
rect 28500 5216 28506 5228
rect 29086 5216 29092 5228
rect 28500 5188 29092 5216
rect 28500 5176 28506 5188
rect 29086 5176 29092 5188
rect 29144 5176 29150 5228
rect 29181 5219 29239 5225
rect 29181 5185 29193 5219
rect 29227 5216 29239 5219
rect 29270 5216 29276 5228
rect 29227 5188 29276 5216
rect 29227 5185 29239 5188
rect 29181 5179 29239 5185
rect 29270 5176 29276 5188
rect 29328 5176 29334 5228
rect 28902 5108 28908 5160
rect 28960 5108 28966 5160
rect 30484 5148 30512 5256
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5216 30619 5219
rect 30760 5216 30788 5324
rect 32140 5284 32168 5324
rect 32309 5321 32321 5355
rect 32355 5352 32367 5355
rect 32674 5352 32680 5364
rect 32355 5324 32680 5352
rect 32355 5321 32367 5324
rect 32309 5315 32367 5321
rect 32674 5312 32680 5324
rect 32732 5312 32738 5364
rect 32950 5312 32956 5364
rect 33008 5352 33014 5364
rect 33502 5352 33508 5364
rect 33008 5324 33508 5352
rect 33008 5312 33014 5324
rect 33502 5312 33508 5324
rect 33560 5312 33566 5364
rect 34606 5312 34612 5364
rect 34664 5312 34670 5364
rect 36170 5312 36176 5364
rect 36228 5312 36234 5364
rect 39390 5312 39396 5364
rect 39448 5312 39454 5364
rect 33042 5284 33048 5296
rect 32140 5256 33048 5284
rect 33042 5244 33048 5256
rect 33100 5244 33106 5296
rect 33812 5287 33870 5293
rect 33812 5253 33824 5287
rect 33858 5284 33870 5287
rect 34330 5284 34336 5296
rect 33858 5256 34336 5284
rect 33858 5253 33870 5256
rect 33812 5247 33870 5253
rect 34330 5244 34336 5256
rect 34388 5244 34394 5296
rect 35894 5244 35900 5296
rect 35952 5244 35958 5296
rect 30607 5188 30788 5216
rect 31021 5219 31079 5225
rect 30607 5185 30619 5188
rect 30561 5179 30619 5185
rect 31021 5185 31033 5219
rect 31067 5216 31079 5219
rect 31113 5219 31171 5225
rect 31113 5216 31125 5219
rect 31067 5188 31125 5216
rect 31067 5185 31079 5188
rect 31021 5179 31079 5185
rect 31113 5185 31125 5188
rect 31159 5185 31171 5219
rect 31113 5179 31171 5185
rect 31386 5176 31392 5228
rect 31444 5216 31450 5228
rect 31481 5219 31539 5225
rect 31481 5216 31493 5219
rect 31444 5188 31493 5216
rect 31444 5176 31450 5188
rect 31481 5185 31493 5188
rect 31527 5185 31539 5219
rect 31481 5179 31539 5185
rect 31662 5176 31668 5228
rect 31720 5216 31726 5228
rect 32125 5219 32183 5225
rect 32125 5216 32137 5219
rect 31720 5188 32137 5216
rect 31720 5176 31726 5188
rect 32125 5185 32137 5188
rect 32171 5185 32183 5219
rect 32125 5179 32183 5185
rect 32214 5176 32220 5228
rect 32272 5216 32278 5228
rect 32401 5220 32459 5225
rect 32324 5219 32459 5220
rect 32324 5216 32413 5219
rect 32272 5192 32413 5216
rect 32272 5188 32352 5192
rect 32272 5176 32278 5188
rect 32401 5185 32413 5192
rect 32447 5185 32459 5219
rect 32401 5179 32459 5185
rect 33060 5188 34008 5216
rect 30484 5120 31800 5148
rect 25700 5052 27844 5080
rect 18288 4984 20024 5012
rect 18288 4972 18294 4984
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 20530 5012 20536 5024
rect 20128 4984 20536 5012
rect 20128 4972 20134 4984
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 20772 4984 21833 5012
rect 20772 4972 20778 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 22281 5015 22339 5021
rect 22281 5012 22293 5015
rect 22244 4984 22293 5012
rect 22244 4972 22250 4984
rect 22281 4981 22293 4984
rect 22327 4981 22339 5015
rect 22281 4975 22339 4981
rect 23750 4972 23756 5024
rect 23808 4972 23814 5024
rect 23934 4972 23940 5024
rect 23992 5012 23998 5024
rect 24486 5012 24492 5024
rect 23992 4984 24492 5012
rect 23992 4972 23998 4984
rect 24486 4972 24492 4984
rect 24544 4972 24550 5024
rect 24762 4972 24768 5024
rect 24820 4972 24826 5024
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25700 5012 25728 5052
rect 30006 5040 30012 5092
rect 30064 5080 30070 5092
rect 30064 5052 30512 5080
rect 30064 5040 30070 5052
rect 25004 4984 25728 5012
rect 25004 4972 25010 4984
rect 25866 4972 25872 5024
rect 25924 5012 25930 5024
rect 26053 5015 26111 5021
rect 26053 5012 26065 5015
rect 25924 4984 26065 5012
rect 25924 4972 25930 4984
rect 26053 4981 26065 4984
rect 26099 4981 26111 5015
rect 26053 4975 26111 4981
rect 26329 5015 26387 5021
rect 26329 4981 26341 5015
rect 26375 5012 26387 5015
rect 26418 5012 26424 5024
rect 26375 4984 26424 5012
rect 26375 4981 26387 4984
rect 26329 4975 26387 4981
rect 26418 4972 26424 4984
rect 26476 4972 26482 5024
rect 26605 5015 26663 5021
rect 26605 4981 26617 5015
rect 26651 5012 26663 5015
rect 26878 5012 26884 5024
rect 26651 4984 26884 5012
rect 26651 4981 26663 4984
rect 26605 4975 26663 4981
rect 26878 4972 26884 4984
rect 26936 4972 26942 5024
rect 27157 5015 27215 5021
rect 27157 4981 27169 5015
rect 27203 5012 27215 5015
rect 27338 5012 27344 5024
rect 27203 4984 27344 5012
rect 27203 4981 27215 4984
rect 27157 4975 27215 4981
rect 27338 4972 27344 4984
rect 27396 4972 27402 5024
rect 27709 5015 27767 5021
rect 27709 4981 27721 5015
rect 27755 5012 27767 5015
rect 28166 5012 28172 5024
rect 27755 4984 28172 5012
rect 27755 4981 27767 4984
rect 27709 4975 27767 4981
rect 28166 4972 28172 4984
rect 28224 4972 28230 5024
rect 28813 5015 28871 5021
rect 28813 4981 28825 5015
rect 28859 5012 28871 5015
rect 29546 5012 29552 5024
rect 28859 4984 29552 5012
rect 28859 4981 28871 4984
rect 28813 4975 28871 4981
rect 29546 4972 29552 4984
rect 29604 4972 29610 5024
rect 30374 4972 30380 5024
rect 30432 4972 30438 5024
rect 30484 5012 30512 5052
rect 30558 5040 30564 5092
rect 30616 5080 30622 5092
rect 30616 5052 31064 5080
rect 30616 5040 30622 5052
rect 30929 5015 30987 5021
rect 30929 5012 30941 5015
rect 30484 4984 30941 5012
rect 30929 4981 30941 4984
rect 30975 4981 30987 5015
rect 31036 5012 31064 5052
rect 31662 5040 31668 5092
rect 31720 5040 31726 5092
rect 31772 5080 31800 5120
rect 32306 5108 32312 5160
rect 32364 5148 32370 5160
rect 33060 5148 33088 5188
rect 32364 5120 33088 5148
rect 33980 5148 34008 5188
rect 34054 5176 34060 5228
rect 34112 5176 34118 5228
rect 34790 5176 34796 5228
rect 34848 5216 34854 5228
rect 35989 5219 36047 5225
rect 35989 5216 36001 5219
rect 34848 5188 36001 5216
rect 34848 5176 34854 5188
rect 35989 5185 36001 5188
rect 36035 5185 36047 5219
rect 35989 5179 36047 5185
rect 38838 5176 38844 5228
rect 38896 5176 38902 5228
rect 38930 5176 38936 5228
rect 38988 5216 38994 5228
rect 39209 5219 39267 5225
rect 39209 5216 39221 5219
rect 38988 5188 39221 5216
rect 38988 5176 38994 5188
rect 39209 5185 39221 5188
rect 39255 5185 39267 5219
rect 39209 5179 39267 5185
rect 36630 5148 36636 5160
rect 33980 5120 36636 5148
rect 32364 5108 32370 5120
rect 36630 5108 36636 5120
rect 36688 5108 36694 5160
rect 31772 5052 33088 5080
rect 31297 5015 31355 5021
rect 31297 5012 31309 5015
rect 31036 4984 31309 5012
rect 30929 4975 30987 4981
rect 31297 4981 31309 4984
rect 31343 4981 31355 5015
rect 31297 4975 31355 4981
rect 31386 4972 31392 5024
rect 31444 5012 31450 5024
rect 32214 5012 32220 5024
rect 31444 4984 32220 5012
rect 31444 4972 31450 4984
rect 32214 4972 32220 4984
rect 32272 4972 32278 5024
rect 32582 4972 32588 5024
rect 32640 4972 32646 5024
rect 32677 5015 32735 5021
rect 32677 4981 32689 5015
rect 32723 5012 32735 5015
rect 32950 5012 32956 5024
rect 32723 4984 32956 5012
rect 32723 4981 32735 4984
rect 32677 4975 32735 4981
rect 32950 4972 32956 4984
rect 33008 4972 33014 5024
rect 33060 5012 33088 5052
rect 35342 5012 35348 5024
rect 33060 4984 35348 5012
rect 35342 4972 35348 4984
rect 35400 4972 35406 5024
rect 39022 4972 39028 5024
rect 39080 4972 39086 5024
rect 1104 4922 39836 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 13950 4922
rect 14002 4870 14014 4922
rect 14066 4870 14078 4922
rect 14130 4870 14142 4922
rect 14194 4870 14206 4922
rect 14258 4870 19950 4922
rect 20002 4870 20014 4922
rect 20066 4870 20078 4922
rect 20130 4870 20142 4922
rect 20194 4870 20206 4922
rect 20258 4870 25950 4922
rect 26002 4870 26014 4922
rect 26066 4870 26078 4922
rect 26130 4870 26142 4922
rect 26194 4870 26206 4922
rect 26258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 37950 4922
rect 38002 4870 38014 4922
rect 38066 4870 38078 4922
rect 38130 4870 38142 4922
rect 38194 4870 38206 4922
rect 38258 4870 39836 4922
rect 1104 4848 39836 4870
rect 1854 4768 1860 4820
rect 1912 4808 1918 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1912 4780 1961 4808
rect 1912 4768 1918 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 1949 4771 2007 4777
rect 2498 4768 2504 4820
rect 2556 4768 2562 4820
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 3878 4808 3884 4820
rect 2915 4780 3884 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4338 4768 4344 4820
rect 4396 4808 4402 4820
rect 4396 4780 6684 4808
rect 4396 4768 4402 4780
rect 3234 4700 3240 4752
rect 3292 4740 3298 4752
rect 3694 4740 3700 4752
rect 3292 4712 3700 4740
rect 3292 4700 3298 4712
rect 3694 4700 3700 4712
rect 3752 4700 3758 4752
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 3602 4672 3608 4684
rect 1728 4644 3608 4672
rect 1728 4632 1734 4644
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 3936 4644 4445 4672
rect 3936 4632 3942 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 4522 4632 4528 4684
rect 4580 4681 4586 4684
rect 4580 4675 4629 4681
rect 4580 4641 4583 4675
rect 4617 4641 4629 4675
rect 4580 4635 4629 4641
rect 4580 4632 4586 4635
rect 4982 4632 4988 4684
rect 5040 4632 5046 4684
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5445 4675 5503 4681
rect 5445 4672 5457 4675
rect 5132 4644 5457 4672
rect 5132 4632 5138 4644
rect 5445 4641 5457 4644
rect 5491 4641 5503 4675
rect 6656 4672 6684 4780
rect 7282 4768 7288 4820
rect 7340 4768 7346 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 8260 4780 8953 4808
rect 8260 4768 8266 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 9088 4780 9137 4808
rect 9088 4768 9094 4780
rect 9125 4777 9137 4780
rect 9171 4777 9183 4811
rect 9125 4771 9183 4777
rect 9585 4811 9643 4817
rect 9585 4777 9597 4811
rect 9631 4808 9643 4811
rect 10318 4808 10324 4820
rect 9631 4780 10324 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 11388 4780 12756 4808
rect 11388 4768 11394 4780
rect 7300 4740 7328 4768
rect 7300 4712 7696 4740
rect 7006 4672 7012 4684
rect 6656 4644 7012 4672
rect 5445 4635 5503 4641
rect 7006 4632 7012 4644
rect 7064 4672 7070 4684
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 7064 4644 7113 4672
rect 7064 4632 7070 4644
rect 7101 4641 7113 4644
rect 7147 4672 7159 4675
rect 7466 4672 7472 4684
rect 7147 4644 7472 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 7558 4632 7564 4684
rect 7616 4632 7622 4684
rect 7668 4672 7696 4712
rect 8496 4712 10941 4740
rect 7954 4675 8012 4681
rect 7954 4672 7966 4675
rect 7668 4644 7966 4672
rect 7954 4641 7966 4644
rect 8000 4641 8012 4675
rect 7954 4635 8012 4641
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8496 4672 8524 4712
rect 8352 4644 8524 4672
rect 8352 4632 8358 4644
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9030 4672 9036 4684
rect 8720 4644 9036 4672
rect 8720 4632 8726 4644
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 9692 4644 10793 4672
rect 1486 4564 1492 4616
rect 1544 4564 1550 4616
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 1964 4576 2789 4604
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 1762 4536 1768 4548
rect 1719 4508 1768 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 1964 4536 1992 4576
rect 2777 4573 2789 4576
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3326 4604 3332 4616
rect 3099 4576 3332 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4604 3479 4607
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3467 4576 3801 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 5767 4576 5856 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 5828 4548 5856 4576
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5960 4576 6009 4604
rect 5960 4564 5966 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 7834 4564 7840 4616
rect 7892 4564 7898 4616
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8812 4576 9137 4604
rect 8812 4564 8818 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 9582 4604 9588 4616
rect 9539 4576 9588 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 9692 4548 9720 4644
rect 10781 4641 10793 4644
rect 10827 4641 10839 4675
rect 10913 4672 10941 4712
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 12728 4740 12756 4780
rect 12986 4768 12992 4820
rect 13044 4808 13050 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 13044 4780 13093 4808
rect 13044 4768 13050 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13725 4811 13783 4817
rect 13725 4808 13737 4811
rect 13228 4780 13737 4808
rect 13228 4768 13234 4780
rect 13725 4777 13737 4780
rect 13771 4808 13783 4811
rect 14366 4808 14372 4820
rect 13771 4780 14372 4808
rect 13771 4777 13783 4780
rect 13725 4771 13783 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 14884 4780 15945 4808
rect 14884 4768 14890 4780
rect 15933 4777 15945 4780
rect 15979 4777 15991 4811
rect 15933 4771 15991 4777
rect 16206 4768 16212 4820
rect 16264 4768 16270 4820
rect 17402 4768 17408 4820
rect 17460 4768 17466 4820
rect 17770 4808 17776 4820
rect 17512 4780 17776 4808
rect 13906 4740 13912 4752
rect 11940 4712 12112 4740
rect 12728 4712 13912 4740
rect 11940 4700 11946 4712
rect 12084 4681 12112 4712
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 17420 4740 17448 4768
rect 14660 4712 14872 4740
rect 12069 4675 12127 4681
rect 10913 4644 12020 4672
rect 10781 4635 10839 4641
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 9858 4604 9864 4616
rect 9815 4576 9864 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 10042 4604 10048 4616
rect 9999 4576 10048 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 10134 4564 10140 4616
rect 10192 4564 10198 4616
rect 10318 4564 10324 4616
rect 10376 4564 10382 4616
rect 11054 4564 11060 4616
rect 11112 4564 11118 4616
rect 11238 4613 11244 4616
rect 11195 4607 11244 4613
rect 11195 4573 11207 4607
rect 11241 4573 11244 4607
rect 11195 4567 11244 4573
rect 11238 4564 11244 4567
rect 11296 4564 11302 4616
rect 11330 4564 11336 4616
rect 11388 4564 11394 4616
rect 11992 4604 12020 4644
rect 12069 4641 12081 4675
rect 12115 4641 12127 4675
rect 14660 4672 14688 4712
rect 12069 4635 12127 4641
rect 12636 4644 14688 4672
rect 12345 4607 12403 4613
rect 11992 4576 12296 4604
rect 1872 4508 1992 4536
rect 2225 4539 2283 4545
rect 474 4428 480 4480
rect 532 4468 538 4480
rect 1872 4468 1900 4508
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 2406 4536 2412 4548
rect 2271 4508 2412 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 5810 4496 5816 4548
rect 5868 4496 5874 4548
rect 7098 4536 7104 4548
rect 5920 4508 7104 4536
rect 532 4440 1900 4468
rect 532 4428 538 4440
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2501 4471 2559 4477
rect 2501 4468 2513 4471
rect 2372 4440 2513 4468
rect 2372 4428 2378 4440
rect 2501 4437 2513 4440
rect 2547 4437 2559 4471
rect 2501 4431 2559 4437
rect 3234 4428 3240 4480
rect 3292 4428 3298 4480
rect 3602 4428 3608 4480
rect 3660 4428 3666 4480
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 5920 4468 5948 4508
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 9674 4536 9680 4548
rect 8588 4508 9680 4536
rect 4764 4440 5948 4468
rect 6733 4471 6791 4477
rect 4764 4428 4770 4440
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 7558 4468 7564 4480
rect 6779 4440 7564 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 7558 4428 7564 4440
rect 7616 4468 7622 4480
rect 8588 4468 8616 4508
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 12268 4536 12296 4576
rect 12345 4573 12357 4607
rect 12391 4604 12403 4607
rect 12434 4604 12440 4616
rect 12391 4576 12440 4604
rect 12391 4573 12403 4576
rect 12345 4567 12403 4573
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 12636 4536 12664 4644
rect 14734 4632 14740 4684
rect 14792 4632 14798 4684
rect 14844 4672 14872 4712
rect 17328 4712 17448 4740
rect 15010 4672 15016 4684
rect 14844 4644 15016 4672
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 15286 4632 15292 4684
rect 15344 4632 15350 4684
rect 17129 4675 17187 4681
rect 17129 4641 17141 4675
rect 17175 4672 17187 4675
rect 17328 4672 17356 4712
rect 17175 4644 17356 4672
rect 17405 4675 17463 4681
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 17405 4641 17417 4675
rect 17451 4672 17463 4675
rect 17512 4672 17540 4780
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 17920 4780 18828 4808
rect 17920 4768 17926 4780
rect 17678 4700 17684 4752
rect 17736 4740 17742 4752
rect 18800 4740 18828 4780
rect 19242 4768 19248 4820
rect 19300 4768 19306 4820
rect 19352 4780 20208 4808
rect 19352 4740 19380 4780
rect 17736 4712 18736 4740
rect 18800 4712 19380 4740
rect 20180 4740 20208 4780
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 22370 4808 22376 4820
rect 20496 4780 22376 4808
rect 20496 4768 20502 4780
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 22554 4768 22560 4820
rect 22612 4808 22618 4820
rect 22612 4780 23704 4808
rect 22612 4768 22618 4780
rect 21542 4740 21548 4752
rect 20180 4712 21548 4740
rect 17736 4700 17742 4712
rect 17451 4644 17540 4672
rect 18049 4675 18107 4681
rect 17451 4641 17463 4644
rect 17405 4635 17463 4641
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18598 4672 18604 4684
rect 18095 4644 18604 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 18708 4672 18736 4712
rect 21542 4700 21548 4712
rect 21600 4700 21606 4752
rect 21634 4700 21640 4752
rect 21692 4700 21698 4752
rect 18708 4644 18828 4672
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 12768 4576 13492 4604
rect 12768 4564 12774 4576
rect 12268 4508 12664 4536
rect 13354 4496 13360 4548
rect 13412 4496 13418 4548
rect 13464 4536 13492 4576
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 13909 4607 13967 4613
rect 13909 4604 13921 4607
rect 13596 4576 13921 4604
rect 13596 4564 13602 4576
rect 13909 4573 13921 4576
rect 13955 4573 13967 4607
rect 13909 4567 13967 4573
rect 14090 4564 14096 4616
rect 14148 4564 14154 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 15102 4564 15108 4616
rect 15160 4613 15166 4616
rect 15160 4607 15188 4613
rect 15176 4573 15188 4607
rect 15160 4567 15188 4573
rect 15160 4564 15166 4567
rect 16850 4564 16856 4616
rect 16908 4564 16914 4616
rect 17034 4613 17040 4616
rect 17012 4607 17040 4613
rect 17012 4573 17024 4607
rect 17012 4567 17040 4573
rect 17034 4564 17040 4567
rect 17092 4564 17098 4616
rect 17678 4564 17684 4616
rect 17736 4604 17742 4616
rect 17865 4607 17923 4613
rect 17865 4604 17877 4607
rect 17736 4576 17877 4604
rect 17736 4564 17742 4576
rect 17865 4573 17877 4576
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 13722 4536 13728 4548
rect 13464 4508 13728 4536
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 7616 4440 8616 4468
rect 8757 4471 8815 4477
rect 7616 4428 7622 4440
rect 8757 4437 8769 4471
rect 8803 4468 8815 4471
rect 10778 4468 10784 4480
rect 8803 4440 10784 4468
rect 8803 4437 8815 4440
rect 8757 4431 8815 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 11882 4468 11888 4480
rect 11480 4440 11888 4468
rect 11480 4428 11486 4440
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 11974 4428 11980 4480
rect 12032 4428 12038 4480
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 12434 4468 12440 4480
rect 12308 4440 12440 4468
rect 12308 4428 12314 4440
rect 12434 4428 12440 4440
rect 12492 4468 12498 4480
rect 13262 4468 13268 4480
rect 12492 4440 13268 4468
rect 12492 4428 12498 4440
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 13449 4471 13507 4477
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13630 4468 13636 4480
rect 13495 4440 13636 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 13906 4428 13912 4480
rect 13964 4468 13970 4480
rect 17402 4468 17408 4480
rect 13964 4440 17408 4468
rect 13964 4428 13970 4440
rect 17402 4428 17408 4440
rect 17460 4428 17466 4480
rect 17494 4428 17500 4480
rect 17552 4468 17558 4480
rect 18156 4468 18184 4567
rect 18690 4564 18696 4616
rect 18748 4564 18754 4616
rect 18800 4613 18828 4644
rect 21082 4632 21088 4684
rect 21140 4632 21146 4684
rect 21192 4644 21772 4672
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 19392 4576 19993 4604
rect 19392 4564 19398 4576
rect 19981 4573 19993 4576
rect 20027 4573 20039 4607
rect 19981 4567 20039 4573
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 19242 4536 19248 4548
rect 18524 4508 19248 4536
rect 17552 4440 18184 4468
rect 17552 4428 17558 4440
rect 18322 4428 18328 4480
rect 18380 4428 18386 4480
rect 18524 4477 18552 4508
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 19702 4496 19708 4548
rect 19760 4536 19766 4548
rect 20272 4536 20300 4567
rect 20714 4564 20720 4616
rect 20772 4564 20778 4616
rect 20806 4564 20812 4616
rect 20864 4604 20870 4616
rect 21192 4604 21220 4644
rect 20864 4576 21220 4604
rect 21269 4607 21327 4613
rect 20864 4564 20870 4576
rect 21269 4573 21281 4607
rect 21315 4604 21327 4607
rect 21358 4604 21364 4616
rect 21315 4576 21364 4604
rect 21315 4573 21327 4576
rect 21269 4567 21327 4573
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 19760 4508 20300 4536
rect 20901 4539 20959 4545
rect 19760 4496 19766 4508
rect 20901 4505 20913 4539
rect 20947 4536 20959 4539
rect 21634 4536 21640 4548
rect 20947 4508 21640 4536
rect 20947 4505 20959 4508
rect 20901 4499 20959 4505
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 21744 4536 21772 4644
rect 22646 4632 22652 4684
rect 22704 4632 22710 4684
rect 23676 4672 23704 4780
rect 27430 4768 27436 4820
rect 27488 4768 27494 4820
rect 31110 4808 31116 4820
rect 27816 4780 31116 4808
rect 23753 4743 23811 4749
rect 23753 4709 23765 4743
rect 23799 4740 23811 4743
rect 24210 4740 24216 4752
rect 23799 4712 24216 4740
rect 23799 4709 23811 4712
rect 23753 4703 23811 4709
rect 24210 4700 24216 4712
rect 24268 4700 24274 4752
rect 25130 4700 25136 4752
rect 25188 4700 25194 4752
rect 25866 4700 25872 4752
rect 25924 4740 25930 4752
rect 26237 4743 26295 4749
rect 26237 4740 26249 4743
rect 25924 4712 26249 4740
rect 25924 4700 25930 4712
rect 26237 4709 26249 4712
rect 26283 4709 26295 4743
rect 26237 4703 26295 4709
rect 23676 4644 24808 4672
rect 21818 4564 21824 4616
rect 21876 4604 21882 4616
rect 22373 4607 22431 4613
rect 21876 4576 22324 4604
rect 21876 4564 21882 4576
rect 22094 4536 22100 4548
rect 21744 4508 22100 4536
rect 22094 4496 22100 4508
rect 22152 4496 22158 4548
rect 22296 4536 22324 4576
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 22419 4576 22692 4604
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 22664 4548 22692 4576
rect 22738 4564 22744 4616
rect 22796 4564 22802 4616
rect 22922 4564 22928 4616
rect 22980 4604 22986 4616
rect 23017 4607 23075 4613
rect 23017 4604 23029 4607
rect 22980 4576 23029 4604
rect 22980 4564 22986 4576
rect 23017 4573 23029 4576
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 22554 4536 22560 4548
rect 22296 4508 22560 4536
rect 22554 4496 22560 4508
rect 22612 4496 22618 4548
rect 22646 4496 22652 4548
rect 22704 4496 22710 4548
rect 23032 4536 23060 4567
rect 23106 4564 23112 4616
rect 23164 4604 23170 4616
rect 23845 4607 23903 4613
rect 23845 4604 23857 4607
rect 23164 4576 23857 4604
rect 23164 4564 23170 4576
rect 23845 4573 23857 4576
rect 23891 4573 23903 4607
rect 23845 4567 23903 4573
rect 24394 4564 24400 4616
rect 24452 4564 24458 4616
rect 24780 4613 24808 4644
rect 25148 4613 25176 4700
rect 25774 4632 25780 4684
rect 25832 4632 25838 4684
rect 26142 4632 26148 4684
rect 26200 4672 26206 4684
rect 26513 4675 26571 4681
rect 26513 4672 26525 4675
rect 26200 4644 26525 4672
rect 26200 4632 26206 4644
rect 26513 4641 26525 4644
rect 26559 4672 26571 4675
rect 27430 4672 27436 4684
rect 26559 4644 27436 4672
rect 26559 4641 26571 4644
rect 26513 4635 26571 4641
rect 27430 4632 27436 4644
rect 27488 4632 27494 4684
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 25593 4607 25651 4613
rect 25593 4573 25605 4607
rect 25639 4573 25651 4607
rect 25593 4567 25651 4573
rect 23382 4536 23388 4548
rect 23032 4508 23388 4536
rect 23382 4496 23388 4508
rect 23440 4496 23446 4548
rect 23934 4536 23940 4548
rect 23492 4508 23940 4536
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4437 18567 4471
rect 18509 4431 18567 4437
rect 18969 4471 19027 4477
rect 18969 4437 18981 4471
rect 19015 4468 19027 4471
rect 19150 4468 19156 4480
rect 19015 4440 19156 4468
rect 19015 4437 19027 4440
rect 18969 4431 19027 4437
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 20438 4468 20444 4480
rect 19668 4440 20444 4468
rect 19668 4428 19674 4440
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 20530 4428 20536 4480
rect 20588 4428 20594 4480
rect 21453 4471 21511 4477
rect 21453 4437 21465 4471
rect 21499 4468 21511 4471
rect 21542 4468 21548 4480
rect 21499 4440 21548 4468
rect 21499 4437 21511 4440
rect 21453 4431 21511 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 22370 4428 22376 4480
rect 22428 4468 22434 4480
rect 23492 4468 23520 4508
rect 23934 4496 23940 4508
rect 23992 4496 23998 4548
rect 24302 4496 24308 4548
rect 24360 4536 24366 4548
rect 25222 4536 25228 4548
rect 24360 4508 25228 4536
rect 24360 4496 24366 4508
rect 25222 4496 25228 4508
rect 25280 4496 25286 4548
rect 25608 4536 25636 4567
rect 26602 4564 26608 4616
rect 26660 4613 26666 4616
rect 26660 4607 26688 4613
rect 26676 4573 26688 4607
rect 26660 4567 26688 4573
rect 26660 4564 26666 4567
rect 26786 4564 26792 4616
rect 26844 4564 26850 4616
rect 27816 4613 27844 4780
rect 31110 4768 31116 4780
rect 31168 4768 31174 4820
rect 32398 4808 32404 4820
rect 31680 4780 32404 4808
rect 29454 4700 29460 4752
rect 29512 4740 29518 4752
rect 29512 4712 29960 4740
rect 29512 4700 29518 4712
rect 27890 4632 27896 4684
rect 27948 4632 27954 4684
rect 29270 4632 29276 4684
rect 29328 4672 29334 4684
rect 29822 4672 29828 4684
rect 29328 4644 29828 4672
rect 29328 4632 29334 4644
rect 29822 4632 29828 4644
rect 29880 4632 29886 4684
rect 29932 4672 29960 4712
rect 30006 4700 30012 4752
rect 30064 4700 30070 4752
rect 31202 4700 31208 4752
rect 31260 4740 31266 4752
rect 31260 4712 31524 4740
rect 31260 4700 31266 4712
rect 29932 4644 30420 4672
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 28166 4564 28172 4616
rect 28224 4564 28230 4616
rect 30006 4604 30012 4616
rect 28966 4576 30012 4604
rect 25774 4536 25780 4548
rect 25608 4508 25780 4536
rect 25774 4496 25780 4508
rect 25832 4496 25838 4548
rect 28966 4536 28994 4576
rect 30006 4564 30012 4576
rect 30064 4564 30070 4616
rect 27540 4508 28994 4536
rect 29181 4539 29239 4545
rect 22428 4440 23520 4468
rect 22428 4428 22434 4440
rect 23566 4428 23572 4480
rect 23624 4468 23630 4480
rect 24029 4471 24087 4477
rect 24029 4468 24041 4471
rect 23624 4440 24041 4468
rect 23624 4428 23630 4440
rect 24029 4437 24041 4440
rect 24075 4437 24087 4471
rect 24029 4431 24087 4437
rect 24118 4428 24124 4480
rect 24176 4468 24182 4480
rect 24581 4471 24639 4477
rect 24581 4468 24593 4471
rect 24176 4440 24593 4468
rect 24176 4428 24182 4440
rect 24581 4437 24593 4440
rect 24627 4437 24639 4471
rect 24581 4431 24639 4437
rect 24946 4428 24952 4480
rect 25004 4428 25010 4480
rect 25314 4428 25320 4480
rect 25372 4428 25378 4480
rect 25590 4428 25596 4480
rect 25648 4468 25654 4480
rect 27540 4468 27568 4508
rect 29181 4505 29193 4539
rect 29227 4536 29239 4539
rect 30282 4536 30288 4548
rect 29227 4508 30288 4536
rect 29227 4505 29239 4508
rect 29181 4499 29239 4505
rect 30282 4496 30288 4508
rect 30340 4496 30346 4548
rect 30392 4536 30420 4644
rect 31386 4632 31392 4684
rect 31444 4632 31450 4684
rect 31496 4672 31524 4712
rect 31573 4675 31631 4681
rect 31573 4672 31585 4675
rect 31496 4644 31585 4672
rect 31573 4641 31585 4644
rect 31619 4641 31631 4675
rect 31573 4635 31631 4641
rect 30742 4564 30748 4616
rect 30800 4564 30806 4616
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4604 31079 4607
rect 31110 4604 31116 4616
rect 31067 4576 31116 4604
rect 31067 4573 31079 4576
rect 31021 4567 31079 4573
rect 31110 4564 31116 4576
rect 31168 4564 31174 4616
rect 31680 4604 31708 4780
rect 32398 4768 32404 4780
rect 32456 4768 32462 4820
rect 32766 4768 32772 4820
rect 32824 4808 32830 4820
rect 33229 4811 33287 4817
rect 33229 4808 33241 4811
rect 32824 4780 33241 4808
rect 32824 4768 32830 4780
rect 33229 4777 33241 4780
rect 33275 4777 33287 4811
rect 33229 4771 33287 4777
rect 33321 4811 33379 4817
rect 33321 4777 33333 4811
rect 33367 4808 33379 4811
rect 33686 4808 33692 4820
rect 33367 4780 33692 4808
rect 33367 4777 33379 4780
rect 33321 4771 33379 4777
rect 33686 4768 33692 4780
rect 33744 4768 33750 4820
rect 33870 4768 33876 4820
rect 33928 4808 33934 4820
rect 34422 4808 34428 4820
rect 33928 4780 34428 4808
rect 33928 4768 33934 4780
rect 34422 4768 34428 4780
rect 34480 4768 34486 4820
rect 34514 4768 34520 4820
rect 34572 4808 34578 4820
rect 35158 4808 35164 4820
rect 34572 4780 35164 4808
rect 34572 4768 34578 4780
rect 35158 4768 35164 4780
rect 35216 4808 35222 4820
rect 35989 4811 36047 4817
rect 35989 4808 36001 4811
rect 35216 4780 36001 4808
rect 35216 4768 35222 4780
rect 35989 4777 36001 4780
rect 36035 4777 36047 4811
rect 35989 4771 36047 4777
rect 36630 4768 36636 4820
rect 36688 4808 36694 4820
rect 36817 4811 36875 4817
rect 36817 4808 36829 4811
rect 36688 4780 36829 4808
rect 36688 4768 36694 4780
rect 36817 4777 36829 4780
rect 36863 4777 36875 4811
rect 36817 4771 36875 4777
rect 39390 4768 39396 4820
rect 39448 4768 39454 4820
rect 31846 4700 31852 4752
rect 31904 4740 31910 4752
rect 32033 4743 32091 4749
rect 32033 4740 32045 4743
rect 31904 4712 32045 4740
rect 31904 4700 31910 4712
rect 32033 4709 32045 4712
rect 32079 4709 32091 4743
rect 32033 4703 32091 4709
rect 32122 4632 32128 4684
rect 32180 4672 32186 4684
rect 32309 4675 32367 4681
rect 32309 4672 32321 4675
rect 32180 4644 32321 4672
rect 32180 4632 32186 4644
rect 32309 4641 32321 4644
rect 32355 4641 32367 4675
rect 32309 4635 32367 4641
rect 32398 4632 32404 4684
rect 32456 4681 32462 4684
rect 32456 4675 32484 4681
rect 32472 4641 32484 4675
rect 34333 4675 34391 4681
rect 32456 4635 32484 4641
rect 32456 4632 32462 4635
rect 31220 4576 31708 4604
rect 32582 4598 32588 4650
rect 32640 4598 32646 4650
rect 34333 4641 34345 4675
rect 34379 4672 34391 4675
rect 34422 4672 34428 4684
rect 34379 4644 34428 4672
rect 34379 4641 34391 4644
rect 34333 4635 34391 4641
rect 34422 4632 34428 4644
rect 34480 4632 34486 4684
rect 34057 4607 34115 4613
rect 31220 4536 31248 4576
rect 32585 4573 32597 4598
rect 32631 4573 32643 4598
rect 32585 4567 32643 4573
rect 34057 4573 34069 4607
rect 34103 4604 34115 4607
rect 34790 4604 34796 4616
rect 34103 4576 34796 4604
rect 34103 4573 34115 4576
rect 34057 4567 34115 4573
rect 34790 4564 34796 4576
rect 34848 4564 34854 4616
rect 36998 4564 37004 4616
rect 37056 4564 37062 4616
rect 37090 4564 37096 4616
rect 37148 4604 37154 4616
rect 38841 4607 38899 4613
rect 38841 4604 38853 4607
rect 37148 4576 38853 4604
rect 37148 4564 37154 4576
rect 38841 4573 38853 4576
rect 38887 4573 38899 4607
rect 38841 4567 38899 4573
rect 39206 4564 39212 4616
rect 39264 4564 39270 4616
rect 30392 4508 31248 4536
rect 34698 4496 34704 4548
rect 34756 4496 34762 4548
rect 25648 4440 27568 4468
rect 25648 4428 25654 4440
rect 27614 4428 27620 4480
rect 27672 4428 27678 4480
rect 28902 4428 28908 4480
rect 28960 4428 28966 4480
rect 29086 4428 29092 4480
rect 29144 4468 29150 4480
rect 31110 4468 31116 4480
rect 29144 4440 31116 4468
rect 29144 4428 29150 4440
rect 31110 4428 31116 4440
rect 31168 4428 31174 4480
rect 31294 4428 31300 4480
rect 31352 4468 31358 4480
rect 32214 4468 32220 4480
rect 31352 4440 32220 4468
rect 31352 4428 31358 4440
rect 32214 4428 32220 4440
rect 32272 4428 32278 4480
rect 36906 4428 36912 4480
rect 36964 4468 36970 4480
rect 38286 4468 38292 4480
rect 36964 4440 38292 4468
rect 36964 4428 36970 4440
rect 38286 4428 38292 4440
rect 38344 4428 38350 4480
rect 39025 4471 39083 4477
rect 39025 4437 39037 4471
rect 39071 4468 39083 4471
rect 39298 4468 39304 4480
rect 39071 4440 39304 4468
rect 39071 4437 39083 4440
rect 39025 4431 39083 4437
rect 39298 4428 39304 4440
rect 39356 4428 39362 4480
rect 1104 4378 39836 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 9010 4378
rect 9062 4326 9074 4378
rect 9126 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 15010 4378
rect 15062 4326 15074 4378
rect 15126 4326 15138 4378
rect 15190 4326 15202 4378
rect 15254 4326 15266 4378
rect 15318 4326 21010 4378
rect 21062 4326 21074 4378
rect 21126 4326 21138 4378
rect 21190 4326 21202 4378
rect 21254 4326 21266 4378
rect 21318 4326 27010 4378
rect 27062 4326 27074 4378
rect 27126 4326 27138 4378
rect 27190 4326 27202 4378
rect 27254 4326 27266 4378
rect 27318 4326 33010 4378
rect 33062 4326 33074 4378
rect 33126 4326 33138 4378
rect 33190 4326 33202 4378
rect 33254 4326 33266 4378
rect 33318 4326 39010 4378
rect 39062 4326 39074 4378
rect 39126 4326 39138 4378
rect 39190 4326 39202 4378
rect 39254 4326 39266 4378
rect 39318 4326 39836 4378
rect 1104 4304 39836 4326
rect 1949 4267 2007 4273
rect 1949 4233 1961 4267
rect 1995 4264 2007 4267
rect 1995 4236 2636 4264
rect 1995 4233 2007 4236
rect 1949 4227 2007 4233
rect 1486 4156 1492 4208
rect 1544 4156 1550 4208
rect 1854 4156 1860 4208
rect 1912 4156 1918 4208
rect 2498 4156 2504 4208
rect 2556 4156 2562 4208
rect 2608 4196 2636 4236
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3326 4264 3332 4276
rect 2740 4236 3332 4264
rect 2740 4224 2746 4236
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3510 4224 3516 4276
rect 3568 4224 3574 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 4488 4236 5396 4264
rect 4488 4224 4494 4236
rect 3142 4196 3148 4208
rect 2608 4168 3148 4196
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 5368 4196 5396 4236
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 5684 4236 7052 4264
rect 5684 4224 5690 4236
rect 5644 4196 5672 4224
rect 5368 4168 5672 4196
rect 5997 4199 6055 4205
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1946 4128 1952 4140
rect 1719 4100 1952 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2516 4128 2544 4156
rect 2179 4100 2544 4128
rect 2685 4131 2743 4137
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 4338 4137 4344 4140
rect 4316 4131 4344 4137
rect 4316 4097 4328 4131
rect 4316 4091 4344 4097
rect 4338 4088 4344 4091
rect 4396 4088 4402 4140
rect 5368 4137 5396 4168
rect 5997 4165 6009 4199
rect 6043 4196 6055 4199
rect 6178 4196 6184 4208
rect 6043 4168 6184 4196
rect 6043 4165 6055 4168
rect 5997 4159 6055 4165
rect 6178 4156 6184 4168
rect 6236 4156 6242 4208
rect 7024 4196 7052 4236
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 7285 4267 7343 4273
rect 7285 4264 7297 4267
rect 7156 4236 7297 4264
rect 7156 4224 7162 4236
rect 7285 4233 7297 4236
rect 7331 4233 7343 4267
rect 7285 4227 7343 4233
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 9030 4264 9036 4276
rect 7432 4236 9036 4264
rect 7432 4224 7438 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10318 4264 10324 4276
rect 10008 4236 10324 4264
rect 10008 4224 10014 4236
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 11793 4267 11851 4273
rect 11793 4233 11805 4267
rect 11839 4264 11851 4267
rect 11974 4264 11980 4276
rect 11839 4236 11980 4264
rect 11839 4233 11851 4236
rect 11793 4227 11851 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 14461 4267 14519 4273
rect 12584 4236 13216 4264
rect 12584 4224 12590 4236
rect 6380 4168 6776 4196
rect 7024 4168 8340 4196
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 5718 4128 5724 4140
rect 5675 4100 5724 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 5718 4088 5724 4100
rect 5776 4128 5782 4140
rect 6380 4128 6408 4168
rect 5776 4100 6408 4128
rect 5776 4088 5782 4100
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 6564 4100 6653 4128
rect 2314 4020 2320 4072
rect 2372 4060 2378 4072
rect 2409 4063 2467 4069
rect 2409 4060 2421 4063
rect 2372 4032 2421 4060
rect 2372 4020 2378 4032
rect 2409 4029 2421 4032
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 4157 4063 4215 4069
rect 4157 4060 4169 4063
rect 3660 4032 4169 4060
rect 3660 4020 3666 4032
rect 4157 4029 4169 4032
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4798 4060 4804 4072
rect 4479 4032 4804 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5132 4032 5181 4060
rect 5132 4020 5138 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 6564 4060 6592 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 5500 4032 6592 4060
rect 5500 4020 5506 4032
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3961 4767 3995
rect 4709 3955 4767 3961
rect 6181 3995 6239 4001
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 6549 3995 6607 4001
rect 6549 3992 6561 3995
rect 6227 3964 6561 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6549 3961 6561 3964
rect 6595 3961 6607 3995
rect 6549 3955 6607 3961
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 3234 3924 3240 3936
rect 2363 3896 3240 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 4724 3924 4752 3955
rect 3467 3896 4752 3924
rect 5997 3927 6055 3933
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6086 3924 6092 3936
rect 6043 3896 6092 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6454 3884 6460 3936
rect 6512 3884 6518 3936
rect 6748 3924 6776 4168
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 6840 4060 6868 4091
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7708 4100 8217 4128
rect 7708 4088 7714 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8312 4128 8340 4168
rect 9122 4156 9128 4208
rect 9180 4156 9186 4208
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 13081 4199 13139 4205
rect 13081 4196 13093 4199
rect 11664 4168 13093 4196
rect 11664 4156 11670 4168
rect 13081 4165 13093 4168
rect 13127 4165 13139 4199
rect 13188 4196 13216 4236
rect 14461 4233 14473 4267
rect 14507 4264 14519 4267
rect 14734 4264 14740 4276
rect 14507 4236 14740 4264
rect 14507 4233 14519 4236
rect 14461 4227 14519 4233
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 15010 4224 15016 4276
rect 15068 4264 15074 4276
rect 16666 4264 16672 4276
rect 15068 4236 16672 4264
rect 15068 4224 15074 4236
rect 16666 4224 16672 4236
rect 16724 4264 16730 4276
rect 22189 4267 22247 4273
rect 16724 4236 21956 4264
rect 16724 4224 16730 4236
rect 17034 4196 17040 4208
rect 13188 4168 17040 4196
rect 13081 4159 13139 4165
rect 17034 4156 17040 4168
rect 17092 4196 17098 4208
rect 20533 4199 20591 4205
rect 17092 4168 18920 4196
rect 17092 4156 17098 4168
rect 9490 4128 9496 4140
rect 8312 4100 9496 4128
rect 8205 4091 8263 4097
rect 9490 4088 9496 4100
rect 9548 4128 9554 4140
rect 9548 4100 9628 4128
rect 9548 4088 9554 4100
rect 6840 4032 6960 4060
rect 6932 4001 6960 4032
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7377 4063 7435 4069
rect 7377 4060 7389 4063
rect 7156 4032 7389 4060
rect 7156 4020 7162 4032
rect 7377 4029 7389 4032
rect 7423 4029 7435 4063
rect 7377 4023 7435 4029
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 6917 3995 6975 4001
rect 6917 3961 6929 3995
rect 6963 3961 6975 3995
rect 7484 3992 7512 4023
rect 7558 3992 7564 4004
rect 6917 3955 6975 3961
rect 7392 3964 7564 3992
rect 7392 3924 7420 3964
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 6748 3896 7420 3924
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7944 3924 7972 4023
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 9398 4060 9404 4072
rect 8996 4032 9404 4060
rect 8996 4020 9002 4032
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 9600 4069 9628 4100
rect 10318 4088 10324 4140
rect 10376 4088 10382 4140
rect 10502 4137 10508 4140
rect 10459 4131 10508 4137
rect 10459 4097 10471 4131
rect 10505 4097 10508 4131
rect 10459 4091 10508 4097
rect 10502 4088 10508 4091
rect 10560 4088 10566 4140
rect 11241 4131 11299 4137
rect 11241 4097 11253 4131
rect 11287 4128 11299 4131
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11287 4100 11897 4128
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 12216 4100 12357 4128
rect 12216 4088 12222 4100
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12618 4088 12624 4140
rect 12676 4088 12682 4140
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12768 4100 12909 4128
rect 12768 4088 12774 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13320 4100 13737 4128
rect 13320 4088 13326 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 15006 4131 15064 4137
rect 15006 4097 15018 4131
rect 15052 4097 15064 4131
rect 15006 4091 15064 4097
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4029 9643 4063
rect 9585 4023 9643 4029
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 9732 4032 10057 4060
rect 9732 4020 9738 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 10045 4023 10103 4029
rect 10594 4020 10600 4072
rect 10652 4020 10658 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 11701 4063 11759 4069
rect 10836 4032 11008 4060
rect 10836 4020 10842 4032
rect 8846 3952 8852 4004
rect 8904 3992 8910 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8904 3964 9321 3992
rect 8904 3952 8910 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 10980 3992 11008 4032
rect 11701 4029 11713 4063
rect 11747 4060 11759 4063
rect 12176 4060 12204 4088
rect 11747 4032 12204 4060
rect 11747 4029 11759 4032
rect 11701 4023 11759 4029
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13412 4032 13461 4060
rect 13412 4020 13418 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13449 4023 13507 4029
rect 12437 3995 12495 4001
rect 12437 3992 12449 3995
rect 10980 3964 12449 3992
rect 9309 3955 9367 3961
rect 12437 3961 12449 3964
rect 12483 3961 12495 3995
rect 12437 3955 12495 3961
rect 7524 3896 7972 3924
rect 7524 3884 7530 3896
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8076 3896 8953 3924
rect 8076 3884 8082 3896
rect 8941 3893 8953 3896
rect 8987 3924 8999 3927
rect 10594 3924 10600 3936
rect 8987 3896 10600 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 10594 3884 10600 3896
rect 10652 3924 10658 3936
rect 11054 3924 11060 3936
rect 10652 3896 11060 3924
rect 10652 3884 10658 3896
rect 11054 3884 11060 3896
rect 11112 3924 11118 3936
rect 11330 3924 11336 3936
rect 11112 3896 11336 3924
rect 11112 3884 11118 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12253 3927 12311 3933
rect 12253 3924 12265 3927
rect 12032 3896 12265 3924
rect 12032 3884 12038 3896
rect 12253 3893 12265 3896
rect 12299 3893 12311 3927
rect 12253 3887 12311 3893
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 12676 3896 12817 3924
rect 12676 3884 12682 3896
rect 12805 3893 12817 3896
rect 12851 3893 12863 3927
rect 12805 3887 12863 3893
rect 13262 3884 13268 3936
rect 13320 3884 13326 3936
rect 14458 3884 14464 3936
rect 14516 3924 14522 3936
rect 14829 3927 14887 3933
rect 14829 3924 14841 3927
rect 14516 3896 14841 3924
rect 14516 3884 14522 3896
rect 14829 3893 14841 3896
rect 14875 3893 14887 3927
rect 15028 3924 15056 4091
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 15304 4100 15761 4128
rect 15102 4020 15108 4072
rect 15160 4060 15166 4072
rect 15304 4060 15332 4100
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 16206 4088 16212 4140
rect 16264 4128 16270 4140
rect 16574 4128 16580 4140
rect 16264 4100 16580 4128
rect 16264 4088 16270 4100
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 17126 4088 17132 4140
rect 17184 4088 17190 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4128 17555 4131
rect 17770 4128 17776 4140
rect 17543 4100 17776 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 18892 4137 18920 4168
rect 20533 4165 20545 4199
rect 20579 4196 20591 4199
rect 20622 4196 20628 4208
rect 20579 4168 20628 4196
rect 20579 4165 20591 4168
rect 20533 4159 20591 4165
rect 20622 4156 20628 4168
rect 20680 4156 20686 4208
rect 20898 4156 20904 4208
rect 20956 4196 20962 4208
rect 20956 4168 21588 4196
rect 20956 4156 20962 4168
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 19610 4088 19616 4140
rect 19668 4088 19674 4140
rect 21450 4088 21456 4140
rect 21508 4088 21514 4140
rect 21560 4128 21588 4168
rect 21634 4156 21640 4208
rect 21692 4156 21698 4208
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21560 4100 21833 4128
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 15160 4032 15332 4060
rect 15381 4063 15439 4069
rect 15160 4020 15166 4032
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 15470 4060 15476 4072
rect 15427 4032 15476 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 17586 4060 17592 4072
rect 16172 4032 17592 4060
rect 16172 4020 16178 4032
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 18690 4020 18696 4072
rect 18748 4020 18754 4072
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19730 4063 19788 4069
rect 19730 4060 19742 4063
rect 19484 4032 19742 4060
rect 19484 4020 19490 4032
rect 19730 4029 19742 4032
rect 19776 4029 19788 4063
rect 19730 4023 19788 4029
rect 19886 4020 19892 4072
rect 19944 4020 19950 4072
rect 21177 4063 21235 4069
rect 21177 4029 21189 4063
rect 21223 4060 21235 4063
rect 21726 4060 21732 4072
rect 21223 4032 21732 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 21928 4060 21956 4236
rect 22189 4233 22201 4267
rect 22235 4264 22247 4267
rect 22462 4264 22468 4276
rect 22235 4236 22468 4264
rect 22235 4233 22247 4236
rect 22189 4227 22247 4233
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 22554 4224 22560 4276
rect 22612 4224 22618 4276
rect 24302 4264 24308 4276
rect 23216 4236 24308 4264
rect 22830 4196 22836 4208
rect 22480 4168 22836 4196
rect 22480 4140 22508 4168
rect 22830 4156 22836 4168
rect 22888 4156 22894 4208
rect 22462 4088 22468 4140
rect 22520 4088 22526 4140
rect 23017 4131 23075 4137
rect 23017 4097 23029 4131
rect 23063 4128 23075 4131
rect 23216 4128 23244 4236
rect 24302 4224 24308 4236
rect 24360 4224 24366 4276
rect 25038 4264 25044 4276
rect 24964 4236 25044 4264
rect 23063 4100 23244 4128
rect 23063 4097 23075 4100
rect 23017 4091 23075 4097
rect 24210 4088 24216 4140
rect 24268 4088 24274 4140
rect 24854 4088 24860 4140
rect 24912 4088 24918 4140
rect 24964 4128 24992 4236
rect 25038 4224 25044 4236
rect 25096 4264 25102 4276
rect 29086 4264 29092 4276
rect 25096 4236 29092 4264
rect 25096 4224 25102 4236
rect 29086 4224 29092 4236
rect 29144 4224 29150 4276
rect 29178 4224 29184 4276
rect 29236 4264 29242 4276
rect 30285 4267 30343 4273
rect 30285 4264 30297 4267
rect 29236 4236 30297 4264
rect 29236 4224 29242 4236
rect 30285 4233 30297 4236
rect 30331 4233 30343 4267
rect 30285 4227 30343 4233
rect 30650 4224 30656 4276
rect 30708 4264 30714 4276
rect 31662 4264 31668 4276
rect 30708 4236 31668 4264
rect 30708 4224 30714 4236
rect 31662 4224 31668 4236
rect 31720 4224 31726 4276
rect 31754 4224 31760 4276
rect 31812 4264 31818 4276
rect 32490 4264 32496 4276
rect 31812 4236 32496 4264
rect 31812 4224 31818 4236
rect 32490 4224 32496 4236
rect 32548 4224 32554 4276
rect 38838 4264 38844 4276
rect 33244 4236 38844 4264
rect 25774 4156 25780 4208
rect 25832 4196 25838 4208
rect 26326 4196 26332 4208
rect 25832 4168 26332 4196
rect 25832 4156 25838 4168
rect 26326 4156 26332 4168
rect 26384 4156 26390 4208
rect 26786 4196 26792 4208
rect 26436 4168 26792 4196
rect 25041 4131 25099 4137
rect 25041 4128 25053 4131
rect 24964 4100 25053 4128
rect 25041 4097 25053 4100
rect 25087 4097 25099 4131
rect 25041 4091 25099 4097
rect 25222 4088 25228 4140
rect 25280 4128 25286 4140
rect 25317 4131 25375 4137
rect 25317 4128 25329 4131
rect 25280 4100 25329 4128
rect 25280 4088 25286 4100
rect 25317 4097 25329 4100
rect 25363 4097 25375 4131
rect 25317 4091 25375 4097
rect 25406 4088 25412 4140
rect 25464 4128 25470 4140
rect 25464 4100 25636 4128
rect 25464 4088 25470 4100
rect 22649 4063 22707 4069
rect 21928 4032 22600 4060
rect 16574 3992 16580 4004
rect 16316 3964 16580 3992
rect 16316 3924 16344 3964
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 16945 3995 17003 4001
rect 16945 3961 16957 3995
rect 16991 3992 17003 3995
rect 18601 3995 18659 4001
rect 16991 3964 17724 3992
rect 16991 3961 17003 3964
rect 16945 3955 17003 3961
rect 15028 3896 16344 3924
rect 14829 3887 14887 3893
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16485 3927 16543 3933
rect 16485 3924 16497 3927
rect 16448 3896 16497 3924
rect 16448 3884 16454 3896
rect 16485 3893 16497 3896
rect 16531 3893 16543 3927
rect 16485 3887 16543 3893
rect 17313 3927 17371 3933
rect 17313 3893 17325 3927
rect 17359 3924 17371 3927
rect 17586 3924 17592 3936
rect 17359 3896 17592 3924
rect 17359 3893 17371 3896
rect 17313 3887 17371 3893
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 17696 3924 17724 3964
rect 18601 3961 18613 3995
rect 18647 3992 18659 3995
rect 19337 3995 19395 4001
rect 19337 3992 19349 3995
rect 18647 3964 19349 3992
rect 18647 3961 18659 3964
rect 18601 3955 18659 3961
rect 19337 3961 19349 3964
rect 19383 3961 19395 3995
rect 19337 3955 19395 3961
rect 20806 3952 20812 4004
rect 20864 3992 20870 4004
rect 22370 3992 22376 4004
rect 20864 3964 22376 3992
rect 20864 3952 20870 3964
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 18414 3924 18420 3936
rect 17696 3896 18420 3924
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 21726 3924 21732 3936
rect 18564 3896 21732 3924
rect 18564 3884 18570 3896
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 21818 3884 21824 3936
rect 21876 3924 21882 3936
rect 22005 3927 22063 3933
rect 22005 3924 22017 3927
rect 21876 3896 22017 3924
rect 21876 3884 21882 3896
rect 22005 3893 22017 3896
rect 22051 3893 22063 3927
rect 22572 3924 22600 4032
rect 22649 4029 22661 4063
rect 22695 4029 22707 4063
rect 22649 4023 22707 4029
rect 22664 3992 22692 4023
rect 22830 4020 22836 4072
rect 22888 4020 22894 4072
rect 23201 4063 23259 4069
rect 23201 4029 23213 4063
rect 23247 4060 23259 4063
rect 23290 4060 23296 4072
rect 23247 4032 23296 4060
rect 23247 4029 23259 4032
rect 23201 4023 23259 4029
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 23658 4020 23664 4072
rect 23716 4020 23722 4072
rect 23934 4060 23940 4072
rect 23768 4032 23940 4060
rect 23768 3992 23796 4032
rect 23934 4020 23940 4032
rect 23992 4020 23998 4072
rect 24026 4020 24032 4072
rect 24084 4069 24090 4072
rect 24084 4063 24112 4069
rect 24100 4029 24112 4063
rect 25608 4060 25636 4100
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 26145 4131 26203 4137
rect 26145 4128 26157 4131
rect 25740 4100 26157 4128
rect 25740 4088 25746 4100
rect 26145 4097 26157 4100
rect 26191 4097 26203 4131
rect 26145 4091 26203 4097
rect 26234 4088 26240 4140
rect 26292 4128 26298 4140
rect 26436 4128 26464 4168
rect 26786 4156 26792 4168
rect 26844 4156 26850 4208
rect 27154 4156 27160 4208
rect 27212 4196 27218 4208
rect 27212 4168 27384 4196
rect 27212 4156 27218 4168
rect 26292 4100 26464 4128
rect 26292 4088 26298 4100
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 26602 4088 26608 4140
rect 26660 4128 26666 4140
rect 27249 4131 27307 4137
rect 27249 4128 27261 4131
rect 26660 4100 27261 4128
rect 26660 4088 26666 4100
rect 27249 4097 27261 4100
rect 27295 4097 27307 4131
rect 27356 4128 27384 4168
rect 30098 4156 30104 4208
rect 30156 4196 30162 4208
rect 30834 4196 30840 4208
rect 30156 4168 30840 4196
rect 30156 4156 30162 4168
rect 30834 4156 30840 4168
rect 30892 4196 30898 4208
rect 30892 4168 31064 4196
rect 30892 4156 30898 4168
rect 27356 4100 27568 4128
rect 27249 4091 27307 4097
rect 26418 4060 26424 4072
rect 25608 4032 26424 4060
rect 24084 4023 24112 4029
rect 24084 4020 24090 4023
rect 26418 4020 26424 4032
rect 26476 4020 26482 4072
rect 26973 4063 27031 4069
rect 26973 4029 26985 4063
rect 27019 4029 27031 4063
rect 27540 4060 27568 4100
rect 27614 4088 27620 4140
rect 27672 4128 27678 4140
rect 28261 4131 28319 4137
rect 28261 4128 28273 4131
rect 27672 4100 28273 4128
rect 27672 4088 27678 4100
rect 28261 4097 28273 4100
rect 28307 4097 28319 4131
rect 28261 4091 28319 4097
rect 29546 4088 29552 4140
rect 29604 4088 29610 4140
rect 30193 4131 30251 4137
rect 30193 4097 30205 4131
rect 30239 4128 30251 4131
rect 30926 4128 30932 4140
rect 30239 4100 30932 4128
rect 30239 4097 30251 4100
rect 30193 4091 30251 4097
rect 30926 4088 30932 4100
rect 30984 4088 30990 4140
rect 31036 4137 31064 4168
rect 31478 4156 31484 4208
rect 31536 4196 31542 4208
rect 33134 4196 33140 4208
rect 31536 4168 33140 4196
rect 31536 4156 31542 4168
rect 33134 4156 33140 4168
rect 33192 4156 33198 4208
rect 31021 4131 31079 4137
rect 31021 4097 31033 4131
rect 31067 4097 31079 4131
rect 31021 4091 31079 4097
rect 31110 4088 31116 4140
rect 31168 4128 31174 4140
rect 31297 4131 31355 4137
rect 31297 4128 31309 4131
rect 31168 4100 31309 4128
rect 31168 4088 31174 4100
rect 31297 4097 31309 4100
rect 31343 4097 31355 4131
rect 31297 4091 31355 4097
rect 31386 4088 31392 4140
rect 31444 4088 31450 4140
rect 31570 4088 31576 4140
rect 31628 4128 31634 4140
rect 32048 4137 32168 4138
rect 32048 4131 32183 4137
rect 32048 4128 32137 4131
rect 31628 4110 32137 4128
rect 31628 4100 32076 4110
rect 31628 4088 31634 4100
rect 32125 4097 32137 4110
rect 32171 4097 32183 4131
rect 32125 4091 32183 4097
rect 32490 4088 32496 4140
rect 32548 4088 32554 4140
rect 28353 4063 28411 4069
rect 27540 4032 27936 4060
rect 26973 4023 27031 4029
rect 22664 3964 23796 3992
rect 26053 3995 26111 4001
rect 26053 3961 26065 3995
rect 26099 3992 26111 3995
rect 26234 3992 26240 4004
rect 26099 3964 26240 3992
rect 26099 3961 26111 3964
rect 26053 3955 26111 3961
rect 26234 3952 26240 3964
rect 26292 3952 26298 4004
rect 24026 3924 24032 3936
rect 22572 3896 24032 3924
rect 22005 3887 22063 3893
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 25682 3924 25688 3936
rect 24268 3896 25688 3924
rect 24268 3884 24274 3896
rect 25682 3884 25688 3896
rect 25740 3924 25746 3936
rect 26142 3924 26148 3936
rect 25740 3896 26148 3924
rect 25740 3884 25746 3896
rect 26142 3884 26148 3896
rect 26200 3884 26206 3936
rect 26326 3884 26332 3936
rect 26384 3884 26390 3936
rect 26694 3884 26700 3936
rect 26752 3884 26758 3936
rect 26988 3924 27016 4023
rect 27798 3924 27804 3936
rect 26988 3896 27804 3924
rect 27798 3884 27804 3896
rect 27856 3884 27862 3936
rect 27908 3924 27936 4032
rect 28353 4029 28365 4063
rect 28399 4029 28411 4063
rect 28353 4023 28411 4029
rect 27985 3995 28043 4001
rect 27985 3961 27997 3995
rect 28031 3992 28043 3995
rect 28166 3992 28172 4004
rect 28031 3964 28172 3992
rect 28031 3961 28043 3964
rect 27985 3955 28043 3961
rect 28166 3952 28172 3964
rect 28224 3952 28230 4004
rect 28258 3952 28264 4004
rect 28316 3992 28322 4004
rect 28368 3992 28396 4023
rect 28442 4020 28448 4072
rect 28500 4060 28506 4072
rect 28537 4063 28595 4069
rect 28537 4060 28549 4063
rect 28500 4032 28549 4060
rect 28500 4020 28506 4032
rect 28537 4029 28549 4032
rect 28583 4029 28595 4063
rect 28537 4023 28595 4029
rect 28902 4020 28908 4072
rect 28960 4060 28966 4072
rect 28997 4063 29055 4069
rect 28997 4060 29009 4063
rect 28960 4032 29009 4060
rect 28960 4020 28966 4032
rect 28997 4029 29009 4032
rect 29043 4029 29055 4063
rect 28997 4023 29055 4029
rect 29086 4020 29092 4072
rect 29144 4060 29150 4072
rect 29273 4063 29331 4069
rect 29273 4060 29285 4063
rect 29144 4032 29285 4060
rect 29144 4020 29150 4032
rect 29273 4029 29285 4032
rect 29319 4029 29331 4063
rect 29273 4023 29331 4029
rect 29411 4063 29469 4069
rect 29411 4029 29423 4063
rect 29457 4060 29469 4063
rect 29914 4060 29920 4072
rect 29457 4032 29920 4060
rect 29457 4029 29469 4032
rect 29411 4023 29469 4029
rect 29914 4020 29920 4032
rect 29972 4020 29978 4072
rect 32214 4020 32220 4072
rect 32272 4060 32278 4072
rect 33244 4060 33272 4236
rect 38838 4224 38844 4236
rect 38896 4224 38902 4276
rect 34330 4156 34336 4208
rect 34388 4196 34394 4208
rect 36081 4199 36139 4205
rect 36081 4196 36093 4199
rect 34388 4168 36093 4196
rect 34388 4156 34394 4168
rect 36081 4165 36093 4168
rect 36127 4165 36139 4199
rect 36081 4159 36139 4165
rect 36354 4156 36360 4208
rect 36412 4196 36418 4208
rect 38286 4196 38292 4208
rect 36412 4168 38292 4196
rect 36412 4156 36418 4168
rect 38286 4156 38292 4168
rect 38344 4156 38350 4208
rect 33318 4088 33324 4140
rect 33376 4128 33382 4140
rect 33686 4128 33692 4140
rect 33376 4100 33692 4128
rect 33376 4088 33382 4100
rect 33686 4088 33692 4100
rect 33744 4128 33750 4140
rect 34066 4131 34124 4137
rect 34066 4128 34078 4131
rect 33744 4100 34078 4128
rect 33744 4088 33750 4100
rect 34066 4097 34078 4100
rect 34112 4097 34124 4131
rect 34066 4091 34124 4097
rect 34238 4088 34244 4140
rect 34296 4128 34302 4140
rect 34609 4131 34667 4137
rect 34609 4128 34621 4131
rect 34296 4100 34621 4128
rect 34296 4088 34302 4100
rect 34609 4097 34621 4100
rect 34655 4097 34667 4131
rect 34609 4091 34667 4097
rect 34977 4131 35035 4137
rect 34977 4097 34989 4131
rect 35023 4128 35035 4131
rect 35066 4128 35072 4140
rect 35023 4100 35072 4128
rect 35023 4097 35035 4100
rect 34977 4091 35035 4097
rect 35066 4088 35072 4100
rect 35124 4088 35130 4140
rect 36170 4088 36176 4140
rect 36228 4088 36234 4140
rect 36817 4131 36875 4137
rect 36817 4128 36829 4131
rect 36464 4100 36829 4128
rect 32272 4032 33272 4060
rect 32272 4020 32278 4032
rect 34330 4020 34336 4072
rect 34388 4020 34394 4072
rect 34514 4020 34520 4072
rect 34572 4060 34578 4072
rect 34701 4063 34759 4069
rect 34701 4060 34713 4063
rect 34572 4032 34713 4060
rect 34572 4020 34578 4032
rect 34701 4029 34713 4032
rect 34747 4029 34759 4063
rect 34701 4023 34759 4029
rect 35897 4063 35955 4069
rect 35897 4029 35909 4063
rect 35943 4029 35955 4063
rect 35897 4023 35955 4029
rect 28316 3964 28396 3992
rect 28316 3952 28322 3964
rect 32122 3952 32128 4004
rect 32180 3992 32186 4004
rect 32582 3992 32588 4004
rect 32180 3964 32588 3992
rect 32180 3952 32186 3964
rect 32582 3952 32588 3964
rect 32640 3992 32646 4004
rect 32953 3995 33011 4001
rect 32953 3992 32965 3995
rect 32640 3964 32965 3992
rect 32640 3952 32646 3964
rect 32953 3961 32965 3964
rect 32999 3961 33011 3995
rect 32953 3955 33011 3961
rect 35713 3995 35771 4001
rect 35713 3961 35725 3995
rect 35759 3992 35771 3995
rect 35912 3992 35940 4023
rect 35759 3964 35940 3992
rect 36464 3992 36492 4100
rect 36817 4097 36829 4100
rect 36863 4097 36875 4131
rect 36817 4091 36875 4097
rect 37182 4088 37188 4140
rect 37240 4128 37246 4140
rect 38746 4128 38752 4140
rect 37240 4100 38752 4128
rect 37240 4088 37246 4100
rect 38746 4088 38752 4100
rect 38804 4088 38810 4140
rect 38841 4131 38899 4137
rect 38841 4097 38853 4131
rect 38887 4097 38899 4131
rect 38841 4091 38899 4097
rect 36541 3995 36599 4001
rect 36541 3992 36553 3995
rect 36464 3964 36553 3992
rect 35759 3961 35771 3964
rect 35713 3955 35771 3961
rect 36541 3961 36553 3964
rect 36587 3961 36599 3995
rect 36541 3955 36599 3961
rect 37274 3952 37280 4004
rect 37332 3992 37338 4004
rect 38856 3992 38884 4091
rect 39114 4088 39120 4140
rect 39172 4128 39178 4140
rect 39209 4131 39267 4137
rect 39209 4128 39221 4131
rect 39172 4100 39221 4128
rect 39172 4088 39178 4100
rect 39209 4097 39221 4100
rect 39255 4097 39267 4131
rect 39209 4091 39267 4097
rect 37332 3964 38884 3992
rect 39393 3995 39451 4001
rect 37332 3952 37338 3964
rect 39393 3961 39405 3995
rect 39439 3992 39451 3995
rect 39482 3992 39488 4004
rect 39439 3964 39488 3992
rect 39439 3961 39451 3964
rect 39393 3955 39451 3961
rect 39482 3952 39488 3964
rect 39540 3952 39546 4004
rect 28077 3927 28135 3933
rect 28077 3924 28089 3927
rect 27908 3896 28089 3924
rect 28077 3893 28089 3896
rect 28123 3893 28135 3927
rect 28077 3887 28135 3893
rect 29638 3884 29644 3936
rect 29696 3924 29702 3936
rect 30466 3924 30472 3936
rect 29696 3896 30472 3924
rect 29696 3884 29702 3896
rect 30466 3884 30472 3896
rect 30524 3924 30530 3936
rect 30834 3924 30840 3936
rect 30524 3896 30840 3924
rect 30524 3884 30530 3896
rect 30834 3884 30840 3896
rect 30892 3884 30898 3936
rect 31570 3884 31576 3936
rect 31628 3884 31634 3936
rect 32306 3884 32312 3936
rect 32364 3884 32370 3936
rect 32674 3884 32680 3936
rect 32732 3884 32738 3936
rect 34054 3884 34060 3936
rect 34112 3924 34118 3936
rect 34425 3927 34483 3933
rect 34425 3924 34437 3927
rect 34112 3896 34437 3924
rect 34112 3884 34118 3896
rect 34425 3893 34437 3896
rect 34471 3893 34483 3927
rect 34425 3887 34483 3893
rect 36630 3884 36636 3936
rect 36688 3884 36694 3936
rect 39022 3884 39028 3936
rect 39080 3884 39086 3936
rect 1104 3834 39836 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 13950 3834
rect 14002 3782 14014 3834
rect 14066 3782 14078 3834
rect 14130 3782 14142 3834
rect 14194 3782 14206 3834
rect 14258 3782 19950 3834
rect 20002 3782 20014 3834
rect 20066 3782 20078 3834
rect 20130 3782 20142 3834
rect 20194 3782 20206 3834
rect 20258 3782 25950 3834
rect 26002 3782 26014 3834
rect 26066 3782 26078 3834
rect 26130 3782 26142 3834
rect 26194 3782 26206 3834
rect 26258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 37950 3834
rect 38002 3782 38014 3834
rect 38066 3782 38078 3834
rect 38130 3782 38142 3834
rect 38194 3782 38206 3834
rect 38258 3782 39836 3834
rect 1104 3760 39836 3782
rect 1118 3680 1124 3732
rect 1176 3720 1182 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 1176 3692 1593 3720
rect 1176 3680 1182 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 1581 3683 1639 3689
rect 3602 3680 3608 3732
rect 3660 3680 3666 3732
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 4663 3692 6776 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 2041 3655 2099 3661
rect 2041 3652 2053 3655
rect 1728 3624 2053 3652
rect 1728 3612 1734 3624
rect 2041 3621 2053 3624
rect 2087 3621 2099 3655
rect 2041 3615 2099 3621
rect 6089 3655 6147 3661
rect 6089 3621 6101 3655
rect 6135 3652 6147 3655
rect 6546 3652 6552 3664
rect 6135 3624 6552 3652
rect 6135 3621 6147 3624
rect 6089 3615 6147 3621
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 6748 3652 6776 3692
rect 6822 3680 6828 3732
rect 6880 3680 6886 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7432 3692 7665 3720
rect 7432 3680 7438 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 7837 3723 7895 3729
rect 7837 3689 7849 3723
rect 7883 3720 7895 3723
rect 7926 3720 7932 3732
rect 7883 3692 7932 3720
rect 7883 3689 7895 3692
rect 7837 3683 7895 3689
rect 7668 3652 7696 3683
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 8444 3692 8585 3720
rect 8444 3680 8450 3692
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 8573 3683 8631 3689
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9306 3720 9312 3732
rect 8904 3692 9312 3720
rect 8904 3680 8910 3692
rect 9306 3680 9312 3692
rect 9364 3720 9370 3732
rect 11701 3723 11759 3729
rect 9364 3692 11468 3720
rect 9364 3680 9370 3692
rect 8662 3652 8668 3664
rect 6748 3624 7512 3652
rect 7668 3624 8668 3652
rect 1302 3544 1308 3596
rect 1360 3584 1366 3596
rect 1360 3556 2268 3584
rect 1360 3544 1366 3556
rect 1486 3476 1492 3528
rect 1544 3476 1550 3528
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2130 3516 2136 3528
rect 1903 3488 2136 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2240 3516 2268 3556
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2593 3587 2651 3593
rect 2593 3584 2605 3587
rect 2372 3556 2605 3584
rect 2372 3544 2378 3556
rect 2593 3553 2605 3556
rect 2639 3553 2651 3587
rect 4890 3584 4896 3596
rect 2593 3547 2651 3553
rect 4264 3556 4896 3584
rect 2869 3519 2927 3525
rect 2240 3488 2820 3516
rect 2222 3408 2228 3460
rect 2280 3408 2286 3460
rect 2409 3451 2467 3457
rect 2409 3417 2421 3451
rect 2455 3448 2467 3451
rect 2682 3448 2688 3460
rect 2455 3420 2688 3448
rect 2455 3417 2467 3420
rect 2409 3411 2467 3417
rect 2682 3408 2688 3420
rect 2740 3408 2746 3460
rect 2792 3448 2820 3488
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 3881 3519 3939 3525
rect 3881 3518 3893 3519
rect 3804 3516 3893 3518
rect 2915 3490 3893 3516
rect 2915 3488 3832 3490
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 3881 3485 3893 3490
rect 3927 3516 3939 3519
rect 3970 3516 3976 3528
rect 3927 3488 3976 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 4264 3525 4292 3556
rect 4890 3544 4896 3556
rect 4948 3584 4954 3596
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 4948 3556 5089 3584
rect 4948 3544 4954 3556
rect 5077 3553 5089 3556
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 6178 3544 6184 3596
rect 6236 3544 6242 3596
rect 6270 3544 6276 3596
rect 6328 3544 6334 3596
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6512 3556 6653 3584
rect 6512 3544 6518 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 7374 3584 7380 3596
rect 7239 3556 7380 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7484 3584 7512 3624
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 8996 3624 9628 3652
rect 8996 3612 9002 3624
rect 9600 3596 9628 3624
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 10505 3655 10563 3661
rect 10505 3652 10517 3655
rect 9732 3624 10517 3652
rect 9732 3612 9738 3624
rect 10505 3621 10517 3624
rect 10551 3621 10563 3655
rect 10505 3615 10563 3621
rect 7929 3587 7987 3593
rect 7484 3573 7788 3584
rect 7929 3573 7941 3587
rect 7484 3556 7941 3573
rect 7760 3553 7941 3556
rect 7975 3584 7987 3587
rect 8754 3584 8760 3596
rect 7975 3553 7997 3584
rect 7760 3545 7997 3553
rect 8036 3556 8760 3584
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4525 3519 4583 3525
rect 4525 3485 4537 3519
rect 4571 3516 4583 3519
rect 4709 3519 4767 3525
rect 4571 3488 4660 3516
rect 4571 3485 4583 3488
rect 4525 3479 4583 3485
rect 4264 3448 4292 3479
rect 2792 3420 4292 3448
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 2130 3380 2136 3392
rect 1452 3352 2136 3380
rect 1452 3340 1458 3352
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 3602 3380 3608 3392
rect 3384 3352 3608 3380
rect 3384 3340 3390 3352
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 3973 3383 4031 3389
rect 3973 3380 3985 3383
rect 3752 3352 3985 3380
rect 3752 3340 3758 3352
rect 3973 3349 3985 3352
rect 4019 3349 4031 3383
rect 3973 3343 4031 3349
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 4632 3380 4660 3488
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4724 3448 4752 3479
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5316 3488 5365 3516
rect 5316 3476 5322 3488
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 6914 3476 6920 3528
rect 6972 3476 6978 3528
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3516 7067 3519
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7055 3488 7297 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 7285 3485 7297 3488
rect 7331 3516 7343 3519
rect 8036 3516 8064 3556
rect 8754 3544 8760 3556
rect 8812 3584 8818 3596
rect 9214 3584 9220 3596
rect 8812 3556 9220 3584
rect 8812 3544 8818 3556
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 10226 3584 10232 3596
rect 9640 3556 10232 3584
rect 9640 3544 9646 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10612 3584 10640 3692
rect 11440 3652 11468 3692
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 12710 3720 12716 3732
rect 11747 3692 12716 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 16482 3720 16488 3732
rect 12820 3692 16488 3720
rect 12158 3652 12164 3664
rect 11440 3624 12164 3652
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 12250 3612 12256 3664
rect 12308 3652 12314 3664
rect 12345 3655 12403 3661
rect 12345 3652 12357 3655
rect 12308 3624 12357 3652
rect 12308 3612 12314 3624
rect 12345 3621 12357 3624
rect 12391 3621 12403 3655
rect 12345 3615 12403 3621
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 12820 3652 12848 3692
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 16666 3680 16672 3732
rect 16724 3720 16730 3732
rect 17586 3720 17592 3732
rect 16724 3692 17172 3720
rect 16724 3680 16730 3692
rect 12492 3624 12848 3652
rect 12492 3612 12498 3624
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 13081 3655 13139 3661
rect 13081 3652 13093 3655
rect 12952 3624 13093 3652
rect 12952 3612 12958 3624
rect 13081 3621 13093 3624
rect 13127 3652 13139 3655
rect 14826 3652 14832 3664
rect 13127 3624 14832 3652
rect 13127 3621 13139 3624
rect 13081 3615 13139 3621
rect 14826 3612 14832 3624
rect 14884 3612 14890 3664
rect 15930 3612 15936 3664
rect 15988 3612 15994 3664
rect 10781 3587 10839 3593
rect 10781 3584 10793 3587
rect 10612 3556 10793 3584
rect 10781 3553 10793 3556
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 11054 3544 11060 3596
rect 11112 3544 11118 3596
rect 13262 3584 13268 3596
rect 12084 3556 13268 3584
rect 7331 3488 8064 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 7024 3448 7052 3479
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8846 3516 8852 3528
rect 8496 3488 8852 3516
rect 4724 3420 7052 3448
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 8021 3451 8079 3457
rect 8021 3448 8033 3451
rect 7239 3420 8033 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 8021 3417 8033 3420
rect 8067 3417 8079 3451
rect 8496 3448 8524 3488
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9674 3516 9680 3528
rect 9355 3488 9680 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9674 3476 9680 3488
rect 9732 3516 9738 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9732 3488 9873 3516
rect 9732 3476 9738 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10042 3476 10048 3528
rect 10100 3476 10106 3528
rect 10870 3476 10876 3528
rect 10928 3525 10934 3528
rect 10928 3519 10956 3525
rect 10944 3485 10956 3519
rect 10928 3479 10956 3485
rect 10928 3476 10934 3479
rect 11790 3476 11796 3528
rect 11848 3476 11854 3528
rect 11974 3476 11980 3528
rect 12032 3476 12038 3528
rect 12084 3525 12112 3556
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 13596 3556 13645 3584
rect 13596 3544 13602 3556
rect 13633 3553 13645 3556
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 13814 3544 13820 3596
rect 13872 3584 13878 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 13872 3556 14749 3584
rect 13872 3544 13878 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15010 3544 15016 3596
rect 15068 3544 15074 3596
rect 15194 3593 15200 3596
rect 15151 3587 15200 3593
rect 15151 3553 15163 3587
rect 15197 3553 15200 3587
rect 15151 3547 15200 3553
rect 15194 3544 15200 3547
rect 15252 3544 15258 3596
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16114 3584 16120 3596
rect 15528 3556 16120 3584
rect 15528 3544 15534 3556
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 16850 3593 16856 3596
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 16540 3556 16681 3584
rect 16540 3544 16546 3556
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 16828 3587 16856 3593
rect 16828 3553 16840 3587
rect 16828 3547 16856 3553
rect 16850 3544 16856 3547
rect 16908 3544 16914 3596
rect 17144 3584 17172 3692
rect 17236 3692 17592 3720
rect 17236 3661 17264 3692
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 18969 3723 19027 3729
rect 18969 3689 18981 3723
rect 19015 3720 19027 3723
rect 19794 3720 19800 3732
rect 19015 3692 19800 3720
rect 19015 3689 19027 3692
rect 18969 3683 19027 3689
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 21821 3723 21879 3729
rect 21821 3720 21833 3723
rect 19904 3692 21833 3720
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3621 17279 3655
rect 17221 3615 17279 3621
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 17460 3624 17724 3652
rect 17460 3612 17466 3624
rect 17696 3593 17724 3624
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 19904 3661 19932 3692
rect 21821 3689 21833 3692
rect 21867 3689 21879 3723
rect 24489 3723 24547 3729
rect 24489 3720 24501 3723
rect 21821 3683 21879 3689
rect 21928 3692 24501 3720
rect 19889 3655 19947 3661
rect 18840 3624 19380 3652
rect 18840 3612 18846 3624
rect 16960 3556 17172 3584
rect 17681 3587 17739 3593
rect 12069 3519 12127 3525
rect 12069 3485 12081 3519
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 12618 3516 12624 3528
rect 12207 3488 12624 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 13228 3488 13369 3516
rect 13228 3476 13234 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13357 3479 13415 3485
rect 13743 3488 14105 3516
rect 8021 3411 8079 3417
rect 8128 3420 8524 3448
rect 4706 3380 4712 3392
rect 4632 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3380 5043 3383
rect 5534 3380 5540 3392
rect 5031 3352 5540 3380
rect 5031 3349 5043 3352
rect 4985 3343 5043 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6454 3340 6460 3392
rect 6512 3340 6518 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7374 3380 7380 3392
rect 6880 3352 7380 3380
rect 6880 3340 6886 3352
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 8128 3380 8156 3420
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9088 3420 9904 3448
rect 9088 3408 9094 3420
rect 7699 3352 8156 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 8202 3340 8208 3392
rect 8260 3340 8266 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 8628 3352 9321 3380
rect 8628 3340 8634 3352
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9309 3343 9367 3349
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9582 3380 9588 3392
rect 9447 3352 9588 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9766 3340 9772 3392
rect 9824 3340 9830 3392
rect 9876 3380 9904 3420
rect 12526 3408 12532 3460
rect 12584 3408 12590 3460
rect 13262 3408 13268 3460
rect 13320 3448 13326 3460
rect 13743 3448 13771 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 13320 3420 13771 3448
rect 13817 3451 13875 3457
rect 13320 3408 13326 3420
rect 13817 3417 13829 3451
rect 13863 3448 13875 3451
rect 13998 3448 14004 3460
rect 13863 3420 14004 3448
rect 13863 3417 13875 3420
rect 13817 3411 13875 3417
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 12434 3380 12440 3392
rect 9876 3352 12440 3380
rect 12434 3340 12440 3352
rect 12492 3340 12498 3392
rect 12618 3340 12624 3392
rect 12676 3340 12682 3392
rect 13538 3340 13544 3392
rect 13596 3340 13602 3392
rect 14108 3380 14136 3479
rect 14182 3476 14188 3528
rect 14240 3516 14246 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14240 3488 14289 3516
rect 14240 3476 14246 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 15286 3476 15292 3528
rect 15344 3476 15350 3528
rect 16960 3525 16988 3556
rect 17681 3553 17693 3587
rect 17727 3553 17739 3587
rect 17681 3547 17739 3553
rect 19352 3528 19380 3624
rect 19889 3621 19901 3655
rect 19935 3621 19947 3655
rect 21928 3652 21956 3692
rect 24489 3689 24501 3692
rect 24535 3689 24547 3723
rect 24489 3683 24547 3689
rect 24762 3680 24768 3732
rect 24820 3720 24826 3732
rect 24820 3692 27568 3720
rect 24820 3680 24826 3692
rect 19889 3615 19947 3621
rect 21284 3624 21956 3652
rect 19426 3544 19432 3596
rect 19484 3544 19490 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 20282 3587 20340 3593
rect 20282 3584 20294 3587
rect 19576 3556 20294 3584
rect 19576 3544 19582 3556
rect 20282 3553 20294 3556
rect 20328 3553 20340 3587
rect 20282 3547 20340 3553
rect 20441 3587 20499 3593
rect 20441 3553 20453 3587
rect 20487 3584 20499 3587
rect 21284 3584 21312 3624
rect 25682 3612 25688 3664
rect 25740 3652 25746 3664
rect 27540 3652 27568 3692
rect 27614 3680 27620 3732
rect 27672 3680 27678 3732
rect 27816 3692 29592 3720
rect 27816 3652 27844 3692
rect 25740 3624 26556 3652
rect 27540 3624 27844 3652
rect 25740 3612 25746 3624
rect 20487 3556 21312 3584
rect 20487 3553 20499 3556
rect 20441 3547 20499 3553
rect 25498 3544 25504 3596
rect 25556 3544 25562 3596
rect 26418 3544 26424 3596
rect 26476 3544 26482 3596
rect 26528 3584 26556 3624
rect 26697 3587 26755 3593
rect 26697 3584 26709 3587
rect 26528 3556 26709 3584
rect 26697 3553 26709 3556
rect 26743 3553 26755 3587
rect 26697 3547 26755 3553
rect 26786 3544 26792 3596
rect 26844 3593 26850 3596
rect 26844 3587 26872 3593
rect 26860 3553 26872 3587
rect 26844 3547 26872 3553
rect 26844 3544 26850 3547
rect 27706 3544 27712 3596
rect 27764 3544 27770 3596
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17865 3519 17923 3525
rect 17865 3485 17877 3519
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18138 3516 18144 3528
rect 18003 3488 18144 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 15948 3420 16252 3448
rect 15948 3380 15976 3420
rect 14108 3352 15976 3380
rect 16022 3340 16028 3392
rect 16080 3340 16086 3392
rect 16224 3380 16252 3420
rect 17880 3380 17908 3479
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 18046 3408 18052 3460
rect 18104 3448 18110 3460
rect 18248 3448 18276 3479
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 18748 3488 19257 3516
rect 18748 3476 18754 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19334 3476 19340 3528
rect 19392 3476 19398 3528
rect 20162 3476 20168 3528
rect 20220 3476 20226 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 21008 3488 21465 3516
rect 21008 3460 21036 3488
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 21726 3476 21732 3528
rect 21784 3516 21790 3528
rect 22557 3519 22615 3525
rect 22557 3516 22569 3519
rect 21784 3488 22569 3516
rect 21784 3476 21790 3488
rect 22557 3485 22569 3488
rect 22603 3516 22615 3519
rect 22646 3516 22652 3528
rect 22603 3488 22652 3516
rect 22603 3485 22615 3488
rect 22557 3479 22615 3485
rect 22646 3476 22652 3488
rect 22704 3476 22710 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 24121 3519 24179 3525
rect 24121 3485 24133 3519
rect 24167 3485 24179 3519
rect 24121 3479 24179 3485
rect 18104 3420 18276 3448
rect 18104 3408 18110 3420
rect 19058 3408 19064 3460
rect 19116 3448 19122 3460
rect 19426 3448 19432 3460
rect 19116 3420 19432 3448
rect 19116 3408 19122 3420
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 20990 3408 20996 3460
rect 21048 3408 21054 3460
rect 21085 3451 21143 3457
rect 21085 3417 21097 3451
rect 21131 3448 21143 3451
rect 21131 3420 21772 3448
rect 21131 3417 21143 3420
rect 21085 3411 21143 3417
rect 20438 3380 20444 3392
rect 16224 3352 20444 3380
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 21637 3383 21695 3389
rect 21637 3380 21649 3383
rect 20956 3352 21649 3380
rect 20956 3340 20962 3352
rect 21637 3349 21649 3352
rect 21683 3349 21695 3383
rect 21744 3380 21772 3420
rect 22094 3408 22100 3460
rect 22152 3448 22158 3460
rect 22848 3448 22876 3479
rect 22152 3420 22876 3448
rect 22152 3408 22158 3420
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 23860 3448 23888 3479
rect 23072 3420 23888 3448
rect 24136 3448 24164 3479
rect 25222 3476 25228 3528
rect 25280 3476 25286 3528
rect 25777 3519 25835 3525
rect 25777 3485 25789 3519
rect 25823 3516 25835 3519
rect 25866 3516 25872 3528
rect 25823 3488 25872 3516
rect 25823 3485 25835 3488
rect 25777 3479 25835 3485
rect 25866 3476 25872 3488
rect 25924 3476 25930 3528
rect 25958 3476 25964 3528
rect 26016 3476 26022 3528
rect 26970 3476 26976 3528
rect 27028 3476 27034 3528
rect 27982 3476 27988 3528
rect 28040 3476 28046 3528
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 28813 3519 28871 3525
rect 28813 3516 28825 3519
rect 28408 3488 28825 3516
rect 28408 3476 28414 3488
rect 28813 3485 28825 3488
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 29564 3525 29592 3692
rect 29914 3680 29920 3732
rect 29972 3720 29978 3732
rect 32030 3720 32036 3732
rect 29972 3692 32036 3720
rect 29972 3680 29978 3692
rect 32030 3680 32036 3692
rect 32088 3680 32094 3732
rect 32122 3680 32128 3732
rect 32180 3720 32186 3732
rect 32861 3723 32919 3729
rect 32180 3692 32812 3720
rect 32180 3680 32186 3692
rect 30929 3655 30987 3661
rect 30929 3621 30941 3655
rect 30975 3652 30987 3655
rect 30975 3624 31800 3652
rect 30975 3621 30987 3624
rect 30929 3615 30987 3621
rect 29638 3544 29644 3596
rect 29696 3584 29702 3596
rect 29917 3587 29975 3593
rect 29917 3584 29929 3587
rect 29696 3556 29929 3584
rect 29696 3544 29702 3556
rect 29917 3553 29929 3556
rect 29963 3553 29975 3587
rect 29917 3547 29975 3553
rect 31018 3544 31024 3596
rect 31076 3544 31082 3596
rect 31662 3544 31668 3596
rect 31720 3544 31726 3596
rect 31772 3584 31800 3624
rect 32217 3587 32275 3593
rect 32217 3584 32229 3587
rect 31772 3556 32229 3584
rect 32217 3553 32229 3556
rect 32263 3553 32275 3587
rect 32217 3547 32275 3553
rect 29181 3519 29239 3525
rect 29181 3516 29193 3519
rect 28960 3488 29193 3516
rect 28960 3476 28966 3488
rect 29181 3485 29193 3488
rect 29227 3485 29239 3519
rect 29181 3479 29239 3485
rect 29549 3519 29607 3525
rect 29549 3485 29561 3519
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 30098 3476 30104 3528
rect 30156 3516 30162 3528
rect 30193 3519 30251 3525
rect 30193 3516 30205 3519
rect 30156 3488 30205 3516
rect 30156 3476 30162 3488
rect 30193 3485 30205 3488
rect 30239 3485 30251 3519
rect 30193 3479 30251 3485
rect 31202 3476 31208 3528
rect 31260 3476 31266 3528
rect 31938 3476 31944 3528
rect 31996 3476 32002 3528
rect 32030 3476 32036 3528
rect 32088 3525 32094 3528
rect 32088 3519 32116 3525
rect 32104 3485 32116 3519
rect 32088 3479 32116 3485
rect 32088 3476 32094 3479
rect 24854 3448 24860 3460
rect 24136 3420 24860 3448
rect 23072 3408 23078 3420
rect 22646 3380 22652 3392
rect 21744 3352 22652 3380
rect 21637 3343 21695 3349
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 23109 3383 23167 3389
rect 23109 3349 23121 3383
rect 23155 3380 23167 3383
rect 23474 3380 23480 3392
rect 23155 3352 23480 3380
rect 23155 3349 23167 3352
rect 23109 3343 23167 3349
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 23860 3380 23888 3420
rect 24854 3408 24860 3420
rect 24912 3408 24918 3460
rect 32784 3448 32812 3692
rect 32861 3689 32873 3723
rect 32907 3720 32919 3723
rect 34238 3720 34244 3732
rect 32907 3692 34244 3720
rect 32907 3689 32919 3692
rect 32861 3683 32919 3689
rect 34238 3680 34244 3692
rect 34296 3680 34302 3732
rect 34330 3680 34336 3732
rect 34388 3720 34394 3732
rect 36449 3723 36507 3729
rect 36449 3720 36461 3723
rect 34388 3692 36461 3720
rect 34388 3680 34394 3692
rect 36449 3689 36461 3692
rect 36495 3689 36507 3723
rect 36449 3683 36507 3689
rect 38286 3680 38292 3732
rect 38344 3720 38350 3732
rect 38473 3723 38531 3729
rect 38473 3720 38485 3723
rect 38344 3692 38485 3720
rect 38344 3680 38350 3692
rect 38473 3689 38485 3692
rect 38519 3689 38531 3723
rect 38473 3683 38531 3689
rect 39390 3680 39396 3732
rect 39448 3680 39454 3732
rect 33137 3655 33195 3661
rect 33137 3621 33149 3655
rect 33183 3652 33195 3655
rect 33502 3652 33508 3664
rect 33183 3624 33508 3652
rect 33183 3621 33195 3624
rect 33137 3615 33195 3621
rect 33502 3612 33508 3624
rect 33560 3612 33566 3664
rect 34606 3612 34612 3664
rect 34664 3652 34670 3664
rect 38010 3652 38016 3664
rect 34664 3624 38016 3652
rect 34664 3612 34670 3624
rect 38010 3612 38016 3624
rect 38068 3612 38074 3664
rect 39025 3655 39083 3661
rect 39025 3621 39037 3655
rect 39071 3652 39083 3655
rect 39942 3652 39948 3664
rect 39071 3624 39948 3652
rect 39071 3621 39083 3624
rect 39025 3615 39083 3621
rect 39942 3612 39948 3624
rect 40000 3612 40006 3664
rect 34333 3587 34391 3593
rect 34333 3553 34345 3587
rect 34379 3584 34391 3587
rect 34422 3584 34428 3596
rect 34379 3556 34428 3584
rect 34379 3553 34391 3556
rect 34333 3547 34391 3553
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35066 3584 35072 3596
rect 34532 3556 35072 3584
rect 32858 3476 32864 3528
rect 32916 3516 32922 3528
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32916 3488 32965 3516
rect 32916 3476 32922 3488
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 34057 3519 34115 3525
rect 34057 3485 34069 3519
rect 34103 3516 34115 3519
rect 34532 3516 34560 3556
rect 35066 3544 35072 3556
rect 35124 3544 35130 3596
rect 34103 3488 34560 3516
rect 34103 3485 34115 3488
rect 34057 3479 34115 3485
rect 34698 3476 34704 3528
rect 34756 3476 34762 3528
rect 35158 3476 35164 3528
rect 35216 3476 35222 3528
rect 35618 3476 35624 3528
rect 35676 3516 35682 3528
rect 38286 3516 38292 3528
rect 35676 3488 38292 3516
rect 35676 3476 35682 3488
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 38657 3519 38715 3525
rect 38657 3485 38669 3519
rect 38703 3516 38715 3519
rect 38746 3516 38752 3528
rect 38703 3488 38752 3516
rect 38703 3485 38715 3488
rect 38657 3479 38715 3485
rect 38746 3476 38752 3488
rect 38804 3476 38810 3528
rect 38838 3476 38844 3528
rect 38896 3476 38902 3528
rect 38930 3476 38936 3528
rect 38988 3516 38994 3528
rect 39209 3519 39267 3525
rect 39209 3516 39221 3519
rect 38988 3488 39221 3516
rect 38988 3476 38994 3488
rect 39209 3485 39221 3488
rect 39255 3485 39267 3519
rect 39209 3479 39267 3485
rect 27448 3420 29868 3448
rect 32784 3420 33916 3448
rect 27448 3380 27476 3420
rect 23860 3352 27476 3380
rect 27614 3340 27620 3392
rect 27672 3380 27678 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 27672 3352 28733 3380
rect 27672 3340 27678 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 28994 3340 29000 3392
rect 29052 3340 29058 3392
rect 29362 3340 29368 3392
rect 29420 3340 29426 3392
rect 29638 3340 29644 3392
rect 29696 3380 29702 3392
rect 29733 3383 29791 3389
rect 29733 3380 29745 3383
rect 29696 3352 29745 3380
rect 29696 3340 29702 3352
rect 29733 3349 29745 3352
rect 29779 3349 29791 3383
rect 29840 3380 29868 3420
rect 31386 3380 31392 3392
rect 29840 3352 31392 3380
rect 29733 3343 29791 3349
rect 31386 3340 31392 3352
rect 31444 3340 31450 3392
rect 33318 3340 33324 3392
rect 33376 3340 33382 3392
rect 33888 3380 33916 3420
rect 35250 3408 35256 3460
rect 35308 3448 35314 3460
rect 39114 3448 39120 3460
rect 35308 3420 39120 3448
rect 35308 3408 35314 3420
rect 39114 3408 39120 3420
rect 39172 3408 39178 3460
rect 34514 3380 34520 3392
rect 33888 3352 34520 3380
rect 34514 3340 34520 3352
rect 34572 3340 34578 3392
rect 34885 3383 34943 3389
rect 34885 3349 34897 3383
rect 34931 3380 34943 3383
rect 34974 3380 34980 3392
rect 34931 3352 34980 3380
rect 34931 3349 34943 3352
rect 34885 3343 34943 3349
rect 34974 3340 34980 3352
rect 35032 3340 35038 3392
rect 35710 3340 35716 3392
rect 35768 3380 35774 3392
rect 37642 3380 37648 3392
rect 35768 3352 37648 3380
rect 35768 3340 35774 3352
rect 37642 3340 37648 3352
rect 37700 3340 37706 3392
rect 1104 3290 39836 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 9010 3290
rect 9062 3238 9074 3290
rect 9126 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 15010 3290
rect 15062 3238 15074 3290
rect 15126 3238 15138 3290
rect 15190 3238 15202 3290
rect 15254 3238 15266 3290
rect 15318 3238 21010 3290
rect 21062 3238 21074 3290
rect 21126 3238 21138 3290
rect 21190 3238 21202 3290
rect 21254 3238 21266 3290
rect 21318 3238 27010 3290
rect 27062 3238 27074 3290
rect 27126 3238 27138 3290
rect 27190 3238 27202 3290
rect 27254 3238 27266 3290
rect 27318 3238 33010 3290
rect 33062 3238 33074 3290
rect 33126 3238 33138 3290
rect 33190 3238 33202 3290
rect 33254 3238 33266 3290
rect 33318 3238 39010 3290
rect 39062 3238 39074 3290
rect 39126 3238 39138 3290
rect 39190 3238 39202 3290
rect 39254 3238 39266 3290
rect 39318 3238 39836 3290
rect 1104 3216 39836 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 1854 3176 1860 3188
rect 1636 3148 1860 3176
rect 1636 3136 1642 3148
rect 1854 3136 1860 3148
rect 1912 3176 1918 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1912 3148 1961 3176
rect 1912 3136 1918 3148
rect 1949 3145 1961 3148
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 3878 3176 3884 3188
rect 3283 3148 3884 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4982 3176 4988 3188
rect 4387 3148 4988 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 7282 3176 7288 3188
rect 5092 3148 7288 3176
rect 1486 3068 1492 3120
rect 1544 3068 1550 3120
rect 4430 3068 4436 3120
rect 4488 3108 4494 3120
rect 5092 3108 5120 3148
rect 7282 3136 7288 3148
rect 7340 3176 7346 3188
rect 7466 3176 7472 3188
rect 7340 3148 7472 3176
rect 7340 3136 7346 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7760 3148 9812 3176
rect 6178 3108 6184 3120
rect 4488 3080 5120 3108
rect 5184 3080 6184 3108
rect 4488 3068 4494 3080
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1452 3012 1869 3040
rect 1452 3000 1458 3012
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2188 3012 2513 3040
rect 2188 3000 2194 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 3602 3040 3608 3052
rect 2501 3003 2559 3009
rect 3252 3012 3608 3040
rect 3252 2984 3280 3012
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4246 3000 4252 3052
rect 4304 3040 4310 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4304 3012 4537 3040
rect 4304 3000 4310 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 5184 3049 5212 3080
rect 6178 3068 6184 3080
rect 6236 3068 6242 3120
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4948 3012 4997 3040
rect 4948 3000 4954 3012
rect 4985 3009 4997 3012
rect 5031 3040 5043 3043
rect 5169 3043 5227 3049
rect 5169 3040 5181 3043
rect 5031 3012 5181 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5169 3009 5181 3012
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5776 3012 6377 3040
rect 5776 3000 5782 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 1670 2864 1676 2916
rect 1728 2864 1734 2916
rect 2240 2836 2268 2935
rect 3234 2932 3240 2984
rect 3292 2932 3298 2984
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3344 2836 3372 2935
rect 5810 2932 5816 2984
rect 5868 2972 5874 2984
rect 7760 2981 7788 3148
rect 9784 3108 9812 3148
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10870 3176 10876 3188
rect 10376 3148 10876 3176
rect 10376 3136 10382 3148
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 11606 3176 11612 3188
rect 11379 3148 11612 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 13814 3136 13820 3188
rect 13872 3136 13878 3188
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 16485 3179 16543 3185
rect 14139 3148 16436 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 9784 3080 9996 3108
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8294 3040 8300 3052
rect 8076 3012 8300 3040
rect 8076 3000 8082 3012
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8904 3012 8953 3040
rect 8904 3000 8910 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 9088 3012 9505 3040
rect 9088 3000 9094 3012
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9968 3040 9996 3080
rect 10042 3068 10048 3120
rect 10100 3108 10106 3120
rect 13262 3108 13268 3120
rect 10100 3080 13268 3108
rect 10100 3068 10106 3080
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 16022 3108 16028 3120
rect 13924 3080 16028 3108
rect 10318 3040 10324 3052
rect 9640 3012 9812 3040
rect 9968 3012 10324 3040
rect 9640 3000 9646 3012
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 5868 2944 7757 2972
rect 5868 2932 5874 2944
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 9180 2944 9229 2972
rect 9180 2932 9186 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9784 2972 9812 3012
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10594 3000 10600 3052
rect 10652 3000 10658 3052
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 12986 3040 12992 3052
rect 12575 3012 12992 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 12986 3000 12992 3012
rect 13044 3000 13050 3052
rect 13924 3049 13952 3080
rect 16022 3068 16028 3080
rect 16080 3068 16086 3120
rect 16408 3108 16436 3148
rect 16485 3145 16497 3179
rect 16531 3176 16543 3179
rect 17586 3176 17592 3188
rect 16531 3148 17592 3176
rect 16531 3145 16543 3148
rect 16485 3139 16543 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 20622 3176 20628 3188
rect 17696 3148 20628 3176
rect 17696 3108 17724 3148
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 28442 3176 28448 3188
rect 20772 3148 22048 3176
rect 20772 3136 20778 3148
rect 16408 3080 17724 3108
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19484 3080 19656 3108
rect 19484 3068 19490 3080
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13909 3043 13967 3049
rect 13127 3012 13584 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 9784 2944 10272 2972
rect 9217 2935 9275 2941
rect 4706 2864 4712 2916
rect 4764 2864 4770 2916
rect 4893 2839 4951 2845
rect 4893 2836 4905 2839
rect 2240 2808 4905 2836
rect 4893 2805 4905 2808
rect 4939 2836 4951 2839
rect 5828 2836 5856 2932
rect 6086 2864 6092 2916
rect 6144 2904 6150 2916
rect 6181 2907 6239 2913
rect 6181 2904 6193 2907
rect 6144 2876 6193 2904
rect 6144 2864 6150 2876
rect 6181 2873 6193 2876
rect 6227 2904 6239 2907
rect 6546 2904 6552 2916
rect 6227 2876 6552 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 10244 2913 10272 2944
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 11572 2944 11621 2972
rect 11572 2932 11578 2944
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11609 2935 11667 2941
rect 11882 2932 11888 2984
rect 11940 2932 11946 2984
rect 12805 2975 12863 2981
rect 12805 2941 12817 2975
rect 12851 2941 12863 2975
rect 12805 2935 12863 2941
rect 10229 2907 10287 2913
rect 8680 2876 9352 2904
rect 4939 2808 5856 2836
rect 7561 2839 7619 2845
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 8680 2836 8708 2876
rect 7607 2808 8708 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 8754 2796 8760 2848
rect 8812 2796 8818 2848
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 9214 2836 9220 2848
rect 9079 2808 9220 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 9324 2836 9352 2876
rect 10229 2873 10241 2907
rect 10275 2873 10287 2907
rect 10229 2867 10287 2873
rect 12710 2864 12716 2916
rect 12768 2864 12774 2916
rect 9582 2836 9588 2848
rect 9324 2808 9588 2836
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 12434 2836 12440 2848
rect 9732 2808 12440 2836
rect 9732 2796 9738 2808
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 12820 2836 12848 2935
rect 13556 2904 13584 3012
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14366 3040 14372 3052
rect 14056 3012 14372 3040
rect 14056 3000 14062 3012
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14461 3043 14519 3049
rect 14461 3009 14473 3043
rect 14507 3040 14519 3043
rect 14734 3040 14740 3052
rect 14507 3012 14740 3040
rect 14507 3009 14519 3012
rect 14461 3003 14519 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15102 3000 15108 3052
rect 15160 3000 15166 3052
rect 15654 3040 15660 3052
rect 15212 3012 15660 3040
rect 13722 2904 13728 2916
rect 13556 2876 13728 2904
rect 13722 2864 13728 2876
rect 13780 2904 13786 2916
rect 15212 2904 15240 3012
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3040 15807 3043
rect 16114 3040 16120 3052
rect 15795 3012 16120 3040
rect 15795 3009 15807 3012
rect 15749 3003 15807 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16758 3000 16764 3052
rect 16816 3000 16822 3052
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3040 17187 3043
rect 17218 3040 17224 3052
rect 17175 3012 17224 3040
rect 17175 3009 17187 3012
rect 17129 3003 17187 3009
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17494 3000 17500 3052
rect 17552 3000 17558 3052
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3040 19395 3043
rect 19518 3040 19524 3052
rect 19383 3012 19524 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19628 3049 19656 3080
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 20346 3000 20352 3052
rect 20404 3000 20410 3052
rect 21361 3043 21419 3049
rect 21361 3009 21373 3043
rect 21407 3040 21419 3043
rect 21910 3040 21916 3052
rect 21407 3012 21916 3040
rect 21407 3009 21419 3012
rect 21361 3003 21419 3009
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 15381 2975 15439 2981
rect 15381 2941 15393 2975
rect 15427 2941 15439 2975
rect 15381 2935 15439 2941
rect 13780 2876 15240 2904
rect 13780 2864 13786 2876
rect 13262 2836 13268 2848
rect 12820 2808 13268 2836
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 14277 2839 14335 2845
rect 14277 2805 14289 2839
rect 14323 2836 14335 2839
rect 14918 2836 14924 2848
rect 14323 2808 14924 2836
rect 14323 2805 14335 2808
rect 14277 2799 14335 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15396 2836 15424 2935
rect 15470 2932 15476 2984
rect 15528 2932 15534 2984
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 18322 2981 18328 2984
rect 18141 2975 18199 2981
rect 18141 2972 18153 2975
rect 17644 2944 18153 2972
rect 17644 2932 17650 2944
rect 18141 2941 18153 2944
rect 18187 2941 18199 2975
rect 18141 2935 18199 2941
rect 18300 2975 18328 2981
rect 18300 2941 18312 2975
rect 18300 2935 18328 2941
rect 18322 2932 18328 2935
rect 18380 2932 18386 2984
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 18598 2972 18604 2984
rect 18463 2944 18604 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 18598 2932 18604 2944
rect 18656 2972 18662 2984
rect 18656 2944 18828 2972
rect 18656 2932 18662 2944
rect 17034 2904 17040 2916
rect 16868 2876 17040 2904
rect 16868 2836 16896 2876
rect 17034 2864 17040 2876
rect 17092 2864 17098 2916
rect 18693 2907 18751 2913
rect 18693 2873 18705 2907
rect 18739 2873 18751 2907
rect 18693 2867 18751 2873
rect 15396 2808 16896 2836
rect 16942 2796 16948 2848
rect 17000 2796 17006 2848
rect 17310 2796 17316 2848
rect 17368 2796 17374 2848
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 17770 2836 17776 2848
rect 17460 2808 17776 2836
rect 17460 2796 17466 2808
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 18708 2836 18736 2867
rect 18012 2808 18736 2836
rect 18800 2836 18828 2944
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19153 2975 19211 2981
rect 19153 2972 19165 2975
rect 19116 2944 19165 2972
rect 19116 2932 19122 2944
rect 19153 2941 19165 2944
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2941 19487 2975
rect 19429 2935 19487 2941
rect 18874 2864 18880 2916
rect 18932 2904 18938 2916
rect 19444 2904 19472 2935
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 20466 2975 20524 2981
rect 20466 2972 20478 2975
rect 19852 2944 20478 2972
rect 19852 2932 19858 2944
rect 20466 2941 20478 2944
rect 20512 2941 20524 2975
rect 20466 2935 20524 2941
rect 20622 2932 20628 2984
rect 20680 2932 20686 2984
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 21821 2975 21879 2981
rect 21821 2972 21833 2975
rect 20864 2944 21833 2972
rect 20864 2932 20870 2944
rect 21821 2941 21833 2944
rect 21867 2941 21879 2975
rect 22020 2972 22048 3148
rect 23032 3148 28448 3176
rect 23032 3052 23060 3148
rect 24673 3111 24731 3117
rect 24673 3077 24685 3111
rect 24719 3108 24731 3111
rect 24719 3080 26656 3108
rect 24719 3077 24731 3080
rect 24673 3071 24731 3077
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 22143 3012 22968 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 22833 2975 22891 2981
rect 22833 2972 22845 2975
rect 22020 2944 22845 2972
rect 21821 2935 21879 2941
rect 22833 2941 22845 2944
rect 22879 2941 22891 2975
rect 22940 2972 22968 3012
rect 23014 3000 23020 3052
rect 23072 3000 23078 3052
rect 23750 3000 23756 3052
rect 23808 3000 23814 3052
rect 24026 3000 24032 3052
rect 24084 3000 24090 3052
rect 25222 3000 25228 3052
rect 25280 3040 25286 3052
rect 25501 3043 25559 3049
rect 25501 3040 25513 3043
rect 25280 3012 25513 3040
rect 25280 3000 25286 3012
rect 25501 3009 25513 3012
rect 25547 3009 25559 3043
rect 25501 3003 25559 3009
rect 25590 3000 25596 3052
rect 25648 3040 25654 3052
rect 25869 3043 25927 3049
rect 25869 3040 25881 3043
rect 25648 3012 25881 3040
rect 25648 3000 25654 3012
rect 25869 3009 25881 3012
rect 25915 3009 25927 3043
rect 25869 3003 25927 3009
rect 26142 3000 26148 3052
rect 26200 3040 26206 3052
rect 26418 3040 26424 3052
rect 26200 3012 26424 3040
rect 26200 3000 26206 3012
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 26628 3050 26656 3080
rect 26620 3049 26656 3050
rect 26513 3043 26571 3049
rect 26513 3009 26525 3043
rect 26559 3009 26571 3043
rect 26513 3003 26571 3009
rect 26605 3043 26663 3049
rect 26605 3009 26617 3043
rect 26651 3009 26663 3043
rect 26605 3003 26663 3009
rect 22940 2944 23428 2972
rect 22833 2935 22891 2941
rect 18932 2876 19472 2904
rect 20073 2907 20131 2913
rect 18932 2864 18938 2876
rect 20073 2873 20085 2907
rect 20119 2873 20131 2907
rect 20073 2867 20131 2873
rect 19978 2836 19984 2848
rect 18800 2808 19984 2836
rect 18012 2796 18018 2808
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 20088 2836 20116 2867
rect 21082 2864 21088 2916
rect 21140 2904 21146 2916
rect 21545 2907 21603 2913
rect 21545 2904 21557 2907
rect 21140 2876 21557 2904
rect 21140 2864 21146 2876
rect 21545 2873 21557 2876
rect 21591 2873 21603 2907
rect 23400 2904 23428 2944
rect 23474 2932 23480 2984
rect 23532 2932 23538 2984
rect 23891 2975 23949 2981
rect 23891 2972 23903 2975
rect 23584 2944 23903 2972
rect 23584 2904 23612 2944
rect 23891 2941 23903 2944
rect 23937 2972 23949 2975
rect 24210 2972 24216 2984
rect 23937 2944 24216 2972
rect 23937 2941 23949 2944
rect 23891 2935 23949 2941
rect 24210 2932 24216 2944
rect 24268 2932 24274 2984
rect 25774 2932 25780 2984
rect 25832 2932 25838 2984
rect 26528 2972 26556 3003
rect 26970 3000 26976 3052
rect 27028 3000 27034 3052
rect 27080 3040 27108 3148
rect 28442 3136 28448 3148
rect 28500 3176 28506 3188
rect 28813 3179 28871 3185
rect 28500 3148 28764 3176
rect 28500 3136 28506 3148
rect 28736 3108 28764 3148
rect 28813 3145 28825 3179
rect 28859 3176 28871 3179
rect 28902 3176 28908 3188
rect 28859 3148 28908 3176
rect 28859 3145 28871 3148
rect 28813 3139 28871 3145
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 29362 3136 29368 3188
rect 29420 3176 29426 3188
rect 29420 3148 31754 3176
rect 29420 3136 29426 3148
rect 31726 3108 31754 3148
rect 31846 3136 31852 3188
rect 31904 3136 31910 3188
rect 31938 3136 31944 3188
rect 31996 3176 32002 3188
rect 33318 3176 33324 3188
rect 31996 3148 33324 3176
rect 31996 3136 32002 3148
rect 33318 3136 33324 3148
rect 33376 3136 33382 3188
rect 33686 3136 33692 3188
rect 33744 3136 33750 3188
rect 33778 3136 33784 3188
rect 33836 3136 33842 3188
rect 34514 3136 34520 3188
rect 34572 3176 34578 3188
rect 35434 3176 35440 3188
rect 34572 3148 35440 3176
rect 34572 3136 34578 3148
rect 35434 3136 35440 3148
rect 35492 3176 35498 3188
rect 35802 3176 35808 3188
rect 35492 3148 35808 3176
rect 35492 3136 35498 3148
rect 35802 3136 35808 3148
rect 35860 3136 35866 3188
rect 35986 3136 35992 3188
rect 36044 3176 36050 3188
rect 36081 3179 36139 3185
rect 36081 3176 36093 3179
rect 36044 3148 36093 3176
rect 36044 3136 36050 3148
rect 36081 3145 36093 3148
rect 36127 3145 36139 3179
rect 36081 3139 36139 3145
rect 36541 3179 36599 3185
rect 36541 3145 36553 3179
rect 36587 3176 36599 3179
rect 37090 3176 37096 3188
rect 36587 3148 37096 3176
rect 36587 3145 36599 3148
rect 36541 3139 36599 3145
rect 37090 3136 37096 3148
rect 37148 3136 37154 3188
rect 37642 3136 37648 3188
rect 37700 3176 37706 3188
rect 37737 3179 37795 3185
rect 37737 3176 37749 3179
rect 37700 3148 37749 3176
rect 37700 3136 37706 3148
rect 37737 3145 37749 3148
rect 37783 3145 37795 3179
rect 37737 3139 37795 3145
rect 38010 3136 38016 3188
rect 38068 3136 38074 3188
rect 39390 3136 39396 3188
rect 39448 3136 39454 3188
rect 38657 3111 38715 3117
rect 38657 3108 38669 3111
rect 28736 3080 28856 3108
rect 31726 3080 34652 3108
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 27080 3012 27169 3040
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 28166 3000 28172 3052
rect 28224 3000 28230 3052
rect 28828 3044 28856 3080
rect 28828 3040 28994 3044
rect 29089 3043 29147 3049
rect 29089 3040 29101 3043
rect 28828 3016 29101 3040
rect 28966 3012 29101 3016
rect 29089 3009 29101 3012
rect 29135 3009 29147 3043
rect 29089 3003 29147 3009
rect 29914 3000 29920 3052
rect 29972 3049 29978 3052
rect 29972 3043 30000 3049
rect 29988 3009 30000 3043
rect 29972 3003 30000 3009
rect 29972 3000 29978 3003
rect 30742 3000 30748 3052
rect 30800 3040 30806 3052
rect 31113 3043 31171 3049
rect 31113 3040 31125 3043
rect 30800 3012 31125 3040
rect 30800 3000 30806 3012
rect 31113 3009 31125 3012
rect 31159 3009 31171 3043
rect 31113 3003 31171 3009
rect 31386 3000 31392 3052
rect 31444 3040 31450 3052
rect 32401 3043 32459 3049
rect 32401 3040 32413 3043
rect 31444 3012 32413 3040
rect 31444 3000 31450 3012
rect 32401 3009 32413 3012
rect 32447 3040 32459 3043
rect 33229 3043 33287 3049
rect 33229 3040 33241 3043
rect 32447 3012 33241 3040
rect 32447 3009 32459 3012
rect 32401 3003 32459 3009
rect 33229 3009 33241 3012
rect 33275 3009 33287 3043
rect 33229 3003 33287 3009
rect 34146 3000 34152 3052
rect 34204 3040 34210 3052
rect 34624 3049 34652 3080
rect 35636 3080 38669 3108
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 34204 3012 34253 3040
rect 34204 3000 34210 3012
rect 34241 3009 34253 3012
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 34609 3043 34667 3049
rect 34609 3009 34621 3043
rect 34655 3009 34667 3043
rect 34609 3003 34667 3009
rect 34790 3000 34796 3052
rect 34848 3040 34854 3052
rect 34977 3043 35035 3049
rect 34977 3040 34989 3043
rect 34848 3012 34989 3040
rect 34848 3000 34854 3012
rect 34977 3009 34989 3012
rect 35023 3009 35035 3043
rect 34977 3003 35035 3009
rect 35342 3000 35348 3052
rect 35400 3000 35406 3052
rect 27522 2972 27528 2984
rect 26528 2944 27528 2972
rect 27522 2932 27528 2944
rect 27580 2932 27586 2984
rect 27614 2932 27620 2984
rect 27672 2932 27678 2984
rect 27893 2975 27951 2981
rect 27893 2972 27905 2975
rect 27724 2944 27905 2972
rect 23400 2876 23612 2904
rect 21545 2867 21603 2873
rect 24486 2864 24492 2916
rect 24544 2904 24550 2916
rect 24765 2907 24823 2913
rect 24765 2904 24777 2907
rect 24544 2876 24777 2904
rect 24544 2864 24550 2876
rect 24765 2873 24777 2876
rect 24811 2873 24823 2907
rect 26602 2904 26608 2916
rect 24765 2867 24823 2873
rect 25700 2876 26608 2904
rect 20346 2836 20352 2848
rect 20088 2808 20352 2836
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 21174 2836 21180 2848
rect 20496 2808 21180 2836
rect 20496 2796 20502 2808
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 21269 2839 21327 2845
rect 21269 2805 21281 2839
rect 21315 2836 21327 2839
rect 21450 2836 21456 2848
rect 21315 2808 21456 2836
rect 21315 2805 21327 2808
rect 21269 2799 21327 2805
rect 21450 2796 21456 2808
rect 21508 2796 21514 2848
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 24854 2836 24860 2848
rect 22796 2808 24860 2836
rect 22796 2796 22802 2808
rect 24854 2796 24860 2808
rect 24912 2796 24918 2848
rect 25498 2796 25504 2848
rect 25556 2836 25562 2848
rect 25700 2836 25728 2876
rect 26602 2864 26608 2876
rect 26660 2864 26666 2916
rect 27724 2904 27752 2944
rect 27893 2941 27905 2944
rect 27939 2941 27951 2975
rect 27893 2935 27951 2941
rect 28031 2975 28089 2981
rect 28031 2941 28043 2975
rect 28077 2972 28089 2975
rect 28350 2972 28356 2984
rect 28077 2944 28356 2972
rect 28077 2941 28089 2944
rect 28031 2935 28089 2941
rect 28350 2932 28356 2944
rect 28408 2932 28414 2984
rect 28810 2932 28816 2984
rect 28868 2972 28874 2984
rect 28905 2975 28963 2981
rect 28905 2972 28917 2975
rect 28868 2944 28917 2972
rect 28868 2932 28874 2944
rect 28905 2941 28917 2944
rect 28951 2941 28963 2975
rect 29822 2972 29828 2984
rect 28905 2935 28963 2941
rect 29288 2944 29828 2972
rect 29288 2904 29316 2944
rect 29822 2932 29828 2944
rect 29880 2932 29886 2984
rect 30101 2975 30159 2981
rect 30101 2941 30113 2975
rect 30147 2972 30159 2975
rect 30466 2972 30472 2984
rect 30147 2944 30472 2972
rect 30147 2941 30159 2944
rect 30101 2935 30159 2941
rect 30466 2932 30472 2944
rect 30524 2932 30530 2984
rect 30834 2932 30840 2984
rect 30892 2932 30898 2984
rect 31478 2932 31484 2984
rect 31536 2972 31542 2984
rect 31536 2944 31754 2972
rect 31536 2932 31542 2944
rect 27586 2876 27752 2904
rect 28828 2876 29316 2904
rect 25556 2808 25728 2836
rect 25556 2796 25562 2808
rect 25774 2796 25780 2848
rect 25832 2836 25838 2848
rect 26053 2839 26111 2845
rect 26053 2836 26065 2839
rect 25832 2808 26065 2836
rect 25832 2796 25838 2808
rect 26053 2805 26065 2808
rect 26099 2805 26111 2839
rect 26053 2799 26111 2805
rect 26329 2839 26387 2845
rect 26329 2805 26341 2839
rect 26375 2836 26387 2839
rect 26418 2836 26424 2848
rect 26375 2808 26424 2836
rect 26375 2805 26387 2808
rect 26329 2799 26387 2805
rect 26418 2796 26424 2808
rect 26476 2796 26482 2848
rect 26786 2796 26792 2848
rect 26844 2796 26850 2848
rect 27062 2796 27068 2848
rect 27120 2836 27126 2848
rect 27586 2836 27614 2876
rect 28828 2836 28856 2876
rect 29362 2864 29368 2916
rect 29420 2904 29426 2916
rect 29549 2907 29607 2913
rect 29549 2904 29561 2907
rect 29420 2876 29561 2904
rect 29420 2864 29426 2876
rect 29549 2873 29561 2876
rect 29595 2873 29607 2907
rect 31726 2904 31754 2944
rect 31846 2932 31852 2984
rect 31904 2972 31910 2984
rect 32122 2972 32128 2984
rect 31904 2944 32128 2972
rect 31904 2932 31910 2944
rect 32122 2932 32128 2944
rect 32180 2932 32186 2984
rect 33505 2975 33563 2981
rect 33505 2941 33517 2975
rect 33551 2941 33563 2975
rect 33505 2935 33563 2941
rect 33137 2907 33195 2913
rect 31726 2876 32168 2904
rect 29549 2867 29607 2873
rect 27120 2808 28856 2836
rect 27120 2796 27126 2808
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 29914 2836 29920 2848
rect 28960 2808 29920 2836
rect 28960 2796 28966 2808
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 30745 2839 30803 2845
rect 30745 2805 30757 2839
rect 30791 2836 30803 2839
rect 31938 2836 31944 2848
rect 30791 2808 31944 2836
rect 30791 2805 30803 2808
rect 30745 2799 30803 2805
rect 31938 2796 31944 2808
rect 31996 2796 32002 2848
rect 32140 2836 32168 2876
rect 33137 2873 33149 2907
rect 33183 2904 33195 2907
rect 33520 2904 33548 2935
rect 33594 2932 33600 2984
rect 33652 2972 33658 2984
rect 35636 2972 35664 3080
rect 38657 3077 38669 3080
rect 38703 3077 38715 3111
rect 38657 3071 38715 3077
rect 35710 3000 35716 3052
rect 35768 3000 35774 3052
rect 35802 3000 35808 3052
rect 35860 3040 35866 3052
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 35860 3012 36277 3040
rect 35860 3000 35866 3012
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 36265 3003 36323 3009
rect 36357 3043 36415 3049
rect 36357 3009 36369 3043
rect 36403 3009 36415 3043
rect 36357 3003 36415 3009
rect 33652 2944 35664 2972
rect 33652 2932 33658 2944
rect 36078 2932 36084 2984
rect 36136 2972 36142 2984
rect 36372 2972 36400 3003
rect 37274 3000 37280 3052
rect 37332 3040 37338 3052
rect 37921 3043 37979 3049
rect 37921 3040 37933 3043
rect 37332 3012 37933 3040
rect 37332 3000 37338 3012
rect 37921 3009 37933 3012
rect 37967 3009 37979 3043
rect 37921 3003 37979 3009
rect 38197 3043 38255 3049
rect 38197 3009 38209 3043
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 36136 2944 36400 2972
rect 36136 2932 36142 2944
rect 37642 2932 37648 2984
rect 37700 2972 37706 2984
rect 38212 2972 38240 3003
rect 38286 3000 38292 3052
rect 38344 3000 38350 3052
rect 38749 3043 38807 3049
rect 38749 3009 38761 3043
rect 38795 3040 38807 3043
rect 38841 3043 38899 3049
rect 38841 3040 38853 3043
rect 38795 3012 38853 3040
rect 38795 3009 38807 3012
rect 38749 3003 38807 3009
rect 38841 3009 38853 3012
rect 38887 3009 38899 3043
rect 38841 3003 38899 3009
rect 39209 3043 39267 3049
rect 39209 3009 39221 3043
rect 39255 3009 39267 3043
rect 39209 3003 39267 3009
rect 39224 2972 39252 3003
rect 37700 2944 38240 2972
rect 38304 2944 39252 2972
rect 37700 2932 37706 2944
rect 34425 2907 34483 2913
rect 34425 2904 34437 2907
rect 33183 2876 33548 2904
rect 33612 2876 34437 2904
rect 33183 2873 33195 2876
rect 33137 2867 33195 2873
rect 33612 2836 33640 2876
rect 34425 2873 34437 2876
rect 34471 2873 34483 2907
rect 36354 2904 36360 2916
rect 34425 2867 34483 2873
rect 34532 2876 36360 2904
rect 32140 2808 33640 2836
rect 34149 2839 34207 2845
rect 34149 2805 34161 2839
rect 34195 2836 34207 2839
rect 34532 2836 34560 2876
rect 36354 2864 36360 2876
rect 36412 2864 36418 2916
rect 36722 2864 36728 2916
rect 36780 2904 36786 2916
rect 38304 2904 38332 2944
rect 36780 2876 38332 2904
rect 38473 2907 38531 2913
rect 36780 2864 36786 2876
rect 38473 2873 38485 2907
rect 38519 2904 38531 2907
rect 39666 2904 39672 2916
rect 38519 2876 39672 2904
rect 38519 2873 38531 2876
rect 38473 2867 38531 2873
rect 39666 2864 39672 2876
rect 39724 2864 39730 2916
rect 34195 2808 34560 2836
rect 34195 2805 34207 2808
rect 34149 2799 34207 2805
rect 34606 2796 34612 2848
rect 34664 2836 34670 2848
rect 34793 2839 34851 2845
rect 34793 2836 34805 2839
rect 34664 2808 34805 2836
rect 34664 2796 34670 2808
rect 34793 2805 34805 2808
rect 34839 2805 34851 2839
rect 34793 2799 34851 2805
rect 35158 2796 35164 2848
rect 35216 2796 35222 2848
rect 35342 2796 35348 2848
rect 35400 2836 35406 2848
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 35400 2808 35541 2836
rect 35400 2796 35406 2808
rect 35529 2805 35541 2808
rect 35575 2805 35587 2839
rect 35529 2799 35587 2805
rect 35897 2839 35955 2845
rect 35897 2805 35909 2839
rect 35943 2836 35955 2839
rect 35986 2836 35992 2848
rect 35943 2808 35992 2836
rect 35943 2805 35955 2808
rect 35897 2799 35955 2805
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 39022 2796 39028 2848
rect 39080 2796 39086 2848
rect 1104 2746 39836 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 13950 2746
rect 14002 2694 14014 2746
rect 14066 2694 14078 2746
rect 14130 2694 14142 2746
rect 14194 2694 14206 2746
rect 14258 2694 19950 2746
rect 20002 2694 20014 2746
rect 20066 2694 20078 2746
rect 20130 2694 20142 2746
rect 20194 2694 20206 2746
rect 20258 2694 25950 2746
rect 26002 2694 26014 2746
rect 26066 2694 26078 2746
rect 26130 2694 26142 2746
rect 26194 2694 26206 2746
rect 26258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 37950 2746
rect 38002 2694 38014 2746
rect 38066 2694 38078 2746
rect 38130 2694 38142 2746
rect 38194 2694 38206 2746
rect 38258 2694 39836 2746
rect 1104 2672 39836 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2774 2632 2780 2644
rect 1627 2604 2780 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 4338 2632 4344 2644
rect 3559 2604 4344 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4663 2604 6408 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 3292 2536 4108 2564
rect 3292 2524 3298 2536
rect 2774 2456 2780 2508
rect 2832 2456 2838 2508
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3970 2496 3976 2508
rect 3191 2468 3976 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3970 2456 3976 2468
rect 4028 2456 4034 2508
rect 1486 2388 1492 2440
rect 1544 2388 1550 2440
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2866 2428 2872 2440
rect 2271 2400 2872 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3050 2428 3056 2440
rect 3007 2400 3056 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3510 2428 3516 2440
rect 3344 2400 3516 2428
rect 1854 2320 1860 2372
rect 1912 2320 1918 2372
rect 2406 2320 2412 2372
rect 2464 2320 2470 2372
rect 2593 2363 2651 2369
rect 2593 2329 2605 2363
rect 2639 2360 2651 2363
rect 3344 2360 3372 2400
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 2639 2332 2774 2360
rect 2639 2329 2651 2332
rect 2593 2323 2651 2329
rect 1946 2252 1952 2304
rect 2004 2252 2010 2304
rect 2746 2292 2774 2332
rect 2976 2332 3372 2360
rect 3421 2363 3479 2369
rect 2976 2292 3004 2332
rect 3421 2329 3433 2363
rect 3467 2360 3479 2363
rect 3878 2360 3884 2372
rect 3467 2332 3884 2360
rect 3467 2329 3479 2332
rect 3421 2323 3479 2329
rect 3878 2320 3884 2332
rect 3936 2320 3942 2372
rect 3973 2363 4031 2369
rect 3973 2329 3985 2363
rect 4019 2360 4031 2363
rect 4080 2360 4108 2536
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 5258 2496 5264 2508
rect 4856 2468 5264 2496
rect 4856 2456 4862 2468
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 6178 2456 6184 2508
rect 6236 2456 6242 2508
rect 6380 2496 6408 2604
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 6604 2604 7481 2632
rect 6604 2592 6610 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 7469 2595 7527 2601
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 11793 2635 11851 2641
rect 11793 2632 11805 2635
rect 7892 2604 11805 2632
rect 7892 2592 7898 2604
rect 11793 2601 11805 2604
rect 11839 2601 11851 2635
rect 13262 2632 13268 2644
rect 11793 2595 11851 2601
rect 12406 2604 13268 2632
rect 6454 2524 6460 2576
rect 6512 2564 6518 2576
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 6512 2536 7297 2564
rect 6512 2524 6518 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 7374 2524 7380 2576
rect 7432 2564 7438 2576
rect 7432 2536 8248 2564
rect 7432 2524 7438 2536
rect 7006 2496 7012 2508
rect 6380 2468 7012 2496
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 7558 2456 7564 2508
rect 7616 2456 7622 2508
rect 8220 2505 8248 2536
rect 8386 2524 8392 2576
rect 8444 2564 8450 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 8444 2536 11989 2564
rect 8444 2524 8450 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 12406 2564 12434 2604
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13630 2592 13636 2644
rect 13688 2632 13694 2644
rect 13725 2635 13783 2641
rect 13725 2632 13737 2635
rect 13688 2604 13737 2632
rect 13688 2592 13694 2604
rect 13725 2601 13737 2604
rect 13771 2632 13783 2635
rect 13906 2632 13912 2644
rect 13771 2604 13912 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 15286 2632 15292 2644
rect 14384 2604 15292 2632
rect 11977 2527 12035 2533
rect 12360 2536 12434 2564
rect 13357 2567 13415 2573
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2465 8263 2499
rect 8205 2459 8263 2465
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 12360 2505 12388 2536
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 14384 2564 14412 2604
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 16114 2632 16120 2644
rect 15804 2604 16120 2632
rect 15804 2592 15810 2604
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 17218 2592 17224 2644
rect 17276 2592 17282 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 18782 2632 18788 2644
rect 17819 2604 18788 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 20257 2635 20315 2641
rect 19306 2604 19932 2632
rect 13403 2536 14412 2564
rect 16485 2567 16543 2573
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 16485 2533 16497 2567
rect 16531 2533 16543 2567
rect 16485 2527 16543 2533
rect 16945 2567 17003 2573
rect 16945 2533 16957 2567
rect 16991 2564 17003 2567
rect 17402 2564 17408 2576
rect 16991 2536 17408 2564
rect 16991 2533 17003 2536
rect 16945 2527 17003 2533
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 8812 2468 11897 2496
rect 8812 2456 8818 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 12345 2499 12403 2505
rect 12345 2465 12357 2499
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 13262 2456 13268 2508
rect 13320 2496 13326 2508
rect 13320 2468 14412 2496
rect 13320 2456 13326 2468
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4571 2400 5856 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 4019 2332 4108 2360
rect 4019 2329 4031 2332
rect 3973 2323 4031 2329
rect 2746 2264 3004 2292
rect 3988 2292 4016 2323
rect 4154 2320 4160 2372
rect 4212 2320 4218 2372
rect 4890 2320 4896 2372
rect 4948 2320 4954 2372
rect 5828 2360 5856 2400
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6328 2400 6377 2428
rect 6328 2388 6334 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 6687 2400 7849 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 6546 2360 6552 2372
rect 5828 2332 6552 2360
rect 6546 2320 6552 2332
rect 6604 2320 6610 2372
rect 7852 2360 7880 2391
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 9214 2428 9220 2440
rect 8536 2400 9220 2428
rect 8536 2388 8542 2400
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9398 2388 9404 2440
rect 9456 2388 9462 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 8662 2360 8668 2372
rect 7852 2332 8668 2360
rect 8662 2320 8668 2332
rect 8720 2320 8726 2372
rect 8754 2320 8760 2372
rect 8812 2360 8818 2372
rect 9030 2360 9036 2372
rect 8812 2332 9036 2360
rect 8812 2320 8818 2332
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 9125 2363 9183 2369
rect 9125 2329 9137 2363
rect 9171 2360 9183 2363
rect 9490 2360 9496 2372
rect 9171 2332 9496 2360
rect 9171 2329 9183 2332
rect 9125 2323 9183 2329
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 9692 2360 9720 2391
rect 11054 2388 11060 2440
rect 11112 2388 11118 2440
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11204 2400 11345 2428
rect 11204 2388 11210 2400
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 11333 2391 11391 2397
rect 11422 2388 11428 2440
rect 11480 2428 11486 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11480 2400 11529 2428
rect 11480 2388 11486 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12158 2428 12164 2440
rect 12115 2400 12164 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 13906 2428 13912 2440
rect 13587 2400 13912 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 14090 2388 14096 2440
rect 14148 2388 14154 2440
rect 14274 2388 14280 2440
rect 14332 2388 14338 2440
rect 14384 2437 14412 2468
rect 15470 2456 15476 2508
rect 15528 2456 15534 2508
rect 16500 2496 16528 2527
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 18874 2564 18880 2576
rect 18380 2536 18880 2564
rect 18380 2524 18386 2536
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 19306 2564 19334 2604
rect 19260 2536 19334 2564
rect 17954 2496 17960 2508
rect 16500 2468 17960 2496
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 19260 2505 19288 2536
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 18104 2468 19257 2496
rect 18104 2456 18110 2468
rect 19245 2465 19257 2468
rect 19291 2465 19303 2499
rect 19904 2496 19932 2604
rect 20257 2601 20269 2635
rect 20303 2632 20315 2635
rect 20346 2632 20352 2644
rect 20303 2604 20352 2632
rect 20303 2601 20315 2604
rect 20257 2595 20315 2601
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 20680 2604 21373 2632
rect 20680 2592 20686 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 32214 2632 32220 2644
rect 22336 2604 32220 2632
rect 22336 2592 22342 2604
rect 32214 2592 32220 2604
rect 32272 2632 32278 2644
rect 33410 2632 33416 2644
rect 32272 2604 33416 2632
rect 32272 2592 32278 2604
rect 33410 2592 33416 2604
rect 33468 2592 33474 2644
rect 33778 2592 33784 2644
rect 33836 2632 33842 2644
rect 33836 2604 37780 2632
rect 33836 2592 33842 2604
rect 22830 2524 22836 2576
rect 22888 2524 22894 2576
rect 23937 2567 23995 2573
rect 23937 2533 23949 2567
rect 23983 2564 23995 2567
rect 24026 2564 24032 2576
rect 23983 2536 24032 2564
rect 23983 2533 23995 2536
rect 23937 2527 23995 2533
rect 24026 2524 24032 2536
rect 24084 2524 24090 2576
rect 26237 2567 26295 2573
rect 26237 2533 26249 2567
rect 26283 2533 26295 2567
rect 26237 2527 26295 2533
rect 20349 2499 20407 2505
rect 20349 2496 20361 2499
rect 19904 2468 20361 2496
rect 19245 2459 19303 2465
rect 20349 2465 20361 2468
rect 20395 2465 20407 2499
rect 20349 2459 20407 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 22796 2468 22937 2496
rect 22796 2456 22802 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 26252 2496 26280 2527
rect 26510 2524 26516 2576
rect 26568 2564 26574 2576
rect 26973 2567 27031 2573
rect 26973 2564 26985 2567
rect 26568 2536 26985 2564
rect 26568 2524 26574 2536
rect 26973 2533 26985 2536
rect 27019 2533 27031 2567
rect 26973 2527 27031 2533
rect 29362 2524 29368 2576
rect 29420 2524 29426 2576
rect 30466 2524 30472 2576
rect 30524 2564 30530 2576
rect 30561 2567 30619 2573
rect 30561 2564 30573 2567
rect 30524 2536 30573 2564
rect 30524 2524 30530 2536
rect 30561 2533 30573 2536
rect 30607 2533 30619 2567
rect 30561 2527 30619 2533
rect 31754 2524 31760 2576
rect 31812 2564 31818 2576
rect 31849 2567 31907 2573
rect 31849 2564 31861 2567
rect 31812 2536 31861 2564
rect 31812 2524 31818 2536
rect 31849 2533 31861 2536
rect 31895 2533 31907 2567
rect 32309 2567 32367 2573
rect 32309 2564 32321 2567
rect 31849 2527 31907 2533
rect 31956 2536 32321 2564
rect 26878 2496 26884 2508
rect 26252 2468 26884 2496
rect 22925 2459 22983 2465
rect 26878 2456 26884 2468
rect 26936 2456 26942 2508
rect 30834 2456 30840 2508
rect 30892 2456 30898 2508
rect 31478 2456 31484 2508
rect 31536 2496 31542 2508
rect 31956 2496 31984 2536
rect 32309 2533 32321 2536
rect 32355 2533 32367 2567
rect 32309 2527 32367 2533
rect 32950 2524 32956 2576
rect 33008 2564 33014 2576
rect 33686 2564 33692 2576
rect 33008 2536 33692 2564
rect 33008 2524 33014 2536
rect 33686 2524 33692 2536
rect 33744 2524 33750 2576
rect 33962 2524 33968 2576
rect 34020 2564 34026 2576
rect 34517 2567 34575 2573
rect 34020 2536 34468 2564
rect 34020 2524 34026 2536
rect 31536 2468 31984 2496
rect 32048 2468 33272 2496
rect 31536 2456 31542 2468
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14292 2360 14320 2388
rect 9692 2332 14320 2360
rect 14384 2360 14412 2391
rect 14642 2388 14648 2440
rect 14700 2428 14706 2440
rect 15010 2428 15016 2440
rect 14700 2400 15016 2428
rect 14700 2388 14706 2400
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15488 2360 15516 2456
rect 15746 2388 15752 2440
rect 15804 2388 15810 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 15948 2400 17049 2428
rect 15948 2372 15976 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 19058 2388 19064 2440
rect 19116 2388 19122 2440
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 20622 2388 20628 2440
rect 20680 2388 20686 2440
rect 21450 2388 21456 2440
rect 21508 2388 21514 2440
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 14384 2332 15516 2360
rect 15930 2320 15936 2372
rect 15988 2320 15994 2372
rect 16574 2320 16580 2372
rect 16632 2360 16638 2372
rect 16761 2363 16819 2369
rect 16761 2360 16773 2363
rect 16632 2332 16773 2360
rect 16632 2320 16638 2332
rect 16761 2329 16773 2332
rect 16807 2329 16819 2363
rect 16761 2323 16819 2329
rect 16850 2320 16856 2372
rect 16908 2360 16914 2372
rect 16908 2332 17724 2360
rect 16908 2320 16914 2332
rect 4246 2292 4252 2304
rect 3988 2264 4252 2292
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 4982 2252 4988 2304
rect 5040 2252 5046 2304
rect 5169 2295 5227 2301
rect 5169 2261 5181 2295
rect 5215 2292 5227 2295
rect 5626 2292 5632 2304
rect 5215 2264 5632 2292
rect 5215 2261 5227 2264
rect 5169 2255 5227 2261
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 8202 2292 8208 2304
rect 6788 2264 8208 2292
rect 6788 2252 6794 2264
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 9217 2295 9275 2301
rect 9217 2261 9229 2295
rect 9263 2292 9275 2295
rect 11238 2292 11244 2304
rect 9263 2264 11244 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11606 2252 11612 2304
rect 11664 2252 11670 2304
rect 12250 2252 12256 2304
rect 12308 2252 12314 2304
rect 14274 2252 14280 2304
rect 14332 2252 14338 2304
rect 15381 2295 15439 2301
rect 15381 2261 15393 2295
rect 15427 2292 15439 2295
rect 17586 2292 17592 2304
rect 15427 2264 17592 2292
rect 15427 2261 15439 2264
rect 15381 2255 15439 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 17696 2292 17724 2332
rect 17770 2320 17776 2372
rect 17828 2360 17834 2372
rect 21836 2360 21864 2391
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 22152 2400 23213 2428
rect 22152 2388 22158 2400
rect 23201 2397 23213 2400
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 24029 2431 24087 2437
rect 24029 2397 24041 2431
rect 24075 2397 24087 2431
rect 24394 2428 24400 2440
rect 24029 2391 24087 2397
rect 24136 2400 24400 2428
rect 21910 2360 21916 2372
rect 17828 2332 21916 2360
rect 17828 2320 17834 2332
rect 21910 2320 21916 2332
rect 21968 2320 21974 2372
rect 22646 2320 22652 2372
rect 22704 2360 22710 2372
rect 24044 2360 24072 2391
rect 22704 2332 24072 2360
rect 22704 2320 22710 2332
rect 20806 2292 20812 2304
rect 17696 2264 20812 2292
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 21637 2295 21695 2301
rect 21637 2261 21649 2295
rect 21683 2292 21695 2295
rect 24136 2292 24164 2400
rect 24394 2388 24400 2400
rect 24452 2388 24458 2440
rect 24670 2388 24676 2440
rect 24728 2388 24734 2440
rect 24762 2388 24768 2440
rect 24820 2388 24826 2440
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 25188 2400 25237 2428
rect 25188 2388 25194 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 25498 2388 25504 2440
rect 25556 2388 25562 2440
rect 26329 2431 26387 2437
rect 26329 2397 26341 2431
rect 26375 2397 26387 2431
rect 26329 2391 26387 2397
rect 26344 2360 26372 2391
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 27709 2431 27767 2437
rect 27709 2428 27721 2431
rect 27672 2400 27721 2428
rect 27672 2388 27678 2400
rect 27709 2397 27721 2400
rect 27755 2397 27767 2431
rect 27709 2391 27767 2397
rect 27985 2431 28043 2437
rect 27985 2397 27997 2431
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 28077 2431 28135 2437
rect 28077 2397 28089 2431
rect 28123 2397 28135 2431
rect 28077 2391 28135 2397
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28399 2424 28488 2428
rect 28534 2424 28540 2440
rect 28399 2400 28540 2424
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28460 2396 28540 2400
rect 28000 2360 28028 2391
rect 24228 2332 26372 2360
rect 26436 2332 28028 2360
rect 28092 2360 28120 2391
rect 28534 2388 28540 2396
rect 28592 2388 28598 2440
rect 28629 2431 28687 2437
rect 28629 2397 28641 2431
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 28644 2390 28675 2391
rect 28644 2360 28672 2390
rect 28718 2388 28724 2440
rect 28776 2428 28782 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 28776 2400 29561 2428
rect 28776 2388 28782 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 29822 2388 29828 2440
rect 29880 2428 29886 2440
rect 31113 2431 31171 2437
rect 31113 2428 31125 2431
rect 29880 2400 31125 2428
rect 29880 2388 29886 2400
rect 31113 2397 31125 2400
rect 31159 2428 31171 2431
rect 31938 2428 31944 2440
rect 31159 2400 31944 2428
rect 31159 2397 31171 2400
rect 31113 2391 31171 2397
rect 31938 2388 31944 2400
rect 31996 2388 32002 2440
rect 28810 2360 28816 2372
rect 28092 2332 28816 2360
rect 24228 2301 24256 2332
rect 21683 2264 24164 2292
rect 24213 2295 24271 2301
rect 21683 2261 21695 2264
rect 21637 2255 21695 2261
rect 24213 2261 24225 2295
rect 24259 2261 24271 2295
rect 24213 2255 24271 2261
rect 24302 2252 24308 2304
rect 24360 2292 24366 2304
rect 24489 2295 24547 2301
rect 24489 2292 24501 2295
rect 24360 2264 24501 2292
rect 24360 2252 24366 2264
rect 24489 2261 24501 2264
rect 24535 2261 24547 2295
rect 24489 2255 24547 2261
rect 24854 2252 24860 2304
rect 24912 2292 24918 2304
rect 24949 2295 25007 2301
rect 24949 2292 24961 2295
rect 24912 2264 24961 2292
rect 24912 2252 24918 2264
rect 24949 2261 24961 2264
rect 24995 2261 25007 2295
rect 24949 2255 25007 2261
rect 25682 2252 25688 2304
rect 25740 2292 25746 2304
rect 26436 2292 26464 2332
rect 25740 2264 26464 2292
rect 25740 2252 25746 2264
rect 26510 2252 26516 2304
rect 26568 2252 26574 2304
rect 26602 2252 26608 2304
rect 26660 2292 26666 2304
rect 28092 2292 28120 2332
rect 28810 2320 28816 2332
rect 28868 2320 28874 2372
rect 28902 2320 28908 2372
rect 28960 2360 28966 2372
rect 29086 2360 29092 2372
rect 28960 2332 29092 2360
rect 28960 2320 28966 2332
rect 29086 2320 29092 2332
rect 29144 2320 29150 2372
rect 29362 2320 29368 2372
rect 29420 2360 29426 2372
rect 32048 2360 32076 2468
rect 32125 2431 32183 2437
rect 32125 2397 32137 2431
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 29420 2332 32076 2360
rect 29420 2320 29426 2332
rect 26660 2264 28120 2292
rect 26660 2252 26666 2264
rect 28258 2252 28264 2304
rect 28316 2252 28322 2304
rect 28442 2252 28448 2304
rect 28500 2292 28506 2304
rect 32140 2292 32168 2391
rect 32398 2388 32404 2440
rect 32456 2428 32462 2440
rect 33244 2437 33272 2468
rect 33318 2456 33324 2508
rect 33376 2496 33382 2508
rect 33376 2468 34376 2496
rect 33376 2456 33382 2468
rect 34348 2437 34376 2468
rect 32493 2431 32551 2437
rect 32493 2428 32505 2431
rect 32456 2400 32505 2428
rect 32456 2388 32462 2400
rect 32493 2397 32505 2400
rect 32539 2397 32551 2431
rect 32493 2391 32551 2397
rect 33137 2431 33195 2437
rect 33137 2397 33149 2431
rect 33183 2397 33195 2431
rect 33137 2391 33195 2397
rect 33229 2431 33287 2437
rect 33229 2397 33241 2431
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 33873 2431 33931 2437
rect 33873 2397 33885 2431
rect 33919 2428 33931 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33919 2400 33977 2428
rect 33919 2397 33931 2400
rect 33873 2391 33931 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 34333 2431 34391 2437
rect 34333 2397 34345 2431
rect 34379 2397 34391 2431
rect 34333 2391 34391 2397
rect 33152 2360 33180 2391
rect 34054 2360 34060 2372
rect 33152 2332 34060 2360
rect 34054 2320 34060 2332
rect 34112 2320 34118 2372
rect 34440 2360 34468 2536
rect 34517 2533 34529 2567
rect 34563 2533 34575 2567
rect 34517 2527 34575 2533
rect 35989 2567 36047 2573
rect 35989 2533 36001 2567
rect 36035 2564 36047 2567
rect 36446 2564 36452 2576
rect 36035 2536 36452 2564
rect 36035 2533 36047 2536
rect 35989 2527 36047 2533
rect 34532 2496 34560 2527
rect 36446 2524 36452 2536
rect 36504 2524 36510 2576
rect 34532 2468 35848 2496
rect 34698 2388 34704 2440
rect 34756 2388 34762 2440
rect 35066 2388 35072 2440
rect 35124 2388 35130 2440
rect 35434 2388 35440 2440
rect 35492 2388 35498 2440
rect 35820 2437 35848 2468
rect 35805 2431 35863 2437
rect 35805 2397 35817 2431
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 36354 2388 36360 2440
rect 36412 2388 36418 2440
rect 37752 2437 37780 2604
rect 39390 2592 39396 2644
rect 39448 2592 39454 2644
rect 38289 2567 38347 2573
rect 38289 2533 38301 2567
rect 38335 2564 38347 2567
rect 39574 2564 39580 2576
rect 38335 2536 39580 2564
rect 38335 2533 38347 2536
rect 38289 2527 38347 2533
rect 39574 2524 39580 2536
rect 39632 2524 39638 2576
rect 37844 2468 38516 2496
rect 37737 2431 37795 2437
rect 37737 2397 37749 2431
rect 37783 2397 37795 2431
rect 37737 2391 37795 2397
rect 37844 2360 37872 2468
rect 38102 2388 38108 2440
rect 38160 2388 38166 2440
rect 38488 2437 38516 2468
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2397 38531 2431
rect 38473 2391 38531 2397
rect 38838 2388 38844 2440
rect 38896 2388 38902 2440
rect 39206 2388 39212 2440
rect 39264 2388 39270 2440
rect 40034 2360 40040 2372
rect 34440 2332 37872 2360
rect 37936 2332 40040 2360
rect 28500 2264 32168 2292
rect 28500 2252 28506 2264
rect 32674 2252 32680 2304
rect 32732 2252 32738 2304
rect 32766 2252 32772 2304
rect 32824 2292 32830 2304
rect 32953 2295 33011 2301
rect 32953 2292 32965 2295
rect 32824 2264 32965 2292
rect 32824 2252 32830 2264
rect 32953 2261 32965 2264
rect 32999 2261 33011 2295
rect 32953 2255 33011 2261
rect 33410 2252 33416 2304
rect 33468 2252 33474 2304
rect 33778 2252 33784 2304
rect 33836 2252 33842 2304
rect 34146 2252 34152 2304
rect 34204 2252 34210 2304
rect 34882 2252 34888 2304
rect 34940 2252 34946 2304
rect 35158 2252 35164 2304
rect 35216 2292 35222 2304
rect 35253 2295 35311 2301
rect 35253 2292 35265 2295
rect 35216 2264 35265 2292
rect 35216 2252 35222 2264
rect 35253 2261 35265 2264
rect 35299 2261 35311 2295
rect 35253 2255 35311 2261
rect 35618 2252 35624 2304
rect 35676 2252 35682 2304
rect 36170 2252 36176 2304
rect 36228 2252 36234 2304
rect 37936 2301 37964 2332
rect 40034 2320 40040 2332
rect 40092 2320 40098 2372
rect 37921 2295 37979 2301
rect 37921 2261 37933 2295
rect 37967 2261 37979 2295
rect 37921 2255 37979 2261
rect 38654 2252 38660 2304
rect 38712 2252 38718 2304
rect 39025 2295 39083 2301
rect 39025 2261 39037 2295
rect 39071 2292 39083 2295
rect 39942 2292 39948 2304
rect 39071 2264 39948 2292
rect 39071 2261 39083 2264
rect 39025 2255 39083 2261
rect 39942 2252 39948 2264
rect 40000 2252 40006 2304
rect 1104 2202 39836 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 9010 2202
rect 9062 2150 9074 2202
rect 9126 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 15010 2202
rect 15062 2150 15074 2202
rect 15126 2150 15138 2202
rect 15190 2150 15202 2202
rect 15254 2150 15266 2202
rect 15318 2150 21010 2202
rect 21062 2150 21074 2202
rect 21126 2150 21138 2202
rect 21190 2150 21202 2202
rect 21254 2150 21266 2202
rect 21318 2150 27010 2202
rect 27062 2150 27074 2202
rect 27126 2150 27138 2202
rect 27190 2150 27202 2202
rect 27254 2150 27266 2202
rect 27318 2150 33010 2202
rect 33062 2150 33074 2202
rect 33126 2150 33138 2202
rect 33190 2150 33202 2202
rect 33254 2150 33266 2202
rect 33318 2150 39010 2202
rect 39062 2150 39074 2202
rect 39126 2150 39138 2202
rect 39190 2150 39202 2202
rect 39254 2150 39266 2202
rect 39318 2150 39836 2202
rect 1104 2128 39836 2150
rect 14274 2048 14280 2100
rect 14332 2088 14338 2100
rect 18322 2088 18328 2100
rect 14332 2060 18328 2088
rect 14332 2048 14338 2060
rect 18322 2048 18328 2060
rect 18380 2048 18386 2100
rect 20806 2048 20812 2100
rect 20864 2088 20870 2100
rect 22002 2088 22008 2100
rect 20864 2060 22008 2088
rect 20864 2048 20870 2060
rect 22002 2048 22008 2060
rect 22060 2048 22066 2100
rect 24670 2048 24676 2100
rect 24728 2088 24734 2100
rect 27430 2088 27436 2100
rect 24728 2060 27436 2088
rect 24728 2048 24734 2060
rect 27430 2048 27436 2060
rect 27488 2048 27494 2100
rect 27522 2048 27528 2100
rect 27580 2088 27586 2100
rect 32490 2088 32496 2100
rect 27580 2060 32496 2088
rect 27580 2048 27586 2060
rect 32490 2048 32496 2060
rect 32548 2048 32554 2100
rect 34422 2048 34428 2100
rect 34480 2088 34486 2100
rect 36538 2088 36544 2100
rect 34480 2060 36544 2088
rect 34480 2048 34486 2060
rect 36538 2048 36544 2060
rect 36596 2048 36602 2100
rect 4982 1980 4988 2032
rect 5040 2020 5046 2032
rect 11330 2020 11336 2032
rect 5040 1992 11336 2020
rect 5040 1980 5046 1992
rect 11330 1980 11336 1992
rect 11388 1980 11394 2032
rect 13906 1980 13912 2032
rect 13964 2020 13970 2032
rect 15194 2020 15200 2032
rect 13964 1992 15200 2020
rect 13964 1980 13970 1992
rect 15194 1980 15200 1992
rect 15252 1980 15258 2032
rect 15654 1980 15660 2032
rect 15712 2020 15718 2032
rect 22094 2020 22100 2032
rect 15712 1992 22100 2020
rect 15712 1980 15718 1992
rect 22094 1980 22100 1992
rect 22152 1980 22158 2032
rect 22554 1980 22560 2032
rect 22612 2020 22618 2032
rect 26602 2020 26608 2032
rect 22612 1992 26608 2020
rect 22612 1980 22618 1992
rect 26602 1980 26608 1992
rect 26660 1980 26666 2032
rect 26786 1980 26792 2032
rect 26844 2020 26850 2032
rect 26844 1992 28488 2020
rect 26844 1980 26850 1992
rect 14274 1952 14280 1964
rect 2746 1924 14280 1952
rect 1946 1776 1952 1828
rect 2004 1816 2010 1828
rect 2746 1816 2774 1924
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 14826 1912 14832 1964
rect 14884 1952 14890 1964
rect 15378 1952 15384 1964
rect 14884 1924 15384 1952
rect 14884 1912 14890 1924
rect 15378 1912 15384 1924
rect 15436 1912 15442 1964
rect 19518 1912 19524 1964
rect 19576 1952 19582 1964
rect 25498 1952 25504 1964
rect 19576 1924 25504 1952
rect 19576 1912 19582 1924
rect 25498 1912 25504 1924
rect 25556 1912 25562 1964
rect 25866 1912 25872 1964
rect 25924 1952 25930 1964
rect 28350 1952 28356 1964
rect 25924 1924 28356 1952
rect 25924 1912 25930 1924
rect 28350 1912 28356 1924
rect 28408 1912 28414 1964
rect 28460 1952 28488 1992
rect 28994 1980 29000 2032
rect 29052 2020 29058 2032
rect 33594 2020 33600 2032
rect 29052 1992 33600 2020
rect 29052 1980 29058 1992
rect 33594 1980 33600 1992
rect 33652 1980 33658 2032
rect 33686 1980 33692 2032
rect 33744 2020 33750 2032
rect 38838 2020 38844 2032
rect 33744 1992 38844 2020
rect 33744 1980 33750 1992
rect 38838 1980 38844 1992
rect 38896 1980 38902 2032
rect 29362 1952 29368 1964
rect 28460 1924 29368 1952
rect 29362 1912 29368 1924
rect 29420 1912 29426 1964
rect 29730 1912 29736 1964
rect 29788 1952 29794 1964
rect 30558 1952 30564 1964
rect 29788 1924 30564 1952
rect 29788 1912 29794 1924
rect 30558 1912 30564 1924
rect 30616 1912 30622 1964
rect 31938 1912 31944 1964
rect 31996 1952 32002 1964
rect 36078 1952 36084 1964
rect 31996 1924 36084 1952
rect 31996 1912 32002 1924
rect 36078 1912 36084 1924
rect 36136 1912 36142 1964
rect 4154 1844 4160 1896
rect 4212 1884 4218 1896
rect 10134 1884 10140 1896
rect 4212 1856 10140 1884
rect 4212 1844 4218 1856
rect 10134 1844 10140 1856
rect 10192 1844 10198 1896
rect 10410 1844 10416 1896
rect 10468 1884 10474 1896
rect 12894 1884 12900 1896
rect 10468 1856 12900 1884
rect 10468 1844 10474 1856
rect 12894 1844 12900 1856
rect 12952 1844 12958 1896
rect 22462 1884 22468 1896
rect 14108 1856 22468 1884
rect 2004 1788 2774 1816
rect 2004 1776 2010 1788
rect 9858 1776 9864 1828
rect 9916 1816 9922 1828
rect 12526 1816 12532 1828
rect 9916 1788 12532 1816
rect 9916 1776 9922 1788
rect 12526 1776 12532 1788
rect 12584 1776 12590 1828
rect 1670 1708 1676 1760
rect 1728 1748 1734 1760
rect 14108 1748 14136 1856
rect 22462 1844 22468 1856
rect 22520 1844 22526 1896
rect 24578 1844 24584 1896
rect 24636 1884 24642 1896
rect 35066 1884 35072 1896
rect 24636 1856 35072 1884
rect 24636 1844 24642 1856
rect 35066 1844 35072 1856
rect 35124 1844 35130 1896
rect 14274 1776 14280 1828
rect 14332 1816 14338 1828
rect 29178 1816 29184 1828
rect 14332 1788 29184 1816
rect 14332 1776 14338 1788
rect 29178 1776 29184 1788
rect 29236 1776 29242 1828
rect 1728 1720 14136 1748
rect 1728 1708 1734 1720
rect 17218 1708 17224 1760
rect 17276 1748 17282 1760
rect 25866 1748 25872 1760
rect 17276 1720 25872 1748
rect 17276 1708 17282 1720
rect 25866 1708 25872 1720
rect 25924 1708 25930 1760
rect 28258 1708 28264 1760
rect 28316 1748 28322 1760
rect 38930 1748 38936 1760
rect 28316 1720 38936 1748
rect 28316 1708 28322 1720
rect 38930 1708 38936 1720
rect 38988 1708 38994 1760
rect 1026 1640 1032 1692
rect 1084 1680 1090 1692
rect 8754 1680 8760 1692
rect 1084 1652 8760 1680
rect 1084 1640 1090 1652
rect 8754 1640 8760 1652
rect 8812 1680 8818 1692
rect 12158 1680 12164 1692
rect 8812 1652 12164 1680
rect 8812 1640 8818 1652
rect 12158 1640 12164 1652
rect 12216 1680 12222 1692
rect 19518 1680 19524 1692
rect 12216 1652 19524 1680
rect 12216 1640 12222 1652
rect 19518 1640 19524 1652
rect 19576 1640 19582 1692
rect 20622 1640 20628 1692
rect 20680 1680 20686 1692
rect 27614 1680 27620 1692
rect 20680 1652 27620 1680
rect 20680 1640 20686 1652
rect 27614 1640 27620 1652
rect 27672 1680 27678 1692
rect 27982 1680 27988 1692
rect 27672 1652 27988 1680
rect 27672 1640 27678 1652
rect 27982 1640 27988 1652
rect 28040 1640 28046 1692
rect 28166 1640 28172 1692
rect 28224 1680 28230 1692
rect 34698 1680 34704 1692
rect 28224 1652 34704 1680
rect 28224 1640 28230 1652
rect 34698 1640 34704 1652
rect 34756 1640 34762 1692
rect 4246 1572 4252 1624
rect 4304 1612 4310 1624
rect 12618 1612 12624 1624
rect 4304 1584 12624 1612
rect 4304 1572 4310 1584
rect 12618 1572 12624 1584
rect 12676 1612 12682 1624
rect 15654 1612 15660 1624
rect 12676 1584 15660 1612
rect 12676 1572 12682 1584
rect 15654 1572 15660 1584
rect 15712 1572 15718 1624
rect 15838 1572 15844 1624
rect 15896 1612 15902 1624
rect 19702 1612 19708 1624
rect 15896 1584 19708 1612
rect 15896 1572 15902 1584
rect 19702 1572 19708 1584
rect 19760 1572 19766 1624
rect 21634 1572 21640 1624
rect 21692 1612 21698 1624
rect 27522 1612 27528 1624
rect 21692 1584 27528 1612
rect 21692 1572 21698 1584
rect 27522 1572 27528 1584
rect 27580 1572 27586 1624
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 17218 1544 17224 1556
rect 8536 1516 17224 1544
rect 8536 1504 8542 1516
rect 17218 1504 17224 1516
rect 17276 1504 17282 1556
rect 20622 1544 20628 1556
rect 17512 1516 20628 1544
rect 11054 1436 11060 1488
rect 11112 1476 11118 1488
rect 16758 1476 16764 1488
rect 11112 1448 16764 1476
rect 11112 1436 11118 1448
rect 16758 1436 16764 1448
rect 16816 1436 16822 1488
rect 16942 1436 16948 1488
rect 17000 1476 17006 1488
rect 17402 1476 17408 1488
rect 17000 1448 17408 1476
rect 17000 1436 17006 1448
rect 17402 1436 17408 1448
rect 17460 1436 17466 1488
rect 7190 1368 7196 1420
rect 7248 1408 7254 1420
rect 9214 1408 9220 1420
rect 7248 1380 9220 1408
rect 7248 1368 7254 1380
rect 9214 1368 9220 1380
rect 9272 1368 9278 1420
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 17512 1408 17540 1516
rect 20622 1504 20628 1516
rect 20680 1504 20686 1556
rect 24670 1504 24676 1556
rect 24728 1544 24734 1556
rect 27890 1544 27896 1556
rect 24728 1516 27896 1544
rect 24728 1504 24734 1516
rect 27890 1504 27896 1516
rect 27948 1504 27954 1556
rect 17586 1436 17592 1488
rect 17644 1476 17650 1488
rect 19242 1476 19248 1488
rect 17644 1448 19248 1476
rect 17644 1436 17650 1448
rect 19242 1436 19248 1448
rect 19300 1436 19306 1488
rect 34606 1436 34612 1488
rect 34664 1476 34670 1488
rect 35250 1476 35256 1488
rect 34664 1448 35256 1476
rect 34664 1436 34670 1448
rect 35250 1436 35256 1448
rect 35308 1436 35314 1488
rect 11388 1380 17540 1408
rect 11388 1368 11394 1380
rect 17678 1368 17684 1420
rect 17736 1408 17742 1420
rect 18690 1408 18696 1420
rect 17736 1380 18696 1408
rect 17736 1368 17742 1380
rect 18690 1368 18696 1380
rect 18748 1368 18754 1420
rect 19150 1368 19156 1420
rect 19208 1408 19214 1420
rect 20346 1408 20352 1420
rect 19208 1380 20352 1408
rect 19208 1368 19214 1380
rect 20346 1368 20352 1380
rect 20404 1368 20410 1420
rect 21910 1368 21916 1420
rect 21968 1408 21974 1420
rect 31846 1408 31852 1420
rect 21968 1380 31852 1408
rect 21968 1368 21974 1380
rect 31846 1368 31852 1380
rect 31904 1368 31910 1420
rect 34238 1368 34244 1420
rect 34296 1408 34302 1420
rect 36814 1408 36820 1420
rect 34296 1380 36820 1408
rect 34296 1368 34302 1380
rect 36814 1368 36820 1380
rect 36872 1368 36878 1420
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 4614 1340 4620 1352
rect 3476 1312 4620 1340
rect 3476 1300 3482 1312
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 4706 1300 4712 1352
rect 4764 1340 4770 1352
rect 7650 1340 7656 1352
rect 4764 1312 7656 1340
rect 4764 1300 4770 1312
rect 7650 1300 7656 1312
rect 7708 1300 7714 1352
rect 8846 1300 8852 1352
rect 8904 1340 8910 1352
rect 10134 1340 10140 1352
rect 8904 1312 10140 1340
rect 8904 1300 8910 1312
rect 10134 1300 10140 1312
rect 10192 1300 10198 1352
rect 12066 1300 12072 1352
rect 12124 1340 12130 1352
rect 12894 1340 12900 1352
rect 12124 1312 12900 1340
rect 12124 1300 12130 1312
rect 12894 1300 12900 1312
rect 12952 1300 12958 1352
rect 13078 1300 13084 1352
rect 13136 1340 13142 1352
rect 15102 1340 15108 1352
rect 13136 1312 15108 1340
rect 13136 1300 13142 1312
rect 15102 1300 15108 1312
rect 15160 1300 15166 1352
rect 17310 1300 17316 1352
rect 17368 1340 17374 1352
rect 19794 1340 19800 1352
rect 17368 1312 19800 1340
rect 17368 1300 17374 1312
rect 19794 1300 19800 1312
rect 19852 1300 19858 1352
rect 20070 1300 20076 1352
rect 20128 1340 20134 1352
rect 21818 1340 21824 1352
rect 20128 1312 21824 1340
rect 20128 1300 20134 1312
rect 21818 1300 21824 1312
rect 21876 1300 21882 1352
rect 24486 1300 24492 1352
rect 24544 1340 24550 1352
rect 25314 1340 25320 1352
rect 24544 1312 25320 1340
rect 24544 1300 24550 1312
rect 25314 1300 25320 1312
rect 25372 1300 25378 1352
rect 33502 1340 33508 1352
rect 30760 1312 33508 1340
rect 3602 1232 3608 1284
rect 3660 1272 3666 1284
rect 5994 1272 6000 1284
rect 3660 1244 6000 1272
rect 3660 1232 3666 1244
rect 5994 1232 6000 1244
rect 6052 1232 6058 1284
rect 12986 1232 12992 1284
rect 13044 1272 13050 1284
rect 16206 1272 16212 1284
rect 13044 1244 16212 1272
rect 13044 1232 13050 1244
rect 16206 1232 16212 1244
rect 16264 1232 16270 1284
rect 16482 1232 16488 1284
rect 16540 1272 16546 1284
rect 20806 1272 20812 1284
rect 16540 1244 20812 1272
rect 16540 1232 16546 1244
rect 20806 1232 20812 1244
rect 20864 1232 20870 1284
rect 22002 1232 22008 1284
rect 22060 1272 22066 1284
rect 24854 1272 24860 1284
rect 22060 1244 24860 1272
rect 22060 1232 22066 1244
rect 24854 1232 24860 1244
rect 24912 1232 24918 1284
rect 25038 1232 25044 1284
rect 25096 1272 25102 1284
rect 26694 1272 26700 1284
rect 25096 1244 26700 1272
rect 25096 1232 25102 1244
rect 26694 1232 26700 1244
rect 26752 1232 26758 1284
rect 30282 1232 30288 1284
rect 30340 1272 30346 1284
rect 30760 1272 30788 1312
rect 33502 1300 33508 1312
rect 33560 1300 33566 1352
rect 36354 1300 36360 1352
rect 36412 1340 36418 1352
rect 37274 1340 37280 1352
rect 36412 1312 37280 1340
rect 36412 1300 36418 1312
rect 37274 1300 37280 1312
rect 37332 1300 37338 1352
rect 32766 1272 32772 1284
rect 30340 1244 30788 1272
rect 30852 1244 32772 1272
rect 30340 1232 30346 1244
rect 2498 1164 2504 1216
rect 2556 1204 2562 1216
rect 2556 1176 2774 1204
rect 2556 1164 2562 1176
rect 2746 1136 2774 1176
rect 4890 1164 4896 1216
rect 4948 1204 4954 1216
rect 8754 1204 8760 1216
rect 4948 1176 8760 1204
rect 4948 1164 4954 1176
rect 8754 1164 8760 1176
rect 8812 1164 8818 1216
rect 9490 1164 9496 1216
rect 9548 1204 9554 1216
rect 10686 1204 10692 1216
rect 9548 1176 10692 1204
rect 9548 1164 9554 1176
rect 10686 1164 10692 1176
rect 10744 1164 10750 1216
rect 13538 1164 13544 1216
rect 13596 1204 13602 1216
rect 13596 1176 17632 1204
rect 13596 1164 13602 1176
rect 6822 1136 6828 1148
rect 2746 1108 6828 1136
rect 6822 1096 6828 1108
rect 6880 1096 6886 1148
rect 7742 1096 7748 1148
rect 7800 1136 7806 1148
rect 11606 1136 11612 1148
rect 7800 1108 11612 1136
rect 7800 1096 7806 1108
rect 11606 1096 11612 1108
rect 11664 1096 11670 1148
rect 17494 1136 17500 1148
rect 12406 1108 17500 1136
rect 3970 1028 3976 1080
rect 4028 1068 4034 1080
rect 12406 1068 12434 1108
rect 17494 1096 17500 1108
rect 17552 1096 17558 1148
rect 4028 1040 12434 1068
rect 4028 1028 4034 1040
rect 16390 1028 16396 1080
rect 16448 1068 16454 1080
rect 17604 1068 17632 1176
rect 21726 1164 21732 1216
rect 21784 1204 21790 1216
rect 24302 1204 24308 1216
rect 21784 1176 24308 1204
rect 21784 1164 21790 1176
rect 24302 1164 24308 1176
rect 24360 1164 24366 1216
rect 30852 1204 30880 1244
rect 32766 1232 32772 1244
rect 32824 1232 32830 1284
rect 35250 1232 35256 1284
rect 35308 1272 35314 1284
rect 37182 1272 37188 1284
rect 35308 1244 37188 1272
rect 35308 1232 35314 1244
rect 37182 1232 37188 1244
rect 37240 1232 37246 1284
rect 26712 1176 30880 1204
rect 26712 1148 26740 1176
rect 31110 1164 31116 1216
rect 31168 1204 31174 1216
rect 36446 1204 36452 1216
rect 31168 1176 36452 1204
rect 31168 1164 31174 1176
rect 36446 1164 36452 1176
rect 36504 1164 36510 1216
rect 17678 1096 17684 1148
rect 17736 1136 17742 1148
rect 23014 1136 23020 1148
rect 17736 1108 23020 1136
rect 17736 1096 17742 1108
rect 23014 1096 23020 1108
rect 23072 1096 23078 1148
rect 23106 1096 23112 1148
rect 23164 1136 23170 1148
rect 26418 1136 26424 1148
rect 23164 1108 26424 1136
rect 23164 1096 23170 1108
rect 26418 1096 26424 1108
rect 26476 1096 26482 1148
rect 26694 1096 26700 1148
rect 26752 1096 26758 1148
rect 29178 1096 29184 1148
rect 29236 1136 29242 1148
rect 34146 1136 34152 1148
rect 29236 1108 34152 1136
rect 29236 1096 29242 1108
rect 34146 1096 34152 1108
rect 34204 1096 34210 1148
rect 34974 1096 34980 1148
rect 35032 1136 35038 1148
rect 36262 1136 36268 1148
rect 35032 1108 36268 1136
rect 35032 1096 35038 1108
rect 36262 1096 36268 1108
rect 36320 1096 36326 1148
rect 24026 1068 24032 1080
rect 16448 1040 17448 1068
rect 17604 1040 24032 1068
rect 16448 1028 16454 1040
rect 8294 960 8300 1012
rect 8352 1000 8358 1012
rect 11330 1000 11336 1012
rect 8352 972 11336 1000
rect 8352 960 8358 972
rect 11330 960 11336 972
rect 11388 960 11394 1012
rect 16482 960 16488 1012
rect 16540 1000 16546 1012
rect 17310 1000 17316 1012
rect 16540 972 17316 1000
rect 16540 960 16546 972
rect 17310 960 17316 972
rect 17368 960 17374 1012
rect 17420 1000 17448 1040
rect 24026 1028 24032 1040
rect 24084 1028 24090 1080
rect 24210 1028 24216 1080
rect 24268 1068 24274 1080
rect 24946 1068 24952 1080
rect 24268 1040 24952 1068
rect 24268 1028 24274 1040
rect 24946 1028 24952 1040
rect 25004 1028 25010 1080
rect 28994 1068 29000 1080
rect 25240 1040 29000 1068
rect 25240 1000 25268 1040
rect 28994 1028 29000 1040
rect 29052 1028 29058 1080
rect 32674 1068 32680 1080
rect 31726 1040 32680 1068
rect 17420 972 25268 1000
rect 26418 960 26424 1012
rect 26476 1000 26482 1012
rect 31726 1000 31754 1040
rect 32674 1028 32680 1040
rect 32732 1028 32738 1080
rect 34698 1028 34704 1080
rect 34756 1068 34762 1080
rect 36998 1068 37004 1080
rect 34756 1040 37004 1068
rect 34756 1028 34762 1040
rect 36998 1028 37004 1040
rect 37056 1028 37062 1080
rect 26476 972 31754 1000
rect 26476 960 26482 972
rect 31938 960 31944 1012
rect 31996 1000 32002 1012
rect 35066 1000 35072 1012
rect 31996 972 35072 1000
rect 31996 960 32002 972
rect 35066 960 35072 972
rect 35124 960 35130 1012
rect 6362 892 6368 944
rect 6420 932 6426 944
rect 6420 904 9168 932
rect 6420 892 6426 904
rect 7466 824 7472 876
rect 7524 864 7530 876
rect 9030 864 9036 876
rect 7524 836 9036 864
rect 7524 824 7530 836
rect 9030 824 9036 836
rect 9088 824 9094 876
rect 9140 864 9168 904
rect 9214 892 9220 944
rect 9272 932 9278 944
rect 11790 932 11796 944
rect 9272 904 11796 932
rect 9272 892 9278 904
rect 11790 892 11796 904
rect 11848 892 11854 944
rect 24762 932 24768 944
rect 16408 904 24768 932
rect 16408 864 16436 904
rect 24762 892 24768 904
rect 24820 892 24826 944
rect 25590 892 25596 944
rect 25648 932 25654 944
rect 27338 932 27344 944
rect 25648 904 27344 932
rect 25648 892 25654 904
rect 27338 892 27344 904
rect 27396 892 27402 944
rect 28902 892 28908 944
rect 28960 932 28966 944
rect 31570 932 31576 944
rect 28960 904 31576 932
rect 28960 892 28966 904
rect 31570 892 31576 904
rect 31628 892 31634 944
rect 31662 892 31668 944
rect 31720 932 31726 944
rect 31720 904 33824 932
rect 31720 892 31726 904
rect 9140 836 16436 864
rect 16482 824 16488 876
rect 16540 864 16546 876
rect 22094 864 22100 876
rect 16540 836 22100 864
rect 16540 824 16546 836
rect 22094 824 22100 836
rect 22152 824 22158 876
rect 22278 824 22284 876
rect 22336 864 22342 876
rect 26510 864 26516 876
rect 22336 836 26516 864
rect 22336 824 22342 836
rect 26510 824 26516 836
rect 26568 824 26574 876
rect 30006 824 30012 876
rect 30064 864 30070 876
rect 32306 864 32312 876
rect 30064 836 32312 864
rect 30064 824 30070 836
rect 32306 824 32312 836
rect 32364 824 32370 876
rect 2682 756 2688 808
rect 2740 796 2746 808
rect 2740 768 7788 796
rect 2740 756 2746 768
rect 2590 688 2596 740
rect 2648 728 2654 740
rect 4890 728 4896 740
rect 2648 700 4896 728
rect 2648 688 2654 700
rect 4890 688 4896 700
rect 4948 688 4954 740
rect 2314 620 2320 672
rect 2372 660 2378 672
rect 7760 660 7788 768
rect 13998 756 14004 808
rect 14056 796 14062 808
rect 14056 768 15792 796
rect 14056 756 14062 768
rect 14550 688 14556 740
rect 14608 728 14614 740
rect 15654 728 15660 740
rect 14608 700 15660 728
rect 14608 688 14614 700
rect 15654 688 15660 700
rect 15712 688 15718 740
rect 15764 728 15792 768
rect 17310 756 17316 808
rect 17368 796 17374 808
rect 27706 796 27712 808
rect 17368 768 27712 796
rect 17368 756 17374 768
rect 27706 756 27712 768
rect 27764 756 27770 808
rect 30374 756 30380 808
rect 30432 796 30438 808
rect 33042 796 33048 808
rect 30432 768 33048 796
rect 30432 756 30438 768
rect 33042 756 33048 768
rect 33100 756 33106 808
rect 33796 796 33824 904
rect 33870 892 33876 944
rect 33928 932 33934 944
rect 34790 932 34796 944
rect 33928 904 34796 932
rect 33928 892 33934 904
rect 34790 892 34796 904
rect 34848 892 34854 944
rect 36078 796 36084 808
rect 33796 768 36084 796
rect 36078 756 36084 768
rect 36136 756 36142 808
rect 24670 728 24676 740
rect 15764 700 24676 728
rect 24670 688 24676 700
rect 24728 688 24734 740
rect 24762 688 24768 740
rect 24820 728 24826 740
rect 26326 728 26332 740
rect 24820 700 26332 728
rect 24820 688 24826 700
rect 26326 688 26332 700
rect 26384 688 26390 740
rect 27798 688 27804 740
rect 27856 728 27862 740
rect 30650 728 30656 740
rect 27856 700 30656 728
rect 27856 688 27862 700
rect 30650 688 30656 700
rect 30708 688 30714 740
rect 22922 660 22928 672
rect 2372 632 2774 660
rect 7760 632 22928 660
rect 2372 620 2378 632
rect 2746 592 2774 632
rect 22922 620 22928 632
rect 22980 620 22986 672
rect 29454 620 29460 672
rect 29512 660 29518 672
rect 35618 660 35624 672
rect 29512 632 35624 660
rect 29512 620 29518 632
rect 35618 620 35624 632
rect 35676 620 35682 672
rect 35802 620 35808 672
rect 35860 660 35866 672
rect 37642 660 37648 672
rect 35860 632 37648 660
rect 35860 620 35866 632
rect 37642 620 37648 632
rect 37700 620 37706 672
rect 9674 592 9680 604
rect 2746 564 9680 592
rect 9674 552 9680 564
rect 9732 552 9738 604
rect 11422 552 11428 604
rect 11480 592 11486 604
rect 23658 592 23664 604
rect 11480 564 23664 592
rect 11480 552 11486 564
rect 23658 552 23664 564
rect 23716 552 23722 604
rect 26970 552 26976 604
rect 27028 592 27034 604
rect 30466 592 30472 604
rect 27028 564 30472 592
rect 27028 552 27034 564
rect 30466 552 30472 564
rect 30524 552 30530 604
rect 31386 552 31392 604
rect 31444 592 31450 604
rect 35342 592 35348 604
rect 31444 564 35348 592
rect 31444 552 31450 564
rect 35342 552 35348 564
rect 35400 552 35406 604
rect 2038 484 2044 536
rect 2096 524 2102 536
rect 13998 524 14004 536
rect 2096 496 14004 524
rect 2096 484 2102 496
rect 13998 484 14004 496
rect 14056 484 14062 536
rect 14090 484 14096 536
rect 14148 524 14154 536
rect 17310 524 17316 536
rect 14148 496 17316 524
rect 14148 484 14154 496
rect 17310 484 17316 496
rect 17368 484 17374 536
rect 17954 484 17960 536
rect 18012 524 18018 536
rect 19426 524 19432 536
rect 18012 496 19432 524
rect 18012 484 18018 496
rect 19426 484 19432 496
rect 19484 484 19490 536
rect 28074 484 28080 536
rect 28132 524 28138 536
rect 34882 524 34888 536
rect 28132 496 34888 524
rect 28132 484 28138 496
rect 34882 484 34888 496
rect 34940 484 34946 536
rect 36078 484 36084 536
rect 36136 524 36142 536
rect 38746 524 38752 536
rect 36136 496 38752 524
rect 36136 484 36142 496
rect 38746 484 38752 496
rect 38804 484 38810 536
rect 5258 416 5264 468
rect 5316 456 5322 468
rect 12066 456 12072 468
rect 5316 428 12072 456
rect 5316 416 5322 428
rect 12066 416 12072 428
rect 12124 416 12130 468
rect 12802 416 12808 468
rect 12860 456 12866 468
rect 14826 456 14832 468
rect 12860 428 14832 456
rect 12860 416 12866 428
rect 14826 416 14832 428
rect 14884 416 14890 468
rect 14918 416 14924 468
rect 14976 456 14982 468
rect 18138 456 18144 468
rect 14976 428 18144 456
rect 14976 416 14982 428
rect 18138 416 18144 428
rect 18196 416 18202 468
rect 23658 416 23664 468
rect 23716 456 23722 468
rect 29086 456 29092 468
rect 23716 428 29092 456
rect 23716 416 23722 428
rect 29086 416 29092 428
rect 29144 416 29150 468
rect 30834 416 30840 468
rect 30892 456 30898 468
rect 32582 456 32588 468
rect 30892 428 32588 456
rect 30892 416 30898 428
rect 32582 416 32588 428
rect 32640 416 32646 468
rect 11698 348 11704 400
rect 11756 388 11762 400
rect 14550 388 14556 400
rect 11756 360 14556 388
rect 11756 348 11762 360
rect 14550 348 14556 360
rect 14608 348 14614 400
rect 14734 348 14740 400
rect 14792 388 14798 400
rect 22186 388 22192 400
rect 14792 360 22192 388
rect 14792 348 14798 360
rect 22186 348 22192 360
rect 22244 348 22250 400
rect 24026 348 24032 400
rect 24084 388 24090 400
rect 24084 360 25912 388
rect 24084 348 24090 360
rect 5902 280 5908 332
rect 5960 320 5966 332
rect 5960 292 14412 320
rect 5960 280 5966 292
rect 8570 212 8576 264
rect 8628 252 8634 264
rect 12250 252 12256 264
rect 8628 224 12256 252
rect 8628 212 8634 224
rect 12250 212 12256 224
rect 12308 212 12314 264
rect 14384 252 14412 292
rect 14458 280 14464 332
rect 14516 320 14522 332
rect 17862 320 17868 332
rect 14516 292 17868 320
rect 14516 280 14522 292
rect 17862 280 17868 292
rect 17920 280 17926 332
rect 20530 280 20536 332
rect 20588 320 20594 332
rect 21174 320 21180 332
rect 20588 292 21180 320
rect 20588 280 20594 292
rect 21174 280 21180 292
rect 21232 280 21238 332
rect 22554 280 22560 332
rect 22612 320 22618 332
rect 25774 320 25780 332
rect 22612 292 25780 320
rect 22612 280 22618 292
rect 25774 280 25780 292
rect 25832 280 25838 332
rect 25884 320 25912 360
rect 26142 348 26148 400
rect 26200 388 26206 400
rect 29638 388 29644 400
rect 26200 360 29644 388
rect 26200 348 26206 360
rect 29638 348 29644 360
rect 29696 348 29702 400
rect 33594 348 33600 400
rect 33652 388 33658 400
rect 37826 388 37832 400
rect 33652 360 37832 388
rect 33652 348 33658 360
rect 37826 348 37832 360
rect 37884 348 37890 400
rect 29270 320 29276 332
rect 25884 292 29276 320
rect 29270 280 29276 292
rect 29328 280 29334 332
rect 30558 280 30564 332
rect 30616 320 30622 332
rect 34606 320 34612 332
rect 30616 292 34612 320
rect 30616 280 30622 292
rect 34606 280 34612 292
rect 34664 280 34670 332
rect 15746 252 15752 264
rect 14384 224 15752 252
rect 15746 212 15752 224
rect 15804 212 15810 264
rect 27246 212 27252 264
rect 27304 252 27310 264
rect 33410 252 33416 264
rect 27304 224 33416 252
rect 27304 212 27310 224
rect 33410 212 33416 224
rect 33468 212 33474 264
rect 11238 144 11244 196
rect 11296 184 11302 196
rect 16022 184 16028 196
rect 11296 156 16028 184
rect 11296 144 11302 156
rect 16022 144 16028 156
rect 16080 144 16086 196
rect 27522 144 27528 196
rect 27580 184 27586 196
rect 31294 184 31300 196
rect 27580 156 31300 184
rect 27580 144 27586 156
rect 31294 144 31300 156
rect 31352 144 31358 196
rect 36630 144 36636 196
rect 36688 184 36694 196
rect 37550 184 37556 196
rect 36688 156 37556 184
rect 36688 144 36694 156
rect 37550 144 37556 156
rect 37608 144 37614 196
rect 22922 8 22928 60
rect 22980 48 22986 60
rect 31478 48 31484 60
rect 22980 20 31484 48
rect 22980 8 22986 20
rect 31478 8 31484 20
rect 31536 8 31542 60
<< via1 >>
rect 5632 10820 5684 10872
rect 16396 10820 16448 10872
rect 2872 10752 2924 10804
rect 18328 10752 18380 10804
rect 7656 10684 7708 10736
rect 19432 10684 19484 10736
rect 12624 10616 12676 10668
rect 13360 10616 13412 10668
rect 28540 10616 28592 10668
rect 14372 10548 14424 10600
rect 23940 10548 23992 10600
rect 9772 10480 9824 10532
rect 17684 10480 17736 10532
rect 17776 10480 17828 10532
rect 6184 10412 6236 10464
rect 17040 10412 17092 10464
rect 17224 10412 17276 10464
rect 22744 10412 22796 10464
rect 33784 10412 33836 10464
rect 9312 10344 9364 10396
rect 32404 10344 32456 10396
rect 1584 10208 1636 10260
rect 28908 10276 28960 10328
rect 2596 10072 2648 10124
rect 31208 10208 31260 10260
rect 9588 10140 9640 10192
rect 17224 10140 17276 10192
rect 17960 10140 18012 10192
rect 26700 10140 26752 10192
rect 12256 10072 12308 10124
rect 21916 10072 21968 10124
rect 35624 10140 35676 10192
rect 16488 10004 16540 10056
rect 27068 10072 27120 10124
rect 36084 10072 36136 10124
rect 26976 10004 27028 10056
rect 34060 10004 34112 10056
rect 1308 9936 1360 9988
rect 21364 9936 21416 9988
rect 22468 9936 22520 9988
rect 34244 9936 34296 9988
rect 2504 9868 2556 9920
rect 12348 9868 12400 9920
rect 21916 9868 21968 9920
rect 34428 9868 34480 9920
rect 2320 9800 2372 9852
rect 9680 9800 9732 9852
rect 16580 9800 16632 9852
rect 7380 9732 7432 9784
rect 3792 9664 3844 9716
rect 15384 9732 15436 9784
rect 20720 9732 20772 9784
rect 15476 9664 15528 9716
rect 20444 9664 20496 9716
rect 21456 9664 21508 9716
rect 22100 9800 22152 9852
rect 35992 9800 36044 9852
rect 22652 9732 22704 9784
rect 23664 9732 23716 9784
rect 24676 9732 24728 9784
rect 26976 9664 27028 9716
rect 28172 9664 28224 9716
rect 29644 9664 29696 9716
rect 33416 9664 33468 9716
rect 16488 9596 16540 9648
rect 22836 9596 22888 9648
rect 6276 9528 6328 9580
rect 8668 9460 8720 9512
rect 13084 9392 13136 9444
rect 3700 9324 3752 9376
rect 12072 9324 12124 9376
rect 2780 9256 2832 9308
rect 4252 9256 4304 9308
rect 9496 9256 9548 9308
rect 13268 9528 13320 9580
rect 15016 9528 15068 9580
rect 23572 9528 23624 9580
rect 31484 9460 31536 9512
rect 13268 9392 13320 9444
rect 20628 9392 20680 9444
rect 22192 9392 22244 9444
rect 30012 9392 30064 9444
rect 35256 9392 35308 9444
rect 16856 9324 16908 9376
rect 25688 9324 25740 9376
rect 25780 9324 25832 9376
rect 36636 9324 36688 9376
rect 26700 9256 26752 9308
rect 37188 9256 37240 9308
rect 38568 9256 38620 9308
rect 6644 9188 6696 9240
rect 10876 9188 10928 9240
rect 12532 9188 12584 9240
rect 15016 9188 15068 9240
rect 15108 9188 15160 9240
rect 17960 9188 18012 9240
rect 19524 9188 19576 9240
rect 24124 9188 24176 9240
rect 24216 9188 24268 9240
rect 36820 9188 36872 9240
rect 8484 9120 8536 9172
rect 20536 9120 20588 9172
rect 20628 9120 20680 9172
rect 22192 9120 22244 9172
rect 22284 9120 22336 9172
rect 26792 9120 26844 9172
rect 2872 9052 2924 9104
rect 4528 9052 4580 9104
rect 5632 9052 5684 9104
rect 8576 9052 8628 9104
rect 31392 9120 31444 9172
rect 4068 8984 4120 9036
rect 10232 8984 10284 9036
rect 2412 8916 2464 8968
rect 12532 8916 12584 8968
rect 1860 8848 1912 8900
rect 5264 8848 5316 8900
rect 14832 8984 14884 9036
rect 15660 8984 15712 9036
rect 14464 8916 14516 8968
rect 22008 8916 22060 8968
rect 23848 8984 23900 9036
rect 35808 8984 35860 9036
rect 24400 8916 24452 8968
rect 26332 8916 26384 8968
rect 37372 8916 37424 8968
rect 12808 8848 12860 8900
rect 19708 8848 19760 8900
rect 20720 8848 20772 8900
rect 24584 8848 24636 8900
rect 25872 8848 25924 8900
rect 32864 8848 32916 8900
rect 33600 8848 33652 8900
rect 36360 8848 36412 8900
rect 7472 8780 7524 8832
rect 8392 8780 8444 8832
rect 16488 8780 16540 8832
rect 19616 8780 19668 8832
rect 22284 8780 22336 8832
rect 22376 8780 22428 8832
rect 28356 8780 28408 8832
rect 28908 8780 28960 8832
rect 30288 8780 30340 8832
rect 30748 8780 30800 8832
rect 37740 8848 37792 8900
rect 36912 8780 36964 8832
rect 38476 8780 38528 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 9010 8678 9062 8730
rect 9074 8678 9126 8730
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 15010 8678 15062 8730
rect 15074 8678 15126 8730
rect 15138 8678 15190 8730
rect 15202 8678 15254 8730
rect 15266 8678 15318 8730
rect 21010 8678 21062 8730
rect 21074 8678 21126 8730
rect 21138 8678 21190 8730
rect 21202 8678 21254 8730
rect 21266 8678 21318 8730
rect 27010 8678 27062 8730
rect 27074 8678 27126 8730
rect 27138 8678 27190 8730
rect 27202 8678 27254 8730
rect 27266 8678 27318 8730
rect 33010 8678 33062 8730
rect 33074 8678 33126 8730
rect 33138 8678 33190 8730
rect 33202 8678 33254 8730
rect 33266 8678 33318 8730
rect 39010 8678 39062 8730
rect 39074 8678 39126 8730
rect 39138 8678 39190 8730
rect 39202 8678 39254 8730
rect 39266 8678 39318 8730
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 2872 8576 2924 8628
rect 1676 8508 1728 8560
rect 3700 8576 3752 8628
rect 4160 8576 4212 8628
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 6000 8576 6052 8628
rect 6092 8576 6144 8628
rect 7196 8576 7248 8628
rect 7472 8576 7524 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 3332 8551 3384 8560
rect 3332 8517 3341 8551
rect 3341 8517 3375 8551
rect 3375 8517 3384 8551
rect 3332 8508 3384 8517
rect 3884 8551 3936 8560
rect 3884 8517 3893 8551
rect 3893 8517 3927 8551
rect 3927 8517 3936 8551
rect 3884 8508 3936 8517
rect 4252 8551 4304 8560
rect 4252 8517 4261 8551
rect 4261 8517 4295 8551
rect 4295 8517 4304 8551
rect 4252 8508 4304 8517
rect 4436 8551 4488 8560
rect 4436 8517 4445 8551
rect 4445 8517 4479 8551
rect 4479 8517 4488 8551
rect 4436 8508 4488 8517
rect 4068 8440 4120 8492
rect 5448 8508 5500 8560
rect 5540 8551 5592 8560
rect 5540 8517 5549 8551
rect 5549 8517 5583 8551
rect 5583 8517 5592 8551
rect 5540 8508 5592 8517
rect 8300 8576 8352 8628
rect 9404 8576 9456 8628
rect 10508 8576 10560 8628
rect 11612 8576 11664 8628
rect 12716 8576 12768 8628
rect 13820 8576 13872 8628
rect 14924 8576 14976 8628
rect 15660 8619 15712 8628
rect 15660 8585 15669 8619
rect 15669 8585 15703 8619
rect 15703 8585 15712 8619
rect 15660 8576 15712 8585
rect 16028 8576 16080 8628
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 17132 8576 17184 8628
rect 18236 8576 18288 8628
rect 19340 8576 19392 8628
rect 19708 8576 19760 8628
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 4988 8440 5040 8492
rect 5264 8440 5316 8492
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 5724 8372 5776 8424
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 8576 8551 8628 8560
rect 8576 8517 8585 8551
rect 8585 8517 8619 8551
rect 8619 8517 8628 8551
rect 8576 8508 8628 8517
rect 9680 8508 9732 8560
rect 9588 8440 9640 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 11152 8508 11204 8560
rect 11244 8551 11296 8560
rect 11244 8517 11253 8551
rect 11253 8517 11287 8551
rect 11287 8517 11296 8551
rect 11244 8508 11296 8517
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 14648 8508 14700 8560
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 14280 8372 14332 8424
rect 15384 8440 15436 8492
rect 15752 8440 15804 8492
rect 16580 8440 16632 8492
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 17500 8440 17552 8492
rect 17316 8415 17368 8424
rect 17316 8381 17325 8415
rect 17325 8381 17359 8415
rect 17359 8381 17368 8415
rect 17316 8372 17368 8381
rect 20904 8508 20956 8560
rect 20444 8440 20496 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 21548 8576 21600 8628
rect 22376 8619 22428 8628
rect 22376 8585 22385 8619
rect 22385 8585 22419 8619
rect 22419 8585 22428 8619
rect 22376 8576 22428 8585
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 23756 8576 23808 8628
rect 24768 8576 24820 8628
rect 25964 8576 26016 8628
rect 29276 8576 29328 8628
rect 30380 8576 30432 8628
rect 31668 8576 31720 8628
rect 31760 8576 31812 8628
rect 32588 8576 32640 8628
rect 33692 8576 33744 8628
rect 34796 8576 34848 8628
rect 35900 8576 35952 8628
rect 36636 8619 36688 8628
rect 36636 8585 36645 8619
rect 36645 8585 36679 8619
rect 36679 8585 36688 8619
rect 36636 8576 36688 8585
rect 20996 8372 21048 8424
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22376 8440 22428 8492
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 24952 8440 25004 8492
rect 26332 8483 26384 8492
rect 26332 8449 26341 8483
rect 26341 8449 26375 8483
rect 26375 8449 26384 8483
rect 26332 8440 26384 8449
rect 27436 8483 27488 8492
rect 27436 8449 27445 8483
rect 27445 8449 27479 8483
rect 27479 8449 27488 8483
rect 27436 8440 27488 8449
rect 8760 8304 8812 8356
rect 9680 8304 9732 8356
rect 4804 8236 4856 8288
rect 8300 8236 8352 8288
rect 8392 8236 8444 8288
rect 11428 8236 11480 8288
rect 14556 8236 14608 8288
rect 18236 8304 18288 8356
rect 18052 8236 18104 8288
rect 19156 8236 19208 8288
rect 21272 8279 21324 8288
rect 21272 8245 21281 8279
rect 21281 8245 21315 8279
rect 21315 8245 21324 8279
rect 21272 8236 21324 8245
rect 21456 8304 21508 8356
rect 22192 8304 22244 8356
rect 23112 8236 23164 8288
rect 23480 8279 23532 8288
rect 23480 8245 23489 8279
rect 23489 8245 23523 8279
rect 23523 8245 23532 8279
rect 23480 8236 23532 8245
rect 26884 8372 26936 8424
rect 24860 8236 24912 8288
rect 26332 8304 26384 8356
rect 25504 8236 25556 8288
rect 29644 8347 29696 8356
rect 29644 8313 29653 8347
rect 29653 8313 29687 8347
rect 29687 8313 29696 8347
rect 29644 8304 29696 8313
rect 28172 8279 28224 8288
rect 28172 8245 28181 8279
rect 28181 8245 28215 8279
rect 28215 8245 28224 8279
rect 28172 8236 28224 8245
rect 29460 8236 29512 8288
rect 30748 8483 30800 8492
rect 30748 8449 30757 8483
rect 30757 8449 30791 8483
rect 30791 8449 30800 8483
rect 30748 8440 30800 8449
rect 36176 8508 36228 8560
rect 37280 8576 37332 8628
rect 38108 8576 38160 8628
rect 39396 8619 39448 8628
rect 39396 8585 39405 8619
rect 39405 8585 39439 8619
rect 39439 8585 39448 8619
rect 39396 8576 39448 8585
rect 38660 8508 38712 8560
rect 31208 8483 31260 8492
rect 31208 8449 31217 8483
rect 31217 8449 31251 8483
rect 31251 8449 31260 8483
rect 31208 8440 31260 8449
rect 32680 8440 32732 8492
rect 33600 8440 33652 8492
rect 33876 8440 33928 8492
rect 35164 8483 35216 8492
rect 35164 8449 35173 8483
rect 35173 8449 35207 8483
rect 35207 8449 35216 8483
rect 35164 8440 35216 8449
rect 36636 8440 36688 8492
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 30748 8304 30800 8356
rect 31668 8372 31720 8424
rect 37096 8372 37148 8424
rect 37648 8372 37700 8424
rect 38476 8440 38528 8492
rect 38844 8483 38896 8492
rect 38844 8449 38853 8483
rect 38853 8449 38887 8483
rect 38887 8449 38896 8483
rect 38844 8440 38896 8449
rect 38936 8440 38988 8492
rect 32312 8304 32364 8356
rect 34428 8236 34480 8288
rect 37832 8236 37884 8288
rect 38476 8304 38528 8356
rect 39028 8347 39080 8356
rect 39028 8313 39037 8347
rect 39037 8313 39071 8347
rect 39071 8313 39080 8347
rect 39028 8304 39080 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 13950 8134 14002 8186
rect 14014 8134 14066 8186
rect 14078 8134 14130 8186
rect 14142 8134 14194 8186
rect 14206 8134 14258 8186
rect 19950 8134 20002 8186
rect 20014 8134 20066 8186
rect 20078 8134 20130 8186
rect 20142 8134 20194 8186
rect 20206 8134 20258 8186
rect 25950 8134 26002 8186
rect 26014 8134 26066 8186
rect 26078 8134 26130 8186
rect 26142 8134 26194 8186
rect 26206 8134 26258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 37950 8134 38002 8186
rect 38014 8134 38066 8186
rect 38078 8134 38130 8186
rect 38142 8134 38194 8186
rect 38206 8134 38258 8186
rect 4528 8032 4580 8084
rect 5264 8032 5316 8084
rect 5356 8032 5408 8084
rect 10784 8032 10836 8084
rect 14464 8032 14516 8084
rect 1400 7964 1452 8016
rect 1400 7828 1452 7880
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 3608 8007 3660 8016
rect 3608 7973 3617 8007
rect 3617 7973 3651 8007
rect 3651 7973 3660 8007
rect 3608 7964 3660 7973
rect 6920 7964 6972 8016
rect 3700 7896 3752 7948
rect 6368 7939 6420 7948
rect 6368 7905 6377 7939
rect 6377 7905 6411 7939
rect 6411 7905 6420 7939
rect 6368 7896 6420 7905
rect 7196 7896 7248 7948
rect 8576 7964 8628 8016
rect 8852 7964 8904 8016
rect 10324 8007 10376 8016
rect 10324 7973 10333 8007
rect 10333 7973 10367 8007
rect 10367 7973 10376 8007
rect 10324 7964 10376 7973
rect 10692 8007 10744 8016
rect 10692 7973 10701 8007
rect 10701 7973 10735 8007
rect 10735 7973 10744 8007
rect 10692 7964 10744 7973
rect 13544 7964 13596 8016
rect 14832 7964 14884 8016
rect 16672 8032 16724 8084
rect 16948 8032 17000 8084
rect 19616 8075 19668 8084
rect 19616 8041 19625 8075
rect 19625 8041 19659 8075
rect 19659 8041 19668 8075
rect 19616 8032 19668 8041
rect 20168 8032 20220 8084
rect 20996 8032 21048 8084
rect 21640 8032 21692 8084
rect 2780 7828 2832 7880
rect 3516 7828 3568 7880
rect 1492 7803 1544 7812
rect 1492 7769 1501 7803
rect 1501 7769 1535 7803
rect 1535 7769 1544 7803
rect 1492 7760 1544 7769
rect 2044 7803 2096 7812
rect 2044 7769 2053 7803
rect 2053 7769 2087 7803
rect 2087 7769 2096 7803
rect 2044 7760 2096 7769
rect 2872 7760 2924 7812
rect 4620 7828 4672 7880
rect 1032 7692 1084 7744
rect 2596 7692 2648 7744
rect 2780 7692 2832 7744
rect 4344 7760 4396 7812
rect 4896 7760 4948 7812
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 5356 7760 5408 7812
rect 5724 7828 5776 7880
rect 7840 7828 7892 7880
rect 6276 7760 6328 7812
rect 8484 7828 8536 7880
rect 10416 7896 10468 7948
rect 11704 7896 11756 7948
rect 4160 7692 4212 7744
rect 8576 7803 8628 7812
rect 8576 7769 8585 7803
rect 8585 7769 8619 7803
rect 8619 7769 8628 7803
rect 8576 7760 8628 7769
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 8208 7692 8260 7744
rect 8852 7692 8904 7744
rect 9588 7828 9640 7880
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 9772 7828 9824 7880
rect 9496 7760 9548 7812
rect 10140 7803 10192 7812
rect 10140 7769 10149 7803
rect 10149 7769 10183 7803
rect 10183 7769 10192 7803
rect 10140 7760 10192 7769
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 11336 7828 11388 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 12440 7896 12492 7948
rect 12624 7896 12676 7948
rect 13636 7896 13688 7948
rect 15568 7896 15620 7948
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 16948 7896 17000 7948
rect 11888 7828 11940 7837
rect 12992 7828 13044 7880
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 14464 7828 14516 7880
rect 14924 7828 14976 7880
rect 16120 7828 16172 7880
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 21272 7964 21324 8016
rect 22376 8032 22428 8084
rect 24308 8032 24360 8084
rect 25044 8032 25096 8084
rect 26148 8032 26200 8084
rect 27344 8032 27396 8084
rect 24124 7964 24176 8016
rect 17960 7896 18012 7948
rect 20996 7896 21048 7948
rect 11980 7692 12032 7744
rect 12532 7692 12584 7744
rect 16304 7692 16356 7744
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 19800 7828 19852 7880
rect 20720 7871 20772 7880
rect 20720 7837 20729 7871
rect 20729 7837 20763 7871
rect 20763 7837 20772 7871
rect 20720 7828 20772 7837
rect 17868 7760 17920 7812
rect 18604 7692 18656 7744
rect 20260 7760 20312 7812
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 21916 7871 21968 7880
rect 21916 7837 21925 7871
rect 21925 7837 21959 7871
rect 21959 7837 21968 7871
rect 21916 7828 21968 7837
rect 23388 7871 23440 7880
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 23756 7828 23808 7880
rect 24032 7871 24084 7880
rect 24032 7837 24041 7871
rect 24041 7837 24075 7871
rect 24075 7837 24084 7871
rect 24032 7828 24084 7837
rect 24492 7828 24544 7880
rect 24952 7896 25004 7948
rect 25044 7939 25096 7948
rect 25044 7905 25053 7939
rect 25053 7905 25087 7939
rect 25087 7905 25096 7939
rect 25044 7896 25096 7905
rect 25504 8007 25556 8016
rect 25504 7973 25513 8007
rect 25513 7973 25547 8007
rect 25547 7973 25556 8007
rect 25504 7964 25556 7973
rect 26884 7964 26936 8016
rect 30748 8032 30800 8084
rect 31576 8032 31628 8084
rect 32128 8032 32180 8084
rect 33968 8032 34020 8084
rect 34428 8032 34480 8084
rect 36176 8032 36228 8084
rect 36820 8075 36872 8084
rect 36820 8041 36829 8075
rect 36829 8041 36863 8075
rect 36863 8041 36872 8075
rect 36820 8032 36872 8041
rect 37648 8075 37700 8084
rect 37648 8041 37657 8075
rect 37657 8041 37691 8075
rect 37691 8041 37700 8075
rect 37648 8032 37700 8041
rect 38292 8075 38344 8084
rect 38292 8041 38301 8075
rect 38301 8041 38335 8075
rect 38335 8041 38344 8075
rect 38292 8032 38344 8041
rect 28172 8007 28224 8016
rect 28172 7973 28181 8007
rect 28181 7973 28215 8007
rect 28215 7973 28224 8007
rect 28172 7964 28224 7973
rect 25412 7896 25464 7948
rect 27344 7896 27396 7948
rect 29092 7896 29144 7948
rect 30288 7896 30340 7948
rect 31300 7939 31352 7948
rect 31300 7905 31309 7939
rect 31309 7905 31343 7939
rect 31343 7905 31352 7939
rect 31300 7896 31352 7905
rect 31760 7939 31812 7948
rect 31760 7905 31769 7939
rect 31769 7905 31803 7939
rect 31803 7905 31812 7939
rect 31760 7896 31812 7905
rect 34152 7964 34204 8016
rect 35808 7964 35860 8016
rect 38384 7964 38436 8016
rect 32312 7939 32364 7948
rect 32312 7905 32321 7939
rect 32321 7905 32355 7939
rect 32355 7905 32364 7939
rect 32312 7896 32364 7905
rect 23112 7760 23164 7812
rect 25780 7871 25832 7880
rect 25780 7837 25789 7871
rect 25789 7837 25823 7871
rect 25823 7837 25832 7871
rect 25780 7828 25832 7837
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 27436 7871 27488 7880
rect 27436 7837 27445 7871
rect 27445 7837 27479 7871
rect 27479 7837 27488 7871
rect 27436 7828 27488 7837
rect 27896 7828 27948 7880
rect 28448 7871 28500 7880
rect 28448 7837 28457 7871
rect 28457 7837 28491 7871
rect 28491 7837 28500 7871
rect 28448 7828 28500 7837
rect 28540 7871 28592 7880
rect 28540 7837 28574 7871
rect 28574 7837 28592 7871
rect 28540 7828 28592 7837
rect 28724 7871 28776 7880
rect 28724 7837 28733 7871
rect 28733 7837 28767 7871
rect 28767 7837 28776 7871
rect 28724 7828 28776 7837
rect 30104 7828 30156 7880
rect 31116 7871 31168 7880
rect 31116 7837 31125 7871
rect 31125 7837 31159 7871
rect 31159 7837 31168 7871
rect 31116 7828 31168 7837
rect 32036 7871 32088 7880
rect 32036 7837 32045 7871
rect 32045 7837 32079 7871
rect 32079 7837 32088 7871
rect 32036 7828 32088 7837
rect 33968 7828 34020 7880
rect 34796 7828 34848 7880
rect 35716 7871 35768 7880
rect 35716 7837 35725 7871
rect 35725 7837 35759 7871
rect 35759 7837 35768 7871
rect 35716 7828 35768 7837
rect 36268 7828 36320 7880
rect 22192 7692 22244 7744
rect 22652 7735 22704 7744
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 23296 7692 23348 7744
rect 24124 7692 24176 7744
rect 24216 7735 24268 7744
rect 24216 7701 24225 7735
rect 24225 7701 24259 7735
rect 24259 7701 24268 7735
rect 24216 7692 24268 7701
rect 25596 7692 25648 7744
rect 25964 7692 26016 7744
rect 26608 7692 26660 7744
rect 29920 7692 29972 7744
rect 31760 7692 31812 7744
rect 32772 7692 32824 7744
rect 33508 7692 33560 7744
rect 34888 7692 34940 7744
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 37832 7896 37884 7948
rect 38660 7939 38712 7948
rect 38660 7905 38669 7939
rect 38669 7905 38703 7939
rect 38703 7905 38712 7939
rect 38660 7896 38712 7905
rect 37832 7760 37884 7812
rect 37280 7692 37332 7744
rect 38936 7692 38988 7744
rect 39396 7735 39448 7744
rect 39396 7701 39405 7735
rect 39405 7701 39439 7735
rect 39439 7701 39448 7735
rect 39396 7692 39448 7701
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 9010 7590 9062 7642
rect 9074 7590 9126 7642
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 15010 7590 15062 7642
rect 15074 7590 15126 7642
rect 15138 7590 15190 7642
rect 15202 7590 15254 7642
rect 15266 7590 15318 7642
rect 21010 7590 21062 7642
rect 21074 7590 21126 7642
rect 21138 7590 21190 7642
rect 21202 7590 21254 7642
rect 21266 7590 21318 7642
rect 27010 7590 27062 7642
rect 27074 7590 27126 7642
rect 27138 7590 27190 7642
rect 27202 7590 27254 7642
rect 27266 7590 27318 7642
rect 33010 7590 33062 7642
rect 33074 7590 33126 7642
rect 33138 7590 33190 7642
rect 33202 7590 33254 7642
rect 33266 7590 33318 7642
rect 39010 7590 39062 7642
rect 39074 7590 39126 7642
rect 39138 7590 39190 7642
rect 39202 7590 39254 7642
rect 39266 7590 39318 7642
rect 9772 7488 9824 7540
rect 9956 7531 10008 7540
rect 9956 7497 9965 7531
rect 9965 7497 9999 7531
rect 9999 7497 10008 7531
rect 9956 7488 10008 7497
rect 11060 7488 11112 7540
rect 11796 7488 11848 7540
rect 11980 7488 12032 7540
rect 756 7420 808 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 1584 7284 1636 7336
rect 1768 7284 1820 7336
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 4896 7420 4948 7472
rect 5816 7463 5868 7472
rect 5816 7429 5825 7463
rect 5825 7429 5859 7463
rect 5859 7429 5868 7463
rect 5816 7420 5868 7429
rect 7380 7420 7432 7472
rect 4252 7352 4304 7404
rect 4620 7352 4672 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 4344 7284 4396 7336
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 7472 7327 7524 7336
rect 7472 7293 7481 7327
rect 7481 7293 7515 7327
rect 7515 7293 7524 7327
rect 7472 7284 7524 7293
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 12348 7420 12400 7472
rect 13084 7488 13136 7540
rect 14464 7488 14516 7540
rect 14740 7488 14792 7540
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 16028 7488 16080 7540
rect 17960 7488 18012 7540
rect 18052 7488 18104 7540
rect 10048 7352 10100 7404
rect 4528 7216 4580 7268
rect 1124 7148 1176 7200
rect 2964 7148 3016 7200
rect 4344 7148 4396 7200
rect 4436 7148 4488 7200
rect 5080 7148 5132 7200
rect 6552 7148 6604 7200
rect 9588 7284 9640 7336
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 16120 7352 16172 7404
rect 17224 7352 17276 7404
rect 17592 7420 17644 7472
rect 19800 7531 19852 7540
rect 19800 7497 19809 7531
rect 19809 7497 19843 7531
rect 19843 7497 19852 7531
rect 19800 7488 19852 7497
rect 19892 7488 19944 7540
rect 20168 7420 20220 7472
rect 21916 7488 21968 7540
rect 24032 7488 24084 7540
rect 24124 7488 24176 7540
rect 17408 7352 17460 7404
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 11060 7284 11112 7336
rect 10416 7148 10468 7200
rect 10968 7148 11020 7200
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 14464 7284 14516 7336
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 14924 7327 14976 7336
rect 14924 7293 14958 7327
rect 14958 7293 14976 7327
rect 14924 7284 14976 7293
rect 15292 7284 15344 7336
rect 16028 7284 16080 7336
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 18236 7284 18288 7336
rect 18604 7327 18656 7336
rect 18604 7293 18613 7327
rect 18613 7293 18647 7327
rect 18647 7293 18656 7327
rect 18604 7284 18656 7293
rect 19064 7284 19116 7336
rect 20168 7284 20220 7336
rect 20444 7352 20496 7404
rect 23296 7420 23348 7472
rect 25136 7488 25188 7540
rect 25964 7488 26016 7540
rect 26056 7488 26108 7540
rect 26792 7488 26844 7540
rect 28080 7488 28132 7540
rect 28724 7488 28776 7540
rect 28816 7488 28868 7540
rect 30104 7531 30156 7540
rect 30104 7497 30113 7531
rect 30113 7497 30147 7531
rect 30147 7497 30156 7531
rect 30104 7488 30156 7497
rect 33048 7488 33100 7540
rect 33416 7488 33468 7540
rect 20628 7352 20680 7404
rect 25136 7352 25188 7404
rect 25872 7352 25924 7404
rect 26884 7352 26936 7404
rect 27436 7395 27488 7404
rect 27436 7361 27445 7395
rect 27445 7361 27479 7395
rect 27479 7361 27488 7395
rect 27436 7352 27488 7361
rect 27712 7352 27764 7404
rect 27896 7352 27948 7404
rect 28264 7395 28316 7404
rect 28264 7361 28273 7395
rect 28273 7361 28307 7395
rect 28307 7361 28316 7395
rect 28264 7352 28316 7361
rect 30380 7420 30432 7472
rect 28632 7352 28684 7404
rect 29460 7395 29512 7404
rect 29460 7361 29469 7395
rect 29469 7361 29503 7395
rect 29503 7361 29512 7395
rect 29460 7352 29512 7361
rect 30656 7395 30708 7404
rect 30656 7361 30665 7395
rect 30665 7361 30699 7395
rect 30699 7361 30708 7395
rect 30656 7352 30708 7361
rect 31024 7420 31076 7472
rect 31116 7420 31168 7472
rect 33968 7531 34020 7540
rect 33968 7497 33977 7531
rect 33977 7497 34011 7531
rect 34011 7497 34020 7531
rect 33968 7488 34020 7497
rect 34244 7488 34296 7540
rect 37280 7488 37332 7540
rect 37372 7488 37424 7540
rect 38752 7488 38804 7540
rect 31300 7352 31352 7404
rect 34336 7420 34388 7472
rect 21272 7284 21324 7336
rect 21548 7284 21600 7336
rect 22192 7284 22244 7336
rect 23480 7284 23532 7336
rect 24124 7284 24176 7336
rect 24308 7327 24360 7336
rect 24308 7293 24317 7327
rect 24317 7293 24351 7327
rect 24351 7293 24360 7327
rect 24308 7284 24360 7293
rect 14648 7216 14700 7268
rect 15936 7216 15988 7268
rect 16764 7216 16816 7268
rect 12900 7148 12952 7200
rect 13176 7148 13228 7200
rect 15108 7148 15160 7200
rect 16028 7191 16080 7200
rect 16028 7157 16037 7191
rect 16037 7157 16071 7191
rect 16071 7157 16080 7191
rect 16028 7148 16080 7157
rect 16396 7148 16448 7200
rect 18512 7148 18564 7200
rect 21180 7216 21232 7268
rect 22100 7216 22152 7268
rect 21272 7148 21324 7200
rect 24952 7284 25004 7336
rect 29184 7327 29236 7336
rect 24860 7216 24912 7268
rect 26332 7216 26384 7268
rect 27160 7216 27212 7268
rect 29184 7293 29193 7327
rect 29193 7293 29227 7327
rect 29227 7293 29236 7327
rect 29184 7284 29236 7293
rect 29276 7327 29328 7336
rect 29276 7293 29310 7327
rect 29310 7293 29328 7327
rect 29276 7284 29328 7293
rect 28908 7259 28960 7268
rect 28908 7225 28917 7259
rect 28917 7225 28951 7259
rect 28951 7225 28960 7259
rect 28908 7216 28960 7225
rect 30748 7216 30800 7268
rect 32404 7284 32456 7336
rect 33048 7395 33100 7404
rect 33048 7361 33057 7395
rect 33057 7361 33091 7395
rect 33091 7361 33100 7395
rect 33048 7352 33100 7361
rect 33968 7352 34020 7404
rect 34612 7352 34664 7404
rect 34980 7352 35032 7404
rect 33508 7284 33560 7336
rect 35440 7395 35492 7404
rect 35440 7361 35449 7395
rect 35449 7361 35483 7395
rect 35483 7361 35492 7395
rect 35440 7352 35492 7361
rect 36544 7352 36596 7404
rect 38476 7395 38528 7404
rect 38476 7361 38485 7395
rect 38485 7361 38519 7395
rect 38519 7361 38528 7395
rect 38476 7352 38528 7361
rect 38660 7352 38712 7404
rect 35716 7284 35768 7336
rect 31852 7216 31904 7268
rect 32036 7216 32088 7268
rect 32496 7216 32548 7268
rect 28632 7148 28684 7200
rect 30564 7148 30616 7200
rect 31576 7148 31628 7200
rect 35256 7259 35308 7268
rect 35256 7225 35265 7259
rect 35265 7225 35299 7259
rect 35299 7225 35308 7259
rect 35256 7216 35308 7225
rect 35348 7216 35400 7268
rect 36728 7216 36780 7268
rect 40040 7216 40092 7268
rect 39396 7191 39448 7200
rect 39396 7157 39405 7191
rect 39405 7157 39439 7191
rect 39439 7157 39448 7191
rect 39396 7148 39448 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 13950 7046 14002 7098
rect 14014 7046 14066 7098
rect 14078 7046 14130 7098
rect 14142 7046 14194 7098
rect 14206 7046 14258 7098
rect 19950 7046 20002 7098
rect 20014 7046 20066 7098
rect 20078 7046 20130 7098
rect 20142 7046 20194 7098
rect 20206 7046 20258 7098
rect 25950 7046 26002 7098
rect 26014 7046 26066 7098
rect 26078 7046 26130 7098
rect 26142 7046 26194 7098
rect 26206 7046 26258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 37950 7046 38002 7098
rect 38014 7046 38066 7098
rect 38078 7046 38130 7098
rect 38142 7046 38194 7098
rect 38206 7046 38258 7098
rect 2044 6944 2096 6996
rect 2412 6944 2464 6996
rect 2688 6944 2740 6996
rect 4252 6944 4304 6996
rect 11060 6944 11112 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 13176 6944 13228 6996
rect 15016 6944 15068 6996
rect 15660 6944 15712 6996
rect 1492 6876 1544 6928
rect 4436 6919 4488 6928
rect 4436 6885 4445 6919
rect 4445 6885 4479 6919
rect 4479 6885 4488 6919
rect 4436 6876 4488 6885
rect 7380 6876 7432 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 3516 6808 3568 6860
rect 4344 6808 4396 6860
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 6368 6851 6420 6860
rect 6368 6817 6377 6851
rect 6377 6817 6411 6851
rect 6411 6817 6420 6851
rect 6368 6808 6420 6817
rect 6552 6851 6604 6860
rect 6552 6817 6570 6851
rect 6570 6817 6604 6851
rect 6552 6808 6604 6817
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 6920 6851 6972 6860
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 7564 6851 7616 6860
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 12716 6876 12768 6928
rect 2320 6740 2372 6792
rect 3700 6740 3752 6792
rect 1860 6672 1912 6724
rect 3240 6672 3292 6724
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 4896 6740 4948 6792
rect 2688 6604 2740 6656
rect 3700 6604 3752 6656
rect 5632 6647 5684 6656
rect 5632 6613 5641 6647
rect 5641 6613 5675 6647
rect 5675 6613 5684 6647
rect 5632 6604 5684 6613
rect 6552 6604 6604 6656
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 14188 6876 14240 6928
rect 16212 6944 16264 6996
rect 16580 6944 16632 6996
rect 19984 6944 20036 6996
rect 20076 6987 20128 6996
rect 20076 6953 20085 6987
rect 20085 6953 20119 6987
rect 20119 6953 20128 6987
rect 20076 6944 20128 6953
rect 20168 6944 20220 6996
rect 24124 6944 24176 6996
rect 17960 6876 18012 6928
rect 20536 6876 20588 6928
rect 8852 6740 8904 6792
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 10600 6715 10652 6724
rect 10600 6681 10609 6715
rect 10609 6681 10643 6715
rect 10643 6681 10652 6715
rect 10600 6672 10652 6681
rect 10692 6715 10744 6724
rect 10692 6681 10701 6715
rect 10701 6681 10735 6715
rect 10735 6681 10744 6715
rect 10692 6672 10744 6681
rect 10784 6672 10836 6724
rect 11612 6740 11664 6792
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 12992 6740 13044 6792
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 13452 6740 13504 6792
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13820 6740 13872 6792
rect 16580 6808 16632 6860
rect 16856 6808 16908 6860
rect 17868 6808 17920 6860
rect 20812 6808 20864 6860
rect 24584 6876 24636 6928
rect 26332 6876 26384 6928
rect 28908 6944 28960 6996
rect 30656 6944 30708 6996
rect 29276 6876 29328 6928
rect 21824 6808 21876 6860
rect 14924 6740 14976 6792
rect 15568 6740 15620 6792
rect 9864 6604 9916 6656
rect 9956 6604 10008 6656
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 10968 6604 11020 6656
rect 11520 6604 11572 6656
rect 11888 6604 11940 6656
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 13544 6647 13596 6656
rect 13544 6613 13553 6647
rect 13553 6613 13587 6647
rect 13587 6613 13596 6647
rect 13544 6604 13596 6613
rect 13728 6672 13780 6724
rect 16764 6740 16816 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 19064 6740 19116 6792
rect 19524 6740 19576 6792
rect 20352 6740 20404 6792
rect 20536 6740 20588 6792
rect 16304 6672 16356 6724
rect 14188 6604 14240 6656
rect 14832 6604 14884 6656
rect 15016 6604 15068 6656
rect 16948 6604 17000 6656
rect 19340 6672 19392 6724
rect 20168 6672 20220 6724
rect 21364 6783 21416 6792
rect 21364 6749 21373 6783
rect 21373 6749 21407 6783
rect 21407 6749 21416 6783
rect 21364 6740 21416 6749
rect 21456 6783 21508 6792
rect 21456 6749 21490 6783
rect 21490 6749 21508 6783
rect 21456 6740 21508 6749
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 23112 6672 23164 6724
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 24768 6740 24820 6792
rect 24860 6783 24912 6792
rect 24860 6749 24869 6783
rect 24869 6749 24903 6783
rect 24903 6749 24912 6783
rect 24860 6740 24912 6749
rect 25136 6740 25188 6792
rect 24032 6672 24084 6724
rect 24492 6672 24544 6724
rect 25872 6740 25924 6792
rect 25964 6783 26016 6792
rect 25964 6749 25973 6783
rect 25973 6749 26007 6783
rect 26007 6749 26016 6783
rect 25964 6740 26016 6749
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 27160 6808 27212 6860
rect 26516 6740 26568 6792
rect 26700 6740 26752 6792
rect 27344 6740 27396 6792
rect 28264 6808 28316 6860
rect 30196 6851 30248 6860
rect 30196 6817 30205 6851
rect 30205 6817 30239 6851
rect 30239 6817 30248 6851
rect 30196 6808 30248 6817
rect 31208 6876 31260 6928
rect 34612 6944 34664 6996
rect 37740 6944 37792 6996
rect 30564 6851 30616 6860
rect 30564 6817 30598 6851
rect 30598 6817 30616 6851
rect 30564 6808 30616 6817
rect 38568 6808 38620 6860
rect 27620 6740 27672 6792
rect 27712 6783 27764 6792
rect 27712 6749 27721 6783
rect 27721 6749 27755 6783
rect 27755 6749 27764 6783
rect 27712 6740 27764 6749
rect 22560 6647 22612 6656
rect 22560 6613 22569 6647
rect 22569 6613 22603 6647
rect 22603 6613 22612 6647
rect 22560 6604 22612 6613
rect 22744 6647 22796 6656
rect 22744 6613 22753 6647
rect 22753 6613 22787 6647
rect 22787 6613 22796 6647
rect 22744 6604 22796 6613
rect 23020 6604 23072 6656
rect 25412 6672 25464 6724
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 31668 6740 31720 6792
rect 32220 6783 32272 6792
rect 32220 6749 32229 6783
rect 32229 6749 32263 6783
rect 32263 6749 32272 6783
rect 32220 6740 32272 6749
rect 33416 6740 33468 6792
rect 34060 6740 34112 6792
rect 34244 6740 34296 6792
rect 34612 6740 34664 6792
rect 25872 6604 25924 6656
rect 27344 6647 27396 6656
rect 27344 6613 27353 6647
rect 27353 6613 27387 6647
rect 27387 6613 27396 6647
rect 27344 6604 27396 6613
rect 27436 6604 27488 6656
rect 28264 6604 28316 6656
rect 32864 6672 32916 6724
rect 32588 6604 32640 6656
rect 32772 6604 32824 6656
rect 33692 6604 33744 6656
rect 35072 6740 35124 6792
rect 37740 6740 37792 6792
rect 34796 6672 34848 6724
rect 35532 6672 35584 6724
rect 38476 6740 38528 6792
rect 35348 6604 35400 6656
rect 35716 6647 35768 6656
rect 35716 6613 35725 6647
rect 35725 6613 35759 6647
rect 35759 6613 35768 6647
rect 35716 6604 35768 6613
rect 35808 6647 35860 6656
rect 35808 6613 35817 6647
rect 35817 6613 35851 6647
rect 35851 6613 35860 6647
rect 35808 6604 35860 6613
rect 38752 6672 38804 6724
rect 38384 6604 38436 6656
rect 38568 6604 38620 6656
rect 39580 6672 39632 6724
rect 39396 6647 39448 6656
rect 39396 6613 39405 6647
rect 39405 6613 39439 6647
rect 39439 6613 39448 6647
rect 39396 6604 39448 6613
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 9010 6502 9062 6554
rect 9074 6502 9126 6554
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 15010 6502 15062 6554
rect 15074 6502 15126 6554
rect 15138 6502 15190 6554
rect 15202 6502 15254 6554
rect 15266 6502 15318 6554
rect 21010 6502 21062 6554
rect 21074 6502 21126 6554
rect 21138 6502 21190 6554
rect 21202 6502 21254 6554
rect 21266 6502 21318 6554
rect 27010 6502 27062 6554
rect 27074 6502 27126 6554
rect 27138 6502 27190 6554
rect 27202 6502 27254 6554
rect 27266 6502 27318 6554
rect 33010 6502 33062 6554
rect 33074 6502 33126 6554
rect 33138 6502 33190 6554
rect 33202 6502 33254 6554
rect 33266 6502 33318 6554
rect 39010 6502 39062 6554
rect 39074 6502 39126 6554
rect 39138 6502 39190 6554
rect 39202 6502 39254 6554
rect 39266 6502 39318 6554
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 7196 6400 7248 6452
rect 9128 6400 9180 6452
rect 9956 6400 10008 6452
rect 10692 6400 10744 6452
rect 11428 6400 11480 6452
rect 1216 6196 1268 6248
rect 2872 6307 2924 6316
rect 2872 6273 2881 6307
rect 2881 6273 2915 6307
rect 2915 6273 2924 6307
rect 2872 6264 2924 6273
rect 3608 6264 3660 6316
rect 6092 6332 6144 6384
rect 4068 6264 4120 6316
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 4804 6264 4856 6316
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 4436 6196 4488 6248
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 6644 6196 6696 6248
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7196 6264 7248 6316
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 10968 6332 11020 6384
rect 8576 6264 8628 6316
rect 9588 6264 9640 6316
rect 10324 6264 10376 6316
rect 10600 6264 10652 6316
rect 11428 6264 11480 6316
rect 6368 6128 6420 6180
rect 8760 6196 8812 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 3516 6060 3568 6112
rect 3976 6060 4028 6112
rect 6184 6060 6236 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8944 6128 8996 6180
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 9864 6196 9916 6248
rect 12256 6400 12308 6452
rect 12440 6400 12492 6452
rect 11980 6264 12032 6316
rect 12072 6264 12124 6316
rect 13728 6332 13780 6384
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 14372 6400 14424 6452
rect 15936 6400 15988 6452
rect 16120 6400 16172 6452
rect 15568 6307 15620 6316
rect 15568 6273 15577 6307
rect 15577 6273 15611 6307
rect 15611 6273 15620 6307
rect 15568 6264 15620 6273
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 16948 6400 17000 6452
rect 20996 6400 21048 6452
rect 21640 6400 21692 6452
rect 21916 6400 21968 6452
rect 23020 6400 23072 6452
rect 24860 6400 24912 6452
rect 25964 6400 26016 6452
rect 19984 6332 20036 6384
rect 21456 6332 21508 6384
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 18052 6264 18104 6316
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 10692 6128 10744 6180
rect 11060 6128 11112 6180
rect 12256 6128 12308 6180
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 14188 6196 14240 6248
rect 14372 6196 14424 6248
rect 14740 6196 14792 6248
rect 15200 6196 15252 6248
rect 16396 6196 16448 6248
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 18512 6196 18564 6248
rect 18880 6196 18932 6248
rect 19156 6239 19208 6248
rect 19156 6205 19190 6239
rect 19190 6205 19208 6239
rect 19156 6196 19208 6205
rect 19524 6196 19576 6248
rect 7840 6060 7892 6112
rect 9588 6060 9640 6112
rect 10048 6060 10100 6112
rect 10508 6060 10560 6112
rect 13176 6060 13228 6112
rect 14464 6060 14516 6112
rect 14740 6060 14792 6112
rect 14924 6128 14976 6180
rect 19892 6196 19944 6248
rect 20076 6239 20128 6248
rect 20076 6205 20085 6239
rect 20085 6205 20119 6239
rect 20119 6205 20128 6239
rect 20076 6196 20128 6205
rect 20720 6264 20772 6316
rect 21916 6239 21968 6248
rect 21916 6205 21925 6239
rect 21925 6205 21959 6239
rect 21959 6205 21968 6239
rect 21916 6196 21968 6205
rect 16580 6060 16632 6112
rect 17868 6060 17920 6112
rect 18144 6060 18196 6112
rect 19156 6060 19208 6112
rect 20720 6060 20772 6112
rect 21364 6060 21416 6112
rect 23020 6239 23072 6248
rect 23020 6205 23029 6239
rect 23029 6205 23063 6239
rect 23063 6205 23072 6239
rect 23020 6196 23072 6205
rect 24124 6171 24176 6180
rect 24124 6137 24133 6171
rect 24133 6137 24167 6171
rect 24167 6137 24176 6171
rect 24124 6128 24176 6137
rect 22928 6103 22980 6112
rect 22928 6069 22937 6103
rect 22937 6069 22971 6103
rect 22971 6069 22980 6103
rect 22928 6060 22980 6069
rect 23664 6060 23716 6112
rect 24308 6264 24360 6316
rect 24952 6264 25004 6316
rect 25504 6264 25556 6316
rect 26516 6332 26568 6384
rect 26700 6332 26752 6384
rect 27436 6332 27488 6384
rect 27804 6264 27856 6316
rect 28540 6332 28592 6384
rect 28080 6307 28132 6316
rect 28080 6273 28089 6307
rect 28089 6273 28123 6307
rect 28123 6273 28132 6307
rect 28080 6264 28132 6273
rect 28264 6264 28316 6316
rect 28448 6264 28500 6316
rect 26424 6196 26476 6248
rect 26516 6196 26568 6248
rect 25412 6128 25464 6180
rect 25596 6060 25648 6112
rect 27160 6128 27212 6180
rect 26884 6060 26936 6112
rect 26976 6103 27028 6112
rect 26976 6069 26985 6103
rect 26985 6069 27019 6103
rect 27019 6069 27028 6103
rect 26976 6060 27028 6069
rect 29184 6239 29236 6248
rect 29184 6205 29193 6239
rect 29193 6205 29227 6239
rect 29227 6205 29236 6239
rect 29184 6196 29236 6205
rect 29276 6196 29328 6248
rect 30288 6264 30340 6316
rect 30380 6307 30432 6316
rect 30380 6273 30389 6307
rect 30389 6273 30423 6307
rect 30423 6273 30432 6307
rect 30380 6264 30432 6273
rect 33416 6400 33468 6452
rect 35072 6400 35124 6452
rect 35440 6400 35492 6452
rect 35900 6400 35952 6452
rect 37556 6400 37608 6452
rect 39488 6400 39540 6452
rect 35716 6332 35768 6384
rect 32312 6307 32364 6316
rect 32312 6273 32321 6307
rect 32321 6273 32355 6307
rect 32355 6273 32364 6307
rect 32312 6264 32364 6273
rect 33416 6307 33468 6316
rect 33416 6273 33425 6307
rect 33425 6273 33459 6307
rect 33459 6273 33468 6307
rect 33416 6264 33468 6273
rect 34520 6264 34572 6316
rect 32404 6196 32456 6248
rect 30840 6128 30892 6180
rect 32772 6196 32824 6248
rect 29000 6060 29052 6112
rect 31116 6103 31168 6112
rect 31116 6069 31125 6103
rect 31125 6069 31159 6103
rect 31159 6069 31168 6103
rect 31116 6060 31168 6069
rect 32312 6060 32364 6112
rect 32588 6128 32640 6180
rect 33692 6239 33744 6248
rect 33692 6205 33701 6239
rect 33701 6205 33735 6239
rect 33735 6205 33744 6239
rect 33692 6196 33744 6205
rect 35440 6239 35492 6248
rect 35440 6205 35449 6239
rect 35449 6205 35483 6239
rect 35483 6205 35492 6239
rect 35440 6196 35492 6205
rect 34244 6060 34296 6112
rect 37372 6264 37424 6316
rect 38752 6307 38804 6316
rect 38752 6273 38761 6307
rect 38761 6273 38795 6307
rect 38795 6273 38804 6307
rect 38752 6264 38804 6273
rect 36176 6196 36228 6248
rect 39212 6307 39264 6316
rect 39212 6273 39221 6307
rect 39221 6273 39255 6307
rect 39255 6273 39264 6307
rect 39212 6264 39264 6273
rect 37096 6128 37148 6180
rect 39028 6103 39080 6112
rect 39028 6069 39037 6103
rect 39037 6069 39071 6103
rect 39071 6069 39080 6103
rect 39028 6060 39080 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 13950 5958 14002 6010
rect 14014 5958 14066 6010
rect 14078 5958 14130 6010
rect 14142 5958 14194 6010
rect 14206 5958 14258 6010
rect 19950 5958 20002 6010
rect 20014 5958 20066 6010
rect 20078 5958 20130 6010
rect 20142 5958 20194 6010
rect 20206 5958 20258 6010
rect 25950 5958 26002 6010
rect 26014 5958 26066 6010
rect 26078 5958 26130 6010
rect 26142 5958 26194 6010
rect 26206 5958 26258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 37950 5958 38002 6010
rect 38014 5958 38066 6010
rect 38078 5958 38130 6010
rect 38142 5958 38194 6010
rect 38206 5958 38258 6010
rect 4068 5856 4120 5908
rect 4896 5856 4948 5908
rect 6092 5856 6144 5908
rect 7104 5856 7156 5908
rect 7196 5856 7248 5908
rect 8208 5856 8260 5908
rect 8668 5856 8720 5908
rect 1768 5788 1820 5840
rect 2504 5788 2556 5840
rect 2780 5831 2832 5840
rect 2780 5797 2789 5831
rect 2789 5797 2823 5831
rect 2823 5797 2832 5831
rect 2780 5788 2832 5797
rect 3148 5831 3200 5840
rect 3148 5797 3157 5831
rect 3157 5797 3191 5831
rect 3191 5797 3200 5831
rect 3148 5788 3200 5797
rect 2964 5720 3016 5772
rect 1400 5652 1452 5704
rect 3608 5720 3660 5772
rect 5908 5720 5960 5772
rect 8576 5788 8628 5840
rect 7472 5720 7524 5772
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 10508 5856 10560 5908
rect 11428 5899 11480 5908
rect 11428 5865 11437 5899
rect 11437 5865 11471 5899
rect 11471 5865 11480 5899
rect 11428 5856 11480 5865
rect 11796 5856 11848 5908
rect 10140 5788 10192 5840
rect 11244 5788 11296 5840
rect 11336 5788 11388 5840
rect 9404 5720 9456 5772
rect 1676 5584 1728 5636
rect 2228 5627 2280 5636
rect 2228 5593 2237 5627
rect 2237 5593 2271 5627
rect 2271 5593 2280 5627
rect 2228 5584 2280 5593
rect 2688 5584 2740 5636
rect 2964 5627 3016 5636
rect 2596 5516 2648 5568
rect 2964 5593 2973 5627
rect 2973 5593 3007 5627
rect 3007 5593 3016 5627
rect 2964 5584 3016 5593
rect 4988 5695 5040 5704
rect 4988 5661 4997 5695
rect 4997 5661 5031 5695
rect 5031 5661 5040 5695
rect 4988 5652 5040 5661
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5632 5652 5684 5704
rect 9680 5720 9732 5772
rect 9956 5720 10008 5772
rect 10508 5763 10560 5772
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 11796 5720 11848 5772
rect 11888 5720 11940 5772
rect 13084 5720 13136 5772
rect 13360 5720 13412 5772
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 8484 5652 8536 5704
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 8852 5652 8904 5704
rect 9496 5652 9548 5704
rect 2872 5516 2924 5568
rect 5908 5584 5960 5636
rect 4068 5516 4120 5568
rect 5080 5516 5132 5568
rect 5540 5516 5592 5568
rect 6552 5516 6604 5568
rect 7288 5516 7340 5568
rect 8392 5516 8444 5568
rect 8668 5516 8720 5568
rect 9496 5516 9548 5568
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11336 5584 11388 5636
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 12532 5695 12584 5704
rect 12532 5661 12566 5695
rect 12566 5661 12584 5695
rect 12532 5652 12584 5661
rect 10140 5516 10192 5568
rect 12440 5516 12492 5568
rect 14464 5788 14516 5840
rect 14832 5788 14884 5840
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 15016 5763 15068 5772
rect 15016 5729 15025 5763
rect 15025 5729 15059 5763
rect 15059 5729 15068 5763
rect 15016 5720 15068 5729
rect 15200 5720 15252 5772
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 14280 5584 14332 5636
rect 16212 5856 16264 5908
rect 16764 5856 16816 5908
rect 17868 5831 17920 5840
rect 17868 5797 17877 5831
rect 17877 5797 17911 5831
rect 17911 5797 17920 5831
rect 17868 5788 17920 5797
rect 19064 5899 19116 5908
rect 19064 5865 19073 5899
rect 19073 5865 19107 5899
rect 19107 5865 19116 5899
rect 19064 5856 19116 5865
rect 19340 5856 19392 5908
rect 20536 5856 20588 5908
rect 20812 5856 20864 5908
rect 20904 5788 20956 5840
rect 19708 5720 19760 5772
rect 20996 5720 21048 5772
rect 22192 5788 22244 5840
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16304 5652 16356 5704
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 18144 5695 18196 5704
rect 18144 5661 18153 5695
rect 18153 5661 18187 5695
rect 18187 5661 18196 5695
rect 18144 5652 18196 5661
rect 18236 5695 18288 5704
rect 18236 5661 18270 5695
rect 18270 5661 18288 5695
rect 18236 5652 18288 5661
rect 19248 5695 19300 5704
rect 19248 5661 19257 5695
rect 19257 5661 19291 5695
rect 19291 5661 19300 5695
rect 19248 5652 19300 5661
rect 14740 5516 14792 5568
rect 14832 5516 14884 5568
rect 15292 5516 15344 5568
rect 15568 5516 15620 5568
rect 19616 5584 19668 5636
rect 20076 5584 20128 5636
rect 20444 5652 20496 5704
rect 21180 5584 21232 5636
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 21548 5652 21600 5704
rect 22376 5788 22428 5840
rect 22928 5788 22980 5840
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 23572 5763 23624 5772
rect 23572 5729 23579 5763
rect 23579 5729 23613 5763
rect 23613 5729 23624 5763
rect 23572 5720 23624 5729
rect 26516 5788 26568 5840
rect 26976 5856 27028 5908
rect 27160 5856 27212 5908
rect 27620 5788 27672 5840
rect 30380 5856 30432 5908
rect 30748 5856 30800 5908
rect 34704 5856 34756 5908
rect 35072 5856 35124 5908
rect 35164 5856 35216 5908
rect 39396 5899 39448 5908
rect 39396 5865 39405 5899
rect 39405 5865 39439 5899
rect 39439 5865 39448 5899
rect 39396 5856 39448 5865
rect 29460 5788 29512 5840
rect 26148 5763 26200 5772
rect 26148 5729 26157 5763
rect 26157 5729 26191 5763
rect 26191 5729 26200 5763
rect 26148 5720 26200 5729
rect 23480 5652 23532 5704
rect 25044 5652 25096 5704
rect 25596 5695 25648 5704
rect 25596 5661 25605 5695
rect 25605 5661 25639 5695
rect 25639 5661 25648 5695
rect 25596 5652 25648 5661
rect 26700 5720 26752 5772
rect 27068 5720 27120 5772
rect 27344 5720 27396 5772
rect 27896 5763 27948 5772
rect 27896 5729 27905 5763
rect 27905 5729 27939 5763
rect 27939 5729 27948 5763
rect 27896 5720 27948 5729
rect 32864 5788 32916 5840
rect 33876 5788 33928 5840
rect 35716 5788 35768 5840
rect 38936 5788 38988 5840
rect 39948 5788 40000 5840
rect 32496 5720 32548 5772
rect 32680 5720 32732 5772
rect 38476 5720 38528 5772
rect 22284 5584 22336 5636
rect 18972 5516 19024 5568
rect 20904 5516 20956 5568
rect 25136 5584 25188 5636
rect 25228 5584 25280 5636
rect 28080 5652 28132 5704
rect 24584 5559 24636 5568
rect 24584 5525 24593 5559
rect 24593 5525 24627 5559
rect 24627 5525 24636 5559
rect 24584 5516 24636 5525
rect 24676 5516 24728 5568
rect 26424 5516 26476 5568
rect 26792 5516 26844 5568
rect 29092 5627 29144 5636
rect 29092 5593 29101 5627
rect 29101 5593 29135 5627
rect 29135 5593 29144 5627
rect 29092 5584 29144 5593
rect 29828 5695 29880 5704
rect 29828 5661 29837 5695
rect 29837 5661 29871 5695
rect 29871 5661 29880 5695
rect 29828 5652 29880 5661
rect 30472 5652 30524 5704
rect 30840 5652 30892 5704
rect 31024 5652 31076 5704
rect 32220 5652 32272 5704
rect 32772 5652 32824 5704
rect 33416 5652 33468 5704
rect 35072 5652 35124 5704
rect 37556 5652 37608 5704
rect 27712 5516 27764 5568
rect 28448 5516 28500 5568
rect 28540 5516 28592 5568
rect 28908 5516 28960 5568
rect 29460 5516 29512 5568
rect 32128 5516 32180 5568
rect 34060 5516 34112 5568
rect 34520 5627 34572 5636
rect 34520 5593 34529 5627
rect 34529 5593 34563 5627
rect 34563 5593 34572 5627
rect 34520 5584 34572 5593
rect 36084 5584 36136 5636
rect 34980 5516 35032 5568
rect 35900 5516 35952 5568
rect 36452 5516 36504 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 9010 5414 9062 5466
rect 9074 5414 9126 5466
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 15010 5414 15062 5466
rect 15074 5414 15126 5466
rect 15138 5414 15190 5466
rect 15202 5414 15254 5466
rect 15266 5414 15318 5466
rect 21010 5414 21062 5466
rect 21074 5414 21126 5466
rect 21138 5414 21190 5466
rect 21202 5414 21254 5466
rect 21266 5414 21318 5466
rect 27010 5414 27062 5466
rect 27074 5414 27126 5466
rect 27138 5414 27190 5466
rect 27202 5414 27254 5466
rect 27266 5414 27318 5466
rect 33010 5414 33062 5466
rect 33074 5414 33126 5466
rect 33138 5414 33190 5466
rect 33202 5414 33254 5466
rect 33266 5414 33318 5466
rect 39010 5414 39062 5466
rect 39074 5414 39126 5466
rect 39138 5414 39190 5466
rect 39202 5414 39254 5466
rect 39266 5414 39318 5466
rect 1400 5312 1452 5364
rect 1952 5355 2004 5364
rect 1952 5321 1961 5355
rect 1961 5321 1995 5355
rect 1995 5321 2004 5355
rect 1952 5312 2004 5321
rect 3424 5355 3476 5364
rect 3424 5321 3433 5355
rect 3433 5321 3467 5355
rect 3467 5321 3476 5355
rect 3424 5312 3476 5321
rect 3884 5312 3936 5364
rect 4804 5312 4856 5364
rect 6092 5312 6144 5364
rect 7564 5312 7616 5364
rect 7748 5312 7800 5364
rect 1492 5287 1544 5296
rect 1492 5253 1501 5287
rect 1501 5253 1535 5287
rect 1535 5253 1544 5287
rect 1492 5244 1544 5253
rect 1676 5287 1728 5296
rect 1676 5253 1685 5287
rect 1685 5253 1719 5287
rect 1719 5253 1728 5287
rect 1676 5244 1728 5253
rect 1860 5287 1912 5296
rect 1860 5253 1869 5287
rect 1869 5253 1903 5287
rect 1903 5253 1912 5287
rect 1860 5244 1912 5253
rect 1584 5176 1636 5228
rect 2320 5244 2372 5296
rect 2412 5176 2464 5228
rect 2596 5176 2648 5228
rect 2872 5176 2924 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 3608 5176 3660 5228
rect 1860 5108 1912 5160
rect 4344 5176 4396 5228
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 4804 5176 4856 5228
rect 5080 5244 5132 5296
rect 6000 5244 6052 5296
rect 6920 5244 6972 5296
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 5724 5176 5776 5228
rect 6184 5176 6236 5228
rect 6552 5176 6604 5228
rect 6736 5176 6788 5228
rect 7196 5176 7248 5228
rect 8392 5219 8444 5228
rect 8392 5185 8426 5219
rect 8426 5185 8444 5219
rect 8392 5176 8444 5185
rect 9404 5312 9456 5364
rect 9312 5244 9364 5296
rect 11520 5312 11572 5364
rect 11704 5312 11756 5364
rect 5080 5108 5132 5160
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 2412 5083 2464 5092
rect 2412 5049 2421 5083
rect 2421 5049 2455 5083
rect 2455 5049 2464 5083
rect 2412 5040 2464 5049
rect 2320 4972 2372 5024
rect 2964 4972 3016 5024
rect 4160 5040 4212 5092
rect 4344 5015 4396 5024
rect 4344 4981 4353 5015
rect 4353 4981 4387 5015
rect 4387 4981 4396 5015
rect 4344 4972 4396 4981
rect 6092 5108 6144 5160
rect 7472 5108 7524 5160
rect 7748 5108 7800 5160
rect 7932 5108 7984 5160
rect 8116 5108 8168 5160
rect 8944 5108 8996 5160
rect 9128 5108 9180 5160
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 9496 5151 9548 5160
rect 9496 5117 9505 5151
rect 9505 5117 9539 5151
rect 9539 5117 9548 5151
rect 9496 5108 9548 5117
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10416 5108 10468 5160
rect 10692 5108 10744 5160
rect 11888 5176 11940 5228
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 12440 5312 12492 5364
rect 12624 5355 12676 5364
rect 12624 5321 12633 5355
rect 12633 5321 12667 5355
rect 12667 5321 12676 5355
rect 12624 5312 12676 5321
rect 12808 5312 12860 5364
rect 14924 5312 14976 5364
rect 15200 5312 15252 5364
rect 21456 5312 21508 5364
rect 22652 5312 22704 5364
rect 23756 5312 23808 5364
rect 24124 5312 24176 5364
rect 25228 5312 25280 5364
rect 25320 5312 25372 5364
rect 26516 5312 26568 5364
rect 26608 5312 26660 5364
rect 27436 5312 27488 5364
rect 12716 5176 12768 5228
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 13084 5176 13136 5228
rect 4896 4972 4948 5024
rect 5172 4972 5224 5024
rect 7012 5083 7064 5092
rect 7012 5049 7021 5083
rect 7021 5049 7055 5083
rect 7055 5049 7064 5083
rect 7012 5040 7064 5049
rect 7104 5040 7156 5092
rect 9956 5083 10008 5092
rect 5448 4972 5500 5024
rect 6276 4972 6328 5024
rect 7656 4972 7708 5024
rect 9956 5049 9965 5083
rect 9965 5049 9999 5083
rect 9999 5049 10008 5083
rect 9956 5040 10008 5049
rect 9036 4972 9088 5024
rect 9588 4972 9640 5024
rect 12624 5108 12676 5160
rect 12992 5108 13044 5160
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 15752 5176 15804 5228
rect 16212 5176 16264 5228
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 16948 5176 17000 5228
rect 18236 5176 18288 5228
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 18880 5219 18932 5228
rect 18880 5185 18914 5219
rect 18914 5185 18932 5219
rect 18880 5176 18932 5185
rect 19892 5176 19944 5228
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 22468 5219 22520 5228
rect 22468 5185 22477 5219
rect 22477 5185 22511 5219
rect 22511 5185 22520 5219
rect 22468 5176 22520 5185
rect 13360 5108 13412 5160
rect 14372 5108 14424 5160
rect 11060 5040 11112 5092
rect 10968 4972 11020 5024
rect 11796 4972 11848 5024
rect 13268 5040 13320 5092
rect 15292 5040 15344 5092
rect 12532 4972 12584 5024
rect 14096 4972 14148 5024
rect 14924 4972 14976 5024
rect 15108 4972 15160 5024
rect 16396 5108 16448 5160
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 18420 5108 18472 5160
rect 19248 5108 19300 5160
rect 16304 4972 16356 5024
rect 17868 4972 17920 5024
rect 18236 4972 18288 5024
rect 22928 5176 22980 5228
rect 24308 5176 24360 5228
rect 24860 5176 24912 5228
rect 22744 5151 22796 5160
rect 22744 5117 22753 5151
rect 22753 5117 22787 5151
rect 22787 5117 22796 5151
rect 22744 5108 22796 5117
rect 23388 5108 23440 5160
rect 24032 5108 24084 5160
rect 25412 5176 25464 5228
rect 26792 5219 26844 5228
rect 26792 5185 26801 5219
rect 26801 5185 26835 5219
rect 26835 5185 26844 5219
rect 26792 5176 26844 5185
rect 25044 5151 25096 5160
rect 25044 5117 25053 5151
rect 25053 5117 25087 5151
rect 25087 5117 25096 5151
rect 25044 5108 25096 5117
rect 27436 5176 27488 5228
rect 27620 5176 27672 5228
rect 27896 5312 27948 5364
rect 29092 5312 29144 5364
rect 29644 5312 29696 5364
rect 30196 5312 30248 5364
rect 28080 5249 28132 5296
rect 28080 5244 28089 5249
rect 28089 5244 28123 5249
rect 28123 5244 28132 5249
rect 28172 5244 28224 5296
rect 27712 5108 27764 5160
rect 20444 5083 20496 5092
rect 20444 5049 20453 5083
rect 20453 5049 20487 5083
rect 20487 5049 20496 5083
rect 20444 5040 20496 5049
rect 21548 5040 21600 5092
rect 22652 5040 22704 5092
rect 28448 5176 28500 5228
rect 29092 5176 29144 5228
rect 29276 5176 29328 5228
rect 28908 5151 28960 5160
rect 28908 5117 28917 5151
rect 28917 5117 28951 5151
rect 28951 5117 28960 5151
rect 28908 5108 28960 5117
rect 32680 5312 32732 5364
rect 32956 5312 33008 5364
rect 33508 5312 33560 5364
rect 34612 5355 34664 5364
rect 34612 5321 34621 5355
rect 34621 5321 34655 5355
rect 34655 5321 34664 5355
rect 34612 5312 34664 5321
rect 36176 5355 36228 5364
rect 36176 5321 36185 5355
rect 36185 5321 36219 5355
rect 36219 5321 36228 5355
rect 36176 5312 36228 5321
rect 39396 5355 39448 5364
rect 39396 5321 39405 5355
rect 39405 5321 39439 5355
rect 39439 5321 39448 5355
rect 39396 5312 39448 5321
rect 33048 5244 33100 5296
rect 34336 5244 34388 5296
rect 35900 5287 35952 5296
rect 35900 5253 35909 5287
rect 35909 5253 35943 5287
rect 35943 5253 35952 5287
rect 35900 5244 35952 5253
rect 31392 5176 31444 5228
rect 31668 5176 31720 5228
rect 32220 5176 32272 5228
rect 20076 4972 20128 5024
rect 20536 4972 20588 5024
rect 20720 4972 20772 5024
rect 22192 4972 22244 5024
rect 23756 5015 23808 5024
rect 23756 4981 23765 5015
rect 23765 4981 23799 5015
rect 23799 4981 23808 5015
rect 23756 4972 23808 4981
rect 23940 4972 23992 5024
rect 24492 4972 24544 5024
rect 24768 5015 24820 5024
rect 24768 4981 24777 5015
rect 24777 4981 24811 5015
rect 24811 4981 24820 5015
rect 24768 4972 24820 4981
rect 24952 4972 25004 5024
rect 30012 5040 30064 5092
rect 25872 4972 25924 5024
rect 26424 4972 26476 5024
rect 26884 4972 26936 5024
rect 27344 4972 27396 5024
rect 28172 4972 28224 5024
rect 29552 4972 29604 5024
rect 30380 5015 30432 5024
rect 30380 4981 30389 5015
rect 30389 4981 30423 5015
rect 30423 4981 30432 5015
rect 30380 4972 30432 4981
rect 30564 5040 30616 5092
rect 31668 5083 31720 5092
rect 31668 5049 31677 5083
rect 31677 5049 31711 5083
rect 31711 5049 31720 5083
rect 31668 5040 31720 5049
rect 32312 5108 32364 5160
rect 34060 5219 34112 5228
rect 34060 5185 34069 5219
rect 34069 5185 34103 5219
rect 34103 5185 34112 5219
rect 34060 5176 34112 5185
rect 34796 5176 34848 5228
rect 38844 5219 38896 5228
rect 38844 5185 38853 5219
rect 38853 5185 38887 5219
rect 38887 5185 38896 5219
rect 38844 5176 38896 5185
rect 38936 5176 38988 5228
rect 36636 5108 36688 5160
rect 31392 4972 31444 5024
rect 32220 4972 32272 5024
rect 32588 5015 32640 5024
rect 32588 4981 32597 5015
rect 32597 4981 32631 5015
rect 32631 4981 32640 5015
rect 32588 4972 32640 4981
rect 32956 4972 33008 5024
rect 35348 4972 35400 5024
rect 39028 5015 39080 5024
rect 39028 4981 39037 5015
rect 39037 4981 39071 5015
rect 39071 4981 39080 5015
rect 39028 4972 39080 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 13950 4870 14002 4922
rect 14014 4870 14066 4922
rect 14078 4870 14130 4922
rect 14142 4870 14194 4922
rect 14206 4870 14258 4922
rect 19950 4870 20002 4922
rect 20014 4870 20066 4922
rect 20078 4870 20130 4922
rect 20142 4870 20194 4922
rect 20206 4870 20258 4922
rect 25950 4870 26002 4922
rect 26014 4870 26066 4922
rect 26078 4870 26130 4922
rect 26142 4870 26194 4922
rect 26206 4870 26258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 37950 4870 38002 4922
rect 38014 4870 38066 4922
rect 38078 4870 38130 4922
rect 38142 4870 38194 4922
rect 38206 4870 38258 4922
rect 1860 4768 1912 4820
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 3884 4768 3936 4820
rect 4344 4768 4396 4820
rect 3240 4700 3292 4752
rect 3700 4700 3752 4752
rect 1676 4632 1728 4684
rect 3608 4632 3660 4684
rect 3884 4632 3936 4684
rect 4528 4632 4580 4684
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 5080 4632 5132 4684
rect 7288 4768 7340 4820
rect 8208 4768 8260 4820
rect 9036 4768 9088 4820
rect 10324 4768 10376 4820
rect 11336 4768 11388 4820
rect 7012 4632 7064 4684
rect 7472 4632 7524 4684
rect 7564 4675 7616 4684
rect 7564 4641 7573 4675
rect 7573 4641 7607 4675
rect 7607 4641 7616 4675
rect 7564 4632 7616 4641
rect 8300 4632 8352 4684
rect 8668 4632 8720 4684
rect 9036 4632 9088 4684
rect 1492 4607 1544 4616
rect 1492 4573 1501 4607
rect 1501 4573 1535 4607
rect 1535 4573 1544 4607
rect 1492 4564 1544 4573
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 1768 4496 1820 4548
rect 3332 4564 3384 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 5908 4564 5960 4616
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 8760 4564 8812 4616
rect 9588 4564 9640 4616
rect 11888 4700 11940 4752
rect 12992 4768 13044 4820
rect 13176 4768 13228 4820
rect 14372 4768 14424 4820
rect 14832 4768 14884 4820
rect 16212 4811 16264 4820
rect 16212 4777 16221 4811
rect 16221 4777 16255 4811
rect 16255 4777 16264 4811
rect 16212 4768 16264 4777
rect 17408 4768 17460 4820
rect 13912 4700 13964 4752
rect 9864 4564 9916 4616
rect 10048 4564 10100 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 11244 4564 11296 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 480 4428 532 4480
rect 2412 4539 2464 4548
rect 2412 4505 2421 4539
rect 2421 4505 2455 4539
rect 2455 4505 2464 4539
rect 2412 4496 2464 4505
rect 5816 4496 5868 4548
rect 2320 4428 2372 4480
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 4712 4428 4764 4480
rect 7104 4496 7156 4548
rect 7564 4428 7616 4480
rect 9680 4496 9732 4548
rect 12440 4564 12492 4616
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 15016 4675 15068 4684
rect 15016 4641 15025 4675
rect 15025 4641 15059 4675
rect 15059 4641 15068 4675
rect 15016 4632 15068 4641
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 17776 4768 17828 4820
rect 17868 4768 17920 4820
rect 17684 4700 17736 4752
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 20444 4768 20496 4820
rect 22376 4768 22428 4820
rect 22560 4768 22612 4820
rect 18604 4632 18656 4684
rect 21548 4700 21600 4752
rect 21640 4743 21692 4752
rect 21640 4709 21649 4743
rect 21649 4709 21683 4743
rect 21683 4709 21692 4743
rect 21640 4700 21692 4709
rect 12716 4564 12768 4616
rect 13360 4539 13412 4548
rect 13360 4505 13369 4539
rect 13369 4505 13403 4539
rect 13403 4505 13412 4539
rect 13360 4496 13412 4505
rect 13544 4564 13596 4616
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15108 4607 15160 4616
rect 15108 4573 15142 4607
rect 15142 4573 15160 4607
rect 15108 4564 15160 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17040 4607 17092 4616
rect 17040 4573 17058 4607
rect 17058 4573 17092 4607
rect 17040 4564 17092 4573
rect 17684 4564 17736 4616
rect 13728 4496 13780 4548
rect 10784 4428 10836 4480
rect 11428 4428 11480 4480
rect 11888 4428 11940 4480
rect 11980 4471 12032 4480
rect 11980 4437 11989 4471
rect 11989 4437 12023 4471
rect 12023 4437 12032 4471
rect 11980 4428 12032 4437
rect 12256 4428 12308 4480
rect 12440 4428 12492 4480
rect 13268 4428 13320 4480
rect 13636 4428 13688 4480
rect 13912 4428 13964 4480
rect 17408 4428 17460 4480
rect 17500 4428 17552 4480
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 21088 4675 21140 4684
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 19340 4564 19392 4616
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 19248 4496 19300 4548
rect 19708 4496 19760 4548
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 20812 4564 20864 4616
rect 21364 4564 21416 4616
rect 21640 4496 21692 4548
rect 22652 4675 22704 4684
rect 22652 4641 22661 4675
rect 22661 4641 22695 4675
rect 22695 4641 22704 4675
rect 22652 4632 22704 4641
rect 27436 4811 27488 4820
rect 27436 4777 27445 4811
rect 27445 4777 27479 4811
rect 27479 4777 27488 4811
rect 27436 4768 27488 4777
rect 24216 4700 24268 4752
rect 25136 4700 25188 4752
rect 25872 4700 25924 4752
rect 21824 4564 21876 4616
rect 22100 4496 22152 4548
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 22928 4564 22980 4616
rect 22560 4496 22612 4548
rect 22652 4496 22704 4548
rect 23112 4564 23164 4616
rect 24400 4607 24452 4616
rect 24400 4573 24409 4607
rect 24409 4573 24443 4607
rect 24443 4573 24452 4607
rect 24400 4564 24452 4573
rect 25780 4675 25832 4684
rect 25780 4641 25789 4675
rect 25789 4641 25823 4675
rect 25823 4641 25832 4675
rect 25780 4632 25832 4641
rect 26148 4632 26200 4684
rect 27436 4632 27488 4684
rect 23388 4496 23440 4548
rect 19156 4428 19208 4480
rect 19616 4428 19668 4480
rect 20444 4428 20496 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 21548 4428 21600 4480
rect 22376 4428 22428 4480
rect 23940 4496 23992 4548
rect 24308 4496 24360 4548
rect 25228 4496 25280 4548
rect 26608 4607 26660 4616
rect 26608 4573 26642 4607
rect 26642 4573 26660 4607
rect 26608 4564 26660 4573
rect 26792 4607 26844 4616
rect 26792 4573 26801 4607
rect 26801 4573 26835 4607
rect 26835 4573 26844 4607
rect 26792 4564 26844 4573
rect 31116 4768 31168 4820
rect 29460 4700 29512 4752
rect 27896 4675 27948 4684
rect 27896 4641 27905 4675
rect 27905 4641 27939 4675
rect 27939 4641 27948 4675
rect 27896 4632 27948 4641
rect 29276 4632 29328 4684
rect 29828 4632 29880 4684
rect 30012 4743 30064 4752
rect 30012 4709 30021 4743
rect 30021 4709 30055 4743
rect 30055 4709 30064 4743
rect 30012 4700 30064 4709
rect 31208 4700 31260 4752
rect 28172 4607 28224 4616
rect 28172 4573 28181 4607
rect 28181 4573 28215 4607
rect 28215 4573 28224 4607
rect 28172 4564 28224 4573
rect 25780 4496 25832 4548
rect 30012 4564 30064 4616
rect 23572 4428 23624 4480
rect 24124 4428 24176 4480
rect 24952 4471 25004 4480
rect 24952 4437 24961 4471
rect 24961 4437 24995 4471
rect 24995 4437 25004 4471
rect 24952 4428 25004 4437
rect 25320 4471 25372 4480
rect 25320 4437 25329 4471
rect 25329 4437 25363 4471
rect 25363 4437 25372 4471
rect 25320 4428 25372 4437
rect 25596 4428 25648 4480
rect 30288 4496 30340 4548
rect 31392 4675 31444 4684
rect 31392 4641 31401 4675
rect 31401 4641 31435 4675
rect 31435 4641 31444 4675
rect 31392 4632 31444 4641
rect 30748 4607 30800 4616
rect 30748 4573 30757 4607
rect 30757 4573 30791 4607
rect 30791 4573 30800 4607
rect 30748 4564 30800 4573
rect 31116 4564 31168 4616
rect 32404 4768 32456 4820
rect 32772 4768 32824 4820
rect 33692 4768 33744 4820
rect 33876 4768 33928 4820
rect 34428 4768 34480 4820
rect 34520 4768 34572 4820
rect 35164 4768 35216 4820
rect 36636 4768 36688 4820
rect 39396 4811 39448 4820
rect 39396 4777 39405 4811
rect 39405 4777 39439 4811
rect 39439 4777 39448 4811
rect 39396 4768 39448 4777
rect 31852 4700 31904 4752
rect 32128 4632 32180 4684
rect 32404 4675 32456 4684
rect 32404 4641 32438 4675
rect 32438 4641 32456 4675
rect 32404 4632 32456 4641
rect 32588 4607 32640 4650
rect 32588 4598 32597 4607
rect 32597 4598 32631 4607
rect 32631 4598 32640 4607
rect 34428 4632 34480 4684
rect 34796 4564 34848 4616
rect 37004 4607 37056 4616
rect 37004 4573 37013 4607
rect 37013 4573 37047 4607
rect 37047 4573 37056 4607
rect 37004 4564 37056 4573
rect 37096 4564 37148 4616
rect 39212 4607 39264 4616
rect 39212 4573 39221 4607
rect 39221 4573 39255 4607
rect 39255 4573 39264 4607
rect 39212 4564 39264 4573
rect 34704 4539 34756 4548
rect 34704 4505 34713 4539
rect 34713 4505 34747 4539
rect 34747 4505 34756 4539
rect 34704 4496 34756 4505
rect 27620 4471 27672 4480
rect 27620 4437 27629 4471
rect 27629 4437 27663 4471
rect 27663 4437 27672 4471
rect 27620 4428 27672 4437
rect 28908 4471 28960 4480
rect 28908 4437 28917 4471
rect 28917 4437 28951 4471
rect 28951 4437 28960 4471
rect 28908 4428 28960 4437
rect 29092 4471 29144 4480
rect 29092 4437 29101 4471
rect 29101 4437 29135 4471
rect 29135 4437 29144 4471
rect 29092 4428 29144 4437
rect 31116 4428 31168 4480
rect 31300 4428 31352 4480
rect 32220 4428 32272 4480
rect 36912 4428 36964 4480
rect 38292 4428 38344 4480
rect 39304 4428 39356 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 9010 4326 9062 4378
rect 9074 4326 9126 4378
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 15010 4326 15062 4378
rect 15074 4326 15126 4378
rect 15138 4326 15190 4378
rect 15202 4326 15254 4378
rect 15266 4326 15318 4378
rect 21010 4326 21062 4378
rect 21074 4326 21126 4378
rect 21138 4326 21190 4378
rect 21202 4326 21254 4378
rect 21266 4326 21318 4378
rect 27010 4326 27062 4378
rect 27074 4326 27126 4378
rect 27138 4326 27190 4378
rect 27202 4326 27254 4378
rect 27266 4326 27318 4378
rect 33010 4326 33062 4378
rect 33074 4326 33126 4378
rect 33138 4326 33190 4378
rect 33202 4326 33254 4378
rect 33266 4326 33318 4378
rect 39010 4326 39062 4378
rect 39074 4326 39126 4378
rect 39138 4326 39190 4378
rect 39202 4326 39254 4378
rect 39266 4326 39318 4378
rect 1492 4199 1544 4208
rect 1492 4165 1501 4199
rect 1501 4165 1535 4199
rect 1535 4165 1544 4199
rect 1492 4156 1544 4165
rect 1860 4199 1912 4208
rect 1860 4165 1869 4199
rect 1869 4165 1903 4199
rect 1903 4165 1912 4199
rect 1860 4156 1912 4165
rect 2504 4156 2556 4208
rect 2688 4224 2740 4276
rect 3332 4224 3384 4276
rect 3516 4267 3568 4276
rect 3516 4233 3525 4267
rect 3525 4233 3559 4267
rect 3559 4233 3568 4267
rect 3516 4224 3568 4233
rect 4436 4224 4488 4276
rect 3148 4156 3200 4208
rect 5632 4224 5684 4276
rect 1952 4088 2004 4140
rect 2964 4088 3016 4140
rect 4344 4131 4396 4140
rect 4344 4097 4362 4131
rect 4362 4097 4396 4131
rect 4344 4088 4396 4097
rect 6184 4156 6236 4208
rect 7104 4224 7156 4276
rect 7380 4224 7432 4276
rect 9036 4224 9088 4276
rect 9956 4224 10008 4276
rect 10324 4224 10376 4276
rect 11980 4224 12032 4276
rect 12532 4224 12584 4276
rect 5724 4088 5776 4140
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 2320 4020 2372 4072
rect 3608 4020 3660 4072
rect 4804 4020 4856 4072
rect 5080 4020 5132 4072
rect 5448 4020 5500 4072
rect 3240 3884 3292 3936
rect 6092 3884 6144 3936
rect 6460 3927 6512 3936
rect 6460 3893 6469 3927
rect 6469 3893 6503 3927
rect 6503 3893 6512 3927
rect 6460 3884 6512 3893
rect 7656 4088 7708 4140
rect 9128 4199 9180 4208
rect 9128 4165 9137 4199
rect 9137 4165 9171 4199
rect 9171 4165 9180 4199
rect 9128 4156 9180 4165
rect 11612 4156 11664 4208
rect 14740 4224 14792 4276
rect 15016 4224 15068 4276
rect 16672 4224 16724 4276
rect 17040 4156 17092 4208
rect 9496 4088 9548 4140
rect 7104 4020 7156 4072
rect 7564 3952 7616 4004
rect 7472 3884 7524 3936
rect 8944 4020 8996 4072
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 10508 4088 10560 4140
rect 12164 4088 12216 4140
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12716 4088 12768 4140
rect 13268 4088 13320 4140
rect 9680 4020 9732 4072
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 10784 4020 10836 4072
rect 8852 3952 8904 4004
rect 13360 4020 13412 4072
rect 8024 3884 8076 3936
rect 10600 3884 10652 3936
rect 11060 3884 11112 3936
rect 11336 3884 11388 3936
rect 11980 3884 12032 3936
rect 12624 3884 12676 3936
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 14464 3884 14516 3936
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 15108 4020 15160 4072
rect 16212 4088 16264 4140
rect 16580 4088 16632 4140
rect 17132 4131 17184 4140
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 17776 4088 17828 4140
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 20628 4156 20680 4208
rect 20904 4156 20956 4208
rect 19616 4131 19668 4140
rect 19616 4097 19625 4131
rect 19625 4097 19659 4131
rect 19659 4097 19668 4131
rect 19616 4088 19668 4097
rect 21456 4131 21508 4140
rect 21456 4097 21465 4131
rect 21465 4097 21499 4131
rect 21499 4097 21508 4131
rect 21456 4088 21508 4097
rect 21640 4199 21692 4208
rect 21640 4165 21649 4199
rect 21649 4165 21683 4199
rect 21683 4165 21692 4199
rect 21640 4156 21692 4165
rect 15476 4063 15528 4072
rect 15476 4029 15485 4063
rect 15485 4029 15519 4063
rect 15519 4029 15528 4063
rect 15476 4020 15528 4029
rect 16120 4020 16172 4072
rect 17592 4063 17644 4072
rect 17592 4029 17601 4063
rect 17601 4029 17635 4063
rect 17635 4029 17644 4063
rect 17592 4020 17644 4029
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19432 4020 19484 4072
rect 19892 4063 19944 4072
rect 19892 4029 19901 4063
rect 19901 4029 19935 4063
rect 19935 4029 19944 4063
rect 19892 4020 19944 4029
rect 21732 4020 21784 4072
rect 22468 4224 22520 4276
rect 22560 4267 22612 4276
rect 22560 4233 22569 4267
rect 22569 4233 22603 4267
rect 22603 4233 22612 4267
rect 22560 4224 22612 4233
rect 22836 4156 22888 4208
rect 22468 4088 22520 4140
rect 24308 4224 24360 4276
rect 24216 4131 24268 4140
rect 24216 4097 24225 4131
rect 24225 4097 24259 4131
rect 24259 4097 24268 4131
rect 24216 4088 24268 4097
rect 24860 4131 24912 4140
rect 24860 4097 24869 4131
rect 24869 4097 24903 4131
rect 24903 4097 24912 4131
rect 24860 4088 24912 4097
rect 25044 4224 25096 4276
rect 29092 4224 29144 4276
rect 29184 4224 29236 4276
rect 30656 4224 30708 4276
rect 31668 4224 31720 4276
rect 31760 4224 31812 4276
rect 32496 4224 32548 4276
rect 25780 4156 25832 4208
rect 26332 4156 26384 4208
rect 25228 4088 25280 4140
rect 25412 4088 25464 4140
rect 16580 3952 16632 4004
rect 16396 3884 16448 3936
rect 17592 3884 17644 3936
rect 20812 3952 20864 4004
rect 22376 3952 22428 4004
rect 18420 3884 18472 3936
rect 18512 3884 18564 3936
rect 21732 3884 21784 3936
rect 21824 3884 21876 3936
rect 22836 4063 22888 4072
rect 22836 4029 22845 4063
rect 22845 4029 22879 4063
rect 22879 4029 22888 4063
rect 22836 4020 22888 4029
rect 23296 4020 23348 4072
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 23940 4063 23992 4072
rect 23940 4029 23949 4063
rect 23949 4029 23983 4063
rect 23983 4029 23992 4063
rect 23940 4020 23992 4029
rect 24032 4063 24084 4072
rect 24032 4029 24066 4063
rect 24066 4029 24084 4063
rect 25688 4088 25740 4140
rect 26240 4088 26292 4140
rect 26792 4156 26844 4208
rect 27160 4156 27212 4208
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 26608 4088 26660 4140
rect 30104 4156 30156 4208
rect 30840 4156 30892 4208
rect 24032 4020 24084 4029
rect 26424 4020 26476 4072
rect 27620 4088 27672 4140
rect 29552 4131 29604 4140
rect 29552 4097 29561 4131
rect 29561 4097 29595 4131
rect 29595 4097 29604 4131
rect 29552 4088 29604 4097
rect 30932 4088 30984 4140
rect 31484 4156 31536 4208
rect 33140 4156 33192 4208
rect 31116 4088 31168 4140
rect 31392 4131 31444 4140
rect 31392 4097 31401 4131
rect 31401 4097 31435 4131
rect 31435 4097 31444 4131
rect 31392 4088 31444 4097
rect 31576 4088 31628 4140
rect 32496 4131 32548 4140
rect 32496 4097 32505 4131
rect 32505 4097 32539 4131
rect 32539 4097 32548 4131
rect 32496 4088 32548 4097
rect 26240 3952 26292 4004
rect 24032 3884 24084 3936
rect 24216 3884 24268 3936
rect 25688 3884 25740 3936
rect 26148 3884 26200 3936
rect 26332 3927 26384 3936
rect 26332 3893 26341 3927
rect 26341 3893 26375 3927
rect 26375 3893 26384 3927
rect 26332 3884 26384 3893
rect 26700 3927 26752 3936
rect 26700 3893 26709 3927
rect 26709 3893 26743 3927
rect 26743 3893 26752 3927
rect 26700 3884 26752 3893
rect 27804 3884 27856 3936
rect 28172 3952 28224 4004
rect 28264 3952 28316 4004
rect 28448 4020 28500 4072
rect 28908 4020 28960 4072
rect 29092 4020 29144 4072
rect 29920 4020 29972 4072
rect 32220 4020 32272 4072
rect 38844 4224 38896 4276
rect 34336 4156 34388 4208
rect 36360 4156 36412 4208
rect 38292 4156 38344 4208
rect 33324 4088 33376 4140
rect 33692 4088 33744 4140
rect 34244 4088 34296 4140
rect 35072 4088 35124 4140
rect 36176 4131 36228 4140
rect 36176 4097 36185 4131
rect 36185 4097 36219 4131
rect 36219 4097 36228 4131
rect 36176 4088 36228 4097
rect 34336 4063 34388 4072
rect 34336 4029 34345 4063
rect 34345 4029 34379 4063
rect 34379 4029 34388 4063
rect 34336 4020 34388 4029
rect 34520 4020 34572 4072
rect 32128 3952 32180 4004
rect 32588 3952 32640 4004
rect 37188 4088 37240 4140
rect 38752 4088 38804 4140
rect 37280 3952 37332 4004
rect 39120 4088 39172 4140
rect 39488 3952 39540 4004
rect 29644 3884 29696 3936
rect 30472 3884 30524 3936
rect 30840 3884 30892 3936
rect 31576 3927 31628 3936
rect 31576 3893 31585 3927
rect 31585 3893 31619 3927
rect 31619 3893 31628 3927
rect 31576 3884 31628 3893
rect 32312 3927 32364 3936
rect 32312 3893 32321 3927
rect 32321 3893 32355 3927
rect 32355 3893 32364 3927
rect 32312 3884 32364 3893
rect 32680 3927 32732 3936
rect 32680 3893 32689 3927
rect 32689 3893 32723 3927
rect 32723 3893 32732 3927
rect 32680 3884 32732 3893
rect 34060 3884 34112 3936
rect 36636 3927 36688 3936
rect 36636 3893 36645 3927
rect 36645 3893 36679 3927
rect 36679 3893 36688 3927
rect 36636 3884 36688 3893
rect 39028 3927 39080 3936
rect 39028 3893 39037 3927
rect 39037 3893 39071 3927
rect 39071 3893 39080 3927
rect 39028 3884 39080 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 13950 3782 14002 3834
rect 14014 3782 14066 3834
rect 14078 3782 14130 3834
rect 14142 3782 14194 3834
rect 14206 3782 14258 3834
rect 19950 3782 20002 3834
rect 20014 3782 20066 3834
rect 20078 3782 20130 3834
rect 20142 3782 20194 3834
rect 20206 3782 20258 3834
rect 25950 3782 26002 3834
rect 26014 3782 26066 3834
rect 26078 3782 26130 3834
rect 26142 3782 26194 3834
rect 26206 3782 26258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 37950 3782 38002 3834
rect 38014 3782 38066 3834
rect 38078 3782 38130 3834
rect 38142 3782 38194 3834
rect 38206 3782 38258 3834
rect 1124 3680 1176 3732
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 1676 3612 1728 3664
rect 6552 3612 6604 3664
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 7380 3680 7432 3732
rect 7932 3680 7984 3732
rect 8392 3680 8444 3732
rect 8852 3680 8904 3732
rect 9312 3680 9364 3732
rect 1308 3544 1360 3596
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 2136 3476 2188 3528
rect 2320 3544 2372 3596
rect 2228 3451 2280 3460
rect 2228 3417 2237 3451
rect 2237 3417 2271 3451
rect 2271 3417 2280 3451
rect 2228 3408 2280 3417
rect 2688 3408 2740 3460
rect 3976 3476 4028 3528
rect 4896 3544 4948 3596
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 6460 3544 6512 3596
rect 7380 3544 7432 3596
rect 8668 3612 8720 3664
rect 8944 3612 8996 3664
rect 9680 3612 9732 3664
rect 1400 3340 1452 3392
rect 2136 3340 2188 3392
rect 3332 3340 3384 3392
rect 3608 3340 3660 3392
rect 3700 3340 3752 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 5264 3476 5316 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 8760 3544 8812 3596
rect 9220 3587 9272 3596
rect 9220 3553 9229 3587
rect 9229 3553 9263 3587
rect 9263 3553 9272 3587
rect 9220 3544 9272 3553
rect 9588 3544 9640 3596
rect 10232 3544 10284 3596
rect 12716 3680 12768 3732
rect 12164 3612 12216 3664
rect 12256 3612 12308 3664
rect 12440 3612 12492 3664
rect 16488 3680 16540 3732
rect 16672 3680 16724 3732
rect 12900 3612 12952 3664
rect 14832 3612 14884 3664
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 11060 3587 11112 3596
rect 11060 3553 11069 3587
rect 11069 3553 11103 3587
rect 11103 3553 11112 3587
rect 11060 3544 11112 3553
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8852 3476 8904 3528
rect 9680 3476 9732 3528
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 10876 3519 10928 3528
rect 10876 3485 10910 3519
rect 10910 3485 10928 3519
rect 10876 3476 10928 3485
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 13268 3544 13320 3596
rect 13544 3544 13596 3596
rect 13820 3544 13872 3596
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 15200 3544 15252 3596
rect 15476 3544 15528 3596
rect 16120 3544 16172 3596
rect 16488 3544 16540 3596
rect 16856 3587 16908 3596
rect 16856 3553 16874 3587
rect 16874 3553 16908 3587
rect 16856 3544 16908 3553
rect 17592 3680 17644 3732
rect 19800 3680 19852 3732
rect 17408 3612 17460 3664
rect 18788 3612 18840 3664
rect 12624 3476 12676 3528
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 13176 3476 13228 3528
rect 4712 3340 4764 3392
rect 5540 3340 5592 3392
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 6828 3340 6880 3392
rect 7380 3340 7432 3392
rect 9036 3408 9088 3460
rect 8208 3383 8260 3392
rect 8208 3349 8217 3383
rect 8217 3349 8251 3383
rect 8251 3349 8260 3383
rect 8208 3340 8260 3349
rect 8576 3340 8628 3392
rect 9588 3340 9640 3392
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 12532 3451 12584 3460
rect 12532 3417 12541 3451
rect 12541 3417 12575 3451
rect 12575 3417 12584 3451
rect 12532 3408 12584 3417
rect 13268 3408 13320 3460
rect 14004 3408 14056 3460
rect 12440 3340 12492 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 13544 3383 13596 3392
rect 13544 3349 13553 3383
rect 13553 3349 13587 3383
rect 13587 3349 13596 3383
rect 13544 3340 13596 3349
rect 14188 3476 14240 3528
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 24768 3680 24820 3732
rect 19432 3587 19484 3596
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 19524 3544 19576 3596
rect 25688 3612 25740 3664
rect 27620 3723 27672 3732
rect 27620 3689 27629 3723
rect 27629 3689 27663 3723
rect 27663 3689 27672 3723
rect 27620 3680 27672 3689
rect 25504 3587 25556 3596
rect 25504 3553 25513 3587
rect 25513 3553 25547 3587
rect 25547 3553 25556 3587
rect 25504 3544 25556 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 26792 3587 26844 3596
rect 26792 3553 26826 3587
rect 26826 3553 26844 3587
rect 26792 3544 26844 3553
rect 27712 3587 27764 3596
rect 27712 3553 27721 3587
rect 27721 3553 27755 3587
rect 27755 3553 27764 3587
rect 27712 3544 27764 3553
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 18144 3476 18196 3528
rect 18052 3408 18104 3460
rect 18696 3476 18748 3528
rect 19340 3476 19392 3528
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 21732 3476 21784 3528
rect 22652 3476 22704 3528
rect 19064 3408 19116 3460
rect 19432 3408 19484 3460
rect 20996 3408 21048 3460
rect 20444 3340 20496 3392
rect 20904 3340 20956 3392
rect 22100 3408 22152 3460
rect 23020 3451 23072 3460
rect 23020 3417 23029 3451
rect 23029 3417 23063 3451
rect 23063 3417 23072 3451
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 25872 3476 25924 3528
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 28356 3476 28408 3528
rect 28908 3476 28960 3528
rect 29920 3680 29972 3732
rect 32036 3680 32088 3732
rect 32128 3680 32180 3732
rect 29644 3544 29696 3596
rect 31024 3587 31076 3596
rect 31024 3553 31033 3587
rect 31033 3553 31067 3587
rect 31067 3553 31076 3587
rect 31024 3544 31076 3553
rect 31668 3587 31720 3596
rect 31668 3553 31677 3587
rect 31677 3553 31711 3587
rect 31711 3553 31720 3587
rect 31668 3544 31720 3553
rect 30104 3476 30156 3528
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31944 3519 31996 3528
rect 31944 3485 31953 3519
rect 31953 3485 31987 3519
rect 31987 3485 31996 3519
rect 31944 3476 31996 3485
rect 32036 3519 32088 3528
rect 32036 3485 32070 3519
rect 32070 3485 32088 3519
rect 32036 3476 32088 3485
rect 23020 3408 23072 3417
rect 22652 3340 22704 3392
rect 23480 3340 23532 3392
rect 24860 3408 24912 3460
rect 34244 3680 34296 3732
rect 34336 3680 34388 3732
rect 38292 3680 38344 3732
rect 39396 3723 39448 3732
rect 39396 3689 39405 3723
rect 39405 3689 39439 3723
rect 39439 3689 39448 3723
rect 39396 3680 39448 3689
rect 33508 3612 33560 3664
rect 34612 3612 34664 3664
rect 38016 3612 38068 3664
rect 39948 3612 40000 3664
rect 34428 3544 34480 3596
rect 32864 3476 32916 3528
rect 35072 3544 35124 3596
rect 34704 3519 34756 3528
rect 34704 3485 34713 3519
rect 34713 3485 34747 3519
rect 34747 3485 34756 3519
rect 34704 3476 34756 3485
rect 35164 3519 35216 3528
rect 35164 3485 35173 3519
rect 35173 3485 35207 3519
rect 35207 3485 35216 3519
rect 35164 3476 35216 3485
rect 35624 3476 35676 3528
rect 38292 3476 38344 3528
rect 38752 3476 38804 3528
rect 38844 3519 38896 3528
rect 38844 3485 38853 3519
rect 38853 3485 38887 3519
rect 38887 3485 38896 3519
rect 38844 3476 38896 3485
rect 38936 3476 38988 3528
rect 27620 3340 27672 3392
rect 29000 3383 29052 3392
rect 29000 3349 29009 3383
rect 29009 3349 29043 3383
rect 29043 3349 29052 3383
rect 29000 3340 29052 3349
rect 29368 3383 29420 3392
rect 29368 3349 29377 3383
rect 29377 3349 29411 3383
rect 29411 3349 29420 3383
rect 29368 3340 29420 3349
rect 29644 3340 29696 3392
rect 31392 3340 31444 3392
rect 33324 3383 33376 3392
rect 33324 3349 33333 3383
rect 33333 3349 33367 3383
rect 33367 3349 33376 3383
rect 33324 3340 33376 3349
rect 35256 3408 35308 3460
rect 39120 3408 39172 3460
rect 34520 3340 34572 3392
rect 34980 3340 35032 3392
rect 35716 3340 35768 3392
rect 37648 3340 37700 3392
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 9010 3238 9062 3290
rect 9074 3238 9126 3290
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 15010 3238 15062 3290
rect 15074 3238 15126 3290
rect 15138 3238 15190 3290
rect 15202 3238 15254 3290
rect 15266 3238 15318 3290
rect 21010 3238 21062 3290
rect 21074 3238 21126 3290
rect 21138 3238 21190 3290
rect 21202 3238 21254 3290
rect 21266 3238 21318 3290
rect 27010 3238 27062 3290
rect 27074 3238 27126 3290
rect 27138 3238 27190 3290
rect 27202 3238 27254 3290
rect 27266 3238 27318 3290
rect 33010 3238 33062 3290
rect 33074 3238 33126 3290
rect 33138 3238 33190 3290
rect 33202 3238 33254 3290
rect 33266 3238 33318 3290
rect 39010 3238 39062 3290
rect 39074 3238 39126 3290
rect 39138 3238 39190 3290
rect 39202 3238 39254 3290
rect 39266 3238 39318 3290
rect 1584 3136 1636 3188
rect 1860 3136 1912 3188
rect 3884 3136 3936 3188
rect 4988 3136 5040 3188
rect 1492 3111 1544 3120
rect 1492 3077 1501 3111
rect 1501 3077 1535 3111
rect 1535 3077 1544 3111
rect 1492 3068 1544 3077
rect 4436 3068 4488 3120
rect 7288 3136 7340 3188
rect 7472 3136 7524 3188
rect 1400 3000 1452 3052
rect 2136 3000 2188 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4252 3000 4304 3052
rect 4896 3000 4948 3052
rect 6184 3068 6236 3120
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 5724 3000 5776 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 1676 2907 1728 2916
rect 1676 2873 1685 2907
rect 1685 2873 1719 2907
rect 1719 2873 1728 2907
rect 1676 2864 1728 2873
rect 3240 2932 3292 2984
rect 5816 2932 5868 2984
rect 10324 3136 10376 3188
rect 10876 3136 10928 3188
rect 11612 3136 11664 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8300 3000 8352 3052
rect 8852 3000 8904 3052
rect 9036 3000 9088 3052
rect 9588 3000 9640 3052
rect 10048 3068 10100 3120
rect 13268 3068 13320 3120
rect 10324 3043 10376 3052
rect 9128 2932 9180 2984
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 12992 3000 13044 3052
rect 16028 3068 16080 3120
rect 17592 3136 17644 3188
rect 20628 3136 20680 3188
rect 20720 3136 20772 3188
rect 19432 3068 19484 3120
rect 4712 2907 4764 2916
rect 4712 2873 4721 2907
rect 4721 2873 4755 2907
rect 4755 2873 4764 2907
rect 4712 2864 4764 2873
rect 6092 2864 6144 2916
rect 6552 2864 6604 2916
rect 11520 2932 11572 2984
rect 11888 2975 11940 2984
rect 11888 2941 11897 2975
rect 11897 2941 11931 2975
rect 11931 2941 11940 2975
rect 11888 2932 11940 2941
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 8760 2796 8812 2805
rect 9220 2796 9272 2848
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 12716 2864 12768 2873
rect 9588 2796 9640 2848
rect 9680 2796 9732 2848
rect 12440 2796 12492 2848
rect 14004 3000 14056 3052
rect 14372 3000 14424 3052
rect 14740 3000 14792 3052
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 13728 2864 13780 2916
rect 15660 3000 15712 3052
rect 16120 3000 16172 3052
rect 16764 3043 16816 3052
rect 16764 3009 16773 3043
rect 16773 3009 16807 3043
rect 16807 3009 16816 3043
rect 16764 3000 16816 3009
rect 17224 3000 17276 3052
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 19524 3000 19576 3052
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 21916 3000 21968 3052
rect 13268 2796 13320 2848
rect 14924 2796 14976 2848
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 17592 2932 17644 2984
rect 18328 2975 18380 2984
rect 18328 2941 18346 2975
rect 18346 2941 18380 2975
rect 18328 2932 18380 2941
rect 18604 2932 18656 2984
rect 17040 2864 17092 2916
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 16948 2796 17000 2805
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17408 2796 17460 2848
rect 17776 2796 17828 2848
rect 17960 2796 18012 2848
rect 19064 2932 19116 2984
rect 18880 2864 18932 2916
rect 19800 2932 19852 2984
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 20812 2932 20864 2984
rect 23020 3043 23072 3052
rect 23020 3009 23029 3043
rect 23029 3009 23063 3043
rect 23063 3009 23072 3043
rect 23020 3000 23072 3009
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 25228 3000 25280 3052
rect 25596 3000 25648 3052
rect 26148 3000 26200 3052
rect 26424 3000 26476 3052
rect 19984 2796 20036 2848
rect 21088 2864 21140 2916
rect 23480 2975 23532 2984
rect 23480 2941 23489 2975
rect 23489 2941 23523 2975
rect 23523 2941 23532 2975
rect 23480 2932 23532 2941
rect 24216 2932 24268 2984
rect 25780 2975 25832 2984
rect 25780 2941 25789 2975
rect 25789 2941 25823 2975
rect 25823 2941 25832 2975
rect 25780 2932 25832 2941
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 28448 3136 28500 3188
rect 28908 3136 28960 3188
rect 29368 3136 29420 3188
rect 31852 3179 31904 3188
rect 31852 3145 31861 3179
rect 31861 3145 31895 3179
rect 31895 3145 31904 3179
rect 31852 3136 31904 3145
rect 31944 3136 31996 3188
rect 33324 3136 33376 3188
rect 33692 3179 33744 3188
rect 33692 3145 33701 3179
rect 33701 3145 33735 3179
rect 33735 3145 33744 3179
rect 33692 3136 33744 3145
rect 33784 3179 33836 3188
rect 33784 3145 33793 3179
rect 33793 3145 33827 3179
rect 33827 3145 33836 3179
rect 33784 3136 33836 3145
rect 34520 3136 34572 3188
rect 35440 3136 35492 3188
rect 35808 3136 35860 3188
rect 35992 3136 36044 3188
rect 37096 3136 37148 3188
rect 37648 3136 37700 3188
rect 38016 3179 38068 3188
rect 38016 3145 38025 3179
rect 38025 3145 38059 3179
rect 38059 3145 38068 3179
rect 38016 3136 38068 3145
rect 39396 3179 39448 3188
rect 39396 3145 39405 3179
rect 39405 3145 39439 3179
rect 39439 3145 39448 3179
rect 39396 3136 39448 3145
rect 28172 3043 28224 3052
rect 28172 3009 28181 3043
rect 28181 3009 28215 3043
rect 28215 3009 28224 3043
rect 28172 3000 28224 3009
rect 29920 3043 29972 3052
rect 29920 3009 29954 3043
rect 29954 3009 29972 3043
rect 29920 3000 29972 3009
rect 30748 3000 30800 3052
rect 31392 3000 31444 3052
rect 34152 3000 34204 3052
rect 34796 3000 34848 3052
rect 35348 3043 35400 3052
rect 35348 3009 35357 3043
rect 35357 3009 35391 3043
rect 35391 3009 35400 3043
rect 35348 3000 35400 3009
rect 27528 2932 27580 2984
rect 27620 2975 27672 2984
rect 27620 2941 27629 2975
rect 27629 2941 27663 2975
rect 27663 2941 27672 2975
rect 27620 2932 27672 2941
rect 24492 2864 24544 2916
rect 20352 2796 20404 2848
rect 20444 2796 20496 2848
rect 21180 2796 21232 2848
rect 21456 2796 21508 2848
rect 22744 2796 22796 2848
rect 24860 2796 24912 2848
rect 25504 2796 25556 2848
rect 26608 2864 26660 2916
rect 28356 2932 28408 2984
rect 28816 2932 28868 2984
rect 29828 2975 29880 2984
rect 29828 2941 29837 2975
rect 29837 2941 29871 2975
rect 29871 2941 29880 2975
rect 29828 2932 29880 2941
rect 30472 2932 30524 2984
rect 30840 2975 30892 2984
rect 30840 2941 30849 2975
rect 30849 2941 30883 2975
rect 30883 2941 30892 2975
rect 30840 2932 30892 2941
rect 31484 2932 31536 2984
rect 25780 2796 25832 2848
rect 26424 2796 26476 2848
rect 26792 2839 26844 2848
rect 26792 2805 26801 2839
rect 26801 2805 26835 2839
rect 26835 2805 26844 2839
rect 26792 2796 26844 2805
rect 27068 2796 27120 2848
rect 29368 2864 29420 2916
rect 31852 2932 31904 2984
rect 32128 2975 32180 2984
rect 32128 2941 32137 2975
rect 32137 2941 32171 2975
rect 32171 2941 32180 2975
rect 32128 2932 32180 2941
rect 28908 2796 28960 2848
rect 29920 2796 29972 2848
rect 31944 2796 31996 2848
rect 33600 2932 33652 2984
rect 35716 3043 35768 3052
rect 35716 3009 35725 3043
rect 35725 3009 35759 3043
rect 35759 3009 35768 3043
rect 35716 3000 35768 3009
rect 35808 3000 35860 3052
rect 36084 2932 36136 2984
rect 37280 3000 37332 3052
rect 37648 2932 37700 2984
rect 38292 3043 38344 3052
rect 38292 3009 38301 3043
rect 38301 3009 38335 3043
rect 38335 3009 38344 3043
rect 38292 3000 38344 3009
rect 36360 2864 36412 2916
rect 36728 2864 36780 2916
rect 39672 2864 39724 2916
rect 34612 2796 34664 2848
rect 35164 2839 35216 2848
rect 35164 2805 35173 2839
rect 35173 2805 35207 2839
rect 35207 2805 35216 2839
rect 35164 2796 35216 2805
rect 35348 2796 35400 2848
rect 35992 2796 36044 2848
rect 39028 2839 39080 2848
rect 39028 2805 39037 2839
rect 39037 2805 39071 2839
rect 39071 2805 39080 2839
rect 39028 2796 39080 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 13950 2694 14002 2746
rect 14014 2694 14066 2746
rect 14078 2694 14130 2746
rect 14142 2694 14194 2746
rect 14206 2694 14258 2746
rect 19950 2694 20002 2746
rect 20014 2694 20066 2746
rect 20078 2694 20130 2746
rect 20142 2694 20194 2746
rect 20206 2694 20258 2746
rect 25950 2694 26002 2746
rect 26014 2694 26066 2746
rect 26078 2694 26130 2746
rect 26142 2694 26194 2746
rect 26206 2694 26258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 37950 2694 38002 2746
rect 38014 2694 38066 2746
rect 38078 2694 38130 2746
rect 38142 2694 38194 2746
rect 38206 2694 38258 2746
rect 2780 2592 2832 2644
rect 4344 2592 4396 2644
rect 3240 2524 3292 2576
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 3976 2456 4028 2508
rect 1492 2431 1544 2440
rect 1492 2397 1501 2431
rect 1501 2397 1535 2431
rect 1535 2397 1544 2431
rect 1492 2388 1544 2397
rect 2872 2388 2924 2440
rect 3056 2388 3108 2440
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 2412 2363 2464 2372
rect 2412 2329 2421 2363
rect 2421 2329 2455 2363
rect 2455 2329 2464 2363
rect 2412 2320 2464 2329
rect 3516 2388 3568 2440
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 3884 2320 3936 2372
rect 4804 2456 4856 2508
rect 5264 2456 5316 2508
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 6552 2592 6604 2644
rect 7840 2592 7892 2644
rect 6460 2524 6512 2576
rect 7380 2524 7432 2576
rect 7012 2456 7064 2508
rect 7564 2499 7616 2508
rect 7564 2465 7573 2499
rect 7573 2465 7607 2499
rect 7607 2465 7616 2499
rect 7564 2456 7616 2465
rect 8392 2524 8444 2576
rect 13268 2592 13320 2644
rect 13636 2592 13688 2644
rect 13912 2592 13964 2644
rect 8760 2456 8812 2508
rect 15292 2592 15344 2644
rect 15752 2592 15804 2644
rect 16120 2592 16172 2644
rect 17224 2635 17276 2644
rect 17224 2601 17233 2635
rect 17233 2601 17267 2635
rect 17267 2601 17276 2635
rect 17224 2592 17276 2601
rect 18788 2592 18840 2644
rect 13268 2456 13320 2508
rect 4160 2363 4212 2372
rect 4160 2329 4169 2363
rect 4169 2329 4203 2363
rect 4203 2329 4212 2363
rect 4160 2320 4212 2329
rect 4896 2363 4948 2372
rect 4896 2329 4905 2363
rect 4905 2329 4939 2363
rect 4939 2329 4948 2363
rect 4896 2320 4948 2329
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6276 2388 6328 2440
rect 6552 2320 6604 2372
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8484 2388 8536 2440
rect 9220 2388 9272 2440
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 8668 2320 8720 2372
rect 8760 2320 8812 2372
rect 9036 2320 9088 2372
rect 9496 2320 9548 2372
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 11152 2388 11204 2440
rect 11428 2388 11480 2440
rect 12164 2388 12216 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14280 2388 14332 2440
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 17408 2524 17460 2576
rect 18328 2524 18380 2576
rect 18880 2524 18932 2576
rect 17960 2456 18012 2508
rect 18052 2456 18104 2508
rect 20352 2592 20404 2644
rect 20628 2592 20680 2644
rect 22284 2592 22336 2644
rect 32220 2592 32272 2644
rect 33416 2592 33468 2644
rect 33784 2592 33836 2644
rect 22836 2567 22888 2576
rect 22836 2533 22845 2567
rect 22845 2533 22879 2567
rect 22879 2533 22888 2567
rect 22836 2524 22888 2533
rect 24032 2524 24084 2576
rect 22744 2456 22796 2508
rect 26516 2524 26568 2576
rect 29368 2567 29420 2576
rect 29368 2533 29377 2567
rect 29377 2533 29411 2567
rect 29411 2533 29420 2567
rect 29368 2524 29420 2533
rect 30472 2524 30524 2576
rect 31760 2524 31812 2576
rect 26884 2456 26936 2508
rect 30840 2499 30892 2508
rect 30840 2465 30849 2499
rect 30849 2465 30883 2499
rect 30883 2465 30892 2499
rect 30840 2456 30892 2465
rect 31484 2456 31536 2508
rect 32956 2524 33008 2576
rect 33692 2524 33744 2576
rect 33968 2524 34020 2576
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 15016 2388 15068 2440
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 19064 2431 19116 2440
rect 19064 2397 19073 2431
rect 19073 2397 19107 2431
rect 19107 2397 19116 2431
rect 19064 2388 19116 2397
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 15936 2320 15988 2372
rect 16580 2320 16632 2372
rect 16856 2320 16908 2372
rect 4252 2252 4304 2304
rect 4988 2295 5040 2304
rect 4988 2261 4997 2295
rect 4997 2261 5031 2295
rect 5031 2261 5040 2295
rect 4988 2252 5040 2261
rect 5632 2252 5684 2304
rect 6736 2252 6788 2304
rect 8208 2252 8260 2304
rect 11244 2252 11296 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12256 2295 12308 2304
rect 12256 2261 12265 2295
rect 12265 2261 12299 2295
rect 12299 2261 12308 2295
rect 12256 2252 12308 2261
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 17592 2252 17644 2304
rect 17776 2320 17828 2372
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 21916 2320 21968 2372
rect 22652 2320 22704 2372
rect 20812 2252 20864 2304
rect 24400 2388 24452 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 25136 2388 25188 2440
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 27620 2388 27672 2440
rect 28540 2388 28592 2440
rect 28724 2388 28776 2440
rect 29828 2431 29880 2440
rect 29828 2397 29837 2431
rect 29837 2397 29871 2431
rect 29871 2397 29880 2431
rect 29828 2388 29880 2397
rect 31944 2388 31996 2440
rect 24308 2252 24360 2304
rect 24860 2252 24912 2304
rect 25688 2252 25740 2304
rect 26516 2295 26568 2304
rect 26516 2261 26525 2295
rect 26525 2261 26559 2295
rect 26559 2261 26568 2295
rect 26516 2252 26568 2261
rect 26608 2252 26660 2304
rect 28816 2320 28868 2372
rect 28908 2320 28960 2372
rect 29092 2320 29144 2372
rect 29368 2320 29420 2372
rect 28264 2295 28316 2304
rect 28264 2261 28273 2295
rect 28273 2261 28307 2295
rect 28307 2261 28316 2295
rect 28264 2252 28316 2261
rect 28448 2252 28500 2304
rect 32404 2388 32456 2440
rect 33324 2456 33376 2508
rect 34060 2320 34112 2372
rect 36452 2524 36504 2576
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 35072 2431 35124 2440
rect 35072 2397 35081 2431
rect 35081 2397 35115 2431
rect 35115 2397 35124 2431
rect 35072 2388 35124 2397
rect 35440 2431 35492 2440
rect 35440 2397 35449 2431
rect 35449 2397 35483 2431
rect 35483 2397 35492 2431
rect 35440 2388 35492 2397
rect 36360 2431 36412 2440
rect 36360 2397 36369 2431
rect 36369 2397 36403 2431
rect 36403 2397 36412 2431
rect 36360 2388 36412 2397
rect 39396 2635 39448 2644
rect 39396 2601 39405 2635
rect 39405 2601 39439 2635
rect 39439 2601 39448 2635
rect 39396 2592 39448 2601
rect 39580 2524 39632 2576
rect 38108 2431 38160 2440
rect 38108 2397 38117 2431
rect 38117 2397 38151 2431
rect 38151 2397 38160 2431
rect 38108 2388 38160 2397
rect 38844 2431 38896 2440
rect 38844 2397 38853 2431
rect 38853 2397 38887 2431
rect 38887 2397 38896 2431
rect 38844 2388 38896 2397
rect 39212 2431 39264 2440
rect 39212 2397 39221 2431
rect 39221 2397 39255 2431
rect 39255 2397 39264 2431
rect 39212 2388 39264 2397
rect 32680 2295 32732 2304
rect 32680 2261 32689 2295
rect 32689 2261 32723 2295
rect 32723 2261 32732 2295
rect 32680 2252 32732 2261
rect 32772 2252 32824 2304
rect 33416 2295 33468 2304
rect 33416 2261 33425 2295
rect 33425 2261 33459 2295
rect 33459 2261 33468 2295
rect 33416 2252 33468 2261
rect 33784 2295 33836 2304
rect 33784 2261 33793 2295
rect 33793 2261 33827 2295
rect 33827 2261 33836 2295
rect 33784 2252 33836 2261
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 34888 2295 34940 2304
rect 34888 2261 34897 2295
rect 34897 2261 34931 2295
rect 34931 2261 34940 2295
rect 34888 2252 34940 2261
rect 35164 2252 35216 2304
rect 35624 2295 35676 2304
rect 35624 2261 35633 2295
rect 35633 2261 35667 2295
rect 35667 2261 35676 2295
rect 35624 2252 35676 2261
rect 36176 2295 36228 2304
rect 36176 2261 36185 2295
rect 36185 2261 36219 2295
rect 36219 2261 36228 2295
rect 36176 2252 36228 2261
rect 40040 2320 40092 2372
rect 38660 2295 38712 2304
rect 38660 2261 38669 2295
rect 38669 2261 38703 2295
rect 38703 2261 38712 2295
rect 38660 2252 38712 2261
rect 39948 2252 40000 2304
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 9010 2150 9062 2202
rect 9074 2150 9126 2202
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 15010 2150 15062 2202
rect 15074 2150 15126 2202
rect 15138 2150 15190 2202
rect 15202 2150 15254 2202
rect 15266 2150 15318 2202
rect 21010 2150 21062 2202
rect 21074 2150 21126 2202
rect 21138 2150 21190 2202
rect 21202 2150 21254 2202
rect 21266 2150 21318 2202
rect 27010 2150 27062 2202
rect 27074 2150 27126 2202
rect 27138 2150 27190 2202
rect 27202 2150 27254 2202
rect 27266 2150 27318 2202
rect 33010 2150 33062 2202
rect 33074 2150 33126 2202
rect 33138 2150 33190 2202
rect 33202 2150 33254 2202
rect 33266 2150 33318 2202
rect 39010 2150 39062 2202
rect 39074 2150 39126 2202
rect 39138 2150 39190 2202
rect 39202 2150 39254 2202
rect 39266 2150 39318 2202
rect 14280 2048 14332 2100
rect 18328 2048 18380 2100
rect 20812 2048 20864 2100
rect 22008 2048 22060 2100
rect 24676 2048 24728 2100
rect 27436 2048 27488 2100
rect 27528 2048 27580 2100
rect 32496 2048 32548 2100
rect 34428 2048 34480 2100
rect 36544 2048 36596 2100
rect 4988 1980 5040 2032
rect 11336 1980 11388 2032
rect 13912 1980 13964 2032
rect 15200 1980 15252 2032
rect 15660 1980 15712 2032
rect 22100 1980 22152 2032
rect 22560 1980 22612 2032
rect 26608 1980 26660 2032
rect 26792 1980 26844 2032
rect 1952 1776 2004 1828
rect 14280 1912 14332 1964
rect 14832 1912 14884 1964
rect 15384 1912 15436 1964
rect 19524 1912 19576 1964
rect 25504 1912 25556 1964
rect 25872 1912 25924 1964
rect 28356 1912 28408 1964
rect 29000 1980 29052 2032
rect 33600 1980 33652 2032
rect 33692 1980 33744 2032
rect 38844 1980 38896 2032
rect 29368 1912 29420 1964
rect 29736 1912 29788 1964
rect 30564 1912 30616 1964
rect 31944 1912 31996 1964
rect 36084 1912 36136 1964
rect 4160 1844 4212 1896
rect 10140 1844 10192 1896
rect 10416 1844 10468 1896
rect 12900 1844 12952 1896
rect 9864 1776 9916 1828
rect 12532 1776 12584 1828
rect 1676 1708 1728 1760
rect 22468 1844 22520 1896
rect 24584 1844 24636 1896
rect 35072 1844 35124 1896
rect 14280 1776 14332 1828
rect 29184 1776 29236 1828
rect 17224 1708 17276 1760
rect 25872 1708 25924 1760
rect 28264 1708 28316 1760
rect 38936 1708 38988 1760
rect 1032 1640 1084 1692
rect 8760 1640 8812 1692
rect 12164 1640 12216 1692
rect 19524 1640 19576 1692
rect 20628 1640 20680 1692
rect 27620 1640 27672 1692
rect 27988 1640 28040 1692
rect 28172 1640 28224 1692
rect 34704 1640 34756 1692
rect 4252 1572 4304 1624
rect 12624 1572 12676 1624
rect 15660 1572 15712 1624
rect 15844 1572 15896 1624
rect 19708 1572 19760 1624
rect 21640 1572 21692 1624
rect 27528 1572 27580 1624
rect 8484 1504 8536 1556
rect 17224 1504 17276 1556
rect 11060 1436 11112 1488
rect 16764 1436 16816 1488
rect 16948 1436 17000 1488
rect 17408 1436 17460 1488
rect 7196 1368 7248 1420
rect 9220 1368 9272 1420
rect 11336 1368 11388 1420
rect 20628 1504 20680 1556
rect 24676 1504 24728 1556
rect 27896 1504 27948 1556
rect 17592 1436 17644 1488
rect 19248 1436 19300 1488
rect 34612 1436 34664 1488
rect 35256 1436 35308 1488
rect 17684 1368 17736 1420
rect 18696 1368 18748 1420
rect 19156 1368 19208 1420
rect 20352 1368 20404 1420
rect 21916 1368 21968 1420
rect 31852 1368 31904 1420
rect 34244 1368 34296 1420
rect 36820 1368 36872 1420
rect 3424 1300 3476 1352
rect 4620 1300 4672 1352
rect 4712 1300 4764 1352
rect 7656 1300 7708 1352
rect 8852 1300 8904 1352
rect 10140 1300 10192 1352
rect 12072 1300 12124 1352
rect 12900 1300 12952 1352
rect 13084 1300 13136 1352
rect 15108 1300 15160 1352
rect 17316 1300 17368 1352
rect 19800 1300 19852 1352
rect 20076 1300 20128 1352
rect 21824 1300 21876 1352
rect 24492 1300 24544 1352
rect 25320 1300 25372 1352
rect 3608 1232 3660 1284
rect 6000 1232 6052 1284
rect 12992 1232 13044 1284
rect 16212 1232 16264 1284
rect 16488 1232 16540 1284
rect 20812 1232 20864 1284
rect 22008 1232 22060 1284
rect 24860 1232 24912 1284
rect 25044 1232 25096 1284
rect 26700 1232 26752 1284
rect 30288 1232 30340 1284
rect 33508 1300 33560 1352
rect 36360 1300 36412 1352
rect 37280 1300 37332 1352
rect 2504 1164 2556 1216
rect 4896 1164 4948 1216
rect 8760 1164 8812 1216
rect 9496 1164 9548 1216
rect 10692 1164 10744 1216
rect 13544 1164 13596 1216
rect 6828 1096 6880 1148
rect 7748 1096 7800 1148
rect 11612 1096 11664 1148
rect 3976 1028 4028 1080
rect 17500 1096 17552 1148
rect 16396 1028 16448 1080
rect 21732 1164 21784 1216
rect 24308 1164 24360 1216
rect 32772 1232 32824 1284
rect 35256 1232 35308 1284
rect 37188 1232 37240 1284
rect 31116 1164 31168 1216
rect 36452 1164 36504 1216
rect 17684 1096 17736 1148
rect 23020 1096 23072 1148
rect 23112 1096 23164 1148
rect 26424 1096 26476 1148
rect 26700 1096 26752 1148
rect 29184 1096 29236 1148
rect 34152 1096 34204 1148
rect 34980 1096 35032 1148
rect 36268 1096 36320 1148
rect 8300 960 8352 1012
rect 11336 960 11388 1012
rect 16488 960 16540 1012
rect 17316 960 17368 1012
rect 24032 1028 24084 1080
rect 24216 1028 24268 1080
rect 24952 1028 25004 1080
rect 29000 1028 29052 1080
rect 26424 960 26476 1012
rect 32680 1028 32732 1080
rect 34704 1028 34756 1080
rect 37004 1028 37056 1080
rect 31944 960 31996 1012
rect 35072 960 35124 1012
rect 6368 892 6420 944
rect 7472 824 7524 876
rect 9036 824 9088 876
rect 9220 892 9272 944
rect 11796 892 11848 944
rect 24768 892 24820 944
rect 25596 892 25648 944
rect 27344 892 27396 944
rect 28908 892 28960 944
rect 31576 892 31628 944
rect 31668 892 31720 944
rect 16488 824 16540 876
rect 22100 824 22152 876
rect 22284 824 22336 876
rect 26516 824 26568 876
rect 30012 824 30064 876
rect 32312 824 32364 876
rect 2688 756 2740 808
rect 2596 688 2648 740
rect 4896 688 4948 740
rect 2320 620 2372 672
rect 14004 756 14056 808
rect 14556 688 14608 740
rect 15660 688 15712 740
rect 17316 756 17368 808
rect 27712 756 27764 808
rect 30380 756 30432 808
rect 33048 756 33100 808
rect 33876 892 33928 944
rect 34796 892 34848 944
rect 36084 756 36136 808
rect 24676 688 24728 740
rect 24768 688 24820 740
rect 26332 688 26384 740
rect 27804 688 27856 740
rect 30656 688 30708 740
rect 22928 620 22980 672
rect 29460 620 29512 672
rect 35624 620 35676 672
rect 35808 620 35860 672
rect 37648 620 37700 672
rect 9680 552 9732 604
rect 11428 552 11480 604
rect 23664 552 23716 604
rect 26976 552 27028 604
rect 30472 552 30524 604
rect 31392 552 31444 604
rect 35348 552 35400 604
rect 2044 484 2096 536
rect 14004 484 14056 536
rect 14096 484 14148 536
rect 17316 484 17368 536
rect 17960 484 18012 536
rect 19432 484 19484 536
rect 28080 484 28132 536
rect 34888 484 34940 536
rect 36084 484 36136 536
rect 38752 484 38804 536
rect 5264 416 5316 468
rect 12072 416 12124 468
rect 12808 416 12860 468
rect 14832 416 14884 468
rect 14924 416 14976 468
rect 18144 416 18196 468
rect 23664 416 23716 468
rect 29092 416 29144 468
rect 30840 416 30892 468
rect 32588 416 32640 468
rect 11704 348 11756 400
rect 14556 348 14608 400
rect 14740 348 14792 400
rect 22192 348 22244 400
rect 24032 348 24084 400
rect 5908 280 5960 332
rect 8576 212 8628 264
rect 12256 212 12308 264
rect 14464 280 14516 332
rect 17868 280 17920 332
rect 20536 280 20588 332
rect 21180 280 21232 332
rect 22560 280 22612 332
rect 25780 280 25832 332
rect 26148 348 26200 400
rect 29644 348 29696 400
rect 33600 348 33652 400
rect 37832 348 37884 400
rect 29276 280 29328 332
rect 30564 280 30616 332
rect 34612 280 34664 332
rect 15752 212 15804 264
rect 27252 212 27304 264
rect 33416 212 33468 264
rect 11244 144 11296 196
rect 16028 144 16080 196
rect 27528 144 27580 196
rect 31300 144 31352 196
rect 36636 144 36688 196
rect 37556 144 37608 196
rect 22928 8 22980 60
rect 31484 8 31536 60
<< metal2 >>
rect 1674 11194 1730 11250
rect 2778 11194 2834 11250
rect 3882 11194 3938 11250
rect 3988 11206 4200 11234
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1308 9988 1360 9994
rect 1308 9930 1360 9936
rect 1032 7744 1084 7750
rect 1032 7686 1084 7692
rect 756 7472 808 7478
rect 756 7414 808 7420
rect 480 4480 532 4486
rect 480 4422 532 4428
rect 492 2009 520 4422
rect 478 2000 534 2009
rect 478 1935 534 1944
rect 768 1465 796 7414
rect 1044 1698 1072 7686
rect 1124 7200 1176 7206
rect 1124 7142 1176 7148
rect 1136 3738 1164 7142
rect 1216 6248 1268 6254
rect 1216 6190 1268 6196
rect 1124 3732 1176 3738
rect 1124 3674 1176 3680
rect 1228 1737 1256 6190
rect 1320 3602 1348 9930
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1412 8498 1440 9007
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1412 8022 1440 8191
rect 1400 8016 1452 8022
rect 1400 7958 1452 7964
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7449 1440 7822
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1504 7721 1532 7754
rect 1490 7712 1546 7721
rect 1490 7647 1546 7656
rect 1398 7440 1454 7449
rect 1596 7426 1624 10202
rect 1688 8566 1716 11194
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2320 9852 2372 9858
rect 2320 9794 2372 9800
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1398 7375 1454 7384
rect 1504 7398 1624 7426
rect 1674 7440 1730 7449
rect 1504 7290 1532 7398
rect 1674 7375 1676 7384
rect 1728 7375 1730 7384
rect 1676 7346 1728 7352
rect 1412 7262 1532 7290
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1412 6746 1440 7262
rect 1490 7168 1546 7177
rect 1490 7103 1546 7112
rect 1504 6934 1532 7103
rect 1492 6928 1544 6934
rect 1492 6870 1544 6876
rect 1412 6718 1532 6746
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1412 6322 1440 6559
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1504 6202 1532 6718
rect 1596 6361 1624 7278
rect 1674 6896 1730 6905
rect 1780 6866 1808 7278
rect 1674 6831 1730 6840
rect 1768 6860 1820 6866
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1504 6174 1624 6202
rect 1398 6080 1454 6089
rect 1398 6015 1454 6024
rect 1412 5710 1440 6015
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1308 3596 1360 3602
rect 1308 3538 1360 3544
rect 1412 3398 1440 5306
rect 1504 5302 1532 5743
rect 1596 5522 1624 6174
rect 1688 5642 1716 6831
rect 1768 6802 1820 6808
rect 1872 6730 1900 8842
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2226 7984 2282 7993
rect 2226 7919 2282 7928
rect 2240 7886 2268 7919
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2044 7812 2096 7818
rect 2044 7754 2096 7760
rect 2056 7313 2084 7754
rect 2042 7304 2098 7313
rect 2042 7239 2098 7248
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1766 6216 1822 6225
rect 1766 6151 1822 6160
rect 1780 5846 1808 6151
rect 2056 6100 2084 6938
rect 2332 6882 2360 9794
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2424 8242 2452 8910
rect 2516 8634 2544 9862
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2424 8214 2544 8242
rect 2516 7936 2544 8214
rect 2424 7908 2544 7936
rect 2424 7002 2452 7908
rect 2608 7834 2636 10066
rect 2792 9314 2820 11194
rect 3896 11098 3924 11194
rect 3988 11098 4016 11206
rect 3896 11070 4016 11098
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2780 9308 2832 9314
rect 2780 9250 2832 9256
rect 2884 9194 2912 10746
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3422 9616 3478 9625
rect 3422 9551 3478 9560
rect 2516 7806 2636 7834
rect 2700 9166 2912 9194
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2332 6854 2452 6882
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 1872 6072 2084 6100
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1596 5494 1716 5522
rect 1688 5302 1716 5494
rect 1872 5386 1900 6072
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 5808 2006 5817
rect 1950 5743 2006 5752
rect 1780 5358 1900 5386
rect 1964 5370 1992 5743
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2240 5545 2268 5578
rect 2226 5536 2282 5545
rect 2226 5471 2282 5480
rect 1952 5364 2004 5370
rect 1492 5296 1544 5302
rect 1492 5238 1544 5244
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1490 4992 1546 5001
rect 1490 4927 1546 4936
rect 1504 4622 1532 4927
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1490 4448 1546 4457
rect 1490 4383 1546 4392
rect 1504 4214 1532 4383
rect 1492 4208 1544 4214
rect 1492 4150 1544 4156
rect 1490 3904 1546 3913
rect 1490 3839 1546 3848
rect 1504 3534 1532 3839
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1490 3360 1546 3369
rect 1490 3295 1546 3304
rect 1504 3126 1532 3295
rect 1596 3194 1624 5170
rect 1780 4706 1808 5358
rect 1952 5306 2004 5312
rect 2332 5302 2360 6734
rect 1860 5296 1912 5302
rect 1858 5264 1860 5273
rect 2320 5296 2372 5302
rect 1912 5264 1914 5273
rect 2320 5238 2372 5244
rect 2424 5234 2452 6854
rect 2516 5846 2544 7806
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2608 5574 2636 7686
rect 2700 7002 2728 9166
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2778 8800 2834 8809
rect 2778 8735 2834 8744
rect 2792 7886 2820 8735
rect 2884 8634 2912 9046
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3332 8560 3384 8566
rect 3330 8528 3332 8537
rect 3384 8528 3386 8537
rect 3330 8463 3386 8472
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7290 2820 7686
rect 2884 7410 2912 7754
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 3436 7528 3464 9551
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3528 7886 3556 8327
rect 3620 8022 3648 9415
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3712 8634 3740 9318
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3698 8256 3754 8265
rect 3698 8191 3754 8200
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3712 7954 3740 8191
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3516 7880 3568 7886
rect 3568 7840 3648 7868
rect 3516 7822 3568 7828
rect 3252 7500 3464 7528
rect 2872 7404 2924 7410
rect 2924 7364 3004 7392
rect 2872 7346 2924 7352
rect 2792 7262 2912 7290
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2686 6896 2742 6905
rect 2686 6831 2742 6840
rect 2700 6662 2728 6831
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2884 6322 2912 7262
rect 2976 7206 3004 7364
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 3252 6730 3280 7500
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 1858 5199 1914 5208
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 2502 5128 2558 5137
rect 1872 4826 1900 5102
rect 2412 5092 2464 5098
rect 2502 5063 2558 5072
rect 2412 5034 2464 5040
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1676 4684 1728 4690
rect 1780 4678 1992 4706
rect 1676 4626 1728 4632
rect 1688 3670 1716 4626
rect 1860 4616 1912 4622
rect 1858 4584 1860 4593
rect 1912 4584 1914 4593
rect 1768 4548 1820 4554
rect 1858 4519 1914 4528
rect 1768 4490 1820 4496
rect 1780 4026 1808 4490
rect 1860 4208 1912 4214
rect 1858 4176 1860 4185
rect 1912 4176 1914 4185
rect 1964 4146 1992 4678
rect 2332 4570 2360 4966
rect 2424 4729 2452 5034
rect 2516 4826 2544 5063
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2410 4720 2466 4729
rect 2410 4655 2466 4664
rect 2240 4542 2360 4570
rect 2412 4548 2464 4554
rect 1858 4111 1914 4120
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2240 4049 2268 4542
rect 2412 4490 2464 4496
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4078 2360 4422
rect 2320 4072 2372 4078
rect 2226 4040 2282 4049
rect 1780 3998 1900 4026
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1872 3618 1900 3998
rect 2320 4014 2372 4020
rect 2226 3975 2282 3984
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2134 3632 2190 3641
rect 1872 3590 2084 3618
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1492 3120 1544 3126
rect 1688 3074 1716 3431
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1492 3062 1544 3068
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1596 3046 1716 3074
rect 1412 2825 1440 2994
rect 1398 2816 1454 2825
rect 1398 2751 1454 2760
rect 1490 2544 1546 2553
rect 1490 2479 1546 2488
rect 1504 2446 1532 2479
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1214 1728 1270 1737
rect 1032 1692 1084 1698
rect 1214 1663 1270 1672
rect 1032 1634 1084 1640
rect 1596 1601 1624 3046
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1688 1766 1716 2858
rect 1872 2530 1900 3130
rect 2056 2938 2084 3590
rect 2332 3602 2360 4014
rect 2134 3567 2190 3576
rect 2320 3596 2372 3602
rect 2148 3534 2176 3567
rect 2320 3538 2372 3544
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2148 3058 2176 3334
rect 2240 3097 2268 3402
rect 2226 3088 2282 3097
rect 2136 3052 2188 3058
rect 2226 3023 2282 3032
rect 2136 2994 2188 3000
rect 2056 2910 2360 2938
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 1872 2502 2084 2530
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 2281 1900 2314
rect 1952 2304 2004 2310
rect 1858 2272 1914 2281
rect 1952 2246 2004 2252
rect 1858 2207 1914 2216
rect 1964 1834 1992 2246
rect 1952 1828 2004 1834
rect 1952 1770 2004 1776
rect 1676 1760 1728 1766
rect 1676 1702 1728 1708
rect 1582 1592 1638 1601
rect 1582 1527 1638 1536
rect 754 1456 810 1465
rect 754 1391 810 1400
rect 2056 542 2084 2502
rect 2332 678 2360 2910
rect 2424 2553 2452 4490
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2410 2544 2466 2553
rect 2410 2479 2466 2488
rect 2410 2408 2466 2417
rect 2410 2343 2412 2352
rect 2464 2343 2466 2352
rect 2412 2314 2464 2320
rect 2516 1222 2544 4150
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 2608 746 2636 5170
rect 2700 4282 2728 5578
rect 2792 5001 2820 5782
rect 2884 5574 2912 6258
rect 3528 6118 3556 6802
rect 3620 6322 3648 7840
rect 3804 6882 3832 9658
rect 3882 9344 3938 9353
rect 3882 9279 3938 9288
rect 3896 8566 3924 9279
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 4080 8498 4108 8978
rect 4172 8634 4200 11206
rect 4986 11194 5042 11250
rect 6090 11194 6146 11250
rect 7194 11194 7250 11250
rect 8298 11194 8354 11250
rect 9402 11194 9458 11250
rect 10506 11194 10562 11250
rect 11610 11194 11666 11250
rect 12714 11194 12770 11250
rect 13818 11194 13874 11250
rect 14922 11194 14978 11250
rect 16026 11194 16082 11250
rect 17130 11194 17186 11250
rect 18234 11194 18290 11250
rect 19338 11194 19394 11250
rect 20442 11194 20498 11250
rect 21546 11194 21602 11250
rect 22650 11194 22706 11250
rect 23754 11194 23810 11250
rect 24858 11194 24914 11250
rect 25962 11194 26018 11250
rect 27066 11194 27122 11250
rect 27172 11206 27384 11234
rect 4252 9308 4304 9314
rect 4252 9250 4304 9256
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4264 8566 4292 9250
rect 4618 9208 4674 9217
rect 4618 9143 4674 9152
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4434 8664 4490 8673
rect 4434 8599 4490 8608
rect 4448 8566 4476 8599
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3804 6854 4108 6882
rect 3700 6792 3752 6798
rect 3976 6792 4028 6798
rect 3752 6752 3832 6780
rect 3700 6734 3752 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3146 5944 3202 5953
rect 3146 5879 3202 5888
rect 3160 5846 3188 5879
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3620 5778 3648 6258
rect 3712 6254 3740 6598
rect 3700 6248 3752 6254
rect 3698 6216 3700 6225
rect 3752 6216 3754 6225
rect 3698 6151 3754 6160
rect 3698 6080 3754 6089
rect 3698 6015 3754 6024
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 2976 5642 3004 5714
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 3422 5400 3478 5409
rect 3422 5335 3424 5344
rect 3476 5335 3478 5344
rect 3424 5306 3476 5312
rect 3606 5264 3662 5273
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3516 5228 3568 5234
rect 3606 5199 3608 5208
rect 3516 5170 3568 5176
rect 3660 5199 3662 5208
rect 3608 5170 3660 5176
rect 2778 4992 2834 5001
rect 2778 4927 2834 4936
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2884 3641 2912 5170
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4729 3004 4966
rect 3252 4758 3280 5170
rect 3240 4752 3292 4758
rect 2962 4720 3018 4729
rect 3240 4694 3292 4700
rect 2962 4655 3018 4664
rect 3332 4616 3384 4622
rect 3238 4584 3294 4593
rect 3384 4576 3464 4604
rect 3332 4558 3384 4564
rect 3238 4519 3294 4528
rect 3252 4486 3280 4519
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 2976 3505 3004 4082
rect 3160 3913 3188 4150
rect 3240 3936 3292 3942
rect 3146 3904 3202 3913
rect 3240 3878 3292 3884
rect 3146 3839 3202 3848
rect 3252 3505 3280 3878
rect 2962 3496 3018 3505
rect 2688 3460 2740 3466
rect 2962 3431 3018 3440
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 2688 3402 2740 3408
rect 2700 814 2728 3402
rect 3344 3398 3372 4218
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 3240 2984 3292 2990
rect 3054 2952 3110 2961
rect 3240 2926 3292 2932
rect 3054 2887 3110 2896
rect 2778 2680 2834 2689
rect 2778 2615 2780 2624
rect 2832 2615 2834 2624
rect 2780 2586 2832 2592
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1737 2820 2450
rect 3068 2446 3096 2887
rect 3252 2582 3280 2926
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2778 1728 2834 1737
rect 2778 1663 2834 1672
rect 2688 808 2740 814
rect 2688 750 2740 756
rect 2596 740 2648 746
rect 2596 682 2648 688
rect 2320 672 2372 678
rect 2320 614 2372 620
rect 2044 536 2096 542
rect 2044 478 2096 484
rect 2884 42 2912 2382
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 3436 1358 3464 4576
rect 3528 4282 3556 5170
rect 3712 4842 3740 6015
rect 3620 4814 3740 4842
rect 3620 4690 3648 4814
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3620 4185 3648 4422
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3620 3738 3648 4014
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3712 3618 3740 4694
rect 3528 3590 3740 3618
rect 3528 2530 3556 3590
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3620 3058 3648 3334
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3528 2502 3648 2530
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3160 56 3280 82
rect 3528 56 3556 2382
rect 3620 1290 3648 2502
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 3712 921 3740 3334
rect 3698 912 3754 921
rect 3698 847 3754 856
rect 3804 56 3832 6752
rect 3896 6752 3976 6780
rect 3896 5370 3924 6752
rect 3976 6734 4028 6740
rect 4080 6440 4108 6854
rect 3988 6412 4108 6440
rect 3988 6202 4016 6412
rect 4068 6316 4120 6322
rect 4172 6304 4200 7686
rect 4264 7410 4292 8502
rect 4540 8090 4568 9046
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4632 7886 4660 9143
rect 5000 8498 5028 11194
rect 5632 10872 5684 10878
rect 5632 10814 5684 10820
rect 5538 9888 5594 9897
rect 5538 9823 5594 9832
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5276 8634 5304 8842
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5552 8566 5580 9823
rect 5644 9110 5672 10814
rect 5814 9344 5870 9353
rect 5814 9279 5870 9288
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 4816 8294 4844 8434
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 5276 8090 5304 8434
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4356 7342 4384 7754
rect 4908 7478 4936 7754
rect 4896 7472 4948 7478
rect 4710 7440 4766 7449
rect 4620 7404 4672 7410
rect 4896 7414 4948 7420
rect 4710 7375 4766 7384
rect 4988 7404 5040 7410
rect 4620 7346 4672 7352
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4120 6276 4200 6304
rect 4068 6258 4120 6264
rect 4264 6202 4292 6938
rect 4356 6866 4384 7142
rect 4448 6934 4476 7142
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4540 6780 4568 7210
rect 4448 6752 4568 6780
rect 4448 6254 4476 6752
rect 4632 6440 4660 7346
rect 4724 6798 4752 7375
rect 4988 7346 5040 7352
rect 5000 7041 5028 7346
rect 5080 7200 5132 7206
rect 5276 7177 5304 7822
rect 5368 7818 5396 8026
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5080 7142 5132 7148
rect 5262 7168 5318 7177
rect 4986 7032 5042 7041
rect 4986 6967 5042 6976
rect 4712 6792 4764 6798
rect 4896 6792 4948 6798
rect 4894 6760 4896 6769
rect 4948 6760 4950 6769
rect 4712 6734 4764 6740
rect 4540 6412 4660 6440
rect 3988 6174 4108 6202
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3896 4826 3924 5199
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3896 3194 3924 4626
rect 3988 3534 4016 6054
rect 4080 5914 4108 6174
rect 4172 6174 4292 6202
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3976 3528 4028 3534
rect 3974 3496 3976 3505
rect 4028 3496 4030 3505
rect 3974 3431 4030 3440
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3160 54 3294 56
rect 3160 42 3188 54
rect 2884 14 3188 42
rect 3238 0 3294 54
rect 3514 0 3570 56
rect 3790 0 3846 56
rect 3896 42 3924 2314
rect 3988 1086 4016 2450
rect 3976 1080 4028 1086
rect 3976 1022 4028 1028
rect 4080 218 4108 5510
rect 4172 5098 4200 6174
rect 4344 5228 4396 5234
rect 4264 5188 4344 5216
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4264 4978 4292 5188
rect 4344 5170 4396 5176
rect 4172 4950 4292 4978
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4172 4049 4200 4950
rect 4250 4856 4306 4865
rect 4356 4826 4384 4966
rect 4250 4791 4306 4800
rect 4344 4820 4396 4826
rect 4158 4040 4214 4049
rect 4158 3975 4214 3984
rect 4264 3058 4292 4791
rect 4344 4762 4396 4768
rect 4342 4720 4398 4729
rect 4342 4655 4398 4664
rect 4356 4146 4384 4655
rect 4448 4282 4476 6190
rect 4540 6089 4568 6412
rect 4620 6316 4672 6322
rect 4724 6304 4752 6734
rect 4816 6718 4894 6746
rect 4816 6322 4844 6718
rect 4894 6695 4950 6704
rect 4672 6276 4752 6304
rect 4804 6316 4856 6322
rect 4620 6258 4672 6264
rect 4804 6258 4856 6264
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4526 6080 4582 6089
rect 4526 6015 4582 6024
rect 4908 5914 4936 6190
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4988 5704 5040 5710
rect 4986 5672 4988 5681
rect 5040 5672 5042 5681
rect 4986 5607 5042 5616
rect 5092 5574 5120 7142
rect 5262 7103 5318 7112
rect 5354 6624 5410 6633
rect 5354 6559 5410 6568
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5080 5568 5132 5574
rect 4986 5536 5042 5545
rect 5080 5510 5132 5516
rect 4986 5471 5042 5480
rect 4710 5400 4766 5409
rect 4894 5400 4950 5409
rect 4710 5335 4766 5344
rect 4804 5364 4856 5370
rect 4528 5228 4580 5234
rect 4580 5188 4660 5216
rect 4528 5170 4580 5176
rect 4526 4720 4582 4729
rect 4526 4655 4528 4664
rect 4580 4655 4582 4664
rect 4528 4626 4580 4632
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3126 4476 3334
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4264 2961 4292 2994
rect 4250 2952 4306 2961
rect 4250 2887 4306 2896
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4172 1902 4200 2314
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4160 1896 4212 1902
rect 4160 1838 4212 1844
rect 4264 1630 4292 2246
rect 4356 2009 4384 2586
rect 4342 2000 4398 2009
rect 4342 1935 4398 1944
rect 4252 1624 4304 1630
rect 4252 1566 4304 1572
rect 4632 1442 4660 5188
rect 4724 4622 4752 5335
rect 4894 5335 4950 5344
rect 4804 5306 4856 5312
rect 4816 5234 4844 5306
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4908 5030 4936 5335
rect 5000 5148 5028 5471
rect 5092 5302 5120 5510
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5080 5160 5132 5166
rect 5000 5120 5080 5148
rect 5172 5160 5224 5166
rect 5080 5102 5132 5108
rect 5170 5128 5172 5137
rect 5276 5148 5304 5646
rect 5224 5128 5304 5148
rect 5226 5120 5304 5128
rect 5170 5063 5226 5072
rect 4896 5024 4948 5030
rect 5172 5024 5224 5030
rect 4896 4966 4948 4972
rect 5078 4992 5134 5001
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4486 4752 4558
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 4060 4752 4422
rect 4804 4072 4856 4078
rect 4724 4032 4804 4060
rect 4804 4014 4856 4020
rect 4908 3720 4936 4966
rect 5172 4966 5224 4972
rect 5078 4927 5134 4936
rect 5092 4690 5120 4927
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 4724 3692 4936 3720
rect 4724 3398 4752 3692
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4724 2122 4752 2858
rect 4816 2514 4844 3470
rect 4908 3058 4936 3538
rect 5000 3194 5028 4626
rect 5092 4078 5120 4626
rect 5184 4321 5212 4966
rect 5276 4457 5304 5120
rect 5262 4448 5318 4457
rect 5262 4383 5318 4392
rect 5170 4312 5226 4321
rect 5368 4298 5396 6559
rect 5460 5234 5488 8502
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8242 5764 8366
rect 5644 8214 5764 8242
rect 5644 7410 5672 8214
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 6746 5672 7346
rect 5736 6866 5764 7822
rect 5828 7478 5856 9279
rect 6104 8634 6132 11194
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5906 8256 5962 8265
rect 5906 8191 5962 8200
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5644 6718 5764 6746
rect 5632 6656 5684 6662
rect 5736 6633 5764 6718
rect 5632 6598 5684 6604
rect 5722 6624 5778 6633
rect 5644 6322 5672 6598
rect 5722 6559 5778 6568
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5814 6080 5870 6089
rect 5814 6015 5870 6024
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5170 4247 5226 4256
rect 5276 4270 5396 4298
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5276 3534 5304 4270
rect 5460 4078 5488 4966
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5552 3777 5580 5510
rect 5644 4865 5672 5646
rect 5722 5536 5778 5545
rect 5722 5471 5778 5480
rect 5736 5234 5764 5471
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5630 4856 5686 4865
rect 5630 4791 5686 4800
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4282 5672 4558
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5736 4146 5764 5170
rect 5828 4554 5856 6015
rect 5920 5778 5948 8191
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 5920 4622 5948 5578
rect 6012 5545 6040 8570
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6104 5914 6132 6326
rect 6196 6118 6224 10406
rect 6366 9752 6422 9761
rect 6366 9687 6422 9696
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 7818 6316 9522
rect 6380 7954 6408 9687
rect 6644 9240 6696 9246
rect 6644 9182 6696 9188
rect 6458 8528 6514 8537
rect 6656 8498 6684 9182
rect 7208 8634 7236 11194
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7286 10160 7342 10169
rect 7286 10095 7342 10104
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 6458 8463 6514 8472
rect 6644 8492 6696 8498
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6366 6896 6422 6905
rect 6366 6831 6368 6840
rect 6420 6831 6422 6840
rect 6368 6802 6420 6808
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5998 5536 6054 5545
rect 5998 5471 6054 5480
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6012 4865 6040 5238
rect 6104 5166 6132 5306
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 5998 4856 6054 4865
rect 5998 4791 6054 4800
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5724 4140 5776 4146
rect 5644 4100 5724 4128
rect 5538 3768 5594 3777
rect 5538 3703 5594 3712
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 4896 2372 4948 2378
rect 4896 2314 4948 2320
rect 4724 2094 4844 2122
rect 4632 1414 4752 1442
rect 4724 1358 4752 1414
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 4080 190 4200 218
rect 3988 56 4108 82
rect 3988 54 4122 56
rect 3988 42 4016 54
rect 3896 14 4016 42
rect 4066 0 4122 54
rect 4172 42 4200 190
rect 4264 56 4384 82
rect 4632 56 4660 1294
rect 4816 1057 4844 2094
rect 4908 1222 4936 2314
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 5000 2038 5028 2246
rect 4988 2032 5040 2038
rect 4988 1974 5040 1980
rect 4896 1216 4948 1222
rect 4896 1158 4948 1164
rect 4802 1048 4858 1057
rect 4802 983 4858 992
rect 4896 740 4948 746
rect 4896 682 4948 688
rect 4908 56 4936 682
rect 5276 474 5304 2450
rect 5264 468 5316 474
rect 5264 410 5316 416
rect 5184 56 5304 82
rect 4264 54 4398 56
rect 4264 42 4292 54
rect 4172 14 4292 42
rect 4342 0 4398 54
rect 4618 0 4674 56
rect 4894 0 4950 56
rect 5170 54 5304 56
rect 5170 0 5226 54
rect 5276 42 5304 54
rect 5368 42 5396 3567
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5446 3088 5502 3097
rect 5446 3023 5448 3032
rect 5500 3023 5502 3032
rect 5448 2994 5500 3000
rect 5446 1320 5502 1329
rect 5446 1255 5502 1264
rect 5460 56 5488 1255
rect 5552 649 5580 3334
rect 5644 2310 5672 4100
rect 5724 4082 5776 4088
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5538 640 5594 649
rect 5538 575 5594 584
rect 5736 56 5764 2994
rect 5828 2990 5856 4490
rect 6104 3942 6132 5102
rect 6196 4214 6224 5170
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6184 4208 6236 4214
rect 6184 4150 6236 4156
rect 6182 4040 6238 4049
rect 6182 3975 6238 3984
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 5906 3496 5962 3505
rect 5906 3431 5962 3440
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5920 2446 5948 3431
rect 6104 2922 6132 3878
rect 6196 3602 6224 3975
rect 6288 3602 6316 4966
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6092 2916 6144 2922
rect 6092 2858 6144 2864
rect 6196 2514 6224 3062
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 5920 338 5948 2382
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 5908 332 5960 338
rect 5908 274 5960 280
rect 6012 56 6040 1226
rect 6288 56 6316 2382
rect 6380 950 6408 6122
rect 6472 5953 6500 8463
rect 6644 8434 6696 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6642 7304 6698 7313
rect 6642 7239 6698 7248
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6866 6592 7142
rect 6656 6866 6684 7239
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6564 6118 6592 6598
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6458 5944 6514 5953
rect 6458 5879 6514 5888
rect 6564 5574 6592 6054
rect 6656 5681 6684 6190
rect 6642 5672 6698 5681
rect 6642 5607 6698 5616
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5234 6592 5510
rect 6748 5352 6776 6258
rect 6656 5324 6776 5352
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6460 4140 6512 4146
rect 6512 4100 6592 4128
rect 6460 4082 6512 4088
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6472 3602 6500 3878
rect 6564 3670 6592 4100
rect 6656 3720 6684 5324
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 4185 6776 5170
rect 6734 4176 6790 4185
rect 6734 4111 6790 4120
rect 6840 3738 6868 8434
rect 7196 8424 7248 8430
rect 7194 8392 7196 8401
rect 7248 8392 7250 8401
rect 7194 8327 7250 8336
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 6866 6960 7958
rect 7208 7954 7236 8327
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7010 7168 7066 7177
rect 7010 7103 7066 7112
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 7024 5681 7052 7103
rect 7208 7041 7236 7686
rect 7194 7032 7250 7041
rect 7194 6967 7250 6976
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7208 6322 7236 6394
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7116 5914 7144 6258
rect 7300 6118 7328 10095
rect 7380 9784 7432 9790
rect 7380 9726 7432 9732
rect 7392 7478 7420 9726
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8634 7512 8774
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7484 8498 7512 8570
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7392 6254 7420 6870
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7010 5672 7066 5681
rect 7010 5607 7066 5616
rect 6918 5536 6974 5545
rect 6918 5471 6974 5480
rect 6932 5302 6960 5471
rect 7208 5409 7236 5850
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7300 5574 7328 5646
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7194 5400 7250 5409
rect 7194 5335 7250 5344
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 4622 6960 5238
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7010 5128 7066 5137
rect 7010 5063 7012 5072
rect 7064 5063 7066 5072
rect 7104 5092 7156 5098
rect 7012 5034 7064 5040
rect 7104 5034 7156 5040
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 3732 6880 3738
rect 6656 3692 6776 3720
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6642 3632 6698 3641
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6564 3534 6592 3606
rect 6642 3567 6698 3576
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 2582 6500 3334
rect 6656 3058 6684 3567
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6564 2650 6592 2858
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6368 944 6420 950
rect 6368 886 6420 892
rect 6564 56 6592 2314
rect 6748 2310 6776 3692
rect 6828 3674 6880 3680
rect 6932 3618 6960 4558
rect 6840 3590 6960 3618
rect 6840 3398 6868 3590
rect 6920 3528 6972 3534
rect 7024 3516 7052 4626
rect 7116 4554 7144 5034
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4282 7144 4490
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6972 3488 7052 3516
rect 7116 3505 7144 4014
rect 7102 3496 7158 3505
rect 6920 3470 6972 3476
rect 7024 3440 7102 3448
rect 7024 3431 7158 3440
rect 7024 3420 7144 3431
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 7024 2514 7052 3420
rect 7102 2816 7158 2825
rect 7102 2751 7158 2760
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6828 1148 6880 1154
rect 6828 1090 6880 1096
rect 6840 56 6868 1090
rect 7116 56 7144 2751
rect 7208 1426 7236 5170
rect 7300 4826 7328 5510
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7392 4706 7420 6190
rect 7484 6089 7512 7278
rect 7576 6905 7604 7278
rect 7562 6896 7618 6905
rect 7562 6831 7564 6840
rect 7616 6831 7618 6840
rect 7564 6802 7616 6808
rect 7668 6474 7696 10678
rect 8312 8634 8340 11194
rect 9312 10396 9364 10402
rect 9312 10338 9364 10344
rect 8850 10024 8906 10033
rect 8850 9959 8906 9968
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8673 8432 8774
rect 8390 8664 8446 8673
rect 8300 8628 8352 8634
rect 8390 8599 8446 8608
rect 8300 8570 8352 8576
rect 8390 8392 8446 8401
rect 8496 8378 8524 9114
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8588 8566 8616 9046
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8496 8350 8616 8378
rect 8390 8327 8446 8336
rect 8404 8294 8432 8327
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7576 6446 7696 6474
rect 7470 6080 7526 6089
rect 7470 6015 7526 6024
rect 7576 5930 7604 6446
rect 7654 6352 7710 6361
rect 7654 6287 7656 6296
rect 7708 6287 7710 6296
rect 7656 6258 7708 6264
rect 7576 5902 7696 5930
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7484 5166 7512 5714
rect 7576 5370 7604 5714
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7300 4678 7420 4706
rect 7484 4690 7512 5102
rect 7668 5030 7696 5902
rect 7760 5370 7788 7278
rect 7852 6780 7880 7822
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7342 8248 7686
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 8024 6792 8076 6798
rect 7852 6752 8024 6780
rect 8024 6734 8076 6740
rect 8036 6497 8064 6734
rect 8022 6488 8078 6497
rect 8022 6423 8078 6432
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 7760 5166 7788 5306
rect 7748 5160 7800 5166
rect 7852 5148 7880 6054
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8220 5710 8248 5850
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7932 5160 7984 5166
rect 7852 5120 7932 5148
rect 7748 5102 7800 5108
rect 7932 5102 7984 5108
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 7656 5024 7708 5030
rect 7944 5012 7972 5102
rect 7656 4966 7708 4972
rect 7760 4984 7972 5012
rect 8128 5012 8156 5102
rect 8312 5080 8340 8230
rect 8588 8022 8616 8350
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8496 7410 8524 7822
rect 8588 7818 8616 7958
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8496 7313 8524 7346
rect 8482 7304 8538 7313
rect 8482 7239 8538 7248
rect 8574 7032 8630 7041
rect 8574 6967 8630 6976
rect 8588 6322 8616 6967
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8588 6089 8616 6258
rect 8574 6080 8630 6089
rect 8574 6015 8630 6024
rect 8588 5846 8616 6015
rect 8680 5914 8708 9454
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8772 7410 8800 8298
rect 8864 8022 8892 9959
rect 9324 8945 9352 10338
rect 9310 8936 9366 8945
rect 9310 8871 9366 8880
rect 9010 8732 9318 8741
rect 9010 8730 9016 8732
rect 9072 8730 9096 8732
rect 9152 8730 9176 8732
rect 9232 8730 9256 8732
rect 9312 8730 9318 8732
rect 9072 8678 9074 8730
rect 9254 8678 9256 8730
rect 9010 8676 9016 8678
rect 9072 8676 9096 8678
rect 9152 8676 9176 8678
rect 9232 8676 9256 8678
rect 9312 8676 9318 8678
rect 9010 8667 9318 8676
rect 9416 8634 9444 11194
rect 9954 10568 10010 10577
rect 9772 10532 9824 10538
rect 9954 10503 10010 10512
rect 9772 10474 9824 10480
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9496 9308 9548 9314
rect 9496 9250 9548 9256
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 8852 8016 8904 8022
rect 9508 7993 9536 9250
rect 9600 8498 9628 10134
rect 9680 9852 9732 9858
rect 9680 9794 9732 9800
rect 9692 9625 9720 9794
rect 9678 9616 9734 9625
rect 9678 9551 9734 9560
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9692 8362 9720 8502
rect 9784 8498 9812 10474
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 8852 7958 8904 7964
rect 9494 7984 9550 7993
rect 9494 7919 9550 7928
rect 9692 7886 9720 8298
rect 9588 7880 9640 7886
rect 9494 7848 9550 7857
rect 9588 7822 9640 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9494 7783 9496 7792
rect 9548 7783 9550 7792
rect 9496 7754 9548 7760
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8864 6798 8892 7686
rect 9010 7644 9318 7653
rect 9010 7642 9016 7644
rect 9072 7642 9096 7644
rect 9152 7642 9176 7644
rect 9232 7642 9256 7644
rect 9312 7642 9318 7644
rect 9072 7590 9074 7642
rect 9254 7590 9256 7642
rect 9010 7588 9016 7590
rect 9072 7588 9096 7590
rect 9152 7588 9176 7590
rect 9232 7588 9256 7590
rect 9312 7588 9318 7590
rect 9010 7579 9318 7588
rect 9508 6798 9536 7754
rect 9600 7342 9628 7822
rect 9784 7546 9812 7822
rect 9968 7546 9996 10503
rect 10322 10432 10378 10441
rect 10322 10367 10378 10376
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7585 10180 7754
rect 10138 7576 10194 7585
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9956 7540 10008 7546
rect 10138 7511 10194 7520
rect 9956 7482 10008 7488
rect 9770 7440 9826 7449
rect 9770 7375 9826 7384
rect 10048 7404 10100 7410
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 7041 9720 7142
rect 9678 7032 9734 7041
rect 9678 6967 9734 6976
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8484 5704 8536 5710
rect 8576 5704 8628 5710
rect 8484 5646 8536 5652
rect 8574 5672 8576 5681
rect 8628 5672 8630 5681
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8404 5234 8432 5510
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8312 5052 8457 5080
rect 8128 4984 8340 5012
rect 7654 4856 7710 4865
rect 7654 4791 7710 4800
rect 7472 4684 7524 4690
rect 7300 3924 7328 4678
rect 7472 4626 7524 4632
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7576 4486 7604 4626
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7392 4049 7420 4218
rect 7668 4146 7696 4791
rect 7760 4604 7788 4984
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7840 4616 7892 4622
rect 7760 4576 7840 4604
rect 7840 4558 7892 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7746 4312 7802 4321
rect 7746 4247 7802 4256
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 4049 7696 4082
rect 7378 4040 7434 4049
rect 7654 4040 7710 4049
rect 7378 3975 7434 3984
rect 7564 4004 7616 4010
rect 7654 3975 7710 3984
rect 7564 3946 7616 3952
rect 7472 3936 7524 3942
rect 7300 3896 7472 3924
rect 7472 3878 7524 3884
rect 7378 3768 7434 3777
rect 7378 3703 7380 3712
rect 7432 3703 7434 3712
rect 7380 3674 7432 3680
rect 7392 3602 7420 3674
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7300 2281 7328 3130
rect 7392 2582 7420 3334
rect 7484 3194 7512 3878
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7286 2272 7342 2281
rect 7286 2207 7342 2216
rect 7196 1420 7248 1426
rect 7196 1362 7248 1368
rect 7378 1184 7434 1193
rect 7378 1119 7434 1128
rect 7392 56 7420 1119
rect 7484 882 7512 2994
rect 7576 2514 7604 3946
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 7472 876 7524 882
rect 7472 818 7524 824
rect 7668 56 7696 1294
rect 7760 1154 7788 4247
rect 8024 3936 8076 3942
rect 8128 3924 8156 4558
rect 8076 3896 8156 3924
rect 8220 3924 8248 4762
rect 8312 4690 8340 4984
rect 8429 4842 8457 5052
rect 8404 4814 8457 4842
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8220 3896 8340 3924
rect 8024 3878 8076 3884
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7932 3732 7984 3738
rect 8312 3720 8340 3896
rect 8404 3738 8432 4814
rect 7932 3674 7984 3680
rect 8220 3692 8340 3720
rect 8392 3732 8444 3738
rect 7944 2836 7972 3674
rect 8220 3398 8248 3692
rect 8392 3674 8444 3680
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8208 3392 8260 3398
rect 8022 3360 8078 3369
rect 8312 3369 8340 3470
rect 8208 3334 8260 3340
rect 8298 3360 8354 3369
rect 8022 3295 8078 3304
rect 8298 3295 8354 3304
rect 8036 3058 8064 3295
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 7852 2808 7972 2836
rect 7852 2650 7880 2808
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7748 1148 7800 1154
rect 7748 1090 7800 1096
rect 7944 56 7972 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 56 8248 2246
rect 8312 1018 8340 2994
rect 8404 2582 8432 3470
rect 8496 2774 8524 5646
rect 8574 5607 8630 5616
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5409 8708 5510
rect 8666 5400 8722 5409
rect 8666 5335 8722 5344
rect 8772 4808 8800 6190
rect 8864 5710 8892 6734
rect 9678 6624 9734 6633
rect 9010 6556 9318 6565
rect 9678 6559 9734 6568
rect 9010 6554 9016 6556
rect 9072 6554 9096 6556
rect 9152 6554 9176 6556
rect 9232 6554 9256 6556
rect 9312 6554 9318 6556
rect 9072 6502 9074 6554
rect 9254 6502 9256 6554
rect 9010 6500 9016 6502
rect 9072 6500 9096 6502
rect 9152 6500 9176 6502
rect 9232 6500 9256 6502
rect 9312 6500 9318 6502
rect 9010 6491 9318 6500
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9140 6254 9168 6394
rect 9692 6338 9720 6559
rect 9600 6322 9720 6338
rect 9588 6316 9720 6322
rect 9508 6276 9588 6304
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8956 5522 8984 6122
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 8864 5494 8984 5522
rect 8864 5250 8892 5494
rect 9010 5468 9318 5477
rect 9010 5466 9016 5468
rect 9072 5466 9096 5468
rect 9152 5466 9176 5468
rect 9232 5466 9256 5468
rect 9312 5466 9318 5468
rect 9072 5414 9074 5466
rect 9254 5414 9256 5466
rect 9010 5412 9016 5414
rect 9072 5412 9096 5414
rect 9152 5412 9176 5414
rect 9232 5412 9256 5414
rect 9312 5412 9318 5414
rect 9010 5403 9318 5412
rect 9416 5370 9444 5714
rect 9508 5710 9536 6276
rect 9640 6310 9720 6316
rect 9588 6258 9640 6264
rect 9680 6248 9732 6254
rect 9600 6196 9680 6202
rect 9600 6190 9732 6196
rect 9600 6174 9720 6190
rect 9600 6118 9628 6174
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5574 9536 5646
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9312 5296 9364 5302
rect 8864 5222 9260 5250
rect 9312 5238 9364 5244
rect 8944 5160 8996 5166
rect 9128 5160 9180 5166
rect 8996 5120 9076 5148
rect 8944 5102 8996 5108
rect 9048 5030 9076 5120
rect 9128 5102 9180 5108
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8588 4780 8800 4808
rect 9036 4820 9088 4826
rect 8588 3398 8616 4780
rect 9036 4762 9088 4768
rect 9048 4690 9076 4762
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 8680 3670 8708 4626
rect 8760 4616 8812 4622
rect 9140 4570 9168 5102
rect 8760 4558 8812 4564
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8772 3602 8800 4558
rect 8956 4542 9168 4570
rect 8956 4434 8984 4542
rect 9232 4536 9260 5222
rect 9324 5166 9352 5238
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9232 4508 9444 4536
rect 8864 4406 8984 4434
rect 8864 4298 8892 4406
rect 9010 4380 9318 4389
rect 9010 4378 9016 4380
rect 9072 4378 9096 4380
rect 9152 4378 9176 4380
rect 9232 4378 9256 4380
rect 9312 4378 9318 4380
rect 9072 4326 9074 4378
rect 9254 4326 9256 4378
rect 9010 4324 9016 4326
rect 9072 4324 9096 4326
rect 9152 4324 9176 4326
rect 9232 4324 9256 4326
rect 9312 4324 9318 4326
rect 9010 4315 9318 4324
rect 8864 4270 8984 4298
rect 8956 4078 8984 4270
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8864 3913 8892 3946
rect 8850 3904 8906 3913
rect 8850 3839 8906 3848
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8864 3534 8892 3674
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8576 3392 8628 3398
rect 8956 3346 8984 3606
rect 9048 3466 9076 4218
rect 9128 4208 9180 4214
rect 9416 4162 9444 4508
rect 9128 4150 9180 4156
rect 9140 3913 9168 4150
rect 9324 4134 9444 4162
rect 9508 4146 9536 5102
rect 9600 5030 9628 6054
rect 9784 5817 9812 7375
rect 10048 7346 10100 7352
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9876 6254 9904 6598
rect 9968 6458 9996 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9770 5808 9826 5817
rect 9680 5772 9732 5778
rect 9770 5743 9826 5752
rect 9680 5714 9732 5720
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9692 4706 9720 5714
rect 9772 5704 9824 5710
rect 9770 5672 9772 5681
rect 9824 5672 9826 5681
rect 9770 5607 9826 5616
rect 9784 5001 9812 5607
rect 9770 4992 9826 5001
rect 9770 4927 9826 4936
rect 9692 4678 9812 4706
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4457 9628 4558
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9586 4448 9642 4457
rect 9586 4383 9642 4392
rect 9496 4140 9548 4146
rect 9126 3904 9182 3913
rect 9126 3839 9182 3848
rect 9324 3738 9352 4134
rect 9496 4082 9548 4088
rect 9692 4078 9720 4490
rect 9784 4128 9812 4678
rect 9876 4622 9904 6190
rect 9968 5778 9996 6394
rect 10060 6361 10088 7346
rect 10244 6644 10272 8978
rect 10336 8022 10364 10367
rect 10520 8634 10548 11194
rect 10876 9240 10928 9246
rect 10876 9182 10928 9188
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10690 8120 10746 8129
rect 10690 8055 10746 8064
rect 10784 8084 10836 8090
rect 10704 8022 10732 8055
rect 10784 8026 10836 8032
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10428 7206 10456 7890
rect 10796 7886 10824 8026
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7721 10824 7822
rect 10782 7712 10838 7721
rect 10782 7647 10838 7656
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10782 6760 10838 6769
rect 10324 6656 10376 6662
rect 10244 6616 10324 6644
rect 10324 6598 10376 6604
rect 10520 6440 10548 6734
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10692 6724 10744 6730
rect 10782 6695 10784 6704
rect 10692 6666 10744 6672
rect 10836 6695 10838 6704
rect 10784 6666 10836 6672
rect 10152 6412 10548 6440
rect 10046 6352 10102 6361
rect 10046 6287 10102 6296
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5098 9996 5714
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9954 4992 10010 5001
rect 9954 4927 10010 4936
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9968 4282 9996 4927
rect 10060 4622 10088 6054
rect 10152 5846 10180 6412
rect 10612 6322 10640 6666
rect 10704 6458 10732 6666
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10230 6080 10286 6089
rect 10230 6015 10286 6024
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 4622 10180 5510
rect 10244 5234 10272 6015
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10048 4616 10100 4622
rect 10140 4616 10192 4622
rect 10048 4558 10100 4564
rect 10138 4584 10140 4593
rect 10192 4584 10194 4593
rect 10138 4519 10194 4528
rect 10046 4312 10102 4321
rect 9956 4276 10008 4282
rect 10046 4247 10102 4256
rect 9956 4218 10008 4224
rect 9784 4100 9996 4128
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9416 3641 9444 4014
rect 9692 3670 9720 4014
rect 9680 3664 9732 3670
rect 9402 3632 9458 3641
rect 9220 3596 9272 3602
rect 9272 3556 9352 3584
rect 9680 3606 9732 3612
rect 9402 3567 9458 3576
rect 9588 3596 9640 3602
rect 9220 3538 9272 3544
rect 9324 3516 9352 3556
rect 9588 3538 9640 3544
rect 9324 3488 9536 3516
rect 9036 3460 9088 3466
rect 9036 3402 9088 3408
rect 8576 3334 8628 3340
rect 8588 3233 8616 3334
rect 8680 3318 8984 3346
rect 8574 3224 8630 3233
rect 8574 3159 8630 3168
rect 8496 2746 8616 2774
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8496 1562 8524 2382
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8482 1320 8538 1329
rect 8482 1255 8538 1264
rect 8300 1012 8352 1018
rect 8300 954 8352 960
rect 8496 56 8524 1255
rect 8588 270 8616 2746
rect 8680 2378 8708 3318
rect 9010 3292 9318 3301
rect 9010 3290 9016 3292
rect 9072 3290 9096 3292
rect 9152 3290 9176 3292
rect 9232 3290 9256 3292
rect 9312 3290 9318 3292
rect 9072 3238 9074 3290
rect 9254 3238 9256 3290
rect 9010 3236 9016 3238
rect 9072 3236 9096 3238
rect 9152 3236 9176 3238
rect 9232 3236 9256 3238
rect 9312 3236 9318 3238
rect 8758 3224 8814 3233
rect 9010 3227 9318 3236
rect 9508 3210 9536 3488
rect 9600 3398 9628 3538
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9508 3182 9628 3210
rect 8758 3159 8814 3168
rect 8772 2854 8800 3159
rect 9600 3058 9628 3182
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2514 8800 2790
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 8772 1698 8800 2314
rect 8760 1692 8812 1698
rect 8760 1634 8812 1640
rect 8864 1358 8892 2994
rect 9048 2378 9076 2994
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9140 2825 9168 2926
rect 9692 2854 9720 3470
rect 9772 3392 9824 3398
rect 9770 3360 9772 3369
rect 9824 3360 9826 3369
rect 9770 3295 9826 3304
rect 9968 3210 9996 4100
rect 10060 3534 10088 4247
rect 10244 4128 10272 5170
rect 10336 4826 10364 6258
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5914 10548 6054
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10704 5794 10732 6122
rect 10520 5778 10732 5794
rect 10508 5772 10732 5778
rect 10560 5766 10732 5772
rect 10508 5714 10560 5720
rect 10784 5704 10836 5710
rect 10704 5664 10784 5692
rect 10704 5166 10732 5664
rect 10784 5646 10836 5652
rect 10416 5160 10468 5166
rect 10692 5160 10744 5166
rect 10468 5120 10548 5148
rect 10416 5102 10468 5108
rect 10414 4992 10470 5001
rect 10414 4927 10470 4936
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4282 10364 4558
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10324 4140 10376 4146
rect 10244 4100 10324 4128
rect 10244 3602 10272 4100
rect 10324 4082 10376 4088
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10048 3528 10100 3534
rect 10046 3496 10048 3505
rect 10100 3496 10102 3505
rect 10046 3431 10102 3440
rect 9968 3194 10364 3210
rect 9968 3188 10376 3194
rect 9968 3182 10324 3188
rect 10324 3130 10376 3136
rect 10048 3120 10100 3126
rect 10048 3062 10100 3068
rect 10322 3088 10378 3097
rect 9220 2848 9272 2854
rect 9126 2816 9182 2825
rect 9220 2790 9272 2796
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9126 2751 9182 2760
rect 9232 2446 9260 2790
rect 9600 2666 9628 2790
rect 10060 2666 10088 3062
rect 10322 3023 10324 3032
rect 10376 3023 10378 3032
rect 10324 2994 10376 3000
rect 10428 2774 10456 4927
rect 10520 4146 10548 5120
rect 10692 5102 10744 5108
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10796 4078 10824 4422
rect 10888 4185 10916 9182
rect 11242 8936 11298 8945
rect 11242 8871 11298 8880
rect 11256 8566 11284 8871
rect 11624 8634 11652 11194
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11072 7546 11100 8434
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11072 7342 11100 7482
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6798 11008 7142
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6662 11008 6734
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10980 5030 11008 6326
rect 11072 6186 11100 6938
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5098 11100 6122
rect 11164 5409 11192 8502
rect 11334 8392 11390 8401
rect 11334 8327 11390 8336
rect 11348 7886 11376 8327
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11336 7880 11388 7886
rect 11256 7840 11336 7868
rect 11256 6798 11284 7840
rect 11336 7822 11388 7828
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11348 5846 11376 7142
rect 11440 6458 11468 8230
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11518 7712 11574 7721
rect 11518 7647 11574 7656
rect 11532 7410 11560 7647
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11440 5914 11468 6258
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11336 5840 11388 5846
rect 11532 5794 11560 6598
rect 11336 5782 11388 5788
rect 11150 5400 11206 5409
rect 11150 5335 11206 5344
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 11072 4622 11100 5034
rect 11256 4865 11284 5782
rect 11440 5766 11560 5794
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11242 4856 11298 4865
rect 11348 4826 11376 5578
rect 11242 4791 11298 4800
rect 11336 4820 11388 4826
rect 11256 4622 11284 4791
rect 11336 4762 11388 4768
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 10874 4176 10930 4185
rect 10874 4111 10930 4120
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10612 3942 10640 4014
rect 11348 3942 11376 4558
rect 11440 4486 11468 5766
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11532 5370 11560 5646
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11532 4321 11560 5306
rect 11518 4312 11574 4321
rect 11518 4247 11574 4256
rect 11624 4214 11652 6734
rect 11716 5681 11744 7890
rect 11888 7880 11940 7886
rect 11886 7848 11888 7857
rect 11940 7848 11942 7857
rect 11886 7783 11942 7792
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 7546 12020 7686
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11808 7410 11836 7482
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11808 5778 11836 5850
rect 11900 5778 11928 6598
rect 12084 6322 12112 9318
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11702 5672 11758 5681
rect 11702 5607 11758 5616
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 10598 3632 10654 3641
rect 11072 3602 11100 3878
rect 10598 3567 10654 3576
rect 11060 3596 11112 3602
rect 10612 3058 10640 3567
rect 11060 3538 11112 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 11334 3496 11390 3505
rect 10888 3194 10916 3470
rect 11334 3431 11390 3440
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10612 2961 10640 2994
rect 10598 2952 10654 2961
rect 10598 2887 10654 2896
rect 9600 2638 10088 2666
rect 10152 2746 10456 2774
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9010 2204 9318 2213
rect 9010 2202 9016 2204
rect 9072 2202 9096 2204
rect 9152 2202 9176 2204
rect 9232 2202 9256 2204
rect 9312 2202 9318 2204
rect 9072 2150 9074 2202
rect 9254 2150 9256 2202
rect 9010 2148 9016 2150
rect 9072 2148 9096 2150
rect 9152 2148 9176 2150
rect 9232 2148 9256 2150
rect 9312 2148 9318 2150
rect 9010 2139 9318 2148
rect 9220 1420 9272 1426
rect 9220 1362 9272 1368
rect 8852 1352 8904 1358
rect 8852 1294 8904 1300
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8576 264 8628 270
rect 8576 206 8628 212
rect 8772 56 8800 1158
rect 9232 950 9260 1362
rect 9416 1204 9444 2382
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 9508 1222 9536 2314
rect 9586 2136 9642 2145
rect 9586 2071 9642 2080
rect 9324 1176 9444 1204
rect 9496 1216 9548 1222
rect 9220 944 9272 950
rect 9220 886 9272 892
rect 9036 876 9088 882
rect 9036 818 9088 824
rect 9048 56 9076 818
rect 9324 56 9352 1176
rect 9496 1158 9548 1164
rect 9600 56 9628 2071
rect 10152 1902 10180 2746
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11072 2009 11100 2382
rect 11058 2000 11114 2009
rect 11058 1935 11114 1944
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 10416 1896 10468 1902
rect 10416 1838 10468 1844
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 9678 1456 9734 1465
rect 9678 1391 9734 1400
rect 9692 610 9720 1391
rect 9680 604 9732 610
rect 9680 546 9732 552
rect 9876 56 9904 1770
rect 10140 1352 10192 1358
rect 10140 1294 10192 1300
rect 10152 56 10180 1294
rect 10428 56 10456 1838
rect 11058 1592 11114 1601
rect 11058 1527 11114 1536
rect 11072 1494 11100 1527
rect 11060 1488 11112 1494
rect 11060 1430 11112 1436
rect 10692 1216 10744 1222
rect 10692 1158 10744 1164
rect 10704 56 10732 1158
rect 10980 56 11100 82
rect 5276 14 5396 42
rect 5446 0 5502 56
rect 5722 0 5778 56
rect 5998 0 6054 56
rect 6274 0 6330 56
rect 6550 0 6606 56
rect 6826 0 6882 56
rect 7102 0 7158 56
rect 7378 0 7434 56
rect 7654 0 7710 56
rect 7930 0 7986 56
rect 8206 0 8262 56
rect 8482 0 8538 56
rect 8758 0 8814 56
rect 9034 0 9090 56
rect 9310 0 9366 56
rect 9586 0 9642 56
rect 9862 0 9918 56
rect 10138 0 10194 56
rect 10414 0 10470 56
rect 10690 0 10746 56
rect 10966 54 11100 56
rect 10966 0 11022 54
rect 11072 42 11100 54
rect 11164 42 11192 2382
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 202 11284 2246
rect 11348 2038 11376 3431
rect 11426 3360 11482 3369
rect 11426 3295 11482 3304
rect 11440 2446 11468 3295
rect 11624 3194 11652 4150
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11426 1864 11482 1873
rect 11426 1799 11482 1808
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11348 1018 11376 1362
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 11440 610 11468 1799
rect 11428 604 11480 610
rect 11428 546 11480 552
rect 11244 196 11296 202
rect 11244 138 11296 144
rect 11072 14 11192 42
rect 11242 96 11298 105
rect 11532 56 11560 2926
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1154 11652 2246
rect 11612 1148 11664 1154
rect 11612 1090 11664 1096
rect 11716 406 11744 5306
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11796 5024 11848 5030
rect 11900 5001 11928 5170
rect 11796 4966 11848 4972
rect 11886 4992 11942 5001
rect 11808 3534 11836 4966
rect 11886 4927 11942 4936
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11900 4486 11928 4694
rect 11992 4672 12020 6258
rect 12084 4865 12112 6258
rect 12070 4856 12126 4865
rect 12070 4791 12126 4800
rect 11992 4644 12112 4672
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11900 3097 11928 4422
rect 11992 4282 12020 4422
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11992 3534 12020 3878
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11886 3088 11942 3097
rect 11886 3023 11942 3032
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11900 1873 11928 2926
rect 11886 1864 11942 1873
rect 11886 1799 11942 1808
rect 12084 1358 12112 4644
rect 12176 4146 12204 6598
rect 12268 6458 12296 10066
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9081 12388 9862
rect 12532 9240 12584 9246
rect 12532 9182 12584 9188
rect 12346 9072 12402 9081
rect 12346 9007 12402 9016
rect 12544 8974 12572 9182
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12530 7984 12586 7993
rect 12452 7954 12530 7970
rect 12440 7948 12530 7954
rect 12492 7942 12530 7948
rect 12636 7954 12664 10610
rect 12728 8634 12756 11194
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 9580 13320 9586
rect 13096 9540 13268 9568
rect 13096 9450 13124 9540
rect 13268 9522 13320 9528
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12530 7919 12586 7928
rect 12624 7948 12676 7954
rect 12440 7890 12492 7896
rect 12624 7890 12676 7896
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12348 7472 12400 7478
rect 12544 7460 12572 7686
rect 12400 7432 12572 7460
rect 12348 7414 12400 7420
rect 12544 6848 12572 7432
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12544 6820 12664 6848
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12530 6760 12586 6769
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12254 6216 12310 6225
rect 12254 6151 12256 6160
rect 12308 6151 12310 6160
rect 12256 6122 12308 6128
rect 12254 5672 12310 5681
rect 12254 5607 12310 5616
rect 12268 5370 12296 5607
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12254 4856 12310 4865
rect 12254 4791 12310 4800
rect 12268 4486 12296 4791
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12254 4176 12310 4185
rect 12164 4140 12216 4146
rect 12254 4111 12310 4120
rect 12164 4082 12216 4088
rect 12162 4040 12218 4049
rect 12162 3975 12218 3984
rect 12176 3670 12204 3975
rect 12268 3670 12296 4111
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12176 1698 12204 2382
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12164 1692 12216 1698
rect 12164 1634 12216 1640
rect 12268 1601 12296 2246
rect 12254 1592 12310 1601
rect 12254 1527 12310 1536
rect 12072 1352 12124 1358
rect 12072 1294 12124 1300
rect 11796 944 11848 950
rect 11796 886 11848 892
rect 11704 400 11756 406
rect 11704 342 11756 348
rect 11808 56 11836 886
rect 12072 468 12124 474
rect 12072 410 12124 416
rect 12084 56 12112 410
rect 12256 264 12308 270
rect 12256 206 12308 212
rect 12268 82 12296 206
rect 12360 184 12388 6734
rect 12530 6695 12586 6704
rect 12544 6662 12572 6695
rect 12532 6656 12584 6662
rect 12438 6624 12494 6633
rect 12532 6598 12584 6604
rect 12438 6559 12494 6568
rect 12452 6458 12480 6559
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12438 6080 12494 6089
rect 12438 6015 12494 6024
rect 12452 5710 12480 6015
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12452 5574 12480 5646
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12452 4865 12480 5306
rect 12544 5030 12572 5646
rect 12636 5370 12664 6820
rect 12728 6361 12756 6870
rect 12820 6662 12848 8842
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 12900 8424 12952 8430
rect 13188 8401 13216 8434
rect 12900 8366 12952 8372
rect 13174 8392 13230 8401
rect 12912 7206 12940 8366
rect 13174 8327 13230 8336
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13004 7290 13032 7822
rect 13096 7546 13124 7822
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13082 7304 13138 7313
rect 13004 7262 13082 7290
rect 13082 7239 13138 7248
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 13096 7002 13124 7239
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 7002 13216 7142
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13280 6882 13308 9386
rect 13096 6854 13308 6882
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12714 6352 12770 6361
rect 12770 6296 12848 6304
rect 12714 6287 12716 6296
rect 12768 6276 12848 6296
rect 12716 6258 12768 6264
rect 12714 5536 12770 5545
rect 12714 5471 12770 5480
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12728 5234 12756 5471
rect 12820 5370 12848 6276
rect 12898 6080 12954 6089
rect 12898 6015 12954 6024
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12452 4486 12480 4558
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12544 4282 12572 4966
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12636 4146 12664 5102
rect 12728 4622 12756 5170
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12452 3398 12480 3606
rect 12636 3534 12664 3878
rect 12728 3738 12756 4082
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12714 3496 12770 3505
rect 12532 3460 12584 3466
rect 12714 3431 12770 3440
rect 12532 3402 12584 3408
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12438 3088 12494 3097
rect 12438 3023 12494 3032
rect 12452 2854 12480 3023
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12544 1834 12572 3402
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 2961 12664 3334
rect 12622 2952 12678 2961
rect 12728 2922 12756 3431
rect 12622 2887 12678 2896
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12532 1828 12584 1834
rect 12532 1770 12584 1776
rect 12636 1630 12664 2382
rect 12624 1624 12676 1630
rect 12624 1566 12676 1572
rect 12820 474 12848 5170
rect 12912 3670 12940 6015
rect 13004 5817 13032 6734
rect 12990 5808 13046 5817
rect 13096 5778 13124 6854
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13280 6361 13308 6734
rect 13266 6352 13322 6361
rect 13266 6287 13322 6296
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12990 5743 13046 5752
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13004 4826 13032 5102
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12912 1902 12940 3470
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 12900 1352 12952 1358
rect 12900 1294 12952 1300
rect 12808 468 12860 474
rect 12808 410 12860 416
rect 12360 156 12480 184
rect 12268 56 12388 82
rect 11242 0 11298 40
rect 11518 0 11574 56
rect 11794 0 11850 56
rect 12070 0 12126 56
rect 12268 54 12402 56
rect 12346 0 12402 54
rect 12452 42 12480 156
rect 12544 56 12664 82
rect 12912 56 12940 1294
rect 13004 1290 13032 2994
rect 13096 1358 13124 5170
rect 13188 4826 13216 6054
rect 13372 5778 13400 10610
rect 13832 8634 13860 11194
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 13910 10296 13966 10305
rect 13910 10231 13966 10240
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13924 8276 13952 10231
rect 14384 8498 14412 10542
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 13832 8248 13952 8276
rect 13542 8120 13598 8129
rect 13832 8106 13860 8248
rect 13950 8188 14258 8197
rect 13950 8186 13956 8188
rect 14012 8186 14036 8188
rect 14092 8186 14116 8188
rect 14172 8186 14196 8188
rect 14252 8186 14258 8188
rect 14012 8134 14014 8186
rect 14194 8134 14196 8186
rect 13950 8132 13956 8134
rect 14012 8132 14036 8134
rect 14092 8132 14116 8134
rect 14172 8132 14196 8134
rect 14252 8132 14258 8134
rect 13950 8123 14258 8132
rect 13598 8078 13860 8106
rect 13542 8055 13598 8064
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13452 6792 13504 6798
rect 13556 6780 13584 7958
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13648 7449 13676 7890
rect 13634 7440 13690 7449
rect 13634 7375 13690 7384
rect 13950 7100 14258 7109
rect 13950 7098 13956 7100
rect 14012 7098 14036 7100
rect 14092 7098 14116 7100
rect 14172 7098 14196 7100
rect 14252 7098 14258 7100
rect 14012 7046 14014 7098
rect 14194 7046 14196 7098
rect 13950 7044 13956 7046
rect 14012 7044 14036 7046
rect 14092 7044 14116 7046
rect 14172 7044 14196 7046
rect 14252 7044 14258 7046
rect 13950 7035 14258 7044
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 13636 6792 13688 6798
rect 13556 6752 13636 6780
rect 13452 6734 13504 6740
rect 13636 6734 13688 6740
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13266 5536 13322 5545
rect 13266 5471 13322 5480
rect 13280 5098 13308 5471
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13372 4593 13400 5102
rect 13358 4584 13414 4593
rect 13358 4519 13360 4528
rect 13412 4519 13414 4528
rect 13360 4490 13412 4496
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13280 4146 13308 4422
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13372 4078 13400 4490
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13268 3936 13320 3942
rect 13174 3904 13230 3913
rect 13268 3878 13320 3884
rect 13174 3839 13230 3848
rect 13188 3641 13216 3839
rect 13174 3632 13230 3641
rect 13280 3602 13308 3878
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 13174 3567 13230 3576
rect 13268 3596 13320 3602
rect 13188 3534 13216 3567
rect 13268 3538 13320 3544
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13280 3126 13308 3402
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13174 2952 13230 2961
rect 13174 2887 13230 2896
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 12992 1284 13044 1290
rect 12992 1226 13044 1232
rect 13188 56 13216 2887
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13280 2650 13308 2790
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13280 2514 13308 2586
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13372 2281 13400 3703
rect 13358 2272 13414 2281
rect 13358 2207 13414 2216
rect 13464 56 13492 6734
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6361 13584 6598
rect 13542 6352 13598 6361
rect 13542 6287 13598 6296
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13556 4622 13584 6190
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 4298 13584 4558
rect 13648 4486 13676 6734
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6390 13768 6666
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13556 4270 13676 4298
rect 13542 3768 13598 3777
rect 13542 3703 13598 3712
rect 13556 3602 13584 3703
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13556 1222 13584 3334
rect 13648 2650 13676 4270
rect 13740 2922 13768 4490
rect 13832 3720 13860 6734
rect 14200 6662 14228 6870
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14200 6254 14228 6598
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 13950 6012 14258 6021
rect 13950 6010 13956 6012
rect 14012 6010 14036 6012
rect 14092 6010 14116 6012
rect 14172 6010 14196 6012
rect 14252 6010 14258 6012
rect 14012 5958 14014 6010
rect 14194 5958 14196 6010
rect 13950 5956 13956 5958
rect 14012 5956 14036 5958
rect 14092 5956 14116 5958
rect 14172 5956 14196 5958
rect 14252 5956 14258 5958
rect 13950 5947 14258 5956
rect 14292 5760 14320 8366
rect 14476 8090 14504 8910
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14384 6458 14412 7822
rect 14476 7546 14504 7822
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14568 7342 14596 8230
rect 14660 7449 14688 8502
rect 14844 8022 14872 8978
rect 14936 8634 14964 11194
rect 15384 9784 15436 9790
rect 15384 9726 15436 9732
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15028 9246 15056 9522
rect 15106 9480 15162 9489
rect 15106 9415 15162 9424
rect 15120 9246 15148 9415
rect 15016 9240 15068 9246
rect 15016 9182 15068 9188
rect 15108 9240 15160 9246
rect 15108 9182 15160 9188
rect 15010 8732 15318 8741
rect 15010 8730 15016 8732
rect 15072 8730 15096 8732
rect 15152 8730 15176 8732
rect 15232 8730 15256 8732
rect 15312 8730 15318 8732
rect 15072 8678 15074 8730
rect 15254 8678 15256 8730
rect 15010 8676 15016 8678
rect 15072 8676 15096 8678
rect 15152 8676 15176 8678
rect 15232 8676 15256 8678
rect 15312 8676 15318 8678
rect 15010 8667 15318 8676
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15396 8498 15424 9726
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14738 7576 14794 7585
rect 14738 7511 14740 7520
rect 14792 7511 14794 7520
rect 14740 7482 14792 7488
rect 14646 7440 14702 7449
rect 14844 7410 14872 7958
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14646 7375 14702 7384
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14936 7342 14964 7822
rect 15010 7644 15318 7653
rect 15010 7642 15016 7644
rect 15072 7642 15096 7644
rect 15152 7642 15176 7644
rect 15232 7642 15256 7644
rect 15312 7642 15318 7644
rect 15072 7590 15074 7642
rect 15254 7590 15256 7642
rect 15010 7588 15016 7590
rect 15072 7588 15096 7590
rect 15152 7588 15176 7590
rect 15232 7588 15256 7590
rect 15312 7588 15318 7590
rect 15010 7579 15318 7588
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14476 7018 14504 7278
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14554 7032 14610 7041
rect 14476 6990 14554 7018
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14372 6248 14424 6254
rect 14476 6236 14504 6990
rect 14554 6967 14610 6976
rect 14554 6896 14610 6905
rect 14554 6831 14610 6840
rect 14568 6633 14596 6831
rect 14554 6624 14610 6633
rect 14554 6559 14610 6568
rect 14424 6208 14504 6236
rect 14660 6236 14688 7210
rect 15120 7206 15148 7346
rect 15292 7336 15344 7342
rect 15344 7296 15424 7324
rect 15292 7278 15344 7284
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14740 6248 14792 6254
rect 14660 6208 14740 6236
rect 14372 6190 14424 6196
rect 14108 5732 14320 5760
rect 14108 5030 14136 5732
rect 14280 5636 14332 5642
rect 14384 5624 14412 6190
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5846 14504 6054
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14332 5596 14412 5624
rect 14280 5578 14332 5584
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 13950 4924 14258 4933
rect 13950 4922 13956 4924
rect 14012 4922 14036 4924
rect 14092 4922 14116 4924
rect 14172 4922 14196 4924
rect 14252 4922 14258 4924
rect 14012 4870 14014 4922
rect 14194 4870 14196 4922
rect 13950 4868 13956 4870
rect 14012 4868 14036 4870
rect 14092 4868 14116 4870
rect 14172 4868 14196 4870
rect 14252 4868 14258 4870
rect 13950 4859 14258 4868
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 14292 4706 14320 5578
rect 14660 5545 14688 6208
rect 14740 6190 14792 6196
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14752 5778 14780 6054
rect 14844 5953 14872 6598
rect 14936 6304 14964 6734
rect 15028 6662 15056 6938
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15010 6556 15318 6565
rect 15010 6554 15016 6556
rect 15072 6554 15096 6556
rect 15152 6554 15176 6556
rect 15232 6554 15256 6556
rect 15312 6554 15318 6556
rect 15072 6502 15074 6554
rect 15254 6502 15256 6554
rect 15010 6500 15016 6502
rect 15072 6500 15096 6502
rect 15152 6500 15176 6502
rect 15232 6500 15256 6502
rect 15312 6500 15318 6502
rect 15010 6491 15318 6500
rect 14936 6276 15056 6304
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14830 5944 14886 5953
rect 14830 5879 14886 5888
rect 14832 5840 14884 5846
rect 14832 5782 14884 5788
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14844 5574 14872 5782
rect 14740 5568 14792 5574
rect 14646 5536 14702 5545
rect 14740 5510 14792 5516
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14646 5471 14702 5480
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14384 4826 14412 5102
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 13924 4486 13952 4694
rect 14292 4678 14412 4706
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 14108 4049 14136 4558
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 13950 3836 14258 3845
rect 13950 3834 13956 3836
rect 14012 3834 14036 3836
rect 14092 3834 14116 3836
rect 14172 3834 14196 3836
rect 14252 3834 14258 3836
rect 14012 3782 14014 3834
rect 14194 3782 14196 3834
rect 13950 3780 13956 3782
rect 14012 3780 14036 3782
rect 14092 3780 14116 3782
rect 14172 3780 14196 3782
rect 14252 3780 14258 3782
rect 13950 3771 14258 3780
rect 13832 3692 13952 3720
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13832 3194 13860 3538
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13924 2836 13952 3692
rect 14188 3528 14240 3534
rect 14292 3516 14320 4558
rect 14240 3488 14320 3516
rect 14188 3470 14240 3476
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 14016 3058 14044 3402
rect 14094 3224 14150 3233
rect 14094 3159 14150 3168
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14108 2961 14136 3159
rect 14200 3097 14228 3470
rect 14384 3448 14412 4678
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14292 3420 14412 3448
rect 14186 3088 14242 3097
rect 14186 3023 14242 3032
rect 14094 2952 14150 2961
rect 14094 2887 14150 2896
rect 13832 2808 13952 2836
rect 13726 2680 13782 2689
rect 13636 2644 13688 2650
rect 13726 2615 13782 2624
rect 13636 2586 13688 2592
rect 13544 1216 13596 1222
rect 13544 1158 13596 1164
rect 13740 56 13768 2615
rect 12544 54 12678 56
rect 12544 42 12572 54
rect 12452 14 12572 42
rect 12622 0 12678 54
rect 12898 0 12954 56
rect 13174 0 13230 56
rect 13450 0 13506 56
rect 13726 0 13782 56
rect 13832 42 13860 2808
rect 13950 2748 14258 2757
rect 13950 2746 13956 2748
rect 14012 2746 14036 2748
rect 14092 2746 14116 2748
rect 14172 2746 14196 2748
rect 14252 2746 14258 2748
rect 14012 2694 14014 2746
rect 14194 2694 14196 2746
rect 13950 2692 13956 2694
rect 14012 2692 14036 2694
rect 14092 2692 14116 2694
rect 14172 2692 14196 2694
rect 14252 2692 14258 2694
rect 13950 2683 14258 2692
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 13924 2553 13952 2586
rect 13910 2544 13966 2553
rect 13910 2479 13966 2488
rect 14292 2446 14320 3420
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 13924 2038 13952 2382
rect 13912 2032 13964 2038
rect 13912 1974 13964 1980
rect 14004 808 14056 814
rect 14004 750 14056 756
rect 14016 542 14044 750
rect 14108 542 14136 2382
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14292 2106 14320 2246
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14292 1834 14320 1906
rect 14280 1828 14332 1834
rect 14280 1770 14332 1776
rect 14384 1442 14412 2994
rect 14292 1414 14412 1442
rect 14004 536 14056 542
rect 14004 478 14056 484
rect 14096 536 14148 542
rect 14096 478 14148 484
rect 13924 56 14044 82
rect 14292 56 14320 1414
rect 14476 338 14504 3878
rect 14568 746 14596 5170
rect 14752 4808 14780 5510
rect 14936 5370 14964 6122
rect 15028 5778 15056 6276
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5778 15240 6190
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15304 5574 15332 5646
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15010 5468 15318 5477
rect 15010 5466 15016 5468
rect 15072 5466 15096 5468
rect 15152 5466 15176 5468
rect 15232 5466 15256 5468
rect 15312 5466 15318 5468
rect 15072 5414 15074 5466
rect 15254 5414 15256 5466
rect 15010 5412 15016 5414
rect 15072 5412 15096 5414
rect 15152 5412 15176 5414
rect 15232 5412 15256 5414
rect 15312 5412 15318 5414
rect 15010 5403 15318 5412
rect 14924 5364 14976 5370
rect 15200 5364 15252 5370
rect 14924 5306 14976 5312
rect 15028 5324 15200 5352
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4826 14872 5170
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14660 4780 14780 4808
rect 14832 4820 14884 4826
rect 14660 3448 14688 4780
rect 14832 4762 14884 4768
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14752 4282 14780 4626
rect 14740 4276 14792 4282
rect 14936 4264 14964 4966
rect 15028 4690 15056 5324
rect 15200 5306 15252 5312
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15108 5024 15160 5030
rect 15106 4992 15108 5001
rect 15160 4992 15162 5001
rect 15106 4927 15162 4936
rect 15304 4690 15332 5034
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15108 4616 15160 4622
rect 15106 4584 15108 4593
rect 15160 4584 15162 4593
rect 15106 4519 15162 4528
rect 15010 4380 15318 4389
rect 15010 4378 15016 4380
rect 15072 4378 15096 4380
rect 15152 4378 15176 4380
rect 15232 4378 15256 4380
rect 15312 4378 15318 4380
rect 15072 4326 15074 4378
rect 15254 4326 15256 4378
rect 15010 4324 15016 4326
rect 15072 4324 15096 4326
rect 15152 4324 15176 4326
rect 15232 4324 15256 4326
rect 15312 4324 15318 4326
rect 15010 4315 15318 4324
rect 15016 4276 15068 4282
rect 14936 4236 15016 4264
rect 14740 4218 14792 4224
rect 15016 4218 15068 4224
rect 14830 3768 14886 3777
rect 14830 3703 14886 3712
rect 14844 3670 14872 3703
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 15028 3602 15056 4218
rect 15396 4162 15424 7296
rect 15488 5556 15516 9658
rect 15842 9616 15898 9625
rect 15842 9551 15898 9560
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8634 15700 8978
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15580 7721 15608 7890
rect 15566 7712 15622 7721
rect 15566 7647 15622 7656
rect 15672 7002 15700 7890
rect 15764 7546 15792 8434
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15856 6905 15884 9551
rect 16040 8634 16068 11194
rect 16396 10872 16448 10878
rect 16396 10814 16448 10820
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16118 8120 16174 8129
rect 16118 8055 16174 8064
rect 16132 7886 16160 8055
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16132 7585 16160 7822
rect 16118 7576 16174 7585
rect 16028 7540 16080 7546
rect 16118 7511 16174 7520
rect 16028 7482 16080 7488
rect 16040 7342 16068 7482
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15948 7041 15976 7210
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15934 7032 15990 7041
rect 15934 6967 15990 6976
rect 15566 6896 15622 6905
rect 15842 6896 15898 6905
rect 15622 6854 15700 6882
rect 15566 6831 15622 6840
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15580 6633 15608 6734
rect 15566 6624 15622 6633
rect 15566 6559 15622 6568
rect 15580 6322 15608 6559
rect 15672 6497 15700 6854
rect 15842 6831 15898 6840
rect 15658 6488 15714 6497
rect 15658 6423 15714 6432
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15568 5568 15620 5574
rect 15488 5528 15568 5556
rect 15568 5510 15620 5516
rect 15474 5400 15530 5409
rect 15474 5335 15530 5344
rect 15488 4593 15516 5335
rect 15752 5228 15804 5234
rect 15856 5216 15884 6831
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15804 5188 15884 5216
rect 15752 5170 15804 5176
rect 15474 4584 15530 4593
rect 15474 4519 15530 4528
rect 15200 4140 15252 4146
rect 15396 4134 15608 4162
rect 15252 4100 15332 4128
rect 15200 4082 15252 4088
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15198 4040 15254 4049
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15120 3506 15148 4014
rect 15198 3975 15254 3984
rect 15212 3602 15240 3975
rect 15304 3777 15332 4100
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15290 3768 15346 3777
rect 15290 3703 15346 3712
rect 15488 3602 15516 4014
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 14936 3478 15148 3506
rect 15292 3528 15344 3534
rect 14660 3420 14872 3448
rect 14646 3360 14702 3369
rect 14646 3295 14702 3304
rect 14660 2961 14688 3295
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14646 2952 14702 2961
rect 14646 2887 14702 2896
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14660 2281 14688 2382
rect 14646 2272 14702 2281
rect 14646 2207 14702 2216
rect 14556 740 14608 746
rect 14556 682 14608 688
rect 14752 406 14780 2994
rect 14844 1970 14872 3420
rect 14936 3176 14964 3478
rect 15344 3488 15424 3516
rect 15292 3470 15344 3476
rect 15010 3292 15318 3301
rect 15010 3290 15016 3292
rect 15072 3290 15096 3292
rect 15152 3290 15176 3292
rect 15232 3290 15256 3292
rect 15312 3290 15318 3292
rect 15072 3238 15074 3290
rect 15254 3238 15256 3290
rect 15010 3236 15016 3238
rect 15072 3236 15096 3238
rect 15152 3236 15176 3238
rect 15232 3236 15256 3238
rect 15312 3236 15318 3238
rect 15010 3227 15318 3236
rect 14936 3148 15056 3176
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 14936 474 14964 2790
rect 15028 2446 15056 3148
rect 15106 3088 15162 3097
rect 15106 3023 15108 3032
rect 15160 3023 15162 3032
rect 15108 2994 15160 3000
rect 15396 2836 15424 3488
rect 15488 2990 15516 3538
rect 15580 3097 15608 4134
rect 15842 3768 15898 3777
rect 15842 3703 15898 3712
rect 15658 3360 15714 3369
rect 15658 3295 15714 3304
rect 15566 3088 15622 3097
rect 15672 3058 15700 3295
rect 15566 3023 15622 3032
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15304 2808 15424 2836
rect 15304 2650 15332 2808
rect 15474 2680 15530 2689
rect 15292 2644 15344 2650
rect 15474 2615 15530 2624
rect 15752 2644 15804 2650
rect 15292 2586 15344 2592
rect 15488 2514 15516 2615
rect 15752 2586 15804 2592
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15764 2446 15792 2586
rect 15856 2553 15884 3703
rect 15948 3670 15976 6394
rect 16040 5681 16068 7142
rect 16132 6610 16160 7346
rect 16224 7002 16252 7822
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7041 16344 7686
rect 16408 7206 16436 10814
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9761 16528 9998
rect 16580 9852 16632 9858
rect 16580 9794 16632 9800
rect 16486 9752 16542 9761
rect 16486 9687 16542 9696
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16500 9489 16528 9590
rect 16486 9480 16542 9489
rect 16486 9415 16542 9424
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8401 16528 8774
rect 16592 8498 16620 9794
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8634 16896 9318
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 17052 8514 17080 10406
rect 17144 8634 17172 11194
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10198 17264 10406
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17590 9072 17646 9081
rect 17590 9007 17646 9016
rect 17604 8809 17632 9007
rect 17590 8800 17646 8809
rect 17590 8735 17646 8744
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16672 8492 16724 8498
rect 17052 8486 17172 8514
rect 16672 8434 16724 8440
rect 16486 8392 16542 8401
rect 16486 8327 16542 8336
rect 16684 8090 16712 8434
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16960 7954 16988 8026
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16670 7168 16726 7177
rect 16670 7103 16726 7112
rect 16302 7032 16358 7041
rect 16212 6996 16264 7002
rect 16302 6967 16358 6976
rect 16408 7002 16620 7018
rect 16408 6996 16632 7002
rect 16408 6990 16580 6996
rect 16212 6938 16264 6944
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16132 6582 16252 6610
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16132 5710 16160 6394
rect 16224 5914 16252 6582
rect 16316 6361 16344 6666
rect 16302 6352 16358 6361
rect 16302 6287 16358 6296
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16316 5710 16344 6287
rect 16408 6254 16436 6990
rect 16580 6938 16632 6944
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16592 6118 16620 6802
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16120 5704 16172 5710
rect 16026 5672 16082 5681
rect 16120 5646 16172 5652
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16026 5607 16082 5616
rect 16026 4584 16082 4593
rect 16026 4519 16082 4528
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 16040 3516 16068 4519
rect 16132 4078 16160 5646
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16224 4826 16252 5170
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16132 3602 16160 4014
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15948 3488 16068 3516
rect 15948 2774 15976 3488
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 3126 16068 3334
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15948 2746 16068 2774
rect 15842 2544 15898 2553
rect 15842 2479 15898 2488
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15010 2204 15318 2213
rect 15010 2202 15016 2204
rect 15072 2202 15096 2204
rect 15152 2202 15176 2204
rect 15232 2202 15256 2204
rect 15312 2202 15318 2204
rect 15072 2150 15074 2202
rect 15254 2150 15256 2202
rect 15010 2148 15016 2150
rect 15072 2148 15096 2150
rect 15152 2148 15176 2150
rect 15232 2148 15256 2150
rect 15312 2148 15318 2150
rect 15010 2139 15318 2148
rect 15200 2032 15252 2038
rect 15200 1974 15252 1980
rect 15660 2032 15712 2038
rect 15660 1974 15712 1980
rect 15108 1352 15160 1358
rect 15108 1294 15160 1300
rect 14832 468 14884 474
rect 14832 410 14884 416
rect 14924 468 14976 474
rect 14924 410 14976 416
rect 14556 400 14608 406
rect 14556 342 14608 348
rect 14740 400 14792 406
rect 14740 342 14792 348
rect 14464 332 14516 338
rect 14464 274 14516 280
rect 14568 56 14596 342
rect 14844 56 14872 410
rect 15120 56 15148 1294
rect 15212 105 15240 1974
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 15198 96 15254 105
rect 13924 54 14058 56
rect 13924 42 13952 54
rect 13832 14 13952 42
rect 14002 0 14058 54
rect 14278 0 14334 56
rect 14554 0 14610 56
rect 14830 0 14886 56
rect 15106 0 15162 56
rect 15396 56 15424 1906
rect 15672 1630 15700 1974
rect 15660 1624 15712 1630
rect 15660 1566 15712 1572
rect 15660 740 15712 746
rect 15660 682 15712 688
rect 15672 56 15700 682
rect 15764 270 15792 2382
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15842 1864 15898 1873
rect 15842 1799 15898 1808
rect 15856 1630 15884 1799
rect 15844 1624 15896 1630
rect 15844 1566 15896 1572
rect 15752 264 15804 270
rect 15752 206 15804 212
rect 15948 56 15976 2314
rect 16040 202 16068 2746
rect 16132 2650 16160 2994
rect 16224 2689 16252 4082
rect 16210 2680 16266 2689
rect 16120 2644 16172 2650
rect 16210 2615 16266 2624
rect 16120 2586 16172 2592
rect 16316 1873 16344 4966
rect 16408 4865 16436 5102
rect 16394 4856 16450 4865
rect 16394 4791 16450 4800
rect 16592 4146 16620 6054
rect 16684 5114 16712 7103
rect 16776 7041 16804 7210
rect 16762 7032 16818 7041
rect 16762 6967 16818 6976
rect 16868 6866 16896 7278
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16776 5914 16804 6734
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6458 16988 6598
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16868 6361 16896 6394
rect 16854 6352 16910 6361
rect 16854 6287 16910 6296
rect 17144 5930 17172 8486
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17236 7993 17264 8434
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17222 7984 17278 7993
rect 17222 7919 17278 7928
rect 17328 7886 17356 8366
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17236 6322 17264 7346
rect 17420 7041 17448 7346
rect 17406 7032 17462 7041
rect 17406 6967 17462 6976
rect 17512 6798 17540 8434
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7478 17632 7822
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17590 7168 17646 7177
rect 17590 7103 17646 7112
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17314 6624 17370 6633
rect 17314 6559 17370 6568
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 17052 5902 17172 5930
rect 16776 5234 16804 5850
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16684 5086 16804 5114
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16408 3584 16436 3878
rect 16486 3768 16542 3777
rect 16486 3703 16488 3712
rect 16540 3703 16542 3712
rect 16488 3674 16540 3680
rect 16488 3596 16540 3602
rect 16408 3556 16488 3584
rect 16488 3538 16540 3544
rect 16592 2530 16620 3946
rect 16684 3738 16712 4218
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16776 3058 16804 5086
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16868 4185 16896 4558
rect 16854 4176 16910 4185
rect 16854 4111 16910 4120
rect 16854 4040 16910 4049
rect 16854 3975 16910 3984
rect 16868 3602 16896 3975
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16868 3233 16896 3538
rect 16854 3224 16910 3233
rect 16854 3159 16910 3168
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16960 2961 16988 5170
rect 17052 4706 17080 5902
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17052 4678 17172 4706
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17052 4214 17080 4558
rect 17144 4468 17172 4678
rect 17236 4593 17264 5646
rect 17222 4584 17278 4593
rect 17222 4519 17278 4528
rect 17144 4440 17264 4468
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 16946 2952 17002 2961
rect 16946 2887 17002 2896
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16592 2502 16712 2530
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16302 1864 16358 1873
rect 16302 1799 16358 1808
rect 16486 1592 16542 1601
rect 16486 1527 16542 1536
rect 16500 1290 16528 1527
rect 16212 1284 16264 1290
rect 16212 1226 16264 1232
rect 16488 1284 16540 1290
rect 16488 1226 16540 1232
rect 16028 196 16080 202
rect 16028 138 16080 144
rect 16224 56 16252 1226
rect 16396 1080 16448 1086
rect 16396 1022 16448 1028
rect 16486 1048 16542 1057
rect 16408 785 16436 1022
rect 16486 983 16488 992
rect 16540 983 16542 992
rect 16488 954 16540 960
rect 16486 912 16542 921
rect 16486 847 16488 856
rect 16540 847 16542 856
rect 16488 818 16540 824
rect 16394 776 16450 785
rect 16592 762 16620 2314
rect 16684 921 16712 2502
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 16764 1488 16816 1494
rect 16762 1456 16764 1465
rect 16816 1456 16818 1465
rect 16762 1391 16818 1400
rect 16868 1306 16896 2314
rect 16960 1494 16988 2790
rect 16948 1488 17000 1494
rect 16948 1430 17000 1436
rect 16776 1278 16896 1306
rect 16670 912 16726 921
rect 16670 847 16726 856
rect 16394 711 16450 720
rect 16500 734 16620 762
rect 16500 56 16528 734
rect 16776 56 16804 1278
rect 17052 56 17080 2858
rect 17144 2281 17172 4082
rect 17236 3058 17264 4440
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17328 2938 17356 6559
rect 17498 6488 17554 6497
rect 17604 6474 17632 7103
rect 17696 6497 17724 10474
rect 17554 6446 17632 6474
rect 17498 6423 17554 6432
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17420 4826 17448 5646
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17408 4480 17460 4486
rect 17406 4448 17408 4457
rect 17500 4480 17552 4486
rect 17460 4448 17462 4457
rect 17500 4422 17552 4428
rect 17406 4383 17462 4392
rect 17420 3670 17448 4383
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17512 3058 17540 4422
rect 17604 4264 17632 6446
rect 17682 6488 17738 6497
rect 17682 6423 17738 6432
rect 17682 5672 17738 5681
rect 17682 5607 17738 5616
rect 17696 4758 17724 5607
rect 17788 4826 17816 10474
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 17972 9897 18000 10134
rect 17958 9888 18014 9897
rect 17958 9823 18014 9832
rect 17960 9240 18012 9246
rect 17960 9182 18012 9188
rect 17972 9081 18000 9182
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 18248 8634 18276 11194
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17880 6866 17908 7754
rect 17972 7721 18000 7890
rect 17958 7712 18014 7721
rect 17958 7647 18014 7656
rect 18064 7546 18092 8230
rect 18142 8120 18198 8129
rect 18142 8055 18198 8064
rect 18156 7721 18184 8055
rect 18142 7712 18198 7721
rect 18142 7647 18198 7656
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17972 6934 18000 7482
rect 18156 7410 18184 7647
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18248 7342 18276 8298
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 18340 6322 18368 10746
rect 18878 8800 18934 8809
rect 18878 8735 18934 8744
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18616 7342 18644 7686
rect 18892 7410 18920 8735
rect 19352 8634 19380 11194
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19156 8288 19208 8294
rect 19062 8256 19118 8265
rect 19156 8230 19208 8236
rect 19062 8191 19118 8200
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5846 17908 6054
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17880 4826 17908 4966
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17696 4457 17724 4558
rect 17972 4457 18000 5743
rect 18064 5166 18092 6258
rect 18144 6248 18196 6254
rect 18142 6216 18144 6225
rect 18196 6216 18198 6225
rect 18142 6151 18198 6160
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5710 18184 6054
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18236 5704 18288 5710
rect 18340 5681 18368 6258
rect 18524 6254 18552 7142
rect 18892 6254 18920 7346
rect 19076 7342 19104 8191
rect 19168 7410 19196 8230
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19076 7041 19104 7278
rect 19062 7032 19118 7041
rect 19062 6967 19118 6976
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18892 5930 18920 6190
rect 18800 5902 18920 5930
rect 19076 5914 19104 6734
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19168 6118 19196 6190
rect 19156 6112 19208 6118
rect 19156 6054 19208 6060
rect 19064 5908 19116 5914
rect 18236 5646 18288 5652
rect 18326 5672 18382 5681
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17682 4448 17738 4457
rect 17682 4383 17738 4392
rect 17958 4448 18014 4457
rect 17958 4383 18014 4392
rect 17604 4236 18000 4264
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17592 4072 17644 4078
rect 17590 4040 17592 4049
rect 17644 4040 17646 4049
rect 17590 3975 17646 3984
rect 17592 3936 17644 3942
rect 17644 3896 17724 3924
rect 17592 3878 17644 3884
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17604 3194 17632 3674
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17236 2910 17356 2938
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17236 2650 17264 2910
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17130 2272 17186 2281
rect 17130 2207 17186 2216
rect 17224 1760 17276 1766
rect 17224 1702 17276 1708
rect 17236 1562 17264 1702
rect 17224 1556 17276 1562
rect 17224 1498 17276 1504
rect 17328 1358 17356 2790
rect 17420 2582 17448 2790
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17604 2310 17632 2926
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17408 1488 17460 1494
rect 17592 1488 17644 1494
rect 17460 1448 17592 1476
rect 17408 1430 17460 1436
rect 17592 1430 17644 1436
rect 17696 1426 17724 3896
rect 17788 2961 17816 4082
rect 17880 3641 17908 4082
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 17972 3516 18000 4236
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 18064 3754 18092 3975
rect 18156 3924 18184 5646
rect 18248 5234 18276 5646
rect 18326 5607 18382 5616
rect 18800 5234 18828 5902
rect 19064 5850 19116 5856
rect 19260 5710 19288 6598
rect 19352 6322 19380 6666
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19444 6066 19472 10678
rect 20456 9722 20484 11194
rect 21364 9988 21416 9994
rect 21364 9930 21416 9936
rect 20720 9784 20772 9790
rect 20720 9726 20772 9732
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 19524 9240 19576 9246
rect 19524 9182 19576 9188
rect 19536 7041 19564 9182
rect 20640 9178 20668 9386
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19628 8090 19656 8774
rect 19720 8634 19748 8842
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 20548 8498 20576 9114
rect 20732 8906 20760 9726
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20810 8800 20866 8809
rect 20810 8735 20866 8744
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20536 8492 20588 8498
rect 20588 8452 20668 8480
rect 20536 8434 20588 8440
rect 19950 8188 20258 8197
rect 19950 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20196 8188
rect 20252 8186 20258 8188
rect 20012 8134 20014 8186
rect 20194 8134 20196 8186
rect 19950 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20196 8134
rect 20252 8132 20258 8134
rect 19950 8123 20258 8132
rect 20350 8120 20406 8129
rect 19616 8084 19668 8090
rect 19616 8026 19668 8032
rect 20168 8084 20220 8090
rect 20350 8055 20406 8064
rect 20168 8026 20220 8032
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19812 7546 19840 7822
rect 19890 7576 19946 7585
rect 19800 7540 19852 7546
rect 19890 7511 19892 7520
rect 19800 7482 19852 7488
rect 19944 7511 19946 7520
rect 20074 7576 20130 7585
rect 20074 7511 20130 7520
rect 19892 7482 19944 7488
rect 19614 7304 19670 7313
rect 20088 7290 20116 7511
rect 20180 7478 20208 8026
rect 20364 7857 20392 8055
rect 20350 7848 20406 7857
rect 20260 7812 20312 7818
rect 20350 7783 20406 7792
rect 20260 7754 20312 7760
rect 20168 7472 20220 7478
rect 20168 7414 20220 7420
rect 19670 7262 20116 7290
rect 20168 7336 20220 7342
rect 20272 7324 20300 7754
rect 20456 7410 20484 8434
rect 20534 8256 20590 8265
rect 20534 8191 20590 8200
rect 20548 7721 20576 8191
rect 20534 7712 20590 7721
rect 20534 7647 20590 7656
rect 20640 7410 20668 8452
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20272 7296 20395 7324
rect 20168 7278 20220 7284
rect 20367 7290 20395 7296
rect 19614 7239 19670 7248
rect 20180 7188 20208 7278
rect 20367 7262 20576 7290
rect 20180 7160 20325 7188
rect 19950 7100 20258 7109
rect 19950 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20196 7100
rect 20252 7098 20258 7100
rect 20012 7046 20014 7098
rect 20194 7046 20196 7098
rect 19950 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20196 7046
rect 20252 7044 20258 7046
rect 19522 7032 19578 7041
rect 19950 7035 20258 7044
rect 19522 6967 19578 6976
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19536 6254 19564 6734
rect 19996 6390 20024 6938
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 20088 6254 20116 6938
rect 20180 6730 20208 6938
rect 20297 6916 20325 7160
rect 20548 6934 20576 7262
rect 20536 6928 20588 6934
rect 20297 6888 20392 6916
rect 20364 6798 20392 6888
rect 20536 6870 20588 6876
rect 20548 6798 20576 6870
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20536 6792 20588 6798
rect 20732 6769 20760 7822
rect 20824 7313 20852 8735
rect 21010 8732 21318 8741
rect 21010 8730 21016 8732
rect 21072 8730 21096 8732
rect 21152 8730 21176 8732
rect 21232 8730 21256 8732
rect 21312 8730 21318 8732
rect 21072 8678 21074 8730
rect 21254 8678 21256 8730
rect 21010 8676 21016 8678
rect 21072 8676 21096 8678
rect 21152 8676 21176 8678
rect 21232 8676 21256 8678
rect 21312 8676 21318 8678
rect 21010 8667 21318 8676
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20810 7304 20866 7313
rect 20810 7239 20866 7248
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20536 6734 20588 6740
rect 20718 6760 20774 6769
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 19524 6248 19576 6254
rect 19892 6248 19944 6254
rect 19524 6190 19576 6196
rect 19628 6196 19892 6202
rect 19628 6190 19944 6196
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19352 6038 19472 6066
rect 19628 6174 19932 6190
rect 19352 5914 19380 6038
rect 19430 5944 19486 5953
rect 19340 5908 19392 5914
rect 19430 5879 19486 5888
rect 19340 5850 19392 5856
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 18972 5568 19024 5574
rect 18878 5536 18934 5545
rect 18972 5510 19024 5516
rect 18878 5471 18934 5480
rect 18892 5234 18920 5471
rect 18236 5228 18288 5234
rect 18788 5228 18840 5234
rect 18236 5170 18288 5176
rect 18524 5188 18788 5216
rect 18248 5030 18276 5170
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18432 4593 18460 5102
rect 18418 4584 18474 4593
rect 18418 4519 18474 4528
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 4049 18368 4422
rect 18326 4040 18382 4049
rect 18524 4026 18552 5188
rect 18788 5170 18840 5176
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18616 4690 18828 4706
rect 18604 4684 18828 4690
rect 18656 4678 18828 4684
rect 18604 4626 18656 4632
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18708 4185 18736 4558
rect 18800 4321 18828 4678
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18694 4176 18750 4185
rect 18694 4111 18750 4120
rect 18696 4072 18748 4078
rect 18524 3998 18644 4026
rect 18696 4014 18748 4020
rect 18326 3975 18382 3984
rect 18420 3936 18472 3942
rect 18156 3896 18368 3924
rect 18064 3726 18184 3754
rect 18156 3534 18184 3726
rect 17880 3488 18000 3516
rect 18144 3528 18196 3534
rect 17774 2952 17830 2961
rect 17774 2887 17830 2896
rect 17776 2848 17828 2854
rect 17880 2802 17908 3488
rect 18144 3470 18196 3476
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 18064 3097 18092 3402
rect 18050 3088 18106 3097
rect 18050 3023 18106 3032
rect 17828 2796 17908 2802
rect 17776 2790 17908 2796
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17788 2774 17908 2790
rect 17774 2544 17830 2553
rect 17972 2514 18000 2790
rect 18050 2680 18106 2689
rect 18050 2615 18106 2624
rect 18064 2514 18092 2615
rect 17774 2479 17830 2488
rect 17960 2508 18012 2514
rect 17788 2378 17816 2479
rect 17960 2450 18012 2456
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 18156 2009 18184 3470
rect 18340 2990 18368 3896
rect 18420 3878 18472 3884
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18340 2582 18368 2926
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18340 2106 18368 2518
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18142 2000 18198 2009
rect 18142 1935 18198 1944
rect 17684 1420 17736 1426
rect 17684 1362 17736 1368
rect 17316 1352 17368 1358
rect 17316 1294 17368 1300
rect 17866 1184 17922 1193
rect 17500 1148 17552 1154
rect 17684 1148 17736 1154
rect 17552 1108 17684 1136
rect 17500 1090 17552 1096
rect 17922 1142 18000 1170
rect 17866 1119 17922 1128
rect 17684 1090 17736 1096
rect 17316 1012 17368 1018
rect 17316 954 17368 960
rect 17328 814 17356 954
rect 17316 808 17368 814
rect 17316 750 17368 756
rect 17972 542 18000 1142
rect 17316 536 17368 542
rect 17316 478 17368 484
rect 17960 536 18012 542
rect 17960 478 18012 484
rect 17328 56 17356 478
rect 18144 468 18196 474
rect 18144 410 18196 416
rect 17868 332 17920 338
rect 17868 274 17920 280
rect 17880 56 17908 274
rect 18156 56 18184 410
rect 18432 56 18460 3878
rect 18524 3777 18552 3878
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18616 2990 18644 3998
rect 18708 3534 18736 4014
rect 18800 3777 18828 4247
rect 18786 3768 18842 3777
rect 18786 3703 18842 3712
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18708 2825 18736 3470
rect 18800 3233 18828 3606
rect 18786 3224 18842 3233
rect 18786 3159 18842 3168
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18694 2816 18750 2825
rect 18694 2751 18750 2760
rect 18786 2680 18842 2689
rect 18786 2615 18788 2624
rect 18840 2615 18842 2624
rect 18788 2586 18840 2592
rect 18892 2582 18920 2858
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18696 1420 18748 1426
rect 18696 1362 18748 1368
rect 18708 56 18736 1362
rect 18984 56 19012 5510
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19260 4826 19288 5102
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19352 4706 19380 5850
rect 19076 4678 19380 4706
rect 19076 3466 19104 4678
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 3460 19116 3466
rect 19064 3402 19116 3408
rect 19062 3088 19118 3097
rect 19062 3023 19118 3032
rect 19076 2990 19104 3023
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19076 2825 19104 2926
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 19062 2544 19118 2553
rect 19062 2479 19118 2488
rect 19076 2446 19104 2479
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19168 1426 19196 4422
rect 19260 2774 19288 4490
rect 19352 3641 19380 4558
rect 19444 4078 19472 5879
rect 19628 5642 19656 6174
rect 20088 6100 20116 6190
rect 19720 6072 20116 6100
rect 20180 6100 20208 6666
rect 20364 6610 20392 6734
rect 20718 6695 20774 6704
rect 20364 6582 20760 6610
rect 20350 6352 20406 6361
rect 20732 6322 20760 6582
rect 20350 6287 20406 6296
rect 20720 6316 20772 6322
rect 20180 6072 20325 6100
rect 19720 5778 19748 6072
rect 19950 6012 20258 6021
rect 19950 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20196 6012
rect 20252 6010 20258 6012
rect 20012 5958 20014 6010
rect 20194 5958 20196 6010
rect 19950 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20196 5958
rect 20252 5956 20258 5958
rect 19950 5947 20258 5956
rect 20297 5896 20325 6072
rect 19812 5868 20325 5896
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19614 4856 19670 4865
rect 19614 4791 19670 4800
rect 19628 4486 19656 4791
rect 19720 4554 19748 5714
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19616 4480 19668 4486
rect 19812 4434 19840 5868
rect 20364 5794 20392 6287
rect 20720 6258 20772 6264
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20534 5944 20590 5953
rect 20534 5879 20536 5888
rect 20588 5879 20590 5888
rect 20536 5850 20588 5856
rect 20180 5766 20392 5794
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 19890 5536 19946 5545
rect 19890 5471 19946 5480
rect 19904 5234 19932 5471
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 20088 5030 20116 5578
rect 20076 5024 20128 5030
rect 20180 5012 20208 5766
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20456 5545 20484 5646
rect 20442 5536 20498 5545
rect 20442 5471 20498 5480
rect 20732 5234 20760 6054
rect 20824 5914 20852 6802
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20916 5846 20944 8502
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21008 8090 21036 8366
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 21376 8242 21404 9930
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21468 8362 21496 9658
rect 21560 8634 21588 11194
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21928 9926 21956 10066
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 22100 9852 22152 9858
rect 22100 9794 22152 9800
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21284 8022 21312 8230
rect 21376 8214 21772 8242
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 20996 7948 21048 7954
rect 21048 7908 21220 7936
rect 20996 7890 21048 7896
rect 21192 7800 21220 7908
rect 21652 7886 21680 8026
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21192 7772 21496 7800
rect 21468 7721 21496 7772
rect 21454 7712 21510 7721
rect 21010 7644 21318 7653
rect 21454 7647 21510 7656
rect 21010 7642 21016 7644
rect 21072 7642 21096 7644
rect 21152 7642 21176 7644
rect 21232 7642 21256 7644
rect 21312 7642 21318 7644
rect 21072 7590 21074 7642
rect 21254 7590 21256 7642
rect 21010 7588 21016 7590
rect 21072 7588 21096 7590
rect 21152 7588 21176 7590
rect 21232 7588 21256 7590
rect 21312 7588 21318 7590
rect 21010 7579 21318 7588
rect 21652 7460 21680 7822
rect 21270 7440 21326 7449
rect 21270 7375 21326 7384
rect 21376 7432 21680 7460
rect 21284 7342 21312 7375
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 21192 6905 21220 7210
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21178 6896 21234 6905
rect 21178 6831 21234 6840
rect 21284 6644 21312 7142
rect 21376 6798 21404 7432
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21364 6792 21416 6798
rect 21456 6792 21508 6798
rect 21364 6734 21416 6740
rect 21454 6760 21456 6769
rect 21508 6760 21510 6769
rect 21454 6695 21510 6704
rect 21284 6616 21404 6644
rect 21010 6556 21318 6565
rect 21010 6554 21016 6556
rect 21072 6554 21096 6556
rect 21152 6554 21176 6556
rect 21232 6554 21256 6556
rect 21312 6554 21318 6556
rect 21072 6502 21074 6554
rect 21254 6502 21256 6554
rect 21010 6500 21016 6502
rect 21072 6500 21096 6502
rect 21152 6500 21176 6502
rect 21232 6500 21256 6502
rect 21312 6500 21318 6502
rect 21010 6491 21318 6500
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 21008 5778 21036 6394
rect 21376 6118 21404 6616
rect 21454 6624 21510 6633
rect 21454 6559 21510 6568
rect 21468 6390 21496 6559
rect 21456 6384 21508 6390
rect 21456 6326 21508 6332
rect 21560 6338 21588 7278
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21652 6458 21680 6734
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21560 6310 21680 6338
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5794 21404 6054
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21192 5766 21404 5794
rect 21192 5642 21220 5766
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 20180 4984 20392 5012
rect 20076 4966 20128 4972
rect 19950 4924 20258 4933
rect 19950 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20196 4924
rect 20252 4922 20258 4924
rect 20012 4870 20014 4922
rect 20194 4870 20196 4922
rect 19950 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20196 4870
rect 20252 4868 20258 4870
rect 19950 4859 20258 4868
rect 19616 4422 19668 4428
rect 19720 4406 19840 4434
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19432 4072 19484 4078
rect 19484 4032 19564 4060
rect 19432 4014 19484 4020
rect 19430 3904 19486 3913
rect 19430 3839 19486 3848
rect 19338 3632 19394 3641
rect 19444 3602 19472 3839
rect 19536 3602 19564 4032
rect 19338 3567 19394 3576
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19352 3233 19380 3470
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19338 3224 19394 3233
rect 19338 3159 19394 3168
rect 19444 3126 19472 3402
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19536 3058 19564 3538
rect 19628 3505 19656 4082
rect 19614 3496 19670 3505
rect 19614 3431 19670 3440
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19260 2746 19380 2774
rect 19248 1488 19300 1494
rect 19248 1430 19300 1436
rect 19156 1420 19208 1426
rect 19156 1362 19208 1368
rect 19260 56 19288 1430
rect 15198 31 15254 40
rect 15382 0 15438 56
rect 15658 0 15714 56
rect 15934 0 15990 56
rect 16210 0 16266 56
rect 16486 0 16542 56
rect 16762 0 16818 56
rect 17038 0 17094 56
rect 17314 0 17370 56
rect 17590 0 17646 56
rect 17866 0 17922 56
rect 18142 0 18198 56
rect 18418 0 18474 56
rect 18694 0 18750 56
rect 18970 0 19026 56
rect 19246 0 19302 56
rect 19352 42 19380 2746
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19536 1970 19564 2382
rect 19524 1964 19576 1970
rect 19524 1906 19576 1912
rect 19536 1698 19564 1906
rect 19524 1692 19576 1698
rect 19524 1634 19576 1640
rect 19720 1630 19748 4406
rect 19892 4072 19944 4078
rect 19812 4032 19892 4060
rect 19812 3738 19840 4032
rect 19892 4014 19944 4020
rect 20364 3913 20392 4984
rect 20456 4826 20484 5034
rect 20536 5024 20588 5030
rect 20720 5024 20772 5030
rect 20588 4984 20668 5012
rect 20536 4966 20588 4972
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20350 3904 20406 3913
rect 19950 3836 20258 3845
rect 20350 3839 20406 3848
rect 19950 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20196 3836
rect 20252 3834 20258 3836
rect 20012 3782 20014 3834
rect 20194 3782 20196 3834
rect 19950 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20196 3782
rect 20252 3780 20258 3782
rect 19950 3771 20258 3780
rect 20456 3777 20484 4422
rect 20442 3768 20498 3777
rect 19800 3732 19852 3738
rect 20442 3703 20498 3712
rect 19800 3674 19852 3680
rect 20442 3632 20498 3641
rect 20364 3590 20442 3618
rect 20168 3528 20220 3534
rect 19798 3496 19854 3505
rect 19798 3431 19854 3440
rect 20166 3496 20168 3505
rect 20220 3496 20222 3505
rect 20166 3431 20222 3440
rect 19812 2990 19840 3431
rect 20364 3369 20392 3590
rect 20442 3567 20498 3576
rect 20444 3392 20496 3398
rect 20350 3360 20406 3369
rect 20444 3334 20496 3340
rect 20350 3295 20406 3304
rect 19996 3058 20392 3074
rect 19996 3052 20404 3058
rect 19996 3046 20352 3052
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19996 2854 20024 3046
rect 20352 2994 20404 3000
rect 20456 2854 20484 3334
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 19950 2748 20258 2757
rect 19950 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20196 2748
rect 20252 2746 20258 2748
rect 20012 2694 20014 2746
rect 20194 2694 20196 2746
rect 19950 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20196 2694
rect 20252 2692 20258 2694
rect 19950 2683 20258 2692
rect 20364 2650 20392 2790
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 19708 1624 19760 1630
rect 19708 1566 19760 1572
rect 20352 1420 20404 1426
rect 20352 1362 20404 1368
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 20076 1352 20128 1358
rect 20076 1294 20128 1300
rect 19432 536 19484 542
rect 19432 478 19484 484
rect 19444 241 19472 478
rect 19430 232 19486 241
rect 19430 167 19486 176
rect 19444 56 19564 82
rect 19812 56 19840 1294
rect 20088 56 20116 1294
rect 20364 56 20392 1362
rect 20548 338 20576 4422
rect 20640 4214 20668 4984
rect 20720 4966 20772 4972
rect 20732 4622 20760 4966
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 4457 20852 4558
rect 20810 4448 20866 4457
rect 20810 4383 20866 4392
rect 20810 4312 20866 4321
rect 20810 4247 20866 4256
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20824 4010 20852 4247
rect 20916 4214 20944 5510
rect 21010 5468 21318 5477
rect 21010 5466 21016 5468
rect 21072 5466 21096 5468
rect 21152 5466 21176 5468
rect 21232 5466 21256 5468
rect 21312 5466 21318 5468
rect 21072 5414 21074 5466
rect 21254 5414 21256 5466
rect 21010 5412 21016 5414
rect 21072 5412 21096 5414
rect 21152 5412 21176 5414
rect 21232 5412 21256 5414
rect 21312 5412 21318 5414
rect 21010 5403 21318 5412
rect 21376 4865 21404 5646
rect 21468 5370 21496 5646
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21560 5250 21588 5646
rect 21468 5222 21588 5250
rect 21468 5001 21496 5222
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21454 4992 21510 5001
rect 21454 4927 21510 4936
rect 21086 4856 21142 4865
rect 21086 4791 21142 4800
rect 21362 4856 21418 4865
rect 21418 4814 21496 4842
rect 21362 4791 21418 4800
rect 21100 4690 21128 4791
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21010 4380 21318 4389
rect 21010 4378 21016 4380
rect 21072 4378 21096 4380
rect 21152 4378 21176 4380
rect 21232 4378 21256 4380
rect 21312 4378 21318 4380
rect 21072 4326 21074 4378
rect 21254 4326 21256 4378
rect 21010 4324 21016 4326
rect 21072 4324 21096 4326
rect 21152 4324 21176 4326
rect 21232 4324 21256 4326
rect 21312 4324 21318 4326
rect 21010 4315 21318 4324
rect 20904 4208 20956 4214
rect 20904 4150 20956 4156
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20640 3726 21036 3754
rect 20640 3194 20668 3726
rect 21008 3466 21036 3726
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20904 3392 20956 3398
rect 20824 3340 20904 3346
rect 20824 3334 20956 3340
rect 20824 3318 20944 3334
rect 20718 3224 20774 3233
rect 20628 3188 20680 3194
rect 20718 3159 20720 3168
rect 20628 3130 20680 3136
rect 20772 3159 20774 3168
rect 20720 3130 20772 3136
rect 20824 3074 20852 3318
rect 21010 3292 21318 3301
rect 21010 3290 21016 3292
rect 21072 3290 21096 3292
rect 21152 3290 21176 3292
rect 21232 3290 21256 3292
rect 21312 3290 21318 3292
rect 21072 3238 21074 3290
rect 21254 3238 21256 3290
rect 21010 3236 21016 3238
rect 21072 3236 21096 3238
rect 21152 3236 21176 3238
rect 21232 3236 21256 3238
rect 21312 3236 21318 3238
rect 21010 3227 21318 3236
rect 20732 3046 20852 3074
rect 20916 3148 21128 3176
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20640 2650 20668 2926
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20640 1698 20668 2382
rect 20628 1692 20680 1698
rect 20628 1634 20680 1640
rect 20640 1562 20668 1634
rect 20628 1556 20680 1562
rect 20628 1498 20680 1504
rect 20732 1306 20760 3046
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20824 2310 20852 2926
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20812 2100 20864 2106
rect 20812 2042 20864 2048
rect 20640 1278 20760 1306
rect 20824 1290 20852 2042
rect 20812 1284 20864 1290
rect 20536 332 20588 338
rect 20536 274 20588 280
rect 20640 56 20668 1278
rect 20812 1226 20864 1232
rect 20916 56 20944 3148
rect 20994 3088 21050 3097
rect 20994 3023 21050 3032
rect 21008 2825 21036 3023
rect 21100 2922 21128 3148
rect 21178 3088 21234 3097
rect 21178 3023 21234 3032
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 21192 2854 21220 3023
rect 21180 2848 21232 2854
rect 20994 2816 21050 2825
rect 21180 2790 21232 2796
rect 20994 2751 21050 2760
rect 21010 2204 21318 2213
rect 21010 2202 21016 2204
rect 21072 2202 21096 2204
rect 21152 2202 21176 2204
rect 21232 2202 21256 2204
rect 21312 2202 21318 2204
rect 21072 2150 21074 2202
rect 21254 2150 21256 2202
rect 21010 2148 21016 2150
rect 21072 2148 21096 2150
rect 21152 2148 21176 2150
rect 21232 2148 21256 2150
rect 21312 2148 21318 2150
rect 21010 2139 21318 2148
rect 21376 513 21404 4558
rect 21468 4146 21496 4814
rect 21560 4758 21588 5034
rect 21652 4758 21680 6310
rect 21548 4752 21600 4758
rect 21548 4694 21600 4700
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21468 2446 21496 2790
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21454 2136 21510 2145
rect 21454 2071 21510 2080
rect 21468 1601 21496 2071
rect 21454 1592 21510 1601
rect 21454 1527 21510 1536
rect 21560 1442 21588 4422
rect 21652 4214 21680 4490
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 21652 1630 21680 4150
rect 21744 4078 21772 8214
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21928 7546 21956 7822
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21824 6860 21876 6866
rect 21876 6820 21956 6848
rect 21824 6802 21876 6808
rect 21928 6458 21956 6820
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21822 6352 21878 6361
rect 21822 6287 21878 6296
rect 21836 6089 21864 6287
rect 21928 6254 21956 6394
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21822 6080 21878 6089
rect 21822 6015 21878 6024
rect 21822 5672 21878 5681
rect 21822 5607 21878 5616
rect 21836 4622 21864 5607
rect 22020 5522 22048 8910
rect 22112 8498 22140 9794
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22204 9178 22232 9386
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22296 8838 22324 9114
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22388 8634 22416 8774
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22204 7750 22232 8298
rect 22388 8090 22416 8434
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 22192 7744 22244 7750
rect 22190 7712 22192 7721
rect 22244 7712 22246 7721
rect 22190 7647 22246 7656
rect 22204 7342 22232 7647
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22112 6769 22140 7210
rect 22098 6760 22154 6769
rect 22098 6695 22154 6704
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22204 5681 22232 5782
rect 22190 5672 22246 5681
rect 22190 5607 22246 5616
rect 22284 5636 22336 5642
rect 22388 5624 22416 5782
rect 22336 5596 22416 5624
rect 22284 5578 22336 5584
rect 22388 5545 22416 5596
rect 21928 5494 22048 5522
rect 22374 5536 22430 5545
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21744 3534 21772 3878
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21640 1624 21692 1630
rect 21640 1566 21692 1572
rect 21468 1414 21588 1442
rect 21362 504 21418 513
rect 21362 439 21418 448
rect 21180 332 21232 338
rect 21180 274 21232 280
rect 21192 56 21220 274
rect 21468 56 21496 1414
rect 21836 1358 21864 3878
rect 21928 3058 21956 5494
rect 22374 5471 22430 5480
rect 22480 5352 22508 9930
rect 22664 9790 22692 11194
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22652 9784 22704 9790
rect 22652 9726 22704 9732
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22020 5324 22508 5352
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 21916 2372 21968 2378
rect 21916 2314 21968 2320
rect 21928 1426 21956 2314
rect 22020 2106 22048 5324
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 22112 4457 22140 4490
rect 22098 4448 22154 4457
rect 22098 4383 22154 4392
rect 22098 3768 22154 3777
rect 22098 3703 22154 3712
rect 22112 3466 22140 3703
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 22112 2038 22140 2382
rect 22100 2032 22152 2038
rect 22100 1974 22152 1980
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 21916 1420 21968 1426
rect 21916 1362 21968 1368
rect 21824 1352 21876 1358
rect 21824 1294 21876 1300
rect 22008 1284 22060 1290
rect 22008 1226 22060 1232
rect 21732 1216 21784 1222
rect 21732 1158 21784 1164
rect 21744 56 21772 1158
rect 22020 56 22048 1226
rect 22112 882 22140 1527
rect 22100 876 22152 882
rect 22100 818 22152 824
rect 22204 406 22232 4966
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22388 4486 22416 4762
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22282 4312 22338 4321
rect 22480 4282 22508 5170
rect 22572 4826 22600 6598
rect 22664 5817 22692 7686
rect 22756 6662 22784 10406
rect 23664 9784 23716 9790
rect 23202 9752 23258 9761
rect 23664 9726 23716 9732
rect 23202 9687 23258 9696
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22650 5808 22706 5817
rect 22650 5743 22706 5752
rect 22742 5672 22798 5681
rect 22742 5607 22798 5616
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22664 5098 22692 5306
rect 22756 5166 22784 5607
rect 22848 5352 22876 9590
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23124 7818 23152 8230
rect 23112 7812 23164 7818
rect 23112 7754 23164 7760
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23032 6458 23060 6598
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23032 6254 23060 6394
rect 23020 6248 23072 6254
rect 23020 6190 23072 6196
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 23018 6080 23074 6089
rect 22940 5846 22968 6054
rect 23018 6015 23074 6024
rect 22928 5840 22980 5846
rect 22928 5782 22980 5788
rect 23032 5681 23060 6015
rect 23018 5672 23074 5681
rect 23018 5607 23074 5616
rect 22848 5324 23060 5352
rect 22928 5228 22980 5234
rect 22848 5188 22928 5216
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22652 5092 22704 5098
rect 22652 5034 22704 5040
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22664 4690 22692 5034
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22756 4622 22784 5102
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 22572 4282 22600 4490
rect 22282 4247 22338 4256
rect 22468 4276 22520 4282
rect 22296 2961 22324 4247
rect 22468 4218 22520 4224
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22376 4004 22428 4010
rect 22376 3946 22428 3952
rect 22282 2952 22338 2961
rect 22282 2887 22338 2896
rect 22284 2644 22336 2650
rect 22388 2632 22416 3946
rect 22336 2604 22416 2632
rect 22284 2586 22336 2592
rect 22480 1902 22508 4082
rect 22664 3534 22692 4490
rect 22652 3528 22704 3534
rect 22572 3488 22652 3516
rect 22572 2038 22600 3488
rect 22652 3470 22704 3476
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22664 2378 22692 3334
rect 22756 2854 22784 4558
rect 22848 4214 22876 5188
rect 22928 5170 22980 5176
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22756 2514 22784 2790
rect 22848 2582 22876 4014
rect 22836 2576 22888 2582
rect 22836 2518 22888 2524
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 22560 2032 22612 2038
rect 22560 1974 22612 1980
rect 22468 1896 22520 1902
rect 22468 1838 22520 1844
rect 22284 876 22336 882
rect 22284 818 22336 824
rect 22192 400 22244 406
rect 22192 342 22244 348
rect 22296 56 22324 818
rect 22940 678 22968 4558
rect 23032 4321 23060 5324
rect 23124 4622 23152 6666
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23018 4312 23074 4321
rect 23018 4247 23074 4256
rect 23018 3632 23074 3641
rect 23018 3567 23074 3576
rect 23032 3466 23060 3567
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23018 3088 23074 3097
rect 23018 3023 23020 3032
rect 23072 3023 23074 3032
rect 23020 2994 23072 3000
rect 23216 2774 23244 9687
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23386 8120 23442 8129
rect 23386 8055 23442 8064
rect 23400 7886 23428 8055
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 7478 23336 7686
rect 23296 7472 23348 7478
rect 23400 7449 23428 7822
rect 23296 7414 23348 7420
rect 23386 7440 23442 7449
rect 23386 7375 23442 7384
rect 23492 7342 23520 8230
rect 23584 7970 23612 9522
rect 23676 8634 23704 9726
rect 23768 8634 23796 11194
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23860 8498 23888 8978
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23584 7942 23888 7970
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23768 6798 23796 7822
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23572 5772 23624 5778
rect 23676 5760 23704 6054
rect 23624 5732 23704 5760
rect 23572 5714 23624 5720
rect 23308 5658 23336 5714
rect 23480 5704 23532 5710
rect 23478 5672 23480 5681
rect 23532 5672 23534 5681
rect 23308 5630 23428 5658
rect 23400 5409 23428 5630
rect 23478 5607 23534 5616
rect 23386 5400 23442 5409
rect 23768 5370 23796 6734
rect 23386 5335 23442 5344
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23294 4992 23350 5001
rect 23294 4927 23350 4936
rect 23308 4078 23336 4927
rect 23400 4554 23428 5102
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2990 23520 3334
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23032 2746 23244 2774
rect 23032 1601 23060 2746
rect 23018 1592 23074 1601
rect 23018 1527 23074 1536
rect 23020 1148 23072 1154
rect 23020 1090 23072 1096
rect 23112 1148 23164 1154
rect 23112 1090 23164 1096
rect 23032 921 23060 1090
rect 23018 912 23074 921
rect 23018 847 23074 856
rect 22928 672 22980 678
rect 22928 614 22980 620
rect 22560 332 22612 338
rect 22560 274 22612 280
rect 22572 56 22600 274
rect 22848 66 22968 82
rect 22848 60 22980 66
rect 22848 56 22928 60
rect 19444 54 19578 56
rect 19444 42 19472 54
rect 19352 14 19472 42
rect 19522 0 19578 54
rect 19798 0 19854 56
rect 20074 0 20130 56
rect 20350 0 20406 56
rect 20626 0 20682 56
rect 20902 0 20958 56
rect 21178 0 21234 56
rect 21454 0 21510 56
rect 21730 0 21786 56
rect 22006 0 22062 56
rect 22282 0 22338 56
rect 22558 0 22614 56
rect 22834 54 22928 56
rect 22834 0 22890 54
rect 23124 56 23152 1090
rect 23400 56 23520 82
rect 22928 2 22980 8
rect 23110 0 23166 56
rect 23386 54 23520 56
rect 23386 0 23442 54
rect 23492 42 23520 54
rect 23584 42 23612 4422
rect 23664 4072 23716 4078
rect 23768 4060 23796 4966
rect 23716 4032 23796 4060
rect 23664 4014 23716 4020
rect 23860 3641 23888 7942
rect 23952 5030 23980 10542
rect 24676 9784 24728 9790
rect 24872 9738 24900 11194
rect 24676 9726 24728 9732
rect 24124 9240 24176 9246
rect 24124 9182 24176 9188
rect 24216 9240 24268 9246
rect 24216 9182 24268 9188
rect 24136 8022 24164 9182
rect 24228 8498 24256 9182
rect 24400 8968 24452 8974
rect 24688 8945 24716 9726
rect 24780 9710 24900 9738
rect 24400 8910 24452 8916
rect 24674 8936 24730 8945
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24044 7546 24072 7822
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24136 7546 24164 7686
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24136 7002 24164 7278
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 24032 6724 24084 6730
rect 24032 6666 24084 6672
rect 24044 5166 24072 6666
rect 24122 6216 24178 6225
rect 24122 6151 24124 6160
rect 24176 6151 24178 6160
rect 24124 6122 24176 6128
rect 24122 5400 24178 5409
rect 24122 5335 24124 5344
rect 24176 5335 24178 5344
rect 24124 5306 24176 5312
rect 24032 5160 24084 5166
rect 24228 5137 24256 7686
rect 24320 7342 24348 8026
rect 24308 7336 24360 7342
rect 24308 7278 24360 7284
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 24320 5234 24348 6258
rect 24412 5409 24440 8910
rect 24584 8900 24636 8906
rect 24674 8871 24730 8880
rect 24584 8842 24636 8848
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24504 6730 24532 7822
rect 24596 6934 24624 8842
rect 24780 8634 24808 9710
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24952 8492 25004 8498
rect 24952 8434 25004 8440
rect 24860 8288 24912 8294
rect 24860 8230 24912 8236
rect 24872 7274 24900 8230
rect 24964 7954 24992 8434
rect 25504 8288 25556 8294
rect 25042 8256 25098 8265
rect 25504 8230 25556 8236
rect 25042 8191 25098 8200
rect 25056 8090 25084 8191
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25056 7954 25084 8026
rect 25516 8022 25544 8230
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 25412 7948 25464 7954
rect 25412 7890 25464 7896
rect 25136 7540 25188 7546
rect 25056 7500 25136 7528
rect 24952 7336 25004 7342
rect 25056 7324 25084 7500
rect 25136 7482 25188 7488
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 25004 7296 25084 7324
rect 24952 7278 25004 7284
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24964 7041 24992 7278
rect 24950 7032 25006 7041
rect 24950 6967 25006 6976
rect 24584 6928 24636 6934
rect 24584 6870 24636 6876
rect 25148 6798 25176 7346
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24492 6724 24544 6730
rect 24492 6666 24544 6672
rect 24780 6338 24808 6734
rect 24872 6458 24900 6734
rect 25424 6730 25452 7890
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25608 7041 25636 7686
rect 25594 7032 25650 7041
rect 25594 6967 25650 6976
rect 25412 6724 25464 6730
rect 25412 6666 25464 6672
rect 25410 6624 25466 6633
rect 25410 6559 25466 6568
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24780 6322 24992 6338
rect 24780 6316 25004 6322
rect 24780 6310 24952 6316
rect 24952 6258 25004 6264
rect 25424 6186 25452 6559
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 25516 5953 25544 6258
rect 25596 6112 25648 6118
rect 25596 6054 25648 6060
rect 25502 5944 25558 5953
rect 25502 5879 25558 5888
rect 25608 5710 25636 6054
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24676 5568 24728 5574
rect 24676 5510 24728 5516
rect 24398 5400 24454 5409
rect 24398 5335 24454 5344
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24032 5102 24084 5108
rect 24214 5128 24270 5137
rect 24214 5063 24270 5072
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 24216 4752 24268 4758
rect 24216 4694 24268 4700
rect 23940 4548 23992 4554
rect 23940 4490 23992 4496
rect 23952 4321 23980 4490
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 23938 4312 23994 4321
rect 23938 4247 23994 4256
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 23846 3632 23902 3641
rect 23846 3567 23902 3576
rect 23662 3224 23718 3233
rect 23662 3159 23718 3168
rect 23676 610 23704 3159
rect 23756 3052 23808 3058
rect 23952 3040 23980 4014
rect 24044 3942 24072 4014
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23808 3012 23980 3040
rect 24032 3052 24084 3058
rect 23756 2994 23808 3000
rect 24032 2994 24084 3000
rect 23768 2281 23796 2994
rect 24044 2582 24072 2994
rect 24032 2576 24084 2582
rect 24032 2518 24084 2524
rect 23754 2272 23810 2281
rect 23754 2207 23810 2216
rect 24032 1080 24084 1086
rect 24032 1022 24084 1028
rect 23664 604 23716 610
rect 23664 546 23716 552
rect 23664 468 23716 474
rect 23664 410 23716 416
rect 23676 56 23704 410
rect 24044 406 24072 1022
rect 24032 400 24084 406
rect 24032 342 24084 348
rect 23952 56 24072 82
rect 23492 14 23612 42
rect 23662 0 23718 56
rect 23938 54 24072 56
rect 23938 0 23994 54
rect 24044 42 24072 54
rect 24136 42 24164 4422
rect 24228 4146 24256 4694
rect 24320 4554 24348 5170
rect 24492 5024 24544 5030
rect 24492 4966 24544 4972
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24216 3936 24268 3942
rect 24320 3924 24348 4218
rect 24268 3896 24348 3924
rect 24216 3878 24268 3884
rect 24228 2990 24256 3878
rect 24216 2984 24268 2990
rect 24216 2926 24268 2932
rect 24412 2446 24440 4558
rect 24504 2922 24532 4966
rect 24492 2916 24544 2922
rect 24492 2858 24544 2864
rect 24400 2440 24452 2446
rect 24400 2382 24452 2388
rect 24308 2304 24360 2310
rect 24308 2246 24360 2252
rect 24320 1222 24348 2246
rect 24596 1902 24624 5510
rect 24688 3777 24716 5510
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24674 3768 24730 3777
rect 24780 3738 24808 4966
rect 24872 4146 24900 5170
rect 25056 5166 25084 5646
rect 25136 5636 25188 5642
rect 25136 5578 25188 5584
rect 25228 5636 25280 5642
rect 25228 5578 25280 5584
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4865 24992 4966
rect 24950 4856 25006 4865
rect 24950 4791 25006 4800
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24674 3703 24730 3712
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24860 3460 24912 3466
rect 24860 3402 24912 3408
rect 24872 3369 24900 3402
rect 24858 3360 24914 3369
rect 24858 3295 24914 3304
rect 24872 2854 24900 3295
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24688 2106 24716 2382
rect 24676 2100 24728 2106
rect 24676 2042 24728 2048
rect 24584 1896 24636 1902
rect 24584 1838 24636 1844
rect 24676 1556 24728 1562
rect 24676 1498 24728 1504
rect 24492 1352 24544 1358
rect 24492 1294 24544 1300
rect 24308 1216 24360 1222
rect 24308 1158 24360 1164
rect 24216 1080 24268 1086
rect 24216 1022 24268 1028
rect 24228 56 24256 1022
rect 24504 56 24532 1294
rect 24688 746 24716 1498
rect 24780 950 24808 2382
rect 24860 2304 24912 2310
rect 24860 2246 24912 2252
rect 24872 1290 24900 2246
rect 24860 1284 24912 1290
rect 24860 1226 24912 1232
rect 24964 1086 24992 4422
rect 25056 4282 25084 5102
rect 25148 4758 25176 5578
rect 25240 5370 25268 5578
rect 25410 5400 25466 5409
rect 25228 5364 25280 5370
rect 25228 5306 25280 5312
rect 25320 5364 25372 5370
rect 25410 5335 25466 5344
rect 25320 5306 25372 5312
rect 25332 5001 25360 5306
rect 25424 5234 25452 5335
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 25318 4992 25374 5001
rect 25318 4927 25374 4936
rect 25136 4752 25188 4758
rect 25136 4694 25188 4700
rect 25228 4548 25280 4554
rect 25228 4490 25280 4496
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 25240 4146 25268 4490
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25596 4480 25648 4486
rect 25596 4422 25648 4428
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 25226 3632 25282 3641
rect 25226 3567 25282 3576
rect 25240 3534 25268 3567
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25042 3088 25098 3097
rect 25240 3058 25268 3470
rect 25042 3023 25098 3032
rect 25228 3052 25280 3058
rect 25056 1442 25084 3023
rect 25228 2994 25280 3000
rect 25134 2952 25190 2961
rect 25134 2887 25190 2896
rect 25148 2446 25176 2887
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25148 2009 25176 2382
rect 25134 2000 25190 2009
rect 25134 1935 25190 1944
rect 25056 1414 25176 1442
rect 25148 1329 25176 1414
rect 25332 1358 25360 4422
rect 25608 4321 25636 4422
rect 25594 4312 25650 4321
rect 25594 4247 25650 4256
rect 25700 4146 25728 9318
rect 25792 8673 25820 9318
rect 25872 8900 25924 8906
rect 25872 8842 25924 8848
rect 25778 8664 25834 8673
rect 25778 8599 25834 8608
rect 25884 7993 25912 8842
rect 25976 8634 26004 11194
rect 27080 11098 27108 11194
rect 27172 11098 27200 11206
rect 27080 11070 27200 11098
rect 26700 10192 26752 10198
rect 26752 10140 27108 10146
rect 26700 10134 27108 10140
rect 26712 10130 27108 10134
rect 26712 10124 27120 10130
rect 26712 10118 27068 10124
rect 27068 10066 27120 10072
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26988 9722 27016 9998
rect 26976 9716 27028 9722
rect 26976 9658 27028 9664
rect 26700 9308 26752 9314
rect 26700 9250 26752 9256
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 26344 8498 26372 8910
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 25950 8188 26258 8197
rect 25950 8186 25956 8188
rect 26012 8186 26036 8188
rect 26092 8186 26116 8188
rect 26172 8186 26196 8188
rect 26252 8186 26258 8188
rect 26012 8134 26014 8186
rect 26194 8134 26196 8186
rect 25950 8132 25956 8134
rect 26012 8132 26036 8134
rect 26092 8132 26116 8134
rect 26172 8132 26196 8134
rect 26252 8132 26258 8134
rect 25950 8123 26258 8132
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26160 7993 26188 8026
rect 25870 7984 25926 7993
rect 25870 7919 25926 7928
rect 26146 7984 26202 7993
rect 26146 7919 26202 7928
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 25792 7585 25820 7822
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25778 7576 25834 7585
rect 25976 7546 26004 7686
rect 26068 7546 26096 7822
rect 25778 7511 25834 7520
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25884 6798 25912 7346
rect 26344 7274 26372 8298
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26422 7576 26478 7585
rect 26422 7511 26478 7520
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 25950 7100 26258 7109
rect 25950 7098 25956 7100
rect 26012 7098 26036 7100
rect 26092 7098 26116 7100
rect 26172 7098 26196 7100
rect 26252 7098 26258 7100
rect 26012 7046 26014 7098
rect 26194 7046 26196 7098
rect 25950 7044 25956 7046
rect 26012 7044 26036 7046
rect 26092 7044 26116 7046
rect 26172 7044 26196 7046
rect 26252 7044 26258 7046
rect 25950 7035 26258 7044
rect 26344 6934 26372 7210
rect 26436 7177 26464 7511
rect 26422 7168 26478 7177
rect 26422 7103 26478 7112
rect 26332 6928 26384 6934
rect 26332 6870 26384 6876
rect 25872 6792 25924 6798
rect 25964 6792 26016 6798
rect 25872 6734 25924 6740
rect 25962 6760 25964 6769
rect 26240 6792 26292 6798
rect 26016 6760 26018 6769
rect 26516 6792 26568 6798
rect 26292 6752 26372 6780
rect 26240 6734 26292 6740
rect 25962 6695 26018 6704
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 25884 5681 25912 6598
rect 25976 6458 26004 6695
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25950 6012 26258 6021
rect 25950 6010 25956 6012
rect 26012 6010 26036 6012
rect 26092 6010 26116 6012
rect 26172 6010 26196 6012
rect 26252 6010 26258 6012
rect 26012 5958 26014 6010
rect 26194 5958 26196 6010
rect 25950 5956 25956 5958
rect 26012 5956 26036 5958
rect 26092 5956 26116 5958
rect 26172 5956 26196 5958
rect 26252 5956 26258 5958
rect 25950 5947 26258 5956
rect 26148 5772 26200 5778
rect 26148 5714 26200 5720
rect 25870 5672 25926 5681
rect 25870 5607 25926 5616
rect 26160 5545 26188 5714
rect 26146 5536 26202 5545
rect 26146 5471 26202 5480
rect 25778 5264 25834 5273
rect 25778 5199 25834 5208
rect 25792 4690 25820 5199
rect 25872 5024 25924 5030
rect 25872 4966 25924 4972
rect 25884 4758 25912 4966
rect 25950 4924 26258 4933
rect 25950 4922 25956 4924
rect 26012 4922 26036 4924
rect 26092 4922 26116 4924
rect 26172 4922 26196 4924
rect 26252 4922 26258 4924
rect 26012 4870 26014 4922
rect 26194 4870 26196 4922
rect 25950 4868 25956 4870
rect 26012 4868 26036 4870
rect 26092 4868 26116 4870
rect 26172 4868 26196 4870
rect 26252 4868 26258 4870
rect 25950 4859 26258 4868
rect 25872 4752 25924 4758
rect 25872 4694 25924 4700
rect 25780 4684 25832 4690
rect 25780 4626 25832 4632
rect 26148 4684 26200 4690
rect 26148 4626 26200 4632
rect 25780 4548 25832 4554
rect 25832 4508 25912 4536
rect 25780 4490 25832 4496
rect 25780 4208 25832 4214
rect 25780 4150 25832 4156
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25320 1352 25372 1358
rect 25134 1320 25190 1329
rect 25044 1284 25096 1290
rect 25320 1294 25372 1300
rect 25134 1255 25190 1264
rect 25044 1226 25096 1232
rect 24952 1080 25004 1086
rect 24952 1022 25004 1028
rect 24768 944 24820 950
rect 24768 886 24820 892
rect 24676 740 24728 746
rect 24676 682 24728 688
rect 24768 740 24820 746
rect 24768 682 24820 688
rect 24780 56 24808 682
rect 25056 56 25084 1226
rect 25424 1204 25452 4082
rect 25688 3936 25740 3942
rect 25594 3904 25650 3913
rect 25688 3878 25740 3884
rect 25594 3839 25650 3848
rect 25502 3768 25558 3777
rect 25502 3703 25558 3712
rect 25516 3602 25544 3703
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25608 3058 25636 3839
rect 25700 3670 25728 3878
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 25792 2990 25820 4150
rect 25884 3534 25912 4508
rect 26160 3942 26188 4626
rect 26344 4214 26372 6752
rect 26514 6760 26516 6769
rect 26568 6760 26570 6769
rect 26514 6695 26570 6704
rect 26528 6390 26556 6695
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 26436 5574 26464 6190
rect 26528 5846 26556 6190
rect 26516 5840 26568 5846
rect 26516 5782 26568 5788
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26620 5370 26648 7686
rect 26712 6798 26740 9250
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 26804 8265 26832 9114
rect 27010 8732 27318 8741
rect 27010 8730 27016 8732
rect 27072 8730 27096 8732
rect 27152 8730 27176 8732
rect 27232 8730 27256 8732
rect 27312 8730 27318 8732
rect 27072 8678 27074 8730
rect 27254 8678 27256 8730
rect 27010 8676 27016 8678
rect 27072 8676 27096 8678
rect 27152 8676 27176 8678
rect 27232 8676 27256 8678
rect 27312 8676 27318 8678
rect 27010 8667 27318 8676
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26790 8256 26846 8265
rect 26790 8191 26846 8200
rect 26896 8022 26924 8366
rect 27356 8090 27384 11206
rect 28170 11194 28226 11250
rect 29274 11194 29330 11250
rect 30378 11194 30434 11250
rect 31482 11194 31538 11250
rect 31588 11206 31800 11234
rect 28184 9722 28212 11194
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 27434 9208 27490 9217
rect 27434 9143 27490 9152
rect 27448 8498 27476 9143
rect 28356 8832 28408 8838
rect 28356 8774 28408 8780
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 27344 8084 27396 8090
rect 27344 8026 27396 8032
rect 28184 8022 28212 8230
rect 26884 8016 26936 8022
rect 26884 7958 26936 7964
rect 28172 8016 28224 8022
rect 28172 7958 28224 7964
rect 26790 7712 26846 7721
rect 26790 7647 26846 7656
rect 26804 7546 26832 7647
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 26896 7410 26924 7958
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 27010 7644 27318 7653
rect 27010 7642 27016 7644
rect 27072 7642 27096 7644
rect 27152 7642 27176 7644
rect 27232 7642 27256 7644
rect 27312 7642 27318 7644
rect 27072 7590 27074 7642
rect 27254 7590 27256 7642
rect 27010 7588 27016 7590
rect 27072 7588 27096 7590
rect 27152 7588 27176 7590
rect 27232 7588 27256 7590
rect 27312 7588 27318 7590
rect 27010 7579 27318 7588
rect 26884 7404 26936 7410
rect 26884 7346 26936 7352
rect 27356 7313 27384 7890
rect 27436 7880 27488 7886
rect 27896 7880 27948 7886
rect 27488 7840 27568 7868
rect 27436 7822 27488 7828
rect 27434 7440 27490 7449
rect 27434 7375 27436 7384
rect 27488 7375 27490 7384
rect 27436 7346 27488 7352
rect 27342 7304 27398 7313
rect 27160 7268 27212 7274
rect 27342 7239 27398 7248
rect 27160 7210 27212 7216
rect 26790 6896 26846 6905
rect 27172 6866 27200 7210
rect 27356 7041 27384 7239
rect 27342 7032 27398 7041
rect 27342 6967 27398 6976
rect 26790 6831 26846 6840
rect 27160 6860 27212 6866
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26698 6488 26754 6497
rect 26698 6423 26754 6432
rect 26712 6390 26740 6423
rect 26700 6384 26752 6390
rect 26700 6326 26752 6332
rect 26698 6216 26754 6225
rect 26698 6151 26754 6160
rect 26712 5778 26740 6151
rect 26804 5817 26832 6831
rect 27160 6802 27212 6808
rect 27344 6792 27396 6798
rect 27396 6752 27476 6780
rect 27344 6734 27396 6740
rect 27448 6662 27476 6752
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27010 6556 27318 6565
rect 27010 6554 27016 6556
rect 27072 6554 27096 6556
rect 27152 6554 27176 6556
rect 27232 6554 27256 6556
rect 27312 6554 27318 6556
rect 27072 6502 27074 6554
rect 27254 6502 27256 6554
rect 27010 6500 27016 6502
rect 27072 6500 27096 6502
rect 27152 6500 27176 6502
rect 27232 6500 27256 6502
rect 27312 6500 27318 6502
rect 27010 6491 27318 6500
rect 27160 6180 27212 6186
rect 27160 6122 27212 6128
rect 26884 6112 26936 6118
rect 26884 6054 26936 6060
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 26790 5808 26846 5817
rect 26700 5772 26752 5778
rect 26790 5743 26846 5752
rect 26700 5714 26752 5720
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26424 5024 26476 5030
rect 26424 4966 26476 4972
rect 26332 4208 26384 4214
rect 26332 4150 26384 4156
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26252 4010 26280 4082
rect 26436 4078 26464 4966
rect 26528 4865 26556 5306
rect 26804 5234 26832 5510
rect 26896 5273 26924 6054
rect 26988 5914 27016 6054
rect 27066 5944 27122 5953
rect 26976 5908 27028 5914
rect 27172 5914 27200 6122
rect 27066 5879 27122 5888
rect 27160 5908 27212 5914
rect 26976 5850 27028 5856
rect 27080 5778 27108 5879
rect 27160 5850 27212 5856
rect 27356 5778 27384 6598
rect 27434 6488 27490 6497
rect 27434 6423 27490 6432
rect 27448 6390 27476 6423
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 27068 5772 27120 5778
rect 27068 5714 27120 5720
rect 27344 5772 27396 5778
rect 27344 5714 27396 5720
rect 27010 5468 27318 5477
rect 27010 5466 27016 5468
rect 27072 5466 27096 5468
rect 27152 5466 27176 5468
rect 27232 5466 27256 5468
rect 27312 5466 27318 5468
rect 27072 5414 27074 5466
rect 27254 5414 27256 5466
rect 27010 5412 27016 5414
rect 27072 5412 27096 5414
rect 27152 5412 27176 5414
rect 27232 5412 27256 5414
rect 27312 5412 27318 5414
rect 27010 5403 27318 5412
rect 27434 5400 27490 5409
rect 27434 5335 27436 5344
rect 27488 5335 27490 5344
rect 27436 5306 27488 5312
rect 26882 5264 26938 5273
rect 26792 5228 26844 5234
rect 26882 5199 26938 5208
rect 27436 5228 27488 5234
rect 26792 5170 26844 5176
rect 27436 5170 27488 5176
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 26514 4856 26570 4865
rect 26514 4791 26570 4800
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26620 4457 26648 4558
rect 26606 4448 26662 4457
rect 26662 4406 26740 4434
rect 26606 4383 26662 4392
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26424 4072 26476 4078
rect 26528 4049 26556 4082
rect 26424 4014 26476 4020
rect 26514 4040 26570 4049
rect 26240 4004 26292 4010
rect 26514 3975 26570 3984
rect 26240 3946 26292 3952
rect 26148 3936 26200 3942
rect 26148 3878 26200 3884
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 25950 3836 26258 3845
rect 25950 3834 25956 3836
rect 26012 3834 26036 3836
rect 26092 3834 26116 3836
rect 26172 3834 26196 3836
rect 26252 3834 26258 3836
rect 26012 3782 26014 3834
rect 26194 3782 26196 3834
rect 25950 3780 25956 3782
rect 26012 3780 26036 3782
rect 26092 3780 26116 3782
rect 26172 3780 26196 3782
rect 26252 3780 26258 3782
rect 25950 3771 26258 3780
rect 25872 3528 25924 3534
rect 25964 3528 26016 3534
rect 25872 3470 25924 3476
rect 25962 3496 25964 3505
rect 26016 3496 26018 3505
rect 25780 2984 25832 2990
rect 25700 2961 25780 2972
rect 25686 2952 25780 2961
rect 25742 2944 25780 2952
rect 25780 2926 25832 2932
rect 25686 2887 25742 2896
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25516 2446 25544 2790
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25516 1970 25544 2382
rect 25700 2310 25728 2887
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 25688 2304 25740 2310
rect 25688 2246 25740 2252
rect 25504 1964 25556 1970
rect 25504 1906 25556 1912
rect 25332 1176 25452 1204
rect 25332 56 25360 1176
rect 25596 944 25648 950
rect 25596 886 25648 892
rect 25608 56 25636 886
rect 25792 338 25820 2790
rect 25884 1970 25912 3470
rect 25962 3431 26018 3440
rect 26146 3088 26202 3097
rect 26146 3023 26148 3032
rect 26200 3023 26202 3032
rect 26148 2994 26200 3000
rect 25950 2748 26258 2757
rect 25950 2746 25956 2748
rect 26012 2746 26036 2748
rect 26092 2746 26116 2748
rect 26172 2746 26196 2748
rect 26252 2746 26258 2748
rect 26012 2694 26014 2746
rect 26194 2694 26196 2746
rect 25950 2692 25956 2694
rect 26012 2692 26036 2694
rect 26092 2692 26116 2694
rect 26172 2692 26196 2694
rect 26252 2692 26258 2694
rect 25950 2683 26258 2692
rect 25872 1964 25924 1970
rect 25872 1906 25924 1912
rect 25884 1766 25912 1906
rect 25872 1760 25924 1766
rect 25872 1702 25924 1708
rect 25870 1320 25926 1329
rect 25870 1255 25926 1264
rect 25780 332 25832 338
rect 25780 274 25832 280
rect 25884 56 25912 1255
rect 26344 746 26372 3878
rect 26424 3596 26476 3602
rect 26476 3556 26556 3584
rect 26424 3538 26476 3544
rect 26422 3496 26478 3505
rect 26422 3431 26478 3440
rect 26436 3058 26464 3431
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26424 2848 26476 2854
rect 26424 2790 26476 2796
rect 26436 1154 26464 2790
rect 26528 2582 26556 3556
rect 26620 2922 26648 4082
rect 26712 4026 26740 4406
rect 26804 4214 26832 4558
rect 26792 4208 26844 4214
rect 26792 4150 26844 4156
rect 26712 3998 26832 4026
rect 26700 3936 26752 3942
rect 26804 3913 26832 3998
rect 26700 3878 26752 3884
rect 26790 3904 26846 3913
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26516 2576 26568 2582
rect 26516 2518 26568 2524
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 26608 2304 26660 2310
rect 26608 2246 26660 2252
rect 26424 1148 26476 1154
rect 26424 1090 26476 1096
rect 26424 1012 26476 1018
rect 26424 954 26476 960
rect 26332 740 26384 746
rect 26332 682 26384 688
rect 26148 400 26200 406
rect 26148 342 26200 348
rect 26160 56 26188 342
rect 26436 56 26464 954
rect 26528 882 26556 2246
rect 26620 2038 26648 2246
rect 26608 2032 26660 2038
rect 26608 1974 26660 1980
rect 26712 1290 26740 3878
rect 26790 3839 26846 3848
rect 26804 3602 26832 3839
rect 26896 3754 26924 4966
rect 27010 4380 27318 4389
rect 27010 4378 27016 4380
rect 27072 4378 27096 4380
rect 27152 4378 27176 4380
rect 27232 4378 27256 4380
rect 27312 4378 27318 4380
rect 27072 4326 27074 4378
rect 27254 4326 27256 4378
rect 27010 4324 27016 4326
rect 27072 4324 27096 4326
rect 27152 4324 27176 4326
rect 27232 4324 27256 4326
rect 27312 4324 27318 4326
rect 27010 4315 27318 4324
rect 27160 4208 27212 4214
rect 27158 4176 27160 4185
rect 27212 4176 27214 4185
rect 27158 4111 27214 4120
rect 27356 3890 27384 4966
rect 27448 4826 27476 5170
rect 27540 5137 27568 7840
rect 27896 7822 27948 7828
rect 27908 7410 27936 7822
rect 28080 7540 28132 7546
rect 28080 7482 28132 7488
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27896 7404 27948 7410
rect 27896 7346 27948 7352
rect 27724 6798 27752 7346
rect 27620 6792 27672 6798
rect 27620 6734 27672 6740
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 27632 6304 27660 6734
rect 28092 6322 28120 7482
rect 28264 7404 28316 7410
rect 28264 7346 28316 7352
rect 28276 6866 28304 7346
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28276 6322 28304 6598
rect 27804 6316 27856 6322
rect 27632 6276 27804 6304
rect 28080 6316 28132 6322
rect 27804 6258 27856 6264
rect 27908 6276 28080 6304
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27632 5234 27660 5782
rect 27908 5778 27936 6276
rect 28080 6258 28132 6264
rect 28264 6316 28316 6322
rect 28264 6258 28316 6264
rect 27896 5772 27948 5778
rect 27816 5732 27896 5760
rect 27712 5568 27764 5574
rect 27712 5510 27764 5516
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 27724 5166 27752 5510
rect 27712 5160 27764 5166
rect 27526 5128 27582 5137
rect 27712 5102 27764 5108
rect 27526 5063 27582 5072
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27448 4457 27476 4626
rect 27620 4480 27672 4486
rect 27434 4448 27490 4457
rect 27620 4422 27672 4428
rect 27434 4383 27490 4392
rect 27632 4321 27660 4422
rect 27618 4312 27674 4321
rect 27618 4247 27674 4256
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27356 3862 27476 3890
rect 26896 3726 27384 3754
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 26976 3528 27028 3534
rect 26896 3488 26976 3516
rect 26790 3360 26846 3369
rect 26790 3295 26846 3304
rect 26804 2961 26832 3295
rect 26790 2952 26846 2961
rect 26790 2887 26846 2896
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26804 2038 26832 2790
rect 26896 2514 26924 3488
rect 26976 3470 27028 3476
rect 27010 3292 27318 3301
rect 27010 3290 27016 3292
rect 27072 3290 27096 3292
rect 27152 3290 27176 3292
rect 27232 3290 27256 3292
rect 27312 3290 27318 3292
rect 27072 3238 27074 3290
rect 27254 3238 27256 3290
rect 27010 3236 27016 3238
rect 27072 3236 27096 3238
rect 27152 3236 27176 3238
rect 27232 3236 27256 3238
rect 27312 3236 27318 3238
rect 27010 3227 27318 3236
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 26988 2825 27016 2994
rect 27068 2848 27120 2854
rect 26974 2816 27030 2825
rect 27068 2790 27120 2796
rect 26974 2751 27030 2760
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 27080 2292 27108 2790
rect 26896 2281 27108 2292
rect 26882 2272 27108 2281
rect 26938 2264 27108 2272
rect 26882 2207 26938 2216
rect 27010 2204 27318 2213
rect 27010 2202 27016 2204
rect 27072 2202 27096 2204
rect 27152 2202 27176 2204
rect 27232 2202 27256 2204
rect 27312 2202 27318 2204
rect 27072 2150 27074 2202
rect 27254 2150 27256 2202
rect 27010 2148 27016 2150
rect 27072 2148 27096 2150
rect 27152 2148 27176 2150
rect 27232 2148 27256 2150
rect 27312 2148 27318 2150
rect 27010 2139 27318 2148
rect 26792 2032 26844 2038
rect 26792 1974 26844 1980
rect 26700 1284 26752 1290
rect 26700 1226 26752 1232
rect 26700 1148 26752 1154
rect 26700 1090 26752 1096
rect 26516 876 26568 882
rect 26516 818 26568 824
rect 26712 56 26740 1090
rect 27356 950 27384 3726
rect 27448 2106 27476 3862
rect 27632 3738 27660 4082
rect 27816 3942 27844 5732
rect 27896 5714 27948 5720
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 27896 5364 27948 5370
rect 27896 5306 27948 5312
rect 27908 4690 27936 5306
rect 28092 5302 28120 5646
rect 28080 5296 28132 5302
rect 28080 5238 28132 5244
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 28092 5080 28120 5238
rect 28000 5052 28120 5080
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27894 4040 27950 4049
rect 27894 3975 27950 3984
rect 27804 3936 27856 3942
rect 27804 3878 27856 3884
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 27712 3596 27764 3602
rect 27816 3584 27844 3878
rect 27908 3777 27936 3975
rect 27894 3768 27950 3777
rect 27894 3703 27950 3712
rect 28000 3652 28028 5052
rect 28184 5030 28212 5238
rect 28172 5024 28224 5030
rect 28078 4992 28134 5001
rect 28172 4966 28224 4972
rect 28078 4927 28134 4936
rect 27764 3556 27844 3584
rect 27908 3624 28028 3652
rect 27712 3538 27764 3544
rect 27620 3392 27672 3398
rect 27526 3360 27582 3369
rect 27620 3334 27672 3340
rect 27526 3295 27582 3304
rect 27540 2990 27568 3295
rect 27632 2990 27660 3334
rect 27710 3224 27766 3233
rect 27710 3159 27766 3168
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27620 2984 27672 2990
rect 27620 2926 27672 2932
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 27436 2100 27488 2106
rect 27436 2042 27488 2048
rect 27528 2100 27580 2106
rect 27528 2042 27580 2048
rect 27540 1630 27568 2042
rect 27632 1698 27660 2382
rect 27620 1692 27672 1698
rect 27620 1634 27672 1640
rect 27528 1624 27580 1630
rect 27528 1566 27580 1572
rect 27344 944 27396 950
rect 27344 886 27396 892
rect 27724 814 27752 3159
rect 27908 1562 27936 3624
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 28000 1698 28028 3470
rect 28092 2938 28120 4927
rect 28172 4616 28224 4622
rect 28276 4604 28304 6258
rect 28224 4576 28304 4604
rect 28172 4558 28224 4564
rect 28172 4004 28224 4010
rect 28172 3946 28224 3952
rect 28264 4004 28316 4010
rect 28264 3946 28316 3952
rect 28184 3058 28212 3946
rect 28172 3052 28224 3058
rect 28172 2994 28224 3000
rect 28092 2910 28212 2938
rect 28184 1698 28212 2910
rect 28276 2689 28304 3946
rect 28368 3534 28396 8774
rect 28552 7970 28580 10610
rect 28908 10328 28960 10334
rect 28908 10270 28960 10276
rect 28920 8838 28948 10270
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 29288 8634 29316 11194
rect 29644 9716 29696 9722
rect 29644 9658 29696 9664
rect 29276 8628 29328 8634
rect 29276 8570 29328 8576
rect 29656 8362 29684 9658
rect 30012 9444 30064 9450
rect 30012 9386 30064 9392
rect 29644 8356 29696 8362
rect 29644 8298 29696 8304
rect 29460 8288 29512 8294
rect 29460 8230 29512 8236
rect 29642 8256 29698 8265
rect 28552 7942 28856 7970
rect 28552 7886 28580 7942
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28540 7880 28592 7886
rect 28540 7822 28592 7828
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28460 6322 28488 7822
rect 28736 7546 28764 7822
rect 28828 7546 28856 7942
rect 29092 7948 29144 7954
rect 29092 7890 29144 7896
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 28632 7404 28684 7410
rect 28632 7346 28684 7352
rect 28644 7206 28672 7346
rect 28908 7268 28960 7274
rect 28908 7210 28960 7216
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28920 7002 28948 7210
rect 29104 7041 29132 7890
rect 29472 7410 29500 8230
rect 29642 8191 29698 8200
rect 29656 7721 29684 8191
rect 29920 7744 29972 7750
rect 29642 7712 29698 7721
rect 29920 7686 29972 7692
rect 29642 7647 29698 7656
rect 29734 7576 29790 7585
rect 29734 7511 29790 7520
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 29366 7304 29422 7313
rect 29090 7032 29146 7041
rect 28908 6996 28960 7002
rect 29090 6967 29146 6976
rect 28908 6938 28960 6944
rect 29196 6905 29224 7278
rect 29288 6934 29316 7278
rect 29366 7239 29422 7248
rect 29276 6928 29328 6934
rect 29182 6896 29238 6905
rect 29276 6870 29328 6876
rect 29182 6831 29238 6840
rect 29274 6488 29330 6497
rect 29274 6423 29330 6432
rect 28540 6384 28592 6390
rect 28540 6326 28592 6332
rect 28448 6316 28500 6322
rect 28448 6258 28500 6264
rect 28460 6225 28488 6258
rect 28446 6216 28502 6225
rect 28446 6151 28502 6160
rect 28552 5574 28580 6326
rect 29288 6254 29316 6423
rect 29184 6248 29236 6254
rect 28814 6216 28870 6225
rect 29184 6190 29236 6196
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 28814 6151 28870 6160
rect 28448 5568 28500 5574
rect 28448 5510 28500 5516
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 28630 5536 28686 5545
rect 28460 5234 28488 5510
rect 28448 5228 28500 5234
rect 28448 5170 28500 5176
rect 28448 4072 28500 4078
rect 28448 4014 28500 4020
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28460 3194 28488 4014
rect 28448 3188 28500 3194
rect 28448 3130 28500 3136
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28368 2825 28396 2926
rect 28354 2816 28410 2825
rect 28354 2751 28410 2760
rect 28262 2680 28318 2689
rect 28262 2615 28318 2624
rect 28264 2304 28316 2310
rect 28264 2246 28316 2252
rect 28276 1766 28304 2246
rect 28368 1970 28396 2751
rect 28552 2446 28580 5510
rect 28630 5471 28686 5480
rect 28644 3233 28672 5471
rect 28828 3618 28856 6151
rect 29000 6112 29052 6118
rect 29196 6089 29224 6190
rect 29000 6054 29052 6060
rect 29182 6080 29238 6089
rect 28908 5568 28960 5574
rect 28908 5510 28960 5516
rect 28920 5166 28948 5510
rect 28908 5160 28960 5166
rect 28908 5102 28960 5108
rect 28908 4480 28960 4486
rect 28908 4422 28960 4428
rect 28920 4078 28948 4422
rect 28908 4072 28960 4078
rect 29012 4060 29040 6054
rect 29182 6015 29238 6024
rect 29092 5636 29144 5642
rect 29092 5578 29144 5584
rect 29104 5370 29132 5578
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29092 5228 29144 5234
rect 29092 5170 29144 5176
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29104 4570 29132 5170
rect 29288 4690 29316 5170
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 29104 4542 29224 4570
rect 29092 4480 29144 4486
rect 29092 4422 29144 4428
rect 29104 4282 29132 4422
rect 29196 4282 29224 4542
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 29288 4162 29316 4626
rect 29196 4134 29316 4162
rect 29092 4072 29144 4078
rect 29012 4032 29092 4060
rect 28908 4014 28960 4020
rect 29092 4014 29144 4020
rect 28828 3590 29040 3618
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 29012 3482 29040 3590
rect 28630 3224 28686 3233
rect 28920 3194 28948 3470
rect 29012 3454 29132 3482
rect 29000 3392 29052 3398
rect 29000 3334 29052 3340
rect 28630 3159 28686 3168
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28816 2984 28868 2990
rect 28644 2944 28816 2972
rect 28644 2689 28672 2944
rect 28816 2926 28868 2932
rect 28908 2848 28960 2854
rect 28828 2825 28908 2836
rect 28814 2816 28908 2825
rect 28870 2808 28908 2816
rect 28908 2790 28960 2796
rect 28814 2751 28870 2760
rect 28630 2680 28686 2689
rect 28630 2615 28686 2624
rect 28814 2680 28870 2689
rect 28814 2615 28870 2624
rect 28540 2440 28592 2446
rect 28724 2440 28776 2446
rect 28592 2400 28724 2428
rect 28540 2382 28592 2388
rect 28724 2382 28776 2388
rect 28828 2378 28856 2615
rect 28816 2372 28868 2378
rect 28816 2314 28868 2320
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 28448 2304 28500 2310
rect 28448 2246 28500 2252
rect 28356 1964 28408 1970
rect 28356 1906 28408 1912
rect 28264 1760 28316 1766
rect 28264 1702 28316 1708
rect 27988 1692 28040 1698
rect 27988 1634 28040 1640
rect 28172 1692 28224 1698
rect 28172 1634 28224 1640
rect 27896 1556 27948 1562
rect 27896 1498 27948 1504
rect 28354 1320 28410 1329
rect 28354 1255 28410 1264
rect 27712 808 27764 814
rect 27712 750 27764 756
rect 27804 740 27856 746
rect 27804 682 27856 688
rect 26976 604 27028 610
rect 26976 546 27028 552
rect 26988 56 27016 546
rect 27252 264 27304 270
rect 27252 206 27304 212
rect 27264 56 27292 206
rect 27528 196 27580 202
rect 27528 138 27580 144
rect 27540 56 27568 138
rect 27816 56 27844 682
rect 28080 536 28132 542
rect 28080 478 28132 484
rect 28092 56 28120 478
rect 28368 56 28396 1255
rect 28460 1193 28488 2246
rect 28446 1184 28502 1193
rect 28446 1119 28502 1128
rect 28630 1048 28686 1057
rect 28920 1034 28948 2314
rect 29012 2122 29040 3334
rect 29104 2378 29132 3454
rect 29092 2372 29144 2378
rect 29092 2314 29144 2320
rect 29012 2094 29132 2122
rect 29000 2032 29052 2038
rect 29000 1974 29052 1980
rect 29012 1086 29040 1974
rect 28630 983 28686 992
rect 28828 1006 28948 1034
rect 29000 1080 29052 1086
rect 29000 1022 29052 1028
rect 28644 56 28672 983
rect 28828 921 28856 1006
rect 28908 944 28960 950
rect 28814 912 28870 921
rect 28908 886 28960 892
rect 28814 847 28870 856
rect 28920 56 28948 886
rect 29104 474 29132 2094
rect 29196 1834 29224 4134
rect 29380 4060 29408 7239
rect 29460 5840 29512 5846
rect 29460 5782 29512 5788
rect 29472 5574 29500 5782
rect 29460 5568 29512 5574
rect 29460 5510 29512 5516
rect 29644 5364 29696 5370
rect 29644 5306 29696 5312
rect 29552 5024 29604 5030
rect 29552 4966 29604 4972
rect 29460 4752 29512 4758
rect 29460 4694 29512 4700
rect 29472 4457 29500 4694
rect 29458 4448 29514 4457
rect 29458 4383 29514 4392
rect 29564 4146 29592 4966
rect 29656 4457 29684 5306
rect 29642 4448 29698 4457
rect 29642 4383 29698 4392
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29288 4032 29408 4060
rect 29458 4040 29514 4049
rect 29184 1828 29236 1834
rect 29184 1770 29236 1776
rect 29184 1148 29236 1154
rect 29184 1090 29236 1096
rect 29092 468 29144 474
rect 29092 410 29144 416
rect 29196 56 29224 1090
rect 29288 338 29316 4032
rect 29458 3975 29514 3984
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29380 3194 29408 3334
rect 29472 3233 29500 3975
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 29656 3602 29684 3878
rect 29644 3596 29696 3602
rect 29644 3538 29696 3544
rect 29656 3482 29684 3538
rect 29564 3454 29684 3482
rect 29458 3224 29514 3233
rect 29368 3188 29420 3194
rect 29458 3159 29514 3168
rect 29368 3130 29420 3136
rect 29564 2961 29592 3454
rect 29644 3392 29696 3398
rect 29748 3369 29776 7511
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 29840 4865 29868 5646
rect 29826 4856 29882 4865
rect 29826 4791 29882 4800
rect 29828 4684 29880 4690
rect 29828 4626 29880 4632
rect 29840 4196 29868 4626
rect 29932 4321 29960 7686
rect 30024 5098 30052 9386
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30300 8072 30328 8774
rect 30392 8634 30420 11194
rect 31496 11098 31524 11194
rect 31588 11098 31616 11206
rect 31496 11070 31616 11098
rect 31208 10260 31260 10266
rect 31208 10202 31260 10208
rect 30748 8832 30800 8838
rect 30748 8774 30800 8780
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30760 8498 30788 8774
rect 31220 8498 31248 10202
rect 31484 9512 31536 9518
rect 31484 9454 31536 9460
rect 31392 9172 31444 9178
rect 31392 9114 31444 9120
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 30748 8356 30800 8362
rect 30748 8298 30800 8304
rect 30760 8090 30788 8298
rect 30748 8084 30800 8090
rect 30300 8044 30420 8072
rect 30288 7948 30340 7954
rect 30288 7890 30340 7896
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30116 7546 30144 7822
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30208 5370 30236 6802
rect 30300 6322 30328 7890
rect 30392 7478 30420 8044
rect 30748 8026 30800 8032
rect 30380 7472 30432 7478
rect 30380 7414 30432 7420
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6866 30604 7142
rect 30668 7002 30696 7346
rect 30760 7274 30788 8026
rect 31116 7880 31168 7886
rect 31114 7848 31116 7857
rect 31168 7848 31170 7857
rect 31114 7783 31170 7792
rect 31128 7478 31156 7783
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 31116 7472 31168 7478
rect 31220 7449 31248 8434
rect 31298 7984 31354 7993
rect 31298 7919 31300 7928
rect 31352 7919 31354 7928
rect 31300 7890 31352 7896
rect 31116 7414 31168 7420
rect 31206 7440 31262 7449
rect 30748 7268 30800 7274
rect 30748 7210 30800 7216
rect 31036 7018 31064 7414
rect 31312 7410 31340 7890
rect 31404 7857 31432 9114
rect 31496 7993 31524 9454
rect 31772 8634 31800 11206
rect 32586 11194 32642 11250
rect 33690 11194 33746 11250
rect 34794 11194 34850 11250
rect 35898 11194 35954 11250
rect 37002 11194 37058 11250
rect 37108 11206 37320 11234
rect 32404 10396 32456 10402
rect 32404 10338 32456 10344
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 31760 8628 31812 8634
rect 31760 8570 31812 8576
rect 31680 8430 31708 8570
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 32312 8356 32364 8362
rect 32312 8298 32364 8304
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 31576 8084 31628 8090
rect 32128 8084 32180 8090
rect 31628 8044 31708 8072
rect 31576 8026 31628 8032
rect 31482 7984 31538 7993
rect 31482 7919 31538 7928
rect 31390 7848 31446 7857
rect 31390 7783 31446 7792
rect 31390 7712 31446 7721
rect 31390 7647 31446 7656
rect 31206 7375 31262 7384
rect 31300 7404 31352 7410
rect 31300 7346 31352 7352
rect 30656 6996 30708 7002
rect 31036 6990 31248 7018
rect 30656 6938 30708 6944
rect 31220 6934 31248 6990
rect 31208 6928 31260 6934
rect 31208 6870 31260 6876
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 30392 5914 30420 6258
rect 30760 5914 30788 6734
rect 30838 6488 30894 6497
rect 30838 6423 30894 6432
rect 30852 6186 30880 6423
rect 30840 6180 30892 6186
rect 30840 6122 30892 6128
rect 31116 6112 31168 6118
rect 31116 6054 31168 6060
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30748 5908 30800 5914
rect 30748 5850 30800 5856
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30840 5704 30892 5710
rect 30840 5646 30892 5652
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 30196 5364 30248 5370
rect 30196 5306 30248 5312
rect 30012 5092 30064 5098
rect 30012 5034 30064 5040
rect 30380 5024 30432 5030
rect 30380 4966 30432 4972
rect 30194 4856 30250 4865
rect 30194 4791 30250 4800
rect 30012 4752 30064 4758
rect 30012 4694 30064 4700
rect 30024 4622 30052 4694
rect 30012 4616 30064 4622
rect 30012 4558 30064 4564
rect 29918 4312 29974 4321
rect 29918 4247 29974 4256
rect 30104 4208 30156 4214
rect 29840 4168 30104 4196
rect 30104 4150 30156 4156
rect 29920 4072 29972 4078
rect 29920 4014 29972 4020
rect 29932 3738 29960 4014
rect 29920 3732 29972 3738
rect 29920 3674 29972 3680
rect 29644 3334 29696 3340
rect 29734 3360 29790 3369
rect 29550 2952 29606 2961
rect 29368 2916 29420 2922
rect 29550 2887 29606 2896
rect 29368 2858 29420 2864
rect 29380 2582 29408 2858
rect 29368 2576 29420 2582
rect 29368 2518 29420 2524
rect 29368 2372 29420 2378
rect 29368 2314 29420 2320
rect 29380 1970 29408 2314
rect 29368 1964 29420 1970
rect 29368 1906 29420 1912
rect 29460 672 29512 678
rect 29460 614 29512 620
rect 29276 332 29328 338
rect 29276 274 29328 280
rect 29472 56 29500 614
rect 29656 406 29684 3334
rect 29734 3295 29790 3304
rect 29734 3224 29790 3233
rect 29734 3159 29790 3168
rect 29748 2774 29776 3159
rect 29932 3058 29960 3674
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30010 3360 30066 3369
rect 30010 3295 30066 3304
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 29828 2984 29880 2990
rect 29826 2952 29828 2961
rect 29880 2952 29882 2961
rect 29826 2887 29882 2896
rect 29932 2854 29960 2994
rect 30024 2961 30052 3295
rect 30010 2952 30066 2961
rect 30010 2887 30066 2896
rect 29920 2848 29972 2854
rect 30116 2825 30144 3470
rect 29920 2790 29972 2796
rect 30102 2816 30158 2825
rect 29748 2746 29868 2774
rect 30102 2751 30158 2760
rect 29840 2446 29868 2746
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 29736 1964 29788 1970
rect 29736 1906 29788 1912
rect 29644 400 29696 406
rect 29644 342 29696 348
rect 29748 56 29776 1906
rect 30012 876 30064 882
rect 30012 818 30064 824
rect 30024 56 30052 818
rect 30208 377 30236 4791
rect 30288 4548 30340 4554
rect 30288 4490 30340 4496
rect 30300 1850 30328 4490
rect 30392 1952 30420 4966
rect 30484 3942 30512 5646
rect 30852 5409 30880 5646
rect 30838 5400 30894 5409
rect 30838 5335 30894 5344
rect 30564 5092 30616 5098
rect 30564 5034 30616 5040
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30472 2984 30524 2990
rect 30472 2926 30524 2932
rect 30484 2582 30512 2926
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30576 1970 30604 5034
rect 30746 4992 30802 5001
rect 30746 4927 30802 4936
rect 30760 4622 30788 4927
rect 30748 4616 30800 4622
rect 30748 4558 30800 4564
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 30564 1964 30616 1970
rect 30392 1924 30512 1952
rect 30300 1822 30420 1850
rect 30288 1284 30340 1290
rect 30288 1226 30340 1232
rect 30194 368 30250 377
rect 30194 303 30250 312
rect 30300 56 30328 1226
rect 30392 814 30420 1822
rect 30380 808 30432 814
rect 30380 750 30432 756
rect 30484 610 30512 1924
rect 30564 1906 30616 1912
rect 30668 746 30696 4218
rect 30760 3058 30788 4558
rect 30852 4214 30880 5335
rect 30840 4208 30892 4214
rect 31036 4162 31064 5646
rect 31128 4826 31156 6054
rect 31298 5672 31354 5681
rect 31298 5607 31354 5616
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31208 4752 31260 4758
rect 31208 4694 31260 4700
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 31128 4486 31156 4558
rect 31116 4480 31168 4486
rect 31116 4422 31168 4428
rect 30840 4150 30892 4156
rect 30944 4146 31064 4162
rect 31128 4146 31156 4422
rect 31220 4185 31248 4694
rect 31312 4486 31340 5607
rect 31404 5234 31432 7647
rect 31576 7200 31628 7206
rect 31482 7168 31538 7177
rect 31576 7142 31628 7148
rect 31482 7103 31538 7112
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 31392 5024 31444 5030
rect 31390 4992 31392 5001
rect 31444 4992 31446 5001
rect 31390 4927 31446 4936
rect 31390 4720 31446 4729
rect 31390 4655 31392 4664
rect 31444 4655 31446 4664
rect 31392 4626 31444 4632
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 31496 4214 31524 7103
rect 31484 4208 31536 4214
rect 31206 4176 31262 4185
rect 30932 4140 31064 4146
rect 30984 4134 31064 4140
rect 31116 4140 31168 4146
rect 30932 4082 30984 4088
rect 31484 4150 31536 4156
rect 31588 4146 31616 7142
rect 31680 6798 31708 8044
rect 32128 8026 32180 8032
rect 31760 7948 31812 7954
rect 31812 7908 31892 7936
rect 31760 7890 31812 7896
rect 31760 7744 31812 7750
rect 31760 7686 31812 7692
rect 31668 6792 31720 6798
rect 31668 6734 31720 6740
rect 31666 5400 31722 5409
rect 31666 5335 31722 5344
rect 31680 5234 31708 5335
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 31668 5092 31720 5098
rect 31668 5034 31720 5040
rect 31680 4282 31708 5034
rect 31772 4282 31800 7686
rect 31864 7274 31892 7908
rect 32036 7880 32088 7886
rect 32036 7822 32088 7828
rect 32048 7274 32076 7822
rect 32140 7585 32168 8026
rect 32324 7954 32352 8298
rect 32312 7948 32364 7954
rect 32312 7890 32364 7896
rect 32126 7576 32182 7585
rect 32126 7511 32182 7520
rect 32416 7342 32444 10338
rect 32600 8634 32628 11194
rect 33416 9716 33468 9722
rect 33416 9658 33468 9664
rect 32770 9344 32826 9353
rect 32770 9279 32826 9288
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32404 7336 32456 7342
rect 32404 7278 32456 7284
rect 31852 7268 31904 7274
rect 31852 7210 31904 7216
rect 32036 7268 32088 7274
rect 32036 7210 32088 7216
rect 32496 7268 32548 7274
rect 32496 7210 32548 7216
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 32220 6792 32272 6798
rect 32218 6760 32220 6769
rect 32272 6760 32274 6769
rect 32218 6695 32274 6704
rect 32508 6361 32536 7210
rect 32588 6656 32640 6662
rect 32588 6598 32640 6604
rect 32310 6352 32366 6361
rect 32310 6287 32312 6296
rect 32364 6287 32366 6296
rect 32494 6352 32550 6361
rect 32494 6287 32550 6296
rect 32312 6258 32364 6264
rect 32404 6248 32456 6254
rect 32508 6236 32536 6287
rect 32456 6208 32536 6236
rect 32404 6190 32456 6196
rect 32600 6186 32628 6598
rect 32588 6180 32640 6186
rect 32588 6122 32640 6128
rect 32312 6112 32364 6118
rect 32312 6054 32364 6060
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 32220 5704 32272 5710
rect 32140 5652 32220 5658
rect 32324 5681 32352 6054
rect 32692 5930 32720 8434
rect 32784 7750 32812 9279
rect 32864 8900 32916 8906
rect 32864 8842 32916 8848
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 32876 6730 32904 8842
rect 33010 8732 33318 8741
rect 33010 8730 33016 8732
rect 33072 8730 33096 8732
rect 33152 8730 33176 8732
rect 33232 8730 33256 8732
rect 33312 8730 33318 8732
rect 33072 8678 33074 8730
rect 33254 8678 33256 8730
rect 33010 8676 33016 8678
rect 33072 8676 33096 8678
rect 33152 8676 33176 8678
rect 33232 8676 33256 8678
rect 33312 8676 33318 8678
rect 33010 8667 33318 8676
rect 33010 7644 33318 7653
rect 33010 7642 33016 7644
rect 33072 7642 33096 7644
rect 33152 7642 33176 7644
rect 33232 7642 33256 7644
rect 33312 7642 33318 7644
rect 33072 7590 33074 7642
rect 33254 7590 33256 7642
rect 33010 7588 33016 7590
rect 33072 7588 33096 7590
rect 33152 7588 33176 7590
rect 33232 7588 33256 7590
rect 33312 7588 33318 7590
rect 33010 7579 33318 7588
rect 33428 7546 33456 9658
rect 33600 8900 33652 8906
rect 33600 8842 33652 8848
rect 33612 8498 33640 8842
rect 33704 8634 33732 11194
rect 33784 10464 33836 10470
rect 33784 10406 33836 10412
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33508 7744 33560 7750
rect 33508 7686 33560 7692
rect 33048 7540 33100 7546
rect 33048 7482 33100 7488
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 33060 7410 33088 7482
rect 33048 7404 33100 7410
rect 33048 7346 33100 7352
rect 33520 7342 33548 7686
rect 33508 7336 33560 7342
rect 33508 7278 33560 7284
rect 33416 6792 33468 6798
rect 33416 6734 33468 6740
rect 32864 6724 32916 6730
rect 32864 6666 32916 6672
rect 32772 6656 32824 6662
rect 32772 6598 32824 6604
rect 32784 6254 32812 6598
rect 33010 6556 33318 6565
rect 33010 6554 33016 6556
rect 33072 6554 33096 6556
rect 33152 6554 33176 6556
rect 33232 6554 33256 6556
rect 33312 6554 33318 6556
rect 33072 6502 33074 6554
rect 33254 6502 33256 6554
rect 33010 6500 33016 6502
rect 33072 6500 33096 6502
rect 33152 6500 33176 6502
rect 33232 6500 33256 6502
rect 33312 6500 33318 6502
rect 33010 6491 33318 6500
rect 33428 6458 33456 6734
rect 33692 6656 33744 6662
rect 33692 6598 33744 6604
rect 33416 6452 33468 6458
rect 33416 6394 33468 6400
rect 33414 6352 33470 6361
rect 33470 6296 33548 6304
rect 33414 6287 33416 6296
rect 33468 6276 33548 6296
rect 33416 6258 33468 6264
rect 32772 6248 32824 6254
rect 32772 6190 32824 6196
rect 32600 5902 32720 5930
rect 32496 5772 32548 5778
rect 32496 5714 32548 5720
rect 32140 5646 32272 5652
rect 32310 5672 32366 5681
rect 32140 5630 32260 5646
rect 32140 5574 32168 5630
rect 32310 5607 32366 5616
rect 32128 5568 32180 5574
rect 32128 5510 32180 5516
rect 32220 5228 32272 5234
rect 32220 5170 32272 5176
rect 32232 5030 32260 5170
rect 32312 5160 32364 5166
rect 32310 5128 32312 5137
rect 32364 5128 32366 5137
rect 32310 5063 32366 5072
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 31760 4276 31812 4282
rect 31760 4218 31812 4224
rect 31206 4111 31262 4120
rect 31392 4140 31444 4146
rect 31116 4082 31168 4088
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 31022 3904 31078 3913
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 30852 2990 30880 3878
rect 31022 3839 31078 3848
rect 31036 3602 31064 3839
rect 31024 3596 31076 3602
rect 31024 3538 31076 3544
rect 31220 3534 31248 4111
rect 31392 4082 31444 4088
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 31404 4049 31432 4082
rect 31390 4040 31446 4049
rect 31390 3975 31446 3984
rect 31576 3936 31628 3942
rect 31576 3878 31628 3884
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 30840 2984 30892 2990
rect 30840 2926 30892 2932
rect 30852 2514 30880 2926
rect 30840 2508 30892 2514
rect 30840 2450 30892 2456
rect 31220 1737 31248 3470
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 31404 3058 31432 3334
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 31496 2774 31524 2926
rect 31312 2746 31524 2774
rect 31206 1728 31262 1737
rect 31206 1663 31262 1672
rect 31116 1216 31168 1222
rect 31116 1158 31168 1164
rect 30656 740 30708 746
rect 30656 682 30708 688
rect 30472 604 30524 610
rect 30472 546 30524 552
rect 30840 468 30892 474
rect 30840 410 30892 416
rect 30564 332 30616 338
rect 30564 274 30616 280
rect 30576 56 30604 274
rect 30852 56 30880 410
rect 31128 56 31156 1158
rect 31312 202 31340 2746
rect 31484 2508 31536 2514
rect 31484 2450 31536 2456
rect 31392 604 31444 610
rect 31392 546 31444 552
rect 31300 196 31352 202
rect 31300 138 31352 144
rect 31404 56 31432 546
rect 31496 66 31524 2450
rect 31588 950 31616 3878
rect 31668 3596 31720 3602
rect 31720 3556 31800 3584
rect 31668 3538 31720 3544
rect 31772 2582 31800 3556
rect 31864 3194 31892 4694
rect 32416 4690 32444 4762
rect 32128 4684 32180 4690
rect 32128 4626 32180 4632
rect 32404 4684 32456 4690
rect 32508 4672 32536 5714
rect 32600 5137 32628 5902
rect 32864 5840 32916 5846
rect 32864 5782 32916 5788
rect 32680 5772 32732 5778
rect 32680 5714 32732 5720
rect 32692 5545 32720 5714
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32678 5536 32734 5545
rect 32678 5471 32734 5480
rect 32680 5364 32732 5370
rect 32680 5306 32732 5312
rect 32586 5128 32642 5137
rect 32586 5063 32642 5072
rect 32588 5024 32640 5030
rect 32588 4966 32640 4972
rect 32600 4865 32628 4966
rect 32586 4856 32642 4865
rect 32586 4791 32642 4800
rect 32508 4656 32628 4672
rect 32508 4650 32640 4656
rect 32508 4644 32588 4650
rect 32404 4626 32456 4632
rect 31942 4448 31998 4457
rect 31942 4383 31998 4392
rect 31956 4049 31984 4383
rect 31942 4040 31998 4049
rect 32140 4010 32168 4626
rect 32588 4592 32640 4598
rect 32220 4480 32272 4486
rect 32220 4422 32272 4428
rect 32232 4078 32260 4422
rect 32402 4312 32458 4321
rect 32402 4247 32458 4256
rect 32496 4276 32548 4282
rect 32220 4072 32272 4078
rect 32220 4014 32272 4020
rect 31942 3975 31998 3984
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 32312 3936 32364 3942
rect 32312 3878 32364 3884
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 32048 3534 32076 3674
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 31956 3369 31984 3470
rect 31942 3360 31998 3369
rect 31942 3295 31998 3304
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31944 3188 31996 3194
rect 31944 3130 31996 3136
rect 31852 2984 31904 2990
rect 31852 2926 31904 2932
rect 31760 2576 31812 2582
rect 31760 2518 31812 2524
rect 31864 1426 31892 2926
rect 31956 2854 31984 3130
rect 32140 2990 32168 3674
rect 32128 2984 32180 2990
rect 32128 2926 32180 2932
rect 31944 2848 31996 2854
rect 31944 2790 31996 2796
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 32220 2644 32272 2650
rect 32220 2586 32272 2592
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 31956 1970 31984 2382
rect 31944 1964 31996 1970
rect 31944 1906 31996 1912
rect 31852 1420 31904 1426
rect 31852 1362 31904 1368
rect 31944 1012 31996 1018
rect 31944 954 31996 960
rect 31576 944 31628 950
rect 31576 886 31628 892
rect 31668 944 31720 950
rect 31668 886 31720 892
rect 31484 60 31536 66
rect 24044 14 24164 42
rect 24214 0 24270 56
rect 24490 0 24546 56
rect 24766 0 24822 56
rect 25042 0 25098 56
rect 25318 0 25374 56
rect 25594 0 25650 56
rect 25870 0 25926 56
rect 26146 0 26202 56
rect 26422 0 26478 56
rect 26698 0 26754 56
rect 26974 0 27030 56
rect 27250 0 27306 56
rect 27526 0 27582 56
rect 27802 0 27858 56
rect 28078 0 28134 56
rect 28354 0 28410 56
rect 28630 0 28686 56
rect 28906 0 28962 56
rect 29182 0 29238 56
rect 29458 0 29514 56
rect 29734 0 29790 56
rect 30010 0 30066 56
rect 30286 0 30342 56
rect 30562 0 30618 56
rect 30838 0 30894 56
rect 31114 0 31170 56
rect 31390 0 31446 56
rect 31680 56 31708 886
rect 31956 56 31984 954
rect 32232 56 32260 2586
rect 32324 882 32352 3878
rect 32416 2446 32444 4247
rect 32496 4218 32548 4224
rect 32508 4146 32536 4218
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32692 4026 32720 5306
rect 32784 4826 32812 5646
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 32588 4004 32640 4010
rect 32692 3998 32812 4026
rect 32588 3946 32640 3952
rect 32600 3369 32628 3946
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32586 3360 32642 3369
rect 32586 3295 32642 3304
rect 32404 2440 32456 2446
rect 32692 2394 32720 3878
rect 32784 2774 32812 3998
rect 32876 3534 32904 5782
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33010 5468 33318 5477
rect 33010 5466 33016 5468
rect 33072 5466 33096 5468
rect 33152 5466 33176 5468
rect 33232 5466 33256 5468
rect 33312 5466 33318 5468
rect 33072 5414 33074 5466
rect 33254 5414 33256 5466
rect 33010 5412 33016 5414
rect 33072 5412 33096 5414
rect 33152 5412 33176 5414
rect 33232 5412 33256 5414
rect 33312 5412 33318 5414
rect 33010 5403 33318 5412
rect 32956 5364 33008 5370
rect 32956 5306 33008 5312
rect 32968 5030 32996 5306
rect 33048 5296 33100 5302
rect 33048 5238 33100 5244
rect 32956 5024 33008 5030
rect 33060 5001 33088 5238
rect 32956 4966 33008 4972
rect 33046 4992 33102 5001
rect 33046 4927 33102 4936
rect 33010 4380 33318 4389
rect 33010 4378 33016 4380
rect 33072 4378 33096 4380
rect 33152 4378 33176 4380
rect 33232 4378 33256 4380
rect 33312 4378 33318 4380
rect 33072 4326 33074 4378
rect 33254 4326 33256 4378
rect 33010 4324 33016 4326
rect 33072 4324 33096 4326
rect 33152 4324 33176 4326
rect 33232 4324 33256 4326
rect 33312 4324 33318 4326
rect 33010 4315 33318 4324
rect 33140 4208 33192 4214
rect 33192 4156 33364 4162
rect 33140 4150 33364 4156
rect 33152 4146 33364 4150
rect 33152 4140 33376 4146
rect 33152 4134 33324 4140
rect 33324 4082 33376 4088
rect 32864 3528 32916 3534
rect 32864 3470 32916 3476
rect 33322 3496 33378 3505
rect 33322 3431 33378 3440
rect 33336 3398 33364 3431
rect 33324 3392 33376 3398
rect 33324 3334 33376 3340
rect 33010 3292 33318 3301
rect 33010 3290 33016 3292
rect 33072 3290 33096 3292
rect 33152 3290 33176 3292
rect 33232 3290 33256 3292
rect 33312 3290 33318 3292
rect 33072 3238 33074 3290
rect 33254 3238 33256 3290
rect 33010 3236 33016 3238
rect 33072 3236 33096 3238
rect 33152 3236 33176 3238
rect 33232 3236 33256 3238
rect 33312 3236 33318 3238
rect 33010 3227 33318 3236
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 32784 2746 32996 2774
rect 32968 2582 32996 2746
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 33336 2514 33364 3130
rect 33428 2650 33456 5646
rect 33520 5370 33548 6276
rect 33704 6254 33732 6598
rect 33692 6248 33744 6254
rect 33692 6190 33744 6196
rect 33796 5930 33824 10406
rect 33966 10296 34022 10305
rect 33966 10231 34022 10240
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33704 5902 33824 5930
rect 33508 5364 33560 5370
rect 33508 5306 33560 5312
rect 33704 4826 33732 5902
rect 33888 5846 33916 8434
rect 33980 8090 34008 10231
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 34334 10024 34390 10033
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33968 7880 34020 7886
rect 33968 7822 34020 7828
rect 33980 7546 34008 7822
rect 33968 7540 34020 7546
rect 33968 7482 34020 7488
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 33876 5840 33928 5846
rect 33782 5808 33838 5817
rect 33876 5782 33928 5788
rect 33782 5743 33838 5752
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 33692 4140 33744 4146
rect 33692 4082 33744 4088
rect 33508 3664 33560 3670
rect 33508 3606 33560 3612
rect 33416 2644 33468 2650
rect 33416 2586 33468 2592
rect 33324 2508 33376 2514
rect 33324 2450 33376 2456
rect 32404 2382 32456 2388
rect 32600 2366 32720 2394
rect 32496 2100 32548 2106
rect 32496 2042 32548 2048
rect 32312 876 32364 882
rect 32312 818 32364 824
rect 32508 56 32536 2042
rect 32600 474 32628 2366
rect 32680 2304 32732 2310
rect 32680 2246 32732 2252
rect 32772 2304 32824 2310
rect 32772 2246 32824 2252
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 32692 1086 32720 2246
rect 32784 1290 32812 2246
rect 33010 2204 33318 2213
rect 33010 2202 33016 2204
rect 33072 2202 33096 2204
rect 33152 2202 33176 2204
rect 33232 2202 33256 2204
rect 33312 2202 33318 2204
rect 33072 2150 33074 2202
rect 33254 2150 33256 2202
rect 33010 2148 33016 2150
rect 33072 2148 33096 2150
rect 33152 2148 33176 2150
rect 33232 2148 33256 2150
rect 33312 2148 33318 2150
rect 33010 2139 33318 2148
rect 32772 1284 32824 1290
rect 32772 1226 32824 1232
rect 32680 1080 32732 1086
rect 32680 1022 32732 1028
rect 33048 808 33100 814
rect 33048 750 33100 756
rect 32588 468 32640 474
rect 32588 410 32640 416
rect 32770 232 32826 241
rect 32770 167 32826 176
rect 32784 56 32812 167
rect 33060 56 33088 750
rect 33428 270 33456 2246
rect 33520 1358 33548 3606
rect 33704 3194 33732 4082
rect 33796 3194 33824 5743
rect 33876 4820 33928 4826
rect 33876 4762 33928 4768
rect 33692 3188 33744 3194
rect 33692 3130 33744 3136
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33612 2038 33640 2926
rect 33888 2774 33916 4762
rect 33796 2746 33916 2774
rect 33796 2650 33824 2746
rect 33784 2644 33836 2650
rect 33784 2586 33836 2592
rect 33980 2582 34008 7346
rect 34072 6798 34100 9998
rect 34244 9988 34296 9994
rect 34334 9959 34390 9968
rect 34244 9930 34296 9936
rect 34152 8016 34204 8022
rect 34152 7958 34204 7964
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 34060 5568 34112 5574
rect 34060 5510 34112 5516
rect 34072 5234 34100 5510
rect 34060 5228 34112 5234
rect 34060 5170 34112 5176
rect 34060 3936 34112 3942
rect 34060 3878 34112 3884
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 33968 2576 34020 2582
rect 33968 2518 34020 2524
rect 33704 2038 33732 2518
rect 34072 2378 34100 3878
rect 34164 3058 34192 7958
rect 34256 7546 34284 9930
rect 34244 7540 34296 7546
rect 34244 7482 34296 7488
rect 34348 7478 34376 9959
rect 34428 9920 34480 9926
rect 34428 9862 34480 9868
rect 34440 8294 34468 9862
rect 34808 8634 34836 11194
rect 35624 10192 35676 10198
rect 35624 10134 35676 10140
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 35164 8492 35216 8498
rect 35164 8434 35216 8440
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34428 8084 34480 8090
rect 34428 8026 34480 8032
rect 34336 7472 34388 7478
rect 34336 7414 34388 7420
rect 34334 6896 34390 6905
rect 34334 6831 34390 6840
rect 34244 6792 34296 6798
rect 34244 6734 34296 6740
rect 34256 6118 34284 6734
rect 34244 6112 34296 6118
rect 34244 6054 34296 6060
rect 34348 5302 34376 6831
rect 34336 5296 34388 5302
rect 34336 5238 34388 5244
rect 34348 4214 34376 5238
rect 34440 4826 34468 8026
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34808 7449 34836 7822
rect 34888 7744 34940 7750
rect 34888 7686 34940 7692
rect 34794 7440 34850 7449
rect 34612 7404 34664 7410
rect 34794 7375 34850 7384
rect 34612 7346 34664 7352
rect 34624 7002 34652 7346
rect 34612 6996 34664 7002
rect 34664 6956 34744 6984
rect 34612 6938 34664 6944
rect 34612 6792 34664 6798
rect 34518 6760 34574 6769
rect 34612 6734 34664 6740
rect 34518 6695 34574 6704
rect 34532 6322 34560 6695
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34532 4826 34560 5578
rect 34624 5370 34652 6734
rect 34716 5914 34744 6956
rect 34808 6730 34836 7375
rect 34796 6724 34848 6730
rect 34796 6666 34848 6672
rect 34704 5908 34756 5914
rect 34704 5850 34756 5856
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 34808 5234 34836 6666
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 34610 5128 34666 5137
rect 34610 5063 34666 5072
rect 34428 4820 34480 4826
rect 34428 4762 34480 4768
rect 34520 4820 34572 4826
rect 34520 4762 34572 4768
rect 34428 4684 34480 4690
rect 34428 4626 34480 4632
rect 34336 4208 34388 4214
rect 34336 4150 34388 4156
rect 34244 4140 34296 4146
rect 34244 4082 34296 4088
rect 34256 3738 34284 4082
rect 34336 4072 34388 4078
rect 34440 4049 34468 4626
rect 34520 4072 34572 4078
rect 34336 4014 34388 4020
rect 34426 4040 34482 4049
rect 34348 3738 34376 4014
rect 34520 4014 34572 4020
rect 34426 3975 34482 3984
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 34336 3732 34388 3738
rect 34336 3674 34388 3680
rect 34440 3602 34468 3975
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34532 3398 34560 4014
rect 34624 3670 34652 5063
rect 34808 4622 34836 5170
rect 34796 4616 34848 4622
rect 34702 4584 34758 4593
rect 34796 4558 34848 4564
rect 34702 4519 34704 4528
rect 34756 4519 34758 4528
rect 34704 4490 34756 4496
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34794 3632 34850 3641
rect 34794 3567 34850 3576
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 34532 3194 34560 3334
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 34612 2848 34664 2854
rect 34612 2790 34664 2796
rect 34624 2666 34652 2790
rect 34532 2638 34652 2666
rect 34060 2372 34112 2378
rect 34060 2314 34112 2320
rect 33784 2304 33836 2310
rect 33784 2246 33836 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 33600 2032 33652 2038
rect 33600 1974 33652 1980
rect 33692 2032 33744 2038
rect 33692 1974 33744 1980
rect 33796 1601 33824 2246
rect 33782 1592 33838 1601
rect 33782 1527 33838 1536
rect 33508 1352 33560 1358
rect 33508 1294 33560 1300
rect 34164 1154 34192 2246
rect 34428 2100 34480 2106
rect 34428 2042 34480 2048
rect 34244 1420 34296 1426
rect 34244 1362 34296 1368
rect 34152 1148 34204 1154
rect 34152 1090 34204 1096
rect 34256 1034 34284 1362
rect 34164 1006 34284 1034
rect 33876 944 33928 950
rect 33876 886 33928 892
rect 33600 400 33652 406
rect 33600 342 33652 348
rect 33416 264 33468 270
rect 33416 206 33468 212
rect 33322 96 33378 105
rect 31484 2 31536 8
rect 31666 0 31722 56
rect 31942 0 31998 56
rect 32218 0 32274 56
rect 32494 0 32550 56
rect 32770 0 32826 56
rect 33046 0 33102 56
rect 33612 56 33640 342
rect 33888 56 33916 886
rect 34164 56 34192 1006
rect 34440 56 34468 2042
rect 34532 1329 34560 2638
rect 34716 2530 34744 3470
rect 34808 3058 34836 3567
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 34900 2774 34928 7686
rect 34980 7404 35032 7410
rect 34980 7346 35032 7352
rect 34992 5574 35020 7346
rect 35072 6792 35124 6798
rect 35072 6734 35124 6740
rect 35084 6458 35112 6734
rect 35072 6452 35124 6458
rect 35072 6394 35124 6400
rect 35176 5914 35204 8434
rect 35268 7274 35296 9386
rect 35346 8392 35402 8401
rect 35346 8327 35402 8336
rect 35360 7274 35388 8327
rect 35440 7404 35492 7410
rect 35440 7346 35492 7352
rect 35256 7268 35308 7274
rect 35256 7210 35308 7216
rect 35348 7268 35400 7274
rect 35348 7210 35400 7216
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 35360 6338 35388 6598
rect 35452 6458 35480 7346
rect 35532 6724 35584 6730
rect 35532 6666 35584 6672
rect 35440 6452 35492 6458
rect 35440 6394 35492 6400
rect 35360 6310 35480 6338
rect 35452 6254 35480 6310
rect 35440 6248 35492 6254
rect 35440 6190 35492 6196
rect 35072 5908 35124 5914
rect 35072 5850 35124 5856
rect 35164 5908 35216 5914
rect 35164 5850 35216 5856
rect 35084 5710 35112 5850
rect 35072 5704 35124 5710
rect 35072 5646 35124 5652
rect 35254 5672 35310 5681
rect 34980 5568 35032 5574
rect 34980 5510 35032 5516
rect 35084 4146 35112 5646
rect 35254 5607 35310 5616
rect 35164 4820 35216 4826
rect 35164 4762 35216 4768
rect 35072 4140 35124 4146
rect 35072 4082 35124 4088
rect 35084 3602 35112 4082
rect 35072 3596 35124 3602
rect 35072 3538 35124 3544
rect 35176 3534 35204 4762
rect 35164 3528 35216 3534
rect 35164 3470 35216 3476
rect 35268 3466 35296 5607
rect 35348 5024 35400 5030
rect 35348 4966 35400 4972
rect 35256 3460 35308 3466
rect 35256 3402 35308 3408
rect 34980 3392 35032 3398
rect 34980 3334 35032 3340
rect 34624 2502 34744 2530
rect 34808 2746 34928 2774
rect 34624 1873 34652 2502
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 34610 1864 34666 1873
rect 34610 1799 34666 1808
rect 34716 1698 34744 2382
rect 34704 1692 34756 1698
rect 34704 1634 34756 1640
rect 34612 1488 34664 1494
rect 34612 1430 34664 1436
rect 34518 1320 34574 1329
rect 34518 1255 34574 1264
rect 34624 338 34652 1430
rect 34704 1080 34756 1086
rect 34704 1022 34756 1028
rect 34612 332 34664 338
rect 34612 274 34664 280
rect 34716 56 34744 1022
rect 34808 950 34836 2746
rect 34888 2304 34940 2310
rect 34888 2246 34940 2252
rect 34796 944 34848 950
rect 34796 886 34848 892
rect 34900 542 34928 2246
rect 34992 1306 35020 3334
rect 35360 3058 35388 4966
rect 35452 3194 35480 6190
rect 35440 3188 35492 3194
rect 35440 3130 35492 3136
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 35164 2848 35216 2854
rect 35164 2790 35216 2796
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 35072 2440 35124 2446
rect 35072 2382 35124 2388
rect 35176 2394 35204 2790
rect 35084 1902 35112 2382
rect 35176 2366 35296 2394
rect 35164 2304 35216 2310
rect 35164 2246 35216 2252
rect 35072 1896 35124 1902
rect 35072 1838 35124 1844
rect 34992 1278 35112 1306
rect 34980 1148 35032 1154
rect 34980 1090 35032 1096
rect 34888 536 34940 542
rect 34888 478 34940 484
rect 34992 56 35020 1090
rect 35084 1018 35112 1278
rect 35176 1057 35204 2246
rect 35268 1494 35296 2366
rect 35256 1488 35308 1494
rect 35256 1430 35308 1436
rect 35256 1284 35308 1290
rect 35256 1226 35308 1232
rect 35162 1048 35218 1057
rect 35072 1012 35124 1018
rect 35162 983 35218 992
rect 35072 954 35124 960
rect 35268 56 35296 1226
rect 35360 610 35388 2790
rect 35440 2440 35492 2446
rect 35440 2382 35492 2388
rect 35452 1465 35480 2382
rect 35438 1456 35494 1465
rect 35438 1391 35494 1400
rect 35348 604 35400 610
rect 35348 546 35400 552
rect 35544 56 35572 6666
rect 35636 3534 35664 10134
rect 35808 9036 35860 9042
rect 35808 8978 35860 8984
rect 35820 8022 35848 8978
rect 35912 8634 35940 11194
rect 37016 11098 37044 11194
rect 37108 11098 37136 11206
rect 37016 11070 37136 11098
rect 37186 10568 37242 10577
rect 37186 10503 37242 10512
rect 36450 10432 36506 10441
rect 36450 10367 36506 10376
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 35992 9852 36044 9858
rect 35992 9794 36044 9800
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 35808 8016 35860 8022
rect 35808 7958 35860 7964
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35728 7342 35756 7822
rect 35716 7336 35768 7342
rect 35716 7278 35768 7284
rect 35716 6656 35768 6662
rect 35716 6598 35768 6604
rect 35808 6656 35860 6662
rect 35808 6598 35860 6604
rect 35728 6390 35756 6598
rect 35716 6384 35768 6390
rect 35716 6326 35768 6332
rect 35716 5840 35768 5846
rect 35716 5782 35768 5788
rect 35624 3528 35676 3534
rect 35624 3470 35676 3476
rect 35728 3398 35756 5782
rect 35820 5001 35848 6598
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 35912 6361 35940 6394
rect 35898 6352 35954 6361
rect 35898 6287 35954 6296
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35912 5302 35940 5510
rect 35900 5296 35952 5302
rect 35900 5238 35952 5244
rect 35806 4992 35862 5001
rect 35806 4927 35862 4936
rect 35898 4856 35954 4865
rect 35898 4791 35954 4800
rect 35716 3392 35768 3398
rect 35716 3334 35768 3340
rect 35808 3188 35860 3194
rect 35808 3130 35860 3136
rect 35714 3088 35770 3097
rect 35820 3058 35848 3130
rect 35714 3023 35716 3032
rect 35768 3023 35770 3032
rect 35808 3052 35860 3058
rect 35716 2994 35768 3000
rect 35808 2994 35860 3000
rect 35912 2553 35940 4791
rect 36004 3194 36032 9794
rect 36096 5642 36124 10066
rect 36360 8900 36412 8906
rect 36360 8842 36412 8848
rect 36176 8560 36228 8566
rect 36176 8502 36228 8508
rect 36188 8090 36216 8502
rect 36176 8084 36228 8090
rect 36176 8026 36228 8032
rect 36268 7880 36320 7886
rect 36268 7822 36320 7828
rect 36176 6248 36228 6254
rect 36176 6190 36228 6196
rect 36084 5636 36136 5642
rect 36084 5578 36136 5584
rect 36188 5370 36216 6190
rect 36176 5364 36228 5370
rect 36176 5306 36228 5312
rect 36174 4176 36230 4185
rect 36174 4111 36176 4120
rect 36228 4111 36230 4120
rect 36176 4082 36228 4088
rect 35992 3188 36044 3194
rect 35992 3130 36044 3136
rect 36084 2984 36136 2990
rect 36084 2926 36136 2932
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 35898 2544 35954 2553
rect 35898 2479 35954 2488
rect 35624 2304 35676 2310
rect 35624 2246 35676 2252
rect 35636 678 35664 2246
rect 36004 1850 36032 2790
rect 36096 1970 36124 2926
rect 36176 2304 36228 2310
rect 36176 2246 36228 2252
rect 36084 1964 36136 1970
rect 36084 1906 36136 1912
rect 36004 1822 36124 1850
rect 36096 814 36124 1822
rect 36084 808 36136 814
rect 36188 785 36216 2246
rect 36280 1154 36308 7822
rect 36372 4214 36400 8842
rect 36464 5574 36492 10367
rect 36636 9376 36688 9382
rect 36636 9318 36688 9324
rect 36648 8634 36676 9318
rect 37200 9314 37228 10503
rect 37188 9308 37240 9314
rect 37188 9250 37240 9256
rect 36820 9240 36872 9246
rect 36820 9182 36872 9188
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 36636 8492 36688 8498
rect 36636 8434 36688 8440
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 36360 2916 36412 2922
rect 36360 2858 36412 2864
rect 36372 2446 36400 2858
rect 36452 2576 36504 2582
rect 36452 2518 36504 2524
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 36360 1352 36412 1358
rect 36360 1294 36412 1300
rect 36268 1148 36320 1154
rect 36268 1090 36320 1096
rect 36084 750 36136 756
rect 36174 776 36230 785
rect 36174 711 36230 720
rect 35624 672 35676 678
rect 35624 614 35676 620
rect 35808 672 35860 678
rect 35808 614 35860 620
rect 35820 56 35848 614
rect 36084 536 36136 542
rect 36084 478 36136 484
rect 36096 56 36124 478
rect 36372 56 36400 1294
rect 36464 1222 36492 2518
rect 36556 2106 36584 7346
rect 36648 6633 36676 8434
rect 36832 8090 36860 9182
rect 37002 9072 37058 9081
rect 37002 9007 37058 9016
rect 36912 8832 36964 8838
rect 36912 8774 36964 8780
rect 36820 8084 36872 8090
rect 36820 8026 36872 8032
rect 36728 7268 36780 7274
rect 36728 7210 36780 7216
rect 36634 6624 36690 6633
rect 36634 6559 36690 6568
rect 36636 5160 36688 5166
rect 36636 5102 36688 5108
rect 36648 4826 36676 5102
rect 36636 4820 36688 4826
rect 36636 4762 36688 4768
rect 36636 3936 36688 3942
rect 36636 3878 36688 3884
rect 36648 2961 36676 3878
rect 36634 2952 36690 2961
rect 36740 2922 36768 7210
rect 36924 6882 36952 8774
rect 36832 6854 36952 6882
rect 36634 2887 36690 2896
rect 36728 2916 36780 2922
rect 36728 2858 36780 2864
rect 36544 2100 36596 2106
rect 36544 2042 36596 2048
rect 36832 1426 36860 6854
rect 37016 6066 37044 9007
rect 37292 8634 37320 11206
rect 38106 11194 38162 11250
rect 39210 11194 39266 11250
rect 37372 8968 37424 8974
rect 37372 8910 37424 8916
rect 37280 8628 37332 8634
rect 37280 8570 37332 8576
rect 37096 8424 37148 8430
rect 37096 8366 37148 8372
rect 37108 6186 37136 8366
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 37292 7546 37320 7686
rect 37384 7546 37412 8910
rect 37740 8900 37792 8906
rect 37740 8842 37792 8848
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37280 7540 37332 7546
rect 37280 7482 37332 7488
rect 37372 7540 37424 7546
rect 37372 7482 37424 7488
rect 37372 6316 37424 6322
rect 37372 6258 37424 6264
rect 37096 6180 37148 6186
rect 37096 6122 37148 6128
rect 37016 6038 37320 6066
rect 37004 4616 37056 4622
rect 37004 4558 37056 4564
rect 37096 4616 37148 4622
rect 37096 4558 37148 4564
rect 36912 4480 36964 4486
rect 36912 4422 36964 4428
rect 36820 1420 36872 1426
rect 36820 1362 36872 1368
rect 36452 1216 36504 1222
rect 36452 1158 36504 1164
rect 36636 196 36688 202
rect 36636 138 36688 144
rect 36648 56 36676 138
rect 36924 56 36952 4422
rect 37016 1086 37044 4558
rect 37108 3194 37136 4558
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 37096 3188 37148 3194
rect 37096 3130 37148 3136
rect 37200 1290 37228 4082
rect 37292 4010 37320 6038
rect 37280 4004 37332 4010
rect 37280 3946 37332 3952
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37292 1358 37320 2994
rect 37280 1352 37332 1358
rect 37280 1294 37332 1300
rect 37188 1284 37240 1290
rect 37188 1226 37240 1232
rect 37004 1080 37056 1086
rect 37004 1022 37056 1028
rect 37200 56 37320 82
rect 33322 0 33378 40
rect 33598 0 33654 56
rect 33874 0 33930 56
rect 34150 0 34206 56
rect 34426 0 34482 56
rect 34702 0 34758 56
rect 34978 0 35034 56
rect 35254 0 35310 56
rect 35530 0 35586 56
rect 35806 0 35862 56
rect 36082 0 36138 56
rect 36358 0 36414 56
rect 36634 0 36690 56
rect 36910 0 36966 56
rect 37186 54 37320 56
rect 37186 0 37242 54
rect 37292 42 37320 54
rect 37384 42 37412 6258
rect 37476 56 37504 7822
rect 37568 6458 37596 8434
rect 37648 8424 37700 8430
rect 37648 8366 37700 8372
rect 37660 8090 37688 8366
rect 37648 8084 37700 8090
rect 37648 8026 37700 8032
rect 37752 7002 37780 8842
rect 38120 8634 38148 11194
rect 39224 9738 39252 11194
rect 39486 9888 39542 9897
rect 39486 9823 39542 9832
rect 39224 9710 39436 9738
rect 38658 9616 38714 9625
rect 38658 9551 38714 9560
rect 38382 9344 38438 9353
rect 38382 9279 38438 9288
rect 38568 9308 38620 9314
rect 38290 9072 38346 9081
rect 38290 9007 38346 9016
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 37830 8528 37886 8537
rect 37830 8463 37832 8472
rect 37884 8463 37886 8472
rect 37832 8434 37884 8440
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 37844 7954 37872 8230
rect 37950 8188 38258 8197
rect 37950 8186 37956 8188
rect 38012 8186 38036 8188
rect 38092 8186 38116 8188
rect 38172 8186 38196 8188
rect 38252 8186 38258 8188
rect 38012 8134 38014 8186
rect 38194 8134 38196 8186
rect 37950 8132 37956 8134
rect 38012 8132 38036 8134
rect 38092 8132 38116 8134
rect 38172 8132 38196 8134
rect 38252 8132 38258 8134
rect 37950 8123 38258 8132
rect 38304 8090 38332 9007
rect 38292 8084 38344 8090
rect 38292 8026 38344 8032
rect 38396 8022 38424 9279
rect 38568 9250 38620 9256
rect 38476 8832 38528 8838
rect 38476 8774 38528 8780
rect 38488 8498 38516 8774
rect 38476 8492 38528 8498
rect 38476 8434 38528 8440
rect 38476 8356 38528 8362
rect 38476 8298 38528 8304
rect 38488 8265 38516 8298
rect 38474 8256 38530 8265
rect 38474 8191 38530 8200
rect 38384 8016 38436 8022
rect 38384 7958 38436 7964
rect 37832 7948 37884 7954
rect 37832 7890 37884 7896
rect 37832 7812 37884 7818
rect 37832 7754 37884 7760
rect 37740 6996 37792 7002
rect 37740 6938 37792 6944
rect 37740 6792 37792 6798
rect 37740 6734 37792 6740
rect 37556 6452 37608 6458
rect 37556 6394 37608 6400
rect 37556 5704 37608 5710
rect 37556 5646 37608 5652
rect 37568 202 37596 5646
rect 37648 3392 37700 3398
rect 37648 3334 37700 3340
rect 37660 3194 37688 3334
rect 37648 3188 37700 3194
rect 37648 3130 37700 3136
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37660 678 37688 2926
rect 37648 672 37700 678
rect 37648 614 37700 620
rect 37556 196 37608 202
rect 37556 138 37608 144
rect 37752 56 37780 6734
rect 37844 406 37872 7754
rect 38476 7404 38528 7410
rect 38476 7346 38528 7352
rect 38488 7313 38516 7346
rect 38474 7304 38530 7313
rect 38474 7239 38530 7248
rect 37950 7100 38258 7109
rect 37950 7098 37956 7100
rect 38012 7098 38036 7100
rect 38092 7098 38116 7100
rect 38172 7098 38196 7100
rect 38252 7098 38258 7100
rect 38012 7046 38014 7098
rect 38194 7046 38196 7098
rect 37950 7044 37956 7046
rect 38012 7044 38036 7046
rect 38092 7044 38116 7046
rect 38172 7044 38196 7046
rect 38252 7044 38258 7046
rect 37950 7035 38258 7044
rect 38580 6866 38608 9250
rect 38672 8566 38700 9551
rect 38842 9480 38898 9489
rect 38842 9415 38898 9424
rect 38660 8560 38712 8566
rect 38660 8502 38712 8508
rect 38750 8528 38806 8537
rect 38856 8498 38884 9415
rect 39010 8732 39318 8741
rect 39010 8730 39016 8732
rect 39072 8730 39096 8732
rect 39152 8730 39176 8732
rect 39232 8730 39256 8732
rect 39312 8730 39318 8732
rect 39072 8678 39074 8730
rect 39254 8678 39256 8730
rect 39010 8676 39016 8678
rect 39072 8676 39096 8678
rect 39152 8676 39176 8678
rect 39232 8676 39256 8678
rect 39312 8676 39318 8678
rect 39010 8667 39318 8676
rect 39408 8634 39436 9710
rect 39396 8628 39448 8634
rect 39396 8570 39448 8576
rect 38750 8463 38806 8472
rect 38844 8492 38896 8498
rect 38658 7984 38714 7993
rect 38658 7919 38660 7928
rect 38712 7919 38714 7928
rect 38660 7890 38712 7896
rect 38658 7848 38714 7857
rect 38658 7783 38714 7792
rect 38672 7410 38700 7783
rect 38764 7546 38792 8463
rect 38844 8434 38896 8440
rect 38936 8492 38988 8498
rect 38936 8434 38988 8440
rect 38948 7834 38976 8434
rect 39028 8356 39080 8362
rect 39028 8298 39080 8304
rect 39040 7993 39068 8298
rect 39026 7984 39082 7993
rect 39026 7919 39082 7928
rect 38856 7806 38976 7834
rect 38752 7540 38804 7546
rect 38752 7482 38804 7488
rect 38660 7404 38712 7410
rect 38660 7346 38712 7352
rect 38568 6860 38620 6866
rect 38568 6802 38620 6808
rect 38476 6792 38528 6798
rect 38304 6752 38476 6780
rect 37950 6012 38258 6021
rect 37950 6010 37956 6012
rect 38012 6010 38036 6012
rect 38092 6010 38116 6012
rect 38172 6010 38196 6012
rect 38252 6010 38258 6012
rect 38012 5958 38014 6010
rect 38194 5958 38196 6010
rect 37950 5956 37956 5958
rect 38012 5956 38036 5958
rect 38092 5956 38116 5958
rect 38172 5956 38196 5958
rect 38252 5956 38258 5958
rect 37950 5947 38258 5956
rect 37950 4924 38258 4933
rect 37950 4922 37956 4924
rect 38012 4922 38036 4924
rect 38092 4922 38116 4924
rect 38172 4922 38196 4924
rect 38252 4922 38258 4924
rect 38012 4870 38014 4922
rect 38194 4870 38196 4922
rect 37950 4868 37956 4870
rect 38012 4868 38036 4870
rect 38092 4868 38116 4870
rect 38172 4868 38196 4870
rect 38252 4868 38258 4870
rect 37950 4859 38258 4868
rect 38304 4486 38332 6752
rect 38856 6746 38884 7806
rect 38936 7744 38988 7750
rect 39396 7744 39448 7750
rect 38936 7686 38988 7692
rect 39394 7712 39396 7721
rect 39448 7712 39450 7721
rect 38948 7449 38976 7686
rect 39010 7644 39318 7653
rect 39394 7647 39450 7656
rect 39010 7642 39016 7644
rect 39072 7642 39096 7644
rect 39152 7642 39176 7644
rect 39232 7642 39256 7644
rect 39312 7642 39318 7644
rect 39072 7590 39074 7642
rect 39254 7590 39256 7642
rect 39010 7588 39016 7590
rect 39072 7588 39096 7590
rect 39152 7588 39176 7590
rect 39232 7588 39256 7590
rect 39312 7588 39318 7590
rect 39010 7579 39318 7588
rect 38934 7440 38990 7449
rect 38934 7375 38990 7384
rect 39396 7200 39448 7206
rect 39394 7168 39396 7177
rect 39448 7168 39450 7177
rect 39394 7103 39450 7112
rect 38476 6734 38528 6740
rect 38764 6730 38884 6746
rect 38752 6724 38884 6730
rect 38804 6718 38884 6724
rect 38752 6666 38804 6672
rect 38384 6656 38436 6662
rect 38382 6624 38384 6633
rect 38568 6656 38620 6662
rect 38436 6624 38438 6633
rect 38382 6559 38438 6568
rect 38488 6616 38568 6644
rect 38488 5778 38516 6616
rect 39396 6656 39448 6662
rect 38568 6598 38620 6604
rect 39394 6624 39396 6633
rect 39448 6624 39450 6633
rect 39010 6556 39318 6565
rect 39394 6559 39450 6568
rect 39010 6554 39016 6556
rect 39072 6554 39096 6556
rect 39152 6554 39176 6556
rect 39232 6554 39256 6556
rect 39312 6554 39318 6556
rect 39072 6502 39074 6554
rect 39254 6502 39256 6554
rect 39010 6500 39016 6502
rect 39072 6500 39096 6502
rect 39152 6500 39176 6502
rect 39232 6500 39256 6502
rect 39312 6500 39318 6502
rect 39010 6491 39318 6500
rect 39500 6458 39528 9823
rect 39578 8800 39634 8809
rect 39578 8735 39634 8744
rect 39592 6730 39620 8735
rect 40040 7268 40092 7274
rect 40040 7210 40092 7216
rect 40052 6905 40080 7210
rect 40038 6896 40094 6905
rect 40038 6831 40094 6840
rect 39580 6724 39632 6730
rect 39580 6666 39632 6672
rect 39488 6452 39540 6458
rect 39488 6394 39540 6400
rect 39394 6352 39450 6361
rect 38752 6316 38804 6322
rect 38752 6258 38804 6264
rect 39212 6316 39264 6322
rect 39394 6287 39450 6296
rect 39212 6258 39264 6264
rect 38476 5772 38528 5778
rect 38476 5714 38528 5720
rect 38292 4480 38344 4486
rect 38292 4422 38344 4428
rect 38292 4208 38344 4214
rect 38292 4150 38344 4156
rect 37950 3836 38258 3845
rect 37950 3834 37956 3836
rect 38012 3834 38036 3836
rect 38092 3834 38116 3836
rect 38172 3834 38196 3836
rect 38252 3834 38258 3836
rect 38012 3782 38014 3834
rect 38194 3782 38196 3834
rect 37950 3780 37956 3782
rect 38012 3780 38036 3782
rect 38092 3780 38116 3782
rect 38172 3780 38196 3782
rect 38252 3780 38258 3782
rect 37950 3771 38258 3780
rect 38304 3738 38332 4150
rect 38764 4146 38792 6258
rect 39224 6225 39252 6258
rect 39210 6216 39266 6225
rect 39210 6151 39266 6160
rect 39028 6112 39080 6118
rect 39026 6080 39028 6089
rect 39080 6080 39082 6089
rect 39026 6015 39082 6024
rect 39408 5914 39436 6287
rect 39396 5908 39448 5914
rect 39396 5850 39448 5856
rect 38936 5840 38988 5846
rect 39948 5840 40000 5846
rect 38936 5782 38988 5788
rect 39394 5808 39450 5817
rect 38842 5264 38898 5273
rect 38948 5234 38976 5782
rect 39948 5782 40000 5788
rect 39394 5743 39450 5752
rect 39010 5468 39318 5477
rect 39010 5466 39016 5468
rect 39072 5466 39096 5468
rect 39152 5466 39176 5468
rect 39232 5466 39256 5468
rect 39312 5466 39318 5468
rect 39072 5414 39074 5466
rect 39254 5414 39256 5466
rect 39010 5412 39016 5414
rect 39072 5412 39096 5414
rect 39152 5412 39176 5414
rect 39232 5412 39256 5414
rect 39312 5412 39318 5414
rect 39010 5403 39318 5412
rect 39408 5370 39436 5743
rect 39960 5545 39988 5782
rect 39946 5536 40002 5545
rect 39946 5471 40002 5480
rect 39396 5364 39448 5370
rect 39396 5306 39448 5312
rect 39394 5264 39450 5273
rect 38842 5199 38844 5208
rect 38896 5199 38898 5208
rect 38936 5228 38988 5234
rect 38844 5170 38896 5176
rect 39394 5199 39450 5208
rect 38936 5170 38988 5176
rect 39028 5024 39080 5030
rect 39026 4992 39028 5001
rect 39080 4992 39082 5001
rect 39026 4927 39082 4936
rect 39408 4826 39436 5199
rect 39396 4820 39448 4826
rect 39396 4762 39448 4768
rect 39210 4720 39266 4729
rect 39210 4655 39266 4664
rect 39486 4720 39542 4729
rect 39486 4655 39542 4664
rect 39224 4622 39252 4655
rect 39212 4616 39264 4622
rect 39212 4558 39264 4564
rect 39304 4480 39356 4486
rect 39356 4457 39436 4468
rect 39356 4448 39450 4457
rect 39356 4440 39394 4448
rect 39304 4422 39356 4428
rect 39010 4380 39318 4389
rect 39394 4383 39450 4392
rect 39010 4378 39016 4380
rect 39072 4378 39096 4380
rect 39152 4378 39176 4380
rect 39232 4378 39256 4380
rect 39312 4378 39318 4380
rect 39072 4326 39074 4378
rect 39254 4326 39256 4378
rect 39010 4324 39016 4326
rect 39072 4324 39096 4326
rect 39152 4324 39176 4326
rect 39232 4324 39256 4326
rect 39312 4324 39318 4326
rect 39010 4315 39318 4324
rect 38844 4276 38896 4282
rect 38844 4218 38896 4224
rect 38752 4140 38804 4146
rect 38752 4082 38804 4088
rect 38292 3732 38344 3738
rect 38292 3674 38344 3680
rect 38016 3664 38068 3670
rect 38016 3606 38068 3612
rect 38028 3194 38056 3606
rect 38856 3534 38884 4218
rect 39394 4176 39450 4185
rect 39120 4140 39172 4146
rect 39394 4111 39450 4120
rect 39120 4082 39172 4088
rect 39028 3936 39080 3942
rect 39026 3904 39028 3913
rect 39080 3904 39082 3913
rect 39026 3839 39082 3848
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 38752 3528 38804 3534
rect 38752 3470 38804 3476
rect 38844 3528 38896 3534
rect 38844 3470 38896 3476
rect 38936 3528 38988 3534
rect 38936 3470 38988 3476
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 38304 3058 38332 3470
rect 38292 3052 38344 3058
rect 38292 2994 38344 3000
rect 37950 2748 38258 2757
rect 37950 2746 37956 2748
rect 38012 2746 38036 2748
rect 38092 2746 38116 2748
rect 38172 2746 38196 2748
rect 38252 2746 38258 2748
rect 38012 2694 38014 2746
rect 38194 2694 38196 2746
rect 37950 2692 37956 2694
rect 38012 2692 38036 2694
rect 38092 2692 38116 2694
rect 38172 2692 38196 2694
rect 38252 2692 38258 2694
rect 37950 2683 38258 2692
rect 38106 2544 38162 2553
rect 38106 2479 38162 2488
rect 38120 2446 38148 2479
rect 38108 2440 38160 2446
rect 38108 2382 38160 2388
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38672 1737 38700 2246
rect 38658 1728 38714 1737
rect 38658 1663 38714 1672
rect 38764 542 38792 3470
rect 38844 2440 38896 2446
rect 38844 2382 38896 2388
rect 38856 2038 38884 2382
rect 38844 2032 38896 2038
rect 38844 1974 38896 1980
rect 38948 1766 38976 3470
rect 39132 3466 39160 4082
rect 39408 3738 39436 4111
rect 39500 4010 39528 4655
rect 39488 4004 39540 4010
rect 39488 3946 39540 3952
rect 39396 3732 39448 3738
rect 39396 3674 39448 3680
rect 39948 3664 40000 3670
rect 39394 3632 39450 3641
rect 39948 3606 40000 3612
rect 39394 3567 39450 3576
rect 39120 3460 39172 3466
rect 39120 3402 39172 3408
rect 39010 3292 39318 3301
rect 39010 3290 39016 3292
rect 39072 3290 39096 3292
rect 39152 3290 39176 3292
rect 39232 3290 39256 3292
rect 39312 3290 39318 3292
rect 39072 3238 39074 3290
rect 39254 3238 39256 3290
rect 39010 3236 39016 3238
rect 39072 3236 39096 3238
rect 39152 3236 39176 3238
rect 39232 3236 39256 3238
rect 39312 3236 39318 3238
rect 39010 3227 39318 3236
rect 39408 3194 39436 3567
rect 39960 3369 39988 3606
rect 39946 3360 40002 3369
rect 39946 3295 40002 3304
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39394 3088 39450 3097
rect 39394 3023 39450 3032
rect 39028 2848 39080 2854
rect 39026 2816 39028 2825
rect 39080 2816 39082 2825
rect 39026 2751 39082 2760
rect 39408 2650 39436 3023
rect 39672 2916 39724 2922
rect 39672 2858 39724 2864
rect 39396 2644 39448 2650
rect 39396 2586 39448 2592
rect 39580 2576 39632 2582
rect 39684 2553 39712 2858
rect 39580 2518 39632 2524
rect 39670 2544 39726 2553
rect 39212 2440 39264 2446
rect 39210 2408 39212 2417
rect 39264 2408 39266 2417
rect 39210 2343 39266 2352
rect 39010 2204 39318 2213
rect 39010 2202 39016 2204
rect 39072 2202 39096 2204
rect 39152 2202 39176 2204
rect 39232 2202 39256 2204
rect 39312 2202 39318 2204
rect 39072 2150 39074 2202
rect 39254 2150 39256 2202
rect 39010 2148 39016 2150
rect 39072 2148 39096 2150
rect 39152 2148 39176 2150
rect 39232 2148 39256 2150
rect 39312 2148 39318 2150
rect 39010 2139 39318 2148
rect 39592 2009 39620 2518
rect 39670 2479 39726 2488
rect 40040 2372 40092 2378
rect 40040 2314 40092 2320
rect 39948 2304 40000 2310
rect 39946 2272 39948 2281
rect 40000 2272 40002 2281
rect 39946 2207 40002 2216
rect 39578 2000 39634 2009
rect 39578 1935 39634 1944
rect 38936 1760 38988 1766
rect 38936 1702 38988 1708
rect 40052 1465 40080 2314
rect 40038 1456 40094 1465
rect 40038 1391 40094 1400
rect 38752 536 38804 542
rect 38752 478 38804 484
rect 37832 400 37884 406
rect 37832 342 37884 348
rect 37292 14 37412 42
rect 37462 0 37518 56
rect 37738 0 37794 56
<< via2 >>
rect 478 1944 534 2000
rect 1398 9016 1454 9072
rect 1398 8200 1454 8256
rect 1490 7656 1546 7712
rect 1398 7384 1454 7440
rect 1674 7404 1730 7440
rect 1674 7384 1676 7404
rect 1676 7384 1728 7404
rect 1728 7384 1730 7404
rect 1490 7112 1546 7168
rect 1398 6568 1454 6624
rect 1674 6840 1730 6896
rect 1582 6296 1638 6352
rect 1398 6024 1454 6080
rect 1490 5752 1546 5808
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2226 7928 2282 7984
rect 2042 7248 2098 7304
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1766 6160 1822 6216
rect 3422 9560 3478 9616
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1950 5752 2006 5808
rect 2226 5480 2282 5536
rect 1490 4936 1546 4992
rect 1490 4392 1546 4448
rect 1490 3848 1546 3904
rect 1490 3304 1546 3360
rect 1858 5244 1860 5264
rect 1860 5244 1912 5264
rect 1912 5244 1914 5264
rect 1858 5208 1914 5244
rect 2778 8744 2834 8800
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 3330 8508 3332 8528
rect 3332 8508 3384 8528
rect 3384 8508 3386 8528
rect 3330 8472 3386 8508
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 3606 9424 3662 9480
rect 3514 8336 3570 8392
rect 3698 8200 3754 8256
rect 2686 6840 2742 6896
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2502 5072 2558 5128
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1858 4564 1860 4584
rect 1860 4564 1912 4584
rect 1912 4564 1914 4584
rect 1858 4528 1914 4564
rect 1858 4156 1860 4176
rect 1860 4156 1912 4176
rect 1912 4156 1914 4176
rect 1858 4120 1914 4156
rect 2410 4664 2466 4720
rect 2226 3984 2282 4040
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 1674 3440 1730 3496
rect 1398 2760 1454 2816
rect 1490 2488 1546 2544
rect 1214 1672 1270 1728
rect 2134 3576 2190 3632
rect 2226 3032 2282 3088
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 1858 2216 1914 2272
rect 1582 1536 1638 1592
rect 754 1400 810 1456
rect 2410 2488 2466 2544
rect 2410 2372 2466 2408
rect 2410 2352 2412 2372
rect 2412 2352 2464 2372
rect 2464 2352 2466 2372
rect 3882 9288 3938 9344
rect 4618 9152 4674 9208
rect 4434 8608 4490 8664
rect 3146 5888 3202 5944
rect 3698 6196 3700 6216
rect 3700 6196 3752 6216
rect 3752 6196 3754 6216
rect 3698 6160 3754 6196
rect 3698 6024 3754 6080
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 3422 5364 3478 5400
rect 3422 5344 3424 5364
rect 3424 5344 3476 5364
rect 3476 5344 3478 5364
rect 3606 5228 3662 5264
rect 3606 5208 3608 5228
rect 3608 5208 3660 5228
rect 3660 5208 3662 5228
rect 2778 4936 2834 4992
rect 2962 4664 3018 4720
rect 3238 4528 3294 4584
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 2870 3576 2926 3632
rect 3146 3848 3202 3904
rect 2962 3440 3018 3496
rect 3238 3440 3294 3496
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 3054 2896 3110 2952
rect 2778 2644 2834 2680
rect 2778 2624 2780 2644
rect 2780 2624 2832 2644
rect 2832 2624 2834 2644
rect 2778 1672 2834 1728
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 3606 4120 3662 4176
rect 3698 856 3754 912
rect 5538 9832 5594 9888
rect 5814 9288 5870 9344
rect 4710 7384 4766 7440
rect 4986 6976 5042 7032
rect 3882 5208 3938 5264
rect 3974 3476 3976 3496
rect 3976 3476 4028 3496
rect 4028 3476 4030 3496
rect 3974 3440 4030 3476
rect 4250 4800 4306 4856
rect 4158 3984 4214 4040
rect 4342 4664 4398 4720
rect 4894 6740 4896 6760
rect 4896 6740 4948 6760
rect 4948 6740 4950 6760
rect 4894 6704 4950 6740
rect 4526 6024 4582 6080
rect 4986 5652 4988 5672
rect 4988 5652 5040 5672
rect 5040 5652 5042 5672
rect 4986 5616 5042 5652
rect 5262 7112 5318 7168
rect 5354 6568 5410 6624
rect 4986 5480 5042 5536
rect 4710 5344 4766 5400
rect 4526 4684 4582 4720
rect 4526 4664 4528 4684
rect 4528 4664 4580 4684
rect 4580 4664 4582 4684
rect 4250 2896 4306 2952
rect 4342 1944 4398 2000
rect 4894 5344 4950 5400
rect 5170 5108 5172 5128
rect 5172 5108 5224 5128
rect 5224 5108 5226 5128
rect 5170 5072 5226 5108
rect 5078 4936 5134 4992
rect 5262 4392 5318 4448
rect 5170 4256 5226 4312
rect 5906 8200 5962 8256
rect 5722 6568 5778 6624
rect 5814 6024 5870 6080
rect 5722 5480 5778 5536
rect 5630 4800 5686 4856
rect 6366 9696 6422 9752
rect 6458 8472 6514 8528
rect 7286 10104 7342 10160
rect 6366 6860 6422 6896
rect 6366 6840 6368 6860
rect 6368 6840 6420 6860
rect 6420 6840 6422 6860
rect 5998 5480 6054 5536
rect 5998 4800 6054 4856
rect 5538 3712 5594 3768
rect 5354 3576 5410 3632
rect 4802 992 4858 1048
rect 5446 3052 5502 3088
rect 5446 3032 5448 3052
rect 5448 3032 5500 3052
rect 5500 3032 5502 3052
rect 5446 1264 5502 1320
rect 5538 584 5594 640
rect 6182 3984 6238 4040
rect 5906 3440 5962 3496
rect 6642 7248 6698 7304
rect 6458 5888 6514 5944
rect 6642 5616 6698 5672
rect 6734 4120 6790 4176
rect 7194 8372 7196 8392
rect 7196 8372 7248 8392
rect 7248 8372 7250 8392
rect 7194 8336 7250 8372
rect 7010 7112 7066 7168
rect 7194 6976 7250 7032
rect 7010 5616 7066 5672
rect 6918 5480 6974 5536
rect 7194 5344 7250 5400
rect 7010 5092 7066 5128
rect 7010 5072 7012 5092
rect 7012 5072 7064 5092
rect 7064 5072 7066 5092
rect 6642 3576 6698 3632
rect 7102 3440 7158 3496
rect 7102 2760 7158 2816
rect 7562 6860 7618 6896
rect 7562 6840 7564 6860
rect 7564 6840 7616 6860
rect 7616 6840 7618 6860
rect 8850 9968 8906 10024
rect 8390 8608 8446 8664
rect 8390 8336 8446 8392
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 7470 6024 7526 6080
rect 7654 6316 7710 6352
rect 7654 6296 7656 6316
rect 7656 6296 7708 6316
rect 7708 6296 7710 6316
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 8022 6432 8078 6488
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 8482 7248 8538 7304
rect 8574 6976 8630 7032
rect 8574 6024 8630 6080
rect 9310 8880 9366 8936
rect 9016 8730 9072 8732
rect 9096 8730 9152 8732
rect 9176 8730 9232 8732
rect 9256 8730 9312 8732
rect 9016 8678 9062 8730
rect 9062 8678 9072 8730
rect 9096 8678 9126 8730
rect 9126 8678 9138 8730
rect 9138 8678 9152 8730
rect 9176 8678 9190 8730
rect 9190 8678 9202 8730
rect 9202 8678 9232 8730
rect 9256 8678 9266 8730
rect 9266 8678 9312 8730
rect 9016 8676 9072 8678
rect 9096 8676 9152 8678
rect 9176 8676 9232 8678
rect 9256 8676 9312 8678
rect 9954 10512 10010 10568
rect 9678 9560 9734 9616
rect 9494 7928 9550 7984
rect 9494 7812 9550 7848
rect 9494 7792 9496 7812
rect 9496 7792 9548 7812
rect 9548 7792 9550 7812
rect 9016 7642 9072 7644
rect 9096 7642 9152 7644
rect 9176 7642 9232 7644
rect 9256 7642 9312 7644
rect 9016 7590 9062 7642
rect 9062 7590 9072 7642
rect 9096 7590 9126 7642
rect 9126 7590 9138 7642
rect 9138 7590 9152 7642
rect 9176 7590 9190 7642
rect 9190 7590 9202 7642
rect 9202 7590 9232 7642
rect 9256 7590 9266 7642
rect 9266 7590 9312 7642
rect 9016 7588 9072 7590
rect 9096 7588 9152 7590
rect 9176 7588 9232 7590
rect 9256 7588 9312 7590
rect 10322 10376 10378 10432
rect 10138 7520 10194 7576
rect 9770 7384 9826 7440
rect 9678 6976 9734 7032
rect 8574 5652 8576 5672
rect 8576 5652 8628 5672
rect 8628 5652 8630 5672
rect 7654 4800 7710 4856
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 7746 4256 7802 4312
rect 7378 3984 7434 4040
rect 7654 3984 7710 4040
rect 7378 3732 7434 3768
rect 7378 3712 7380 3732
rect 7380 3712 7432 3732
rect 7432 3712 7434 3732
rect 7286 2216 7342 2272
rect 7378 1128 7434 1184
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 8022 3304 8078 3360
rect 8298 3304 8354 3360
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 8574 5616 8630 5652
rect 8666 5344 8722 5400
rect 9678 6568 9734 6624
rect 9016 6554 9072 6556
rect 9096 6554 9152 6556
rect 9176 6554 9232 6556
rect 9256 6554 9312 6556
rect 9016 6502 9062 6554
rect 9062 6502 9072 6554
rect 9096 6502 9126 6554
rect 9126 6502 9138 6554
rect 9138 6502 9152 6554
rect 9176 6502 9190 6554
rect 9190 6502 9202 6554
rect 9202 6502 9232 6554
rect 9256 6502 9266 6554
rect 9266 6502 9312 6554
rect 9016 6500 9072 6502
rect 9096 6500 9152 6502
rect 9176 6500 9232 6502
rect 9256 6500 9312 6502
rect 9016 5466 9072 5468
rect 9096 5466 9152 5468
rect 9176 5466 9232 5468
rect 9256 5466 9312 5468
rect 9016 5414 9062 5466
rect 9062 5414 9072 5466
rect 9096 5414 9126 5466
rect 9126 5414 9138 5466
rect 9138 5414 9152 5466
rect 9176 5414 9190 5466
rect 9190 5414 9202 5466
rect 9202 5414 9232 5466
rect 9256 5414 9266 5466
rect 9266 5414 9312 5466
rect 9016 5412 9072 5414
rect 9096 5412 9152 5414
rect 9176 5412 9232 5414
rect 9256 5412 9312 5414
rect 9016 4378 9072 4380
rect 9096 4378 9152 4380
rect 9176 4378 9232 4380
rect 9256 4378 9312 4380
rect 9016 4326 9062 4378
rect 9062 4326 9072 4378
rect 9096 4326 9126 4378
rect 9126 4326 9138 4378
rect 9138 4326 9152 4378
rect 9176 4326 9190 4378
rect 9190 4326 9202 4378
rect 9202 4326 9232 4378
rect 9256 4326 9266 4378
rect 9266 4326 9312 4378
rect 9016 4324 9072 4326
rect 9096 4324 9152 4326
rect 9176 4324 9232 4326
rect 9256 4324 9312 4326
rect 8850 3848 8906 3904
rect 9770 5752 9826 5808
rect 9770 5652 9772 5672
rect 9772 5652 9824 5672
rect 9824 5652 9826 5672
rect 9770 5616 9826 5652
rect 9770 4936 9826 4992
rect 9586 4392 9642 4448
rect 9126 3848 9182 3904
rect 10690 8064 10746 8120
rect 10782 7656 10838 7712
rect 10782 6724 10838 6760
rect 10782 6704 10784 6724
rect 10784 6704 10836 6724
rect 10836 6704 10838 6724
rect 10046 6296 10102 6352
rect 9954 4936 10010 4992
rect 10230 6024 10286 6080
rect 10138 4564 10140 4584
rect 10140 4564 10192 4584
rect 10192 4564 10194 4584
rect 10138 4528 10194 4564
rect 10046 4256 10102 4312
rect 9402 3576 9458 3632
rect 8574 3168 8630 3224
rect 8482 1264 8538 1320
rect 9016 3290 9072 3292
rect 9096 3290 9152 3292
rect 9176 3290 9232 3292
rect 9256 3290 9312 3292
rect 9016 3238 9062 3290
rect 9062 3238 9072 3290
rect 9096 3238 9126 3290
rect 9126 3238 9138 3290
rect 9138 3238 9152 3290
rect 9176 3238 9190 3290
rect 9190 3238 9202 3290
rect 9202 3238 9232 3290
rect 9256 3238 9266 3290
rect 9266 3238 9312 3290
rect 9016 3236 9072 3238
rect 9096 3236 9152 3238
rect 9176 3236 9232 3238
rect 9256 3236 9312 3238
rect 8758 3168 8814 3224
rect 9770 3340 9772 3360
rect 9772 3340 9824 3360
rect 9824 3340 9826 3360
rect 9770 3304 9826 3340
rect 10414 4936 10470 4992
rect 10046 3476 10048 3496
rect 10048 3476 10100 3496
rect 10100 3476 10102 3496
rect 10046 3440 10102 3476
rect 9126 2760 9182 2816
rect 10322 3052 10378 3088
rect 10322 3032 10324 3052
rect 10324 3032 10376 3052
rect 10376 3032 10378 3052
rect 11242 8880 11298 8936
rect 11334 8336 11390 8392
rect 11518 7656 11574 7712
rect 11150 5344 11206 5400
rect 11242 4800 11298 4856
rect 10874 4120 10930 4176
rect 11518 4256 11574 4312
rect 11886 7828 11888 7848
rect 11888 7828 11940 7848
rect 11940 7828 11942 7848
rect 11886 7792 11942 7828
rect 11702 5616 11758 5672
rect 10598 3576 10654 3632
rect 11334 3440 11390 3496
rect 10598 2896 10654 2952
rect 9016 2202 9072 2204
rect 9096 2202 9152 2204
rect 9176 2202 9232 2204
rect 9256 2202 9312 2204
rect 9016 2150 9062 2202
rect 9062 2150 9072 2202
rect 9096 2150 9126 2202
rect 9126 2150 9138 2202
rect 9138 2150 9152 2202
rect 9176 2150 9190 2202
rect 9190 2150 9202 2202
rect 9202 2150 9232 2202
rect 9256 2150 9266 2202
rect 9266 2150 9312 2202
rect 9016 2148 9072 2150
rect 9096 2148 9152 2150
rect 9176 2148 9232 2150
rect 9256 2148 9312 2150
rect 9586 2080 9642 2136
rect 11058 1944 11114 2000
rect 9678 1400 9734 1456
rect 11058 1536 11114 1592
rect 11426 3304 11482 3360
rect 11426 1808 11482 1864
rect 11242 40 11298 96
rect 11886 4936 11942 4992
rect 12070 4800 12126 4856
rect 11886 3032 11942 3088
rect 11886 1808 11942 1864
rect 12346 9016 12402 9072
rect 12530 7928 12586 7984
rect 12254 6180 12310 6216
rect 12254 6160 12256 6180
rect 12256 6160 12308 6180
rect 12308 6160 12310 6180
rect 12254 5616 12310 5672
rect 12254 4800 12310 4856
rect 12254 4120 12310 4176
rect 12162 3984 12218 4040
rect 12254 1536 12310 1592
rect 12530 6704 12586 6760
rect 12438 6568 12494 6624
rect 12438 6024 12494 6080
rect 13174 8336 13230 8392
rect 13082 7248 13138 7304
rect 12714 6316 12770 6352
rect 12714 6296 12716 6316
rect 12716 6296 12768 6316
rect 12768 6296 12770 6316
rect 12714 5480 12770 5536
rect 12898 6024 12954 6080
rect 12438 4800 12494 4856
rect 12714 3440 12770 3496
rect 12438 3032 12494 3088
rect 12622 2896 12678 2952
rect 12990 5752 13046 5808
rect 13266 6296 13322 6352
rect 13910 10240 13966 10296
rect 13542 8064 13598 8120
rect 13956 8186 14012 8188
rect 14036 8186 14092 8188
rect 14116 8186 14172 8188
rect 14196 8186 14252 8188
rect 13956 8134 14002 8186
rect 14002 8134 14012 8186
rect 14036 8134 14066 8186
rect 14066 8134 14078 8186
rect 14078 8134 14092 8186
rect 14116 8134 14130 8186
rect 14130 8134 14142 8186
rect 14142 8134 14172 8186
rect 14196 8134 14206 8186
rect 14206 8134 14252 8186
rect 13956 8132 14012 8134
rect 14036 8132 14092 8134
rect 14116 8132 14172 8134
rect 14196 8132 14252 8134
rect 13634 7384 13690 7440
rect 13956 7098 14012 7100
rect 14036 7098 14092 7100
rect 14116 7098 14172 7100
rect 14196 7098 14252 7100
rect 13956 7046 14002 7098
rect 14002 7046 14012 7098
rect 14036 7046 14066 7098
rect 14066 7046 14078 7098
rect 14078 7046 14092 7098
rect 14116 7046 14130 7098
rect 14130 7046 14142 7098
rect 14142 7046 14172 7098
rect 14196 7046 14206 7098
rect 14206 7046 14252 7098
rect 13956 7044 14012 7046
rect 14036 7044 14092 7046
rect 14116 7044 14172 7046
rect 14196 7044 14252 7046
rect 13266 5480 13322 5536
rect 13358 4548 13414 4584
rect 13358 4528 13360 4548
rect 13360 4528 13412 4548
rect 13412 4528 13414 4548
rect 13174 3848 13230 3904
rect 13174 3576 13230 3632
rect 13358 3712 13414 3768
rect 13174 2896 13230 2952
rect 13358 2216 13414 2272
rect 13542 6296 13598 6352
rect 13542 3712 13598 3768
rect 13956 6010 14012 6012
rect 14036 6010 14092 6012
rect 14116 6010 14172 6012
rect 14196 6010 14252 6012
rect 13956 5958 14002 6010
rect 14002 5958 14012 6010
rect 14036 5958 14066 6010
rect 14066 5958 14078 6010
rect 14078 5958 14092 6010
rect 14116 5958 14130 6010
rect 14130 5958 14142 6010
rect 14142 5958 14172 6010
rect 14196 5958 14206 6010
rect 14206 5958 14252 6010
rect 13956 5956 14012 5958
rect 14036 5956 14092 5958
rect 14116 5956 14172 5958
rect 14196 5956 14252 5958
rect 15106 9424 15162 9480
rect 15016 8730 15072 8732
rect 15096 8730 15152 8732
rect 15176 8730 15232 8732
rect 15256 8730 15312 8732
rect 15016 8678 15062 8730
rect 15062 8678 15072 8730
rect 15096 8678 15126 8730
rect 15126 8678 15138 8730
rect 15138 8678 15152 8730
rect 15176 8678 15190 8730
rect 15190 8678 15202 8730
rect 15202 8678 15232 8730
rect 15256 8678 15266 8730
rect 15266 8678 15312 8730
rect 15016 8676 15072 8678
rect 15096 8676 15152 8678
rect 15176 8676 15232 8678
rect 15256 8676 15312 8678
rect 14738 7540 14794 7576
rect 14738 7520 14740 7540
rect 14740 7520 14792 7540
rect 14792 7520 14794 7540
rect 14646 7384 14702 7440
rect 15016 7642 15072 7644
rect 15096 7642 15152 7644
rect 15176 7642 15232 7644
rect 15256 7642 15312 7644
rect 15016 7590 15062 7642
rect 15062 7590 15072 7642
rect 15096 7590 15126 7642
rect 15126 7590 15138 7642
rect 15138 7590 15152 7642
rect 15176 7590 15190 7642
rect 15190 7590 15202 7642
rect 15202 7590 15232 7642
rect 15256 7590 15266 7642
rect 15266 7590 15312 7642
rect 15016 7588 15072 7590
rect 15096 7588 15152 7590
rect 15176 7588 15232 7590
rect 15256 7588 15312 7590
rect 14554 6976 14610 7032
rect 14554 6840 14610 6896
rect 14554 6568 14610 6624
rect 13956 4922 14012 4924
rect 14036 4922 14092 4924
rect 14116 4922 14172 4924
rect 14196 4922 14252 4924
rect 13956 4870 14002 4922
rect 14002 4870 14012 4922
rect 14036 4870 14066 4922
rect 14066 4870 14078 4922
rect 14078 4870 14092 4922
rect 14116 4870 14130 4922
rect 14130 4870 14142 4922
rect 14142 4870 14172 4922
rect 14196 4870 14206 4922
rect 14206 4870 14252 4922
rect 13956 4868 14012 4870
rect 14036 4868 14092 4870
rect 14116 4868 14172 4870
rect 14196 4868 14252 4870
rect 15016 6554 15072 6556
rect 15096 6554 15152 6556
rect 15176 6554 15232 6556
rect 15256 6554 15312 6556
rect 15016 6502 15062 6554
rect 15062 6502 15072 6554
rect 15096 6502 15126 6554
rect 15126 6502 15138 6554
rect 15138 6502 15152 6554
rect 15176 6502 15190 6554
rect 15190 6502 15202 6554
rect 15202 6502 15232 6554
rect 15256 6502 15266 6554
rect 15266 6502 15312 6554
rect 15016 6500 15072 6502
rect 15096 6500 15152 6502
rect 15176 6500 15232 6502
rect 15256 6500 15312 6502
rect 14830 5888 14886 5944
rect 14646 5480 14702 5536
rect 14094 3984 14150 4040
rect 13956 3834 14012 3836
rect 14036 3834 14092 3836
rect 14116 3834 14172 3836
rect 14196 3834 14252 3836
rect 13956 3782 14002 3834
rect 14002 3782 14012 3834
rect 14036 3782 14066 3834
rect 14066 3782 14078 3834
rect 14078 3782 14092 3834
rect 14116 3782 14130 3834
rect 14130 3782 14142 3834
rect 14142 3782 14172 3834
rect 14196 3782 14206 3834
rect 14206 3782 14252 3834
rect 13956 3780 14012 3782
rect 14036 3780 14092 3782
rect 14116 3780 14172 3782
rect 14196 3780 14252 3782
rect 14094 3168 14150 3224
rect 14186 3032 14242 3088
rect 14094 2896 14150 2952
rect 13726 2624 13782 2680
rect 13956 2746 14012 2748
rect 14036 2746 14092 2748
rect 14116 2746 14172 2748
rect 14196 2746 14252 2748
rect 13956 2694 14002 2746
rect 14002 2694 14012 2746
rect 14036 2694 14066 2746
rect 14066 2694 14078 2746
rect 14078 2694 14092 2746
rect 14116 2694 14130 2746
rect 14130 2694 14142 2746
rect 14142 2694 14172 2746
rect 14196 2694 14206 2746
rect 14206 2694 14252 2746
rect 13956 2692 14012 2694
rect 14036 2692 14092 2694
rect 14116 2692 14172 2694
rect 14196 2692 14252 2694
rect 13910 2488 13966 2544
rect 15016 5466 15072 5468
rect 15096 5466 15152 5468
rect 15176 5466 15232 5468
rect 15256 5466 15312 5468
rect 15016 5414 15062 5466
rect 15062 5414 15072 5466
rect 15096 5414 15126 5466
rect 15126 5414 15138 5466
rect 15138 5414 15152 5466
rect 15176 5414 15190 5466
rect 15190 5414 15202 5466
rect 15202 5414 15232 5466
rect 15256 5414 15266 5466
rect 15266 5414 15312 5466
rect 15016 5412 15072 5414
rect 15096 5412 15152 5414
rect 15176 5412 15232 5414
rect 15256 5412 15312 5414
rect 15106 4972 15108 4992
rect 15108 4972 15160 4992
rect 15160 4972 15162 4992
rect 15106 4936 15162 4972
rect 15106 4564 15108 4584
rect 15108 4564 15160 4584
rect 15160 4564 15162 4584
rect 15106 4528 15162 4564
rect 15016 4378 15072 4380
rect 15096 4378 15152 4380
rect 15176 4378 15232 4380
rect 15256 4378 15312 4380
rect 15016 4326 15062 4378
rect 15062 4326 15072 4378
rect 15096 4326 15126 4378
rect 15126 4326 15138 4378
rect 15138 4326 15152 4378
rect 15176 4326 15190 4378
rect 15190 4326 15202 4378
rect 15202 4326 15232 4378
rect 15256 4326 15266 4378
rect 15266 4326 15312 4378
rect 15016 4324 15072 4326
rect 15096 4324 15152 4326
rect 15176 4324 15232 4326
rect 15256 4324 15312 4326
rect 14830 3712 14886 3768
rect 15842 9560 15898 9616
rect 15566 7656 15622 7712
rect 16118 8064 16174 8120
rect 16118 7520 16174 7576
rect 15934 6976 15990 7032
rect 15566 6840 15622 6896
rect 15566 6568 15622 6624
rect 15842 6840 15898 6896
rect 15658 6432 15714 6488
rect 15474 5344 15530 5400
rect 15474 4528 15530 4584
rect 15198 3984 15254 4040
rect 15290 3712 15346 3768
rect 14646 3304 14702 3360
rect 14646 2896 14702 2952
rect 14646 2216 14702 2272
rect 15016 3290 15072 3292
rect 15096 3290 15152 3292
rect 15176 3290 15232 3292
rect 15256 3290 15312 3292
rect 15016 3238 15062 3290
rect 15062 3238 15072 3290
rect 15096 3238 15126 3290
rect 15126 3238 15138 3290
rect 15138 3238 15152 3290
rect 15176 3238 15190 3290
rect 15190 3238 15202 3290
rect 15202 3238 15232 3290
rect 15256 3238 15266 3290
rect 15266 3238 15312 3290
rect 15016 3236 15072 3238
rect 15096 3236 15152 3238
rect 15176 3236 15232 3238
rect 15256 3236 15312 3238
rect 15106 3052 15162 3088
rect 15106 3032 15108 3052
rect 15108 3032 15160 3052
rect 15160 3032 15162 3052
rect 15842 3712 15898 3768
rect 15658 3304 15714 3360
rect 15566 3032 15622 3088
rect 15474 2624 15530 2680
rect 16486 9696 16542 9752
rect 16486 9424 16542 9480
rect 17590 9016 17646 9072
rect 17590 8744 17646 8800
rect 16486 8336 16542 8392
rect 16670 7112 16726 7168
rect 16302 6976 16358 7032
rect 16302 6296 16358 6352
rect 16026 5616 16082 5672
rect 16026 4528 16082 4584
rect 15842 2488 15898 2544
rect 15016 2202 15072 2204
rect 15096 2202 15152 2204
rect 15176 2202 15232 2204
rect 15256 2202 15312 2204
rect 15016 2150 15062 2202
rect 15062 2150 15072 2202
rect 15096 2150 15126 2202
rect 15126 2150 15138 2202
rect 15138 2150 15152 2202
rect 15176 2150 15190 2202
rect 15190 2150 15202 2202
rect 15202 2150 15232 2202
rect 15256 2150 15266 2202
rect 15266 2150 15312 2202
rect 15016 2148 15072 2150
rect 15096 2148 15152 2150
rect 15176 2148 15232 2150
rect 15256 2148 15312 2150
rect 15198 40 15254 96
rect 15842 1808 15898 1864
rect 16210 2624 16266 2680
rect 16394 4800 16450 4856
rect 16762 6976 16818 7032
rect 16854 6296 16910 6352
rect 17222 7928 17278 7984
rect 17406 6976 17462 7032
rect 17590 7112 17646 7168
rect 17314 6568 17370 6624
rect 16486 3732 16542 3768
rect 16486 3712 16488 3732
rect 16488 3712 16540 3732
rect 16540 3712 16542 3732
rect 16854 4120 16910 4176
rect 16854 3984 16910 4040
rect 16854 3168 16910 3224
rect 17222 4528 17278 4584
rect 16946 2896 17002 2952
rect 16302 1808 16358 1864
rect 16486 1536 16542 1592
rect 16486 1012 16542 1048
rect 16486 992 16488 1012
rect 16488 992 16540 1012
rect 16540 992 16542 1012
rect 16486 876 16542 912
rect 16486 856 16488 876
rect 16488 856 16540 876
rect 16540 856 16542 876
rect 16394 720 16450 776
rect 16762 1436 16764 1456
rect 16764 1436 16816 1456
rect 16816 1436 16818 1456
rect 16762 1400 16818 1436
rect 16670 856 16726 912
rect 17498 6432 17554 6488
rect 17406 4428 17408 4448
rect 17408 4428 17460 4448
rect 17460 4428 17462 4448
rect 17406 4392 17462 4428
rect 17682 6432 17738 6488
rect 17682 5616 17738 5672
rect 17958 9832 18014 9888
rect 17958 9016 18014 9072
rect 17958 7656 18014 7712
rect 18142 8064 18198 8120
rect 18142 7656 18198 7712
rect 18878 8744 18934 8800
rect 19062 8200 19118 8256
rect 17958 5752 18014 5808
rect 18142 6196 18144 6216
rect 18144 6196 18196 6216
rect 18196 6196 18198 6216
rect 18142 6160 18198 6196
rect 19062 6976 19118 7032
rect 17682 4392 17738 4448
rect 17958 4392 18014 4448
rect 17590 4020 17592 4040
rect 17592 4020 17644 4040
rect 17644 4020 17646 4040
rect 17590 3984 17646 4020
rect 17130 2216 17186 2272
rect 17866 3576 17922 3632
rect 18050 3984 18106 4040
rect 18326 5616 18382 5672
rect 20810 8744 20866 8800
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 20196 8186 20252 8188
rect 19956 8134 20002 8186
rect 20002 8134 20012 8186
rect 20036 8134 20066 8186
rect 20066 8134 20078 8186
rect 20078 8134 20092 8186
rect 20116 8134 20130 8186
rect 20130 8134 20142 8186
rect 20142 8134 20172 8186
rect 20196 8134 20206 8186
rect 20206 8134 20252 8186
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 20196 8132 20252 8134
rect 20350 8064 20406 8120
rect 19890 7540 19946 7576
rect 19890 7520 19892 7540
rect 19892 7520 19944 7540
rect 19944 7520 19946 7540
rect 20074 7520 20130 7576
rect 19614 7248 19670 7304
rect 20350 7792 20406 7848
rect 20534 8200 20590 8256
rect 20534 7656 20590 7712
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 20196 7098 20252 7100
rect 19956 7046 20002 7098
rect 20002 7046 20012 7098
rect 20036 7046 20066 7098
rect 20066 7046 20078 7098
rect 20078 7046 20092 7098
rect 20116 7046 20130 7098
rect 20130 7046 20142 7098
rect 20142 7046 20172 7098
rect 20196 7046 20206 7098
rect 20206 7046 20252 7098
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 20196 7044 20252 7046
rect 19522 6976 19578 7032
rect 21016 8730 21072 8732
rect 21096 8730 21152 8732
rect 21176 8730 21232 8732
rect 21256 8730 21312 8732
rect 21016 8678 21062 8730
rect 21062 8678 21072 8730
rect 21096 8678 21126 8730
rect 21126 8678 21138 8730
rect 21138 8678 21152 8730
rect 21176 8678 21190 8730
rect 21190 8678 21202 8730
rect 21202 8678 21232 8730
rect 21256 8678 21266 8730
rect 21266 8678 21312 8730
rect 21016 8676 21072 8678
rect 21096 8676 21152 8678
rect 21176 8676 21232 8678
rect 21256 8676 21312 8678
rect 20810 7248 20866 7304
rect 19430 5888 19486 5944
rect 18878 5480 18934 5536
rect 18418 4528 18474 4584
rect 18326 3984 18382 4040
rect 18786 4256 18842 4312
rect 18694 4120 18750 4176
rect 17774 2896 17830 2952
rect 18050 3032 18106 3088
rect 17774 2488 17830 2544
rect 18050 2624 18106 2680
rect 18142 1944 18198 2000
rect 17866 1128 17922 1184
rect 18510 3712 18566 3768
rect 18786 3712 18842 3768
rect 18786 3168 18842 3224
rect 18694 2760 18750 2816
rect 18786 2644 18842 2680
rect 18786 2624 18788 2644
rect 18788 2624 18840 2644
rect 18840 2624 18842 2644
rect 19062 3032 19118 3088
rect 19062 2760 19118 2816
rect 19062 2488 19118 2544
rect 20718 6704 20774 6760
rect 20350 6296 20406 6352
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 20196 6010 20252 6012
rect 19956 5958 20002 6010
rect 20002 5958 20012 6010
rect 20036 5958 20066 6010
rect 20066 5958 20078 6010
rect 20078 5958 20092 6010
rect 20116 5958 20130 6010
rect 20130 5958 20142 6010
rect 20142 5958 20172 6010
rect 20196 5958 20206 6010
rect 20206 5958 20252 6010
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 20196 5956 20252 5958
rect 19614 4800 19670 4856
rect 20534 5908 20590 5944
rect 20534 5888 20536 5908
rect 20536 5888 20588 5908
rect 20588 5888 20590 5908
rect 19890 5480 19946 5536
rect 20442 5480 20498 5536
rect 21454 7656 21510 7712
rect 21016 7642 21072 7644
rect 21096 7642 21152 7644
rect 21176 7642 21232 7644
rect 21256 7642 21312 7644
rect 21016 7590 21062 7642
rect 21062 7590 21072 7642
rect 21096 7590 21126 7642
rect 21126 7590 21138 7642
rect 21138 7590 21152 7642
rect 21176 7590 21190 7642
rect 21190 7590 21202 7642
rect 21202 7590 21232 7642
rect 21256 7590 21266 7642
rect 21266 7590 21312 7642
rect 21016 7588 21072 7590
rect 21096 7588 21152 7590
rect 21176 7588 21232 7590
rect 21256 7588 21312 7590
rect 21270 7384 21326 7440
rect 21178 6840 21234 6896
rect 21454 6740 21456 6760
rect 21456 6740 21508 6760
rect 21508 6740 21510 6760
rect 21454 6704 21510 6740
rect 21016 6554 21072 6556
rect 21096 6554 21152 6556
rect 21176 6554 21232 6556
rect 21256 6554 21312 6556
rect 21016 6502 21062 6554
rect 21062 6502 21072 6554
rect 21096 6502 21126 6554
rect 21126 6502 21138 6554
rect 21138 6502 21152 6554
rect 21176 6502 21190 6554
rect 21190 6502 21202 6554
rect 21202 6502 21232 6554
rect 21256 6502 21266 6554
rect 21266 6502 21312 6554
rect 21016 6500 21072 6502
rect 21096 6500 21152 6502
rect 21176 6500 21232 6502
rect 21256 6500 21312 6502
rect 21454 6568 21510 6624
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 20196 4922 20252 4924
rect 19956 4870 20002 4922
rect 20002 4870 20012 4922
rect 20036 4870 20066 4922
rect 20066 4870 20078 4922
rect 20078 4870 20092 4922
rect 20116 4870 20130 4922
rect 20130 4870 20142 4922
rect 20142 4870 20172 4922
rect 20196 4870 20206 4922
rect 20206 4870 20252 4922
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 20196 4868 20252 4870
rect 19430 3848 19486 3904
rect 19338 3576 19394 3632
rect 19338 3168 19394 3224
rect 19614 3440 19670 3496
rect 20350 3848 20406 3904
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 20196 3834 20252 3836
rect 19956 3782 20002 3834
rect 20002 3782 20012 3834
rect 20036 3782 20066 3834
rect 20066 3782 20078 3834
rect 20078 3782 20092 3834
rect 20116 3782 20130 3834
rect 20130 3782 20142 3834
rect 20142 3782 20172 3834
rect 20196 3782 20206 3834
rect 20206 3782 20252 3834
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 20196 3780 20252 3782
rect 20442 3712 20498 3768
rect 19798 3440 19854 3496
rect 20166 3476 20168 3496
rect 20168 3476 20220 3496
rect 20220 3476 20222 3496
rect 20166 3440 20222 3476
rect 20442 3576 20498 3632
rect 20350 3304 20406 3360
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 20196 2746 20252 2748
rect 19956 2694 20002 2746
rect 20002 2694 20012 2746
rect 20036 2694 20066 2746
rect 20066 2694 20078 2746
rect 20078 2694 20092 2746
rect 20116 2694 20130 2746
rect 20130 2694 20142 2746
rect 20142 2694 20172 2746
rect 20196 2694 20206 2746
rect 20206 2694 20252 2746
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 20196 2692 20252 2694
rect 19430 176 19486 232
rect 20810 4392 20866 4448
rect 20810 4256 20866 4312
rect 21016 5466 21072 5468
rect 21096 5466 21152 5468
rect 21176 5466 21232 5468
rect 21256 5466 21312 5468
rect 21016 5414 21062 5466
rect 21062 5414 21072 5466
rect 21096 5414 21126 5466
rect 21126 5414 21138 5466
rect 21138 5414 21152 5466
rect 21176 5414 21190 5466
rect 21190 5414 21202 5466
rect 21202 5414 21232 5466
rect 21256 5414 21266 5466
rect 21266 5414 21312 5466
rect 21016 5412 21072 5414
rect 21096 5412 21152 5414
rect 21176 5412 21232 5414
rect 21256 5412 21312 5414
rect 21454 4936 21510 4992
rect 21086 4800 21142 4856
rect 21362 4800 21418 4856
rect 21016 4378 21072 4380
rect 21096 4378 21152 4380
rect 21176 4378 21232 4380
rect 21256 4378 21312 4380
rect 21016 4326 21062 4378
rect 21062 4326 21072 4378
rect 21096 4326 21126 4378
rect 21126 4326 21138 4378
rect 21138 4326 21152 4378
rect 21176 4326 21190 4378
rect 21190 4326 21202 4378
rect 21202 4326 21232 4378
rect 21256 4326 21266 4378
rect 21266 4326 21312 4378
rect 21016 4324 21072 4326
rect 21096 4324 21152 4326
rect 21176 4324 21232 4326
rect 21256 4324 21312 4326
rect 20718 3188 20774 3224
rect 20718 3168 20720 3188
rect 20720 3168 20772 3188
rect 20772 3168 20774 3188
rect 21016 3290 21072 3292
rect 21096 3290 21152 3292
rect 21176 3290 21232 3292
rect 21256 3290 21312 3292
rect 21016 3238 21062 3290
rect 21062 3238 21072 3290
rect 21096 3238 21126 3290
rect 21126 3238 21138 3290
rect 21138 3238 21152 3290
rect 21176 3238 21190 3290
rect 21190 3238 21202 3290
rect 21202 3238 21232 3290
rect 21256 3238 21266 3290
rect 21266 3238 21312 3290
rect 21016 3236 21072 3238
rect 21096 3236 21152 3238
rect 21176 3236 21232 3238
rect 21256 3236 21312 3238
rect 20994 3032 21050 3088
rect 21178 3032 21234 3088
rect 20994 2760 21050 2816
rect 21016 2202 21072 2204
rect 21096 2202 21152 2204
rect 21176 2202 21232 2204
rect 21256 2202 21312 2204
rect 21016 2150 21062 2202
rect 21062 2150 21072 2202
rect 21096 2150 21126 2202
rect 21126 2150 21138 2202
rect 21138 2150 21152 2202
rect 21176 2150 21190 2202
rect 21190 2150 21202 2202
rect 21202 2150 21232 2202
rect 21256 2150 21266 2202
rect 21266 2150 21312 2202
rect 21016 2148 21072 2150
rect 21096 2148 21152 2150
rect 21176 2148 21232 2150
rect 21256 2148 21312 2150
rect 21454 2080 21510 2136
rect 21454 1536 21510 1592
rect 21822 6296 21878 6352
rect 21822 6024 21878 6080
rect 21822 5616 21878 5672
rect 22190 7692 22192 7712
rect 22192 7692 22244 7712
rect 22244 7692 22246 7712
rect 22190 7656 22246 7692
rect 22098 6704 22154 6760
rect 22190 5616 22246 5672
rect 21362 448 21418 504
rect 22374 5480 22430 5536
rect 22098 4392 22154 4448
rect 22098 3712 22154 3768
rect 22098 1536 22154 1592
rect 22282 4256 22338 4312
rect 23202 9696 23258 9752
rect 22650 5752 22706 5808
rect 22742 5616 22798 5672
rect 23018 6024 23074 6080
rect 23018 5616 23074 5672
rect 22282 2896 22338 2952
rect 23018 4256 23074 4312
rect 23018 3576 23074 3632
rect 23018 3052 23074 3088
rect 23018 3032 23020 3052
rect 23020 3032 23072 3052
rect 23072 3032 23074 3052
rect 23386 8064 23442 8120
rect 23386 7384 23442 7440
rect 23478 5652 23480 5672
rect 23480 5652 23532 5672
rect 23532 5652 23534 5672
rect 23478 5616 23534 5652
rect 23386 5344 23442 5400
rect 23294 4936 23350 4992
rect 23018 1536 23074 1592
rect 23018 856 23074 912
rect 24122 6180 24178 6216
rect 24122 6160 24124 6180
rect 24124 6160 24176 6180
rect 24176 6160 24178 6180
rect 24122 5364 24178 5400
rect 24122 5344 24124 5364
rect 24124 5344 24176 5364
rect 24176 5344 24178 5364
rect 24674 8880 24730 8936
rect 25042 8200 25098 8256
rect 24950 6976 25006 7032
rect 25594 6976 25650 7032
rect 25410 6568 25466 6624
rect 25502 5888 25558 5944
rect 24398 5344 24454 5400
rect 24214 5072 24270 5128
rect 23938 4256 23994 4312
rect 23846 3576 23902 3632
rect 23662 3168 23718 3224
rect 23754 2216 23810 2272
rect 24674 3712 24730 3768
rect 24950 4800 25006 4856
rect 24858 3304 24914 3360
rect 25410 5344 25466 5400
rect 25318 4936 25374 4992
rect 25226 3576 25282 3632
rect 25042 3032 25098 3088
rect 25134 2896 25190 2952
rect 25134 1944 25190 2000
rect 25594 4256 25650 4312
rect 25778 8608 25834 8664
rect 25956 8186 26012 8188
rect 26036 8186 26092 8188
rect 26116 8186 26172 8188
rect 26196 8186 26252 8188
rect 25956 8134 26002 8186
rect 26002 8134 26012 8186
rect 26036 8134 26066 8186
rect 26066 8134 26078 8186
rect 26078 8134 26092 8186
rect 26116 8134 26130 8186
rect 26130 8134 26142 8186
rect 26142 8134 26172 8186
rect 26196 8134 26206 8186
rect 26206 8134 26252 8186
rect 25956 8132 26012 8134
rect 26036 8132 26092 8134
rect 26116 8132 26172 8134
rect 26196 8132 26252 8134
rect 25870 7928 25926 7984
rect 26146 7928 26202 7984
rect 25778 7520 25834 7576
rect 26422 7520 26478 7576
rect 25956 7098 26012 7100
rect 26036 7098 26092 7100
rect 26116 7098 26172 7100
rect 26196 7098 26252 7100
rect 25956 7046 26002 7098
rect 26002 7046 26012 7098
rect 26036 7046 26066 7098
rect 26066 7046 26078 7098
rect 26078 7046 26092 7098
rect 26116 7046 26130 7098
rect 26130 7046 26142 7098
rect 26142 7046 26172 7098
rect 26196 7046 26206 7098
rect 26206 7046 26252 7098
rect 25956 7044 26012 7046
rect 26036 7044 26092 7046
rect 26116 7044 26172 7046
rect 26196 7044 26252 7046
rect 26422 7112 26478 7168
rect 25962 6740 25964 6760
rect 25964 6740 26016 6760
rect 26016 6740 26018 6760
rect 25962 6704 26018 6740
rect 25956 6010 26012 6012
rect 26036 6010 26092 6012
rect 26116 6010 26172 6012
rect 26196 6010 26252 6012
rect 25956 5958 26002 6010
rect 26002 5958 26012 6010
rect 26036 5958 26066 6010
rect 26066 5958 26078 6010
rect 26078 5958 26092 6010
rect 26116 5958 26130 6010
rect 26130 5958 26142 6010
rect 26142 5958 26172 6010
rect 26196 5958 26206 6010
rect 26206 5958 26252 6010
rect 25956 5956 26012 5958
rect 26036 5956 26092 5958
rect 26116 5956 26172 5958
rect 26196 5956 26252 5958
rect 25870 5616 25926 5672
rect 26146 5480 26202 5536
rect 25778 5208 25834 5264
rect 25956 4922 26012 4924
rect 26036 4922 26092 4924
rect 26116 4922 26172 4924
rect 26196 4922 26252 4924
rect 25956 4870 26002 4922
rect 26002 4870 26012 4922
rect 26036 4870 26066 4922
rect 26066 4870 26078 4922
rect 26078 4870 26092 4922
rect 26116 4870 26130 4922
rect 26130 4870 26142 4922
rect 26142 4870 26172 4922
rect 26196 4870 26206 4922
rect 26206 4870 26252 4922
rect 25956 4868 26012 4870
rect 26036 4868 26092 4870
rect 26116 4868 26172 4870
rect 26196 4868 26252 4870
rect 25134 1264 25190 1320
rect 25594 3848 25650 3904
rect 25502 3712 25558 3768
rect 26514 6740 26516 6760
rect 26516 6740 26568 6760
rect 26568 6740 26570 6760
rect 26514 6704 26570 6740
rect 27016 8730 27072 8732
rect 27096 8730 27152 8732
rect 27176 8730 27232 8732
rect 27256 8730 27312 8732
rect 27016 8678 27062 8730
rect 27062 8678 27072 8730
rect 27096 8678 27126 8730
rect 27126 8678 27138 8730
rect 27138 8678 27152 8730
rect 27176 8678 27190 8730
rect 27190 8678 27202 8730
rect 27202 8678 27232 8730
rect 27256 8678 27266 8730
rect 27266 8678 27312 8730
rect 27016 8676 27072 8678
rect 27096 8676 27152 8678
rect 27176 8676 27232 8678
rect 27256 8676 27312 8678
rect 26790 8200 26846 8256
rect 27434 9152 27490 9208
rect 26790 7656 26846 7712
rect 27016 7642 27072 7644
rect 27096 7642 27152 7644
rect 27176 7642 27232 7644
rect 27256 7642 27312 7644
rect 27016 7590 27062 7642
rect 27062 7590 27072 7642
rect 27096 7590 27126 7642
rect 27126 7590 27138 7642
rect 27138 7590 27152 7642
rect 27176 7590 27190 7642
rect 27190 7590 27202 7642
rect 27202 7590 27232 7642
rect 27256 7590 27266 7642
rect 27266 7590 27312 7642
rect 27016 7588 27072 7590
rect 27096 7588 27152 7590
rect 27176 7588 27232 7590
rect 27256 7588 27312 7590
rect 27434 7404 27490 7440
rect 27434 7384 27436 7404
rect 27436 7384 27488 7404
rect 27488 7384 27490 7404
rect 27342 7248 27398 7304
rect 26790 6840 26846 6896
rect 27342 6976 27398 7032
rect 26698 6432 26754 6488
rect 26698 6160 26754 6216
rect 27016 6554 27072 6556
rect 27096 6554 27152 6556
rect 27176 6554 27232 6556
rect 27256 6554 27312 6556
rect 27016 6502 27062 6554
rect 27062 6502 27072 6554
rect 27096 6502 27126 6554
rect 27126 6502 27138 6554
rect 27138 6502 27152 6554
rect 27176 6502 27190 6554
rect 27190 6502 27202 6554
rect 27202 6502 27232 6554
rect 27256 6502 27266 6554
rect 27266 6502 27312 6554
rect 27016 6500 27072 6502
rect 27096 6500 27152 6502
rect 27176 6500 27232 6502
rect 27256 6500 27312 6502
rect 26790 5752 26846 5808
rect 27066 5888 27122 5944
rect 27434 6432 27490 6488
rect 27016 5466 27072 5468
rect 27096 5466 27152 5468
rect 27176 5466 27232 5468
rect 27256 5466 27312 5468
rect 27016 5414 27062 5466
rect 27062 5414 27072 5466
rect 27096 5414 27126 5466
rect 27126 5414 27138 5466
rect 27138 5414 27152 5466
rect 27176 5414 27190 5466
rect 27190 5414 27202 5466
rect 27202 5414 27232 5466
rect 27256 5414 27266 5466
rect 27266 5414 27312 5466
rect 27016 5412 27072 5414
rect 27096 5412 27152 5414
rect 27176 5412 27232 5414
rect 27256 5412 27312 5414
rect 27434 5364 27490 5400
rect 27434 5344 27436 5364
rect 27436 5344 27488 5364
rect 27488 5344 27490 5364
rect 26882 5208 26938 5264
rect 26514 4800 26570 4856
rect 26606 4392 26662 4448
rect 26514 3984 26570 4040
rect 25956 3834 26012 3836
rect 26036 3834 26092 3836
rect 26116 3834 26172 3836
rect 26196 3834 26252 3836
rect 25956 3782 26002 3834
rect 26002 3782 26012 3834
rect 26036 3782 26066 3834
rect 26066 3782 26078 3834
rect 26078 3782 26092 3834
rect 26116 3782 26130 3834
rect 26130 3782 26142 3834
rect 26142 3782 26172 3834
rect 26196 3782 26206 3834
rect 26206 3782 26252 3834
rect 25956 3780 26012 3782
rect 26036 3780 26092 3782
rect 26116 3780 26172 3782
rect 26196 3780 26252 3782
rect 25962 3476 25964 3496
rect 25964 3476 26016 3496
rect 26016 3476 26018 3496
rect 25686 2896 25742 2952
rect 25962 3440 26018 3476
rect 26146 3052 26202 3088
rect 26146 3032 26148 3052
rect 26148 3032 26200 3052
rect 26200 3032 26202 3052
rect 25956 2746 26012 2748
rect 26036 2746 26092 2748
rect 26116 2746 26172 2748
rect 26196 2746 26252 2748
rect 25956 2694 26002 2746
rect 26002 2694 26012 2746
rect 26036 2694 26066 2746
rect 26066 2694 26078 2746
rect 26078 2694 26092 2746
rect 26116 2694 26130 2746
rect 26130 2694 26142 2746
rect 26142 2694 26172 2746
rect 26196 2694 26206 2746
rect 26206 2694 26252 2746
rect 25956 2692 26012 2694
rect 26036 2692 26092 2694
rect 26116 2692 26172 2694
rect 26196 2692 26252 2694
rect 25870 1264 25926 1320
rect 26422 3440 26478 3496
rect 26790 3848 26846 3904
rect 27016 4378 27072 4380
rect 27096 4378 27152 4380
rect 27176 4378 27232 4380
rect 27256 4378 27312 4380
rect 27016 4326 27062 4378
rect 27062 4326 27072 4378
rect 27096 4326 27126 4378
rect 27126 4326 27138 4378
rect 27138 4326 27152 4378
rect 27176 4326 27190 4378
rect 27190 4326 27202 4378
rect 27202 4326 27232 4378
rect 27256 4326 27266 4378
rect 27266 4326 27312 4378
rect 27016 4324 27072 4326
rect 27096 4324 27152 4326
rect 27176 4324 27232 4326
rect 27256 4324 27312 4326
rect 27158 4156 27160 4176
rect 27160 4156 27212 4176
rect 27212 4156 27214 4176
rect 27158 4120 27214 4156
rect 27526 5072 27582 5128
rect 27434 4392 27490 4448
rect 27618 4256 27674 4312
rect 26790 3304 26846 3360
rect 26790 2896 26846 2952
rect 27016 3290 27072 3292
rect 27096 3290 27152 3292
rect 27176 3290 27232 3292
rect 27256 3290 27312 3292
rect 27016 3238 27062 3290
rect 27062 3238 27072 3290
rect 27096 3238 27126 3290
rect 27126 3238 27138 3290
rect 27138 3238 27152 3290
rect 27176 3238 27190 3290
rect 27190 3238 27202 3290
rect 27202 3238 27232 3290
rect 27256 3238 27266 3290
rect 27266 3238 27312 3290
rect 27016 3236 27072 3238
rect 27096 3236 27152 3238
rect 27176 3236 27232 3238
rect 27256 3236 27312 3238
rect 26974 2760 27030 2816
rect 26882 2216 26938 2272
rect 27016 2202 27072 2204
rect 27096 2202 27152 2204
rect 27176 2202 27232 2204
rect 27256 2202 27312 2204
rect 27016 2150 27062 2202
rect 27062 2150 27072 2202
rect 27096 2150 27126 2202
rect 27126 2150 27138 2202
rect 27138 2150 27152 2202
rect 27176 2150 27190 2202
rect 27190 2150 27202 2202
rect 27202 2150 27232 2202
rect 27256 2150 27266 2202
rect 27266 2150 27312 2202
rect 27016 2148 27072 2150
rect 27096 2148 27152 2150
rect 27176 2148 27232 2150
rect 27256 2148 27312 2150
rect 27894 3984 27950 4040
rect 27894 3712 27950 3768
rect 28078 4936 28134 4992
rect 27526 3304 27582 3360
rect 27710 3168 27766 3224
rect 29642 8200 29698 8256
rect 29642 7656 29698 7712
rect 29734 7520 29790 7576
rect 29090 6976 29146 7032
rect 29366 7248 29422 7304
rect 29182 6840 29238 6896
rect 29274 6432 29330 6488
rect 28446 6160 28502 6216
rect 28814 6160 28870 6216
rect 28354 2760 28410 2816
rect 28262 2624 28318 2680
rect 28630 5480 28686 5536
rect 29182 6024 29238 6080
rect 28630 3168 28686 3224
rect 28814 2760 28870 2816
rect 28630 2624 28686 2680
rect 28814 2624 28870 2680
rect 28354 1264 28410 1320
rect 28446 1128 28502 1184
rect 28630 992 28686 1048
rect 28814 856 28870 912
rect 29458 4392 29514 4448
rect 29642 4392 29698 4448
rect 29458 3984 29514 4040
rect 29458 3168 29514 3224
rect 29826 4800 29882 4856
rect 31114 7828 31116 7848
rect 31116 7828 31168 7848
rect 31168 7828 31170 7848
rect 31114 7792 31170 7828
rect 31298 7948 31354 7984
rect 31298 7928 31300 7948
rect 31300 7928 31352 7948
rect 31352 7928 31354 7948
rect 31206 7384 31262 7440
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 31482 7928 31538 7984
rect 31390 7792 31446 7848
rect 31390 7656 31446 7712
rect 30838 6432 30894 6488
rect 30194 4800 30250 4856
rect 29918 4256 29974 4312
rect 29550 2896 29606 2952
rect 29734 3304 29790 3360
rect 29734 3168 29790 3224
rect 30010 3304 30066 3360
rect 29826 2932 29828 2952
rect 29828 2932 29880 2952
rect 29880 2932 29882 2952
rect 29826 2896 29882 2932
rect 30010 2896 30066 2952
rect 30102 2760 30158 2816
rect 30838 5344 30894 5400
rect 30746 4936 30802 4992
rect 30194 312 30250 368
rect 31298 5616 31354 5672
rect 31482 7112 31538 7168
rect 31390 4972 31392 4992
rect 31392 4972 31444 4992
rect 31444 4972 31446 4992
rect 31390 4936 31446 4972
rect 31390 4684 31446 4720
rect 31390 4664 31392 4684
rect 31392 4664 31444 4684
rect 31444 4664 31446 4684
rect 31206 4120 31262 4176
rect 31666 5344 31722 5400
rect 32126 7520 32182 7576
rect 32770 9288 32826 9344
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 32218 6740 32220 6760
rect 32220 6740 32272 6760
rect 32272 6740 32274 6760
rect 32218 6704 32274 6740
rect 32310 6316 32366 6352
rect 32310 6296 32312 6316
rect 32312 6296 32364 6316
rect 32364 6296 32366 6316
rect 32494 6296 32550 6352
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 33016 8730 33072 8732
rect 33096 8730 33152 8732
rect 33176 8730 33232 8732
rect 33256 8730 33312 8732
rect 33016 8678 33062 8730
rect 33062 8678 33072 8730
rect 33096 8678 33126 8730
rect 33126 8678 33138 8730
rect 33138 8678 33152 8730
rect 33176 8678 33190 8730
rect 33190 8678 33202 8730
rect 33202 8678 33232 8730
rect 33256 8678 33266 8730
rect 33266 8678 33312 8730
rect 33016 8676 33072 8678
rect 33096 8676 33152 8678
rect 33176 8676 33232 8678
rect 33256 8676 33312 8678
rect 33016 7642 33072 7644
rect 33096 7642 33152 7644
rect 33176 7642 33232 7644
rect 33256 7642 33312 7644
rect 33016 7590 33062 7642
rect 33062 7590 33072 7642
rect 33096 7590 33126 7642
rect 33126 7590 33138 7642
rect 33138 7590 33152 7642
rect 33176 7590 33190 7642
rect 33190 7590 33202 7642
rect 33202 7590 33232 7642
rect 33256 7590 33266 7642
rect 33266 7590 33312 7642
rect 33016 7588 33072 7590
rect 33096 7588 33152 7590
rect 33176 7588 33232 7590
rect 33256 7588 33312 7590
rect 33016 6554 33072 6556
rect 33096 6554 33152 6556
rect 33176 6554 33232 6556
rect 33256 6554 33312 6556
rect 33016 6502 33062 6554
rect 33062 6502 33072 6554
rect 33096 6502 33126 6554
rect 33126 6502 33138 6554
rect 33138 6502 33152 6554
rect 33176 6502 33190 6554
rect 33190 6502 33202 6554
rect 33202 6502 33232 6554
rect 33256 6502 33266 6554
rect 33266 6502 33312 6554
rect 33016 6500 33072 6502
rect 33096 6500 33152 6502
rect 33176 6500 33232 6502
rect 33256 6500 33312 6502
rect 33414 6316 33470 6352
rect 33414 6296 33416 6316
rect 33416 6296 33468 6316
rect 33468 6296 33470 6316
rect 32310 5616 32366 5672
rect 32310 5108 32312 5128
rect 32312 5108 32364 5128
rect 32364 5108 32366 5128
rect 32310 5072 32366 5108
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 31022 3848 31078 3904
rect 31390 3984 31446 4040
rect 31206 1672 31262 1728
rect 32678 5480 32734 5536
rect 32586 5072 32642 5128
rect 32586 4800 32642 4856
rect 31942 4392 31998 4448
rect 31942 3984 31998 4040
rect 32402 4256 32458 4312
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 31942 3304 31998 3360
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 32586 3304 32642 3360
rect 33016 5466 33072 5468
rect 33096 5466 33152 5468
rect 33176 5466 33232 5468
rect 33256 5466 33312 5468
rect 33016 5414 33062 5466
rect 33062 5414 33072 5466
rect 33096 5414 33126 5466
rect 33126 5414 33138 5466
rect 33138 5414 33152 5466
rect 33176 5414 33190 5466
rect 33190 5414 33202 5466
rect 33202 5414 33232 5466
rect 33256 5414 33266 5466
rect 33266 5414 33312 5466
rect 33016 5412 33072 5414
rect 33096 5412 33152 5414
rect 33176 5412 33232 5414
rect 33256 5412 33312 5414
rect 33046 4936 33102 4992
rect 33016 4378 33072 4380
rect 33096 4378 33152 4380
rect 33176 4378 33232 4380
rect 33256 4378 33312 4380
rect 33016 4326 33062 4378
rect 33062 4326 33072 4378
rect 33096 4326 33126 4378
rect 33126 4326 33138 4378
rect 33138 4326 33152 4378
rect 33176 4326 33190 4378
rect 33190 4326 33202 4378
rect 33202 4326 33232 4378
rect 33256 4326 33266 4378
rect 33266 4326 33312 4378
rect 33016 4324 33072 4326
rect 33096 4324 33152 4326
rect 33176 4324 33232 4326
rect 33256 4324 33312 4326
rect 33322 3440 33378 3496
rect 33016 3290 33072 3292
rect 33096 3290 33152 3292
rect 33176 3290 33232 3292
rect 33256 3290 33312 3292
rect 33016 3238 33062 3290
rect 33062 3238 33072 3290
rect 33096 3238 33126 3290
rect 33126 3238 33138 3290
rect 33138 3238 33152 3290
rect 33176 3238 33190 3290
rect 33190 3238 33202 3290
rect 33202 3238 33232 3290
rect 33256 3238 33266 3290
rect 33266 3238 33312 3290
rect 33016 3236 33072 3238
rect 33096 3236 33152 3238
rect 33176 3236 33232 3238
rect 33256 3236 33312 3238
rect 33966 10240 34022 10296
rect 33782 5752 33838 5808
rect 33016 2202 33072 2204
rect 33096 2202 33152 2204
rect 33176 2202 33232 2204
rect 33256 2202 33312 2204
rect 33016 2150 33062 2202
rect 33062 2150 33072 2202
rect 33096 2150 33126 2202
rect 33126 2150 33138 2202
rect 33138 2150 33152 2202
rect 33176 2150 33190 2202
rect 33190 2150 33202 2202
rect 33202 2150 33232 2202
rect 33256 2150 33266 2202
rect 33266 2150 33312 2202
rect 33016 2148 33072 2150
rect 33096 2148 33152 2150
rect 33176 2148 33232 2150
rect 33256 2148 33312 2150
rect 32770 176 32826 232
rect 34334 9968 34390 10024
rect 34334 6840 34390 6896
rect 34794 7384 34850 7440
rect 34518 6704 34574 6760
rect 34610 5072 34666 5128
rect 34426 3984 34482 4040
rect 34702 4548 34758 4584
rect 34702 4528 34704 4548
rect 34704 4528 34756 4548
rect 34756 4528 34758 4548
rect 34794 3576 34850 3632
rect 33782 1536 33838 1592
rect 33322 40 33378 96
rect 35346 8336 35402 8392
rect 35254 5616 35310 5672
rect 34610 1808 34666 1864
rect 34518 1264 34574 1320
rect 35162 992 35218 1048
rect 35438 1400 35494 1456
rect 37186 10512 37242 10568
rect 36450 10376 36506 10432
rect 35898 6296 35954 6352
rect 35806 4936 35862 4992
rect 35898 4800 35954 4856
rect 35714 3052 35770 3088
rect 35714 3032 35716 3052
rect 35716 3032 35768 3052
rect 35768 3032 35770 3052
rect 36174 4140 36230 4176
rect 36174 4120 36176 4140
rect 36176 4120 36228 4140
rect 36228 4120 36230 4140
rect 35898 2488 35954 2544
rect 36174 720 36230 776
rect 37002 9016 37058 9072
rect 36634 6568 36690 6624
rect 36634 2896 36690 2952
rect 39486 9832 39542 9888
rect 38658 9560 38714 9616
rect 38382 9288 38438 9344
rect 38290 9016 38346 9072
rect 37830 8492 37886 8528
rect 37830 8472 37832 8492
rect 37832 8472 37884 8492
rect 37884 8472 37886 8492
rect 37956 8186 38012 8188
rect 38036 8186 38092 8188
rect 38116 8186 38172 8188
rect 38196 8186 38252 8188
rect 37956 8134 38002 8186
rect 38002 8134 38012 8186
rect 38036 8134 38066 8186
rect 38066 8134 38078 8186
rect 38078 8134 38092 8186
rect 38116 8134 38130 8186
rect 38130 8134 38142 8186
rect 38142 8134 38172 8186
rect 38196 8134 38206 8186
rect 38206 8134 38252 8186
rect 37956 8132 38012 8134
rect 38036 8132 38092 8134
rect 38116 8132 38172 8134
rect 38196 8132 38252 8134
rect 38474 8200 38530 8256
rect 38474 7248 38530 7304
rect 37956 7098 38012 7100
rect 38036 7098 38092 7100
rect 38116 7098 38172 7100
rect 38196 7098 38252 7100
rect 37956 7046 38002 7098
rect 38002 7046 38012 7098
rect 38036 7046 38066 7098
rect 38066 7046 38078 7098
rect 38078 7046 38092 7098
rect 38116 7046 38130 7098
rect 38130 7046 38142 7098
rect 38142 7046 38172 7098
rect 38196 7046 38206 7098
rect 38206 7046 38252 7098
rect 37956 7044 38012 7046
rect 38036 7044 38092 7046
rect 38116 7044 38172 7046
rect 38196 7044 38252 7046
rect 38842 9424 38898 9480
rect 38750 8472 38806 8528
rect 39016 8730 39072 8732
rect 39096 8730 39152 8732
rect 39176 8730 39232 8732
rect 39256 8730 39312 8732
rect 39016 8678 39062 8730
rect 39062 8678 39072 8730
rect 39096 8678 39126 8730
rect 39126 8678 39138 8730
rect 39138 8678 39152 8730
rect 39176 8678 39190 8730
rect 39190 8678 39202 8730
rect 39202 8678 39232 8730
rect 39256 8678 39266 8730
rect 39266 8678 39312 8730
rect 39016 8676 39072 8678
rect 39096 8676 39152 8678
rect 39176 8676 39232 8678
rect 39256 8676 39312 8678
rect 38658 7948 38714 7984
rect 38658 7928 38660 7948
rect 38660 7928 38712 7948
rect 38712 7928 38714 7948
rect 38658 7792 38714 7848
rect 39026 7928 39082 7984
rect 37956 6010 38012 6012
rect 38036 6010 38092 6012
rect 38116 6010 38172 6012
rect 38196 6010 38252 6012
rect 37956 5958 38002 6010
rect 38002 5958 38012 6010
rect 38036 5958 38066 6010
rect 38066 5958 38078 6010
rect 38078 5958 38092 6010
rect 38116 5958 38130 6010
rect 38130 5958 38142 6010
rect 38142 5958 38172 6010
rect 38196 5958 38206 6010
rect 38206 5958 38252 6010
rect 37956 5956 38012 5958
rect 38036 5956 38092 5958
rect 38116 5956 38172 5958
rect 38196 5956 38252 5958
rect 37956 4922 38012 4924
rect 38036 4922 38092 4924
rect 38116 4922 38172 4924
rect 38196 4922 38252 4924
rect 37956 4870 38002 4922
rect 38002 4870 38012 4922
rect 38036 4870 38066 4922
rect 38066 4870 38078 4922
rect 38078 4870 38092 4922
rect 38116 4870 38130 4922
rect 38130 4870 38142 4922
rect 38142 4870 38172 4922
rect 38196 4870 38206 4922
rect 38206 4870 38252 4922
rect 37956 4868 38012 4870
rect 38036 4868 38092 4870
rect 38116 4868 38172 4870
rect 38196 4868 38252 4870
rect 39394 7692 39396 7712
rect 39396 7692 39448 7712
rect 39448 7692 39450 7712
rect 39394 7656 39450 7692
rect 39016 7642 39072 7644
rect 39096 7642 39152 7644
rect 39176 7642 39232 7644
rect 39256 7642 39312 7644
rect 39016 7590 39062 7642
rect 39062 7590 39072 7642
rect 39096 7590 39126 7642
rect 39126 7590 39138 7642
rect 39138 7590 39152 7642
rect 39176 7590 39190 7642
rect 39190 7590 39202 7642
rect 39202 7590 39232 7642
rect 39256 7590 39266 7642
rect 39266 7590 39312 7642
rect 39016 7588 39072 7590
rect 39096 7588 39152 7590
rect 39176 7588 39232 7590
rect 39256 7588 39312 7590
rect 38934 7384 38990 7440
rect 39394 7148 39396 7168
rect 39396 7148 39448 7168
rect 39448 7148 39450 7168
rect 39394 7112 39450 7148
rect 38382 6604 38384 6624
rect 38384 6604 38436 6624
rect 38436 6604 38438 6624
rect 38382 6568 38438 6604
rect 39394 6604 39396 6624
rect 39396 6604 39448 6624
rect 39448 6604 39450 6624
rect 39394 6568 39450 6604
rect 39016 6554 39072 6556
rect 39096 6554 39152 6556
rect 39176 6554 39232 6556
rect 39256 6554 39312 6556
rect 39016 6502 39062 6554
rect 39062 6502 39072 6554
rect 39096 6502 39126 6554
rect 39126 6502 39138 6554
rect 39138 6502 39152 6554
rect 39176 6502 39190 6554
rect 39190 6502 39202 6554
rect 39202 6502 39232 6554
rect 39256 6502 39266 6554
rect 39266 6502 39312 6554
rect 39016 6500 39072 6502
rect 39096 6500 39152 6502
rect 39176 6500 39232 6502
rect 39256 6500 39312 6502
rect 39578 8744 39634 8800
rect 40038 6840 40094 6896
rect 39394 6296 39450 6352
rect 37956 3834 38012 3836
rect 38036 3834 38092 3836
rect 38116 3834 38172 3836
rect 38196 3834 38252 3836
rect 37956 3782 38002 3834
rect 38002 3782 38012 3834
rect 38036 3782 38066 3834
rect 38066 3782 38078 3834
rect 38078 3782 38092 3834
rect 38116 3782 38130 3834
rect 38130 3782 38142 3834
rect 38142 3782 38172 3834
rect 38196 3782 38206 3834
rect 38206 3782 38252 3834
rect 37956 3780 38012 3782
rect 38036 3780 38092 3782
rect 38116 3780 38172 3782
rect 38196 3780 38252 3782
rect 39210 6160 39266 6216
rect 39026 6060 39028 6080
rect 39028 6060 39080 6080
rect 39080 6060 39082 6080
rect 39026 6024 39082 6060
rect 38842 5228 38898 5264
rect 39394 5752 39450 5808
rect 39016 5466 39072 5468
rect 39096 5466 39152 5468
rect 39176 5466 39232 5468
rect 39256 5466 39312 5468
rect 39016 5414 39062 5466
rect 39062 5414 39072 5466
rect 39096 5414 39126 5466
rect 39126 5414 39138 5466
rect 39138 5414 39152 5466
rect 39176 5414 39190 5466
rect 39190 5414 39202 5466
rect 39202 5414 39232 5466
rect 39256 5414 39266 5466
rect 39266 5414 39312 5466
rect 39016 5412 39072 5414
rect 39096 5412 39152 5414
rect 39176 5412 39232 5414
rect 39256 5412 39312 5414
rect 39946 5480 40002 5536
rect 38842 5208 38844 5228
rect 38844 5208 38896 5228
rect 38896 5208 38898 5228
rect 39394 5208 39450 5264
rect 39026 4972 39028 4992
rect 39028 4972 39080 4992
rect 39080 4972 39082 4992
rect 39026 4936 39082 4972
rect 39210 4664 39266 4720
rect 39486 4664 39542 4720
rect 39394 4392 39450 4448
rect 39016 4378 39072 4380
rect 39096 4378 39152 4380
rect 39176 4378 39232 4380
rect 39256 4378 39312 4380
rect 39016 4326 39062 4378
rect 39062 4326 39072 4378
rect 39096 4326 39126 4378
rect 39126 4326 39138 4378
rect 39138 4326 39152 4378
rect 39176 4326 39190 4378
rect 39190 4326 39202 4378
rect 39202 4326 39232 4378
rect 39256 4326 39266 4378
rect 39266 4326 39312 4378
rect 39016 4324 39072 4326
rect 39096 4324 39152 4326
rect 39176 4324 39232 4326
rect 39256 4324 39312 4326
rect 39394 4120 39450 4176
rect 39026 3884 39028 3904
rect 39028 3884 39080 3904
rect 39080 3884 39082 3904
rect 39026 3848 39082 3884
rect 37956 2746 38012 2748
rect 38036 2746 38092 2748
rect 38116 2746 38172 2748
rect 38196 2746 38252 2748
rect 37956 2694 38002 2746
rect 38002 2694 38012 2746
rect 38036 2694 38066 2746
rect 38066 2694 38078 2746
rect 38078 2694 38092 2746
rect 38116 2694 38130 2746
rect 38130 2694 38142 2746
rect 38142 2694 38172 2746
rect 38196 2694 38206 2746
rect 38206 2694 38252 2746
rect 37956 2692 38012 2694
rect 38036 2692 38092 2694
rect 38116 2692 38172 2694
rect 38196 2692 38252 2694
rect 38106 2488 38162 2544
rect 38658 1672 38714 1728
rect 39394 3576 39450 3632
rect 39016 3290 39072 3292
rect 39096 3290 39152 3292
rect 39176 3290 39232 3292
rect 39256 3290 39312 3292
rect 39016 3238 39062 3290
rect 39062 3238 39072 3290
rect 39096 3238 39126 3290
rect 39126 3238 39138 3290
rect 39138 3238 39152 3290
rect 39176 3238 39190 3290
rect 39190 3238 39202 3290
rect 39202 3238 39232 3290
rect 39256 3238 39266 3290
rect 39266 3238 39312 3290
rect 39016 3236 39072 3238
rect 39096 3236 39152 3238
rect 39176 3236 39232 3238
rect 39256 3236 39312 3238
rect 39946 3304 40002 3360
rect 39394 3032 39450 3088
rect 39026 2796 39028 2816
rect 39028 2796 39080 2816
rect 39080 2796 39082 2816
rect 39026 2760 39082 2796
rect 39210 2388 39212 2408
rect 39212 2388 39264 2408
rect 39264 2388 39266 2408
rect 39210 2352 39266 2388
rect 39016 2202 39072 2204
rect 39096 2202 39152 2204
rect 39176 2202 39232 2204
rect 39256 2202 39312 2204
rect 39016 2150 39062 2202
rect 39062 2150 39072 2202
rect 39096 2150 39126 2202
rect 39126 2150 39138 2202
rect 39138 2150 39152 2202
rect 39176 2150 39190 2202
rect 39190 2150 39202 2202
rect 39202 2150 39232 2202
rect 39256 2150 39266 2202
rect 39266 2150 39312 2202
rect 39016 2148 39072 2150
rect 39096 2148 39152 2150
rect 39176 2148 39232 2150
rect 39256 2148 39312 2150
rect 39670 2488 39726 2544
rect 39946 2252 39948 2272
rect 39948 2252 40000 2272
rect 40000 2252 40002 2272
rect 39946 2216 40002 2252
rect 39578 1944 39634 2000
rect 40038 1400 40094 1456
<< metal3 >>
rect 9949 10570 10015 10573
rect 37181 10570 37247 10573
rect 9949 10568 37247 10570
rect 9949 10512 9954 10568
rect 10010 10512 37186 10568
rect 37242 10512 37247 10568
rect 9949 10510 37247 10512
rect 9949 10507 10015 10510
rect 37181 10507 37247 10510
rect 10317 10434 10383 10437
rect 36445 10434 36511 10437
rect 10317 10432 36511 10434
rect 10317 10376 10322 10432
rect 10378 10376 36450 10432
rect 36506 10376 36511 10432
rect 10317 10374 36511 10376
rect 10317 10371 10383 10374
rect 36445 10371 36511 10374
rect 13905 10298 13971 10301
rect 33961 10298 34027 10301
rect 13905 10296 34027 10298
rect 13905 10240 13910 10296
rect 13966 10240 33966 10296
rect 34022 10240 34027 10296
rect 13905 10238 34027 10240
rect 13905 10235 13971 10238
rect 33961 10235 34027 10238
rect 7281 10162 7347 10165
rect 30414 10162 30420 10164
rect 7281 10160 30420 10162
rect 7281 10104 7286 10160
rect 7342 10104 30420 10160
rect 7281 10102 30420 10104
rect 7281 10099 7347 10102
rect 30414 10100 30420 10102
rect 30484 10100 30490 10164
rect 8845 10026 8911 10029
rect 34329 10026 34395 10029
rect 8845 10024 34395 10026
rect 8845 9968 8850 10024
rect 8906 9968 34334 10024
rect 34390 9968 34395 10024
rect 8845 9966 34395 9968
rect 8845 9963 8911 9966
rect 34329 9963 34395 9966
rect 0 9890 120 9920
rect 5533 9890 5599 9893
rect 0 9888 5599 9890
rect 0 9832 5538 9888
rect 5594 9832 5599 9888
rect 0 9830 5599 9832
rect 0 9800 120 9830
rect 5533 9827 5599 9830
rect 11094 9828 11100 9892
rect 11164 9890 11170 9892
rect 17953 9890 18019 9893
rect 11164 9888 18019 9890
rect 11164 9832 17958 9888
rect 18014 9832 18019 9888
rect 11164 9830 18019 9832
rect 11164 9828 11170 9830
rect 17953 9827 18019 9830
rect 39481 9890 39547 9893
rect 40880 9890 41000 9920
rect 39481 9888 41000 9890
rect 39481 9832 39486 9888
rect 39542 9832 41000 9888
rect 39481 9830 41000 9832
rect 39481 9827 39547 9830
rect 40880 9800 41000 9830
rect 6361 9754 6427 9757
rect 16481 9754 16547 9757
rect 6361 9752 16547 9754
rect 6361 9696 6366 9752
rect 6422 9696 16486 9752
rect 16542 9696 16547 9752
rect 6361 9694 16547 9696
rect 6361 9691 6427 9694
rect 16481 9691 16547 9694
rect 16614 9692 16620 9756
rect 16684 9754 16690 9756
rect 23197 9754 23263 9757
rect 16684 9752 23263 9754
rect 16684 9696 23202 9752
rect 23258 9696 23263 9752
rect 16684 9694 23263 9696
rect 16684 9692 16690 9694
rect 23197 9691 23263 9694
rect 0 9618 120 9648
rect 3417 9618 3483 9621
rect 0 9616 3483 9618
rect 0 9560 3422 9616
rect 3478 9560 3483 9616
rect 0 9558 3483 9560
rect 0 9528 120 9558
rect 3417 9555 3483 9558
rect 9673 9618 9739 9621
rect 15837 9618 15903 9621
rect 9673 9616 15903 9618
rect 9673 9560 9678 9616
rect 9734 9560 15842 9616
rect 15898 9560 15903 9616
rect 9673 9558 15903 9560
rect 9673 9555 9739 9558
rect 15837 9555 15903 9558
rect 38653 9618 38719 9621
rect 40880 9618 41000 9648
rect 38653 9616 41000 9618
rect 38653 9560 38658 9616
rect 38714 9560 41000 9616
rect 38653 9558 41000 9560
rect 38653 9555 38719 9558
rect 40880 9528 41000 9558
rect 3601 9482 3667 9485
rect 15101 9482 15167 9485
rect 3601 9480 15167 9482
rect 3601 9424 3606 9480
rect 3662 9424 15106 9480
rect 15162 9424 15167 9480
rect 3601 9422 15167 9424
rect 3601 9419 3667 9422
rect 15101 9419 15167 9422
rect 16481 9482 16547 9485
rect 38837 9482 38903 9485
rect 16481 9480 38903 9482
rect 16481 9424 16486 9480
rect 16542 9424 38842 9480
rect 38898 9424 38903 9480
rect 16481 9422 38903 9424
rect 16481 9419 16547 9422
rect 38837 9419 38903 9422
rect 0 9346 120 9376
rect 3877 9346 3943 9349
rect 0 9344 3943 9346
rect 0 9288 3882 9344
rect 3938 9288 3943 9344
rect 0 9286 3943 9288
rect 0 9256 120 9286
rect 3877 9283 3943 9286
rect 5809 9346 5875 9349
rect 32765 9346 32831 9349
rect 5809 9344 32831 9346
rect 5809 9288 5814 9344
rect 5870 9288 32770 9344
rect 32826 9288 32831 9344
rect 5809 9286 32831 9288
rect 5809 9283 5875 9286
rect 32765 9283 32831 9286
rect 38377 9346 38443 9349
rect 40880 9346 41000 9376
rect 38377 9344 41000 9346
rect 38377 9288 38382 9344
rect 38438 9288 41000 9344
rect 38377 9286 41000 9288
rect 38377 9283 38443 9286
rect 40880 9256 41000 9286
rect 4613 9210 4679 9213
rect 27429 9210 27495 9213
rect 4613 9208 27495 9210
rect 4613 9152 4618 9208
rect 4674 9152 27434 9208
rect 27490 9152 27495 9208
rect 4613 9150 27495 9152
rect 4613 9147 4679 9150
rect 27429 9147 27495 9150
rect 0 9074 120 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 120 9014
rect 1393 9011 1459 9014
rect 12341 9074 12407 9077
rect 17585 9074 17651 9077
rect 12341 9072 17651 9074
rect 12341 9016 12346 9072
rect 12402 9016 17590 9072
rect 17646 9016 17651 9072
rect 12341 9014 17651 9016
rect 12341 9011 12407 9014
rect 17585 9011 17651 9014
rect 17953 9074 18019 9077
rect 36997 9074 37063 9077
rect 17953 9072 37063 9074
rect 17953 9016 17958 9072
rect 18014 9016 37002 9072
rect 37058 9016 37063 9072
rect 17953 9014 37063 9016
rect 17953 9011 18019 9014
rect 36997 9011 37063 9014
rect 38285 9074 38351 9077
rect 40880 9074 41000 9104
rect 38285 9072 41000 9074
rect 38285 9016 38290 9072
rect 38346 9016 41000 9072
rect 38285 9014 41000 9016
rect 38285 9011 38351 9014
rect 40880 8984 41000 9014
rect 8518 8876 8524 8940
rect 8588 8938 8594 8940
rect 9305 8938 9371 8941
rect 8588 8936 9371 8938
rect 8588 8880 9310 8936
rect 9366 8880 9371 8936
rect 8588 8878 9371 8880
rect 8588 8876 8594 8878
rect 9305 8875 9371 8878
rect 11237 8938 11303 8941
rect 24669 8938 24735 8941
rect 11237 8936 24735 8938
rect 11237 8880 11242 8936
rect 11298 8880 24674 8936
rect 24730 8880 24735 8936
rect 11237 8878 24735 8880
rect 11237 8875 11303 8878
rect 24669 8875 24735 8878
rect 0 8802 120 8832
rect 2773 8802 2839 8805
rect 0 8800 2839 8802
rect 0 8744 2778 8800
rect 2834 8744 2839 8800
rect 0 8742 2839 8744
rect 0 8712 120 8742
rect 2773 8739 2839 8742
rect 17585 8802 17651 8805
rect 18873 8802 18939 8805
rect 20805 8802 20871 8805
rect 17585 8800 20871 8802
rect 17585 8744 17590 8800
rect 17646 8744 18878 8800
rect 18934 8744 20810 8800
rect 20866 8744 20871 8800
rect 17585 8742 20871 8744
rect 17585 8739 17651 8742
rect 18873 8739 18939 8742
rect 20805 8739 20871 8742
rect 39573 8802 39639 8805
rect 40880 8802 41000 8832
rect 39573 8800 41000 8802
rect 39573 8744 39578 8800
rect 39634 8744 41000 8800
rect 39573 8742 41000 8744
rect 39573 8739 39639 8742
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 9006 8736 9322 8737
rect 9006 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9322 8736
rect 9006 8671 9322 8672
rect 15006 8736 15322 8737
rect 15006 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15322 8736
rect 15006 8671 15322 8672
rect 21006 8736 21322 8737
rect 21006 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21322 8736
rect 21006 8671 21322 8672
rect 27006 8736 27322 8737
rect 27006 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27322 8736
rect 27006 8671 27322 8672
rect 33006 8736 33322 8737
rect 33006 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33322 8736
rect 33006 8671 33322 8672
rect 39006 8736 39322 8737
rect 39006 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39322 8736
rect 40880 8712 41000 8742
rect 39006 8671 39322 8672
rect 4429 8666 4495 8669
rect 8385 8666 8451 8669
rect 4429 8664 8451 8666
rect 4429 8608 4434 8664
rect 4490 8608 8390 8664
rect 8446 8608 8451 8664
rect 4429 8606 8451 8608
rect 4429 8603 4495 8606
rect 8385 8603 8451 8606
rect 22502 8604 22508 8668
rect 22572 8666 22578 8668
rect 25773 8666 25839 8669
rect 22572 8664 25839 8666
rect 22572 8608 25778 8664
rect 25834 8608 25839 8664
rect 22572 8606 25839 8608
rect 22572 8604 22578 8606
rect 25773 8603 25839 8606
rect 0 8530 120 8560
rect 3325 8530 3391 8533
rect 0 8528 3391 8530
rect 0 8472 3330 8528
rect 3386 8472 3391 8528
rect 0 8470 3391 8472
rect 0 8440 120 8470
rect 3325 8467 3391 8470
rect 6453 8530 6519 8533
rect 37825 8530 37891 8533
rect 6453 8528 37891 8530
rect 6453 8472 6458 8528
rect 6514 8472 37830 8528
rect 37886 8472 37891 8528
rect 6453 8470 37891 8472
rect 6453 8467 6519 8470
rect 37825 8467 37891 8470
rect 38745 8530 38811 8533
rect 40880 8530 41000 8560
rect 38745 8528 41000 8530
rect 38745 8472 38750 8528
rect 38806 8472 41000 8528
rect 38745 8470 41000 8472
rect 38745 8467 38811 8470
rect 40880 8440 41000 8470
rect 3509 8394 3575 8397
rect 7189 8394 7255 8397
rect 8385 8394 8451 8397
rect 3509 8392 8451 8394
rect 3509 8336 3514 8392
rect 3570 8336 7194 8392
rect 7250 8336 8390 8392
rect 8446 8336 8451 8392
rect 3509 8334 8451 8336
rect 3509 8331 3575 8334
rect 7189 8331 7255 8334
rect 8385 8331 8451 8334
rect 11329 8394 11395 8397
rect 13169 8394 13235 8397
rect 11329 8392 13235 8394
rect 11329 8336 11334 8392
rect 11390 8336 13174 8392
rect 13230 8336 13235 8392
rect 11329 8334 13235 8336
rect 11329 8331 11395 8334
rect 13169 8331 13235 8334
rect 13670 8332 13676 8396
rect 13740 8394 13746 8396
rect 16481 8394 16547 8397
rect 35341 8394 35407 8397
rect 13740 8334 14474 8394
rect 13740 8332 13746 8334
rect 0 8258 120 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 120 8198
rect 1393 8195 1459 8198
rect 3693 8258 3759 8261
rect 5901 8258 5967 8261
rect 3693 8256 5967 8258
rect 3693 8200 3698 8256
rect 3754 8200 5906 8256
rect 5962 8200 5967 8256
rect 3693 8198 5967 8200
rect 14414 8258 14474 8334
rect 16481 8392 35407 8394
rect 16481 8336 16486 8392
rect 16542 8336 35346 8392
rect 35402 8336 35407 8392
rect 16481 8334 35407 8336
rect 16481 8331 16547 8334
rect 35341 8331 35407 8334
rect 19057 8258 19123 8261
rect 14414 8256 19123 8258
rect 14414 8200 19062 8256
rect 19118 8200 19123 8256
rect 14414 8198 19123 8200
rect 3693 8195 3759 8198
rect 5901 8195 5967 8198
rect 19057 8195 19123 8198
rect 20529 8258 20595 8261
rect 25037 8258 25103 8261
rect 20529 8256 25103 8258
rect 20529 8200 20534 8256
rect 20590 8200 25042 8256
rect 25098 8200 25103 8256
rect 20529 8198 25103 8200
rect 20529 8195 20595 8198
rect 25037 8195 25103 8198
rect 26785 8258 26851 8261
rect 29637 8258 29703 8261
rect 26785 8256 29703 8258
rect 26785 8200 26790 8256
rect 26846 8200 29642 8256
rect 29698 8200 29703 8256
rect 26785 8198 29703 8200
rect 26785 8195 26851 8198
rect 29637 8195 29703 8198
rect 38469 8258 38535 8261
rect 40880 8258 41000 8288
rect 38469 8256 41000 8258
rect 38469 8200 38474 8256
rect 38530 8200 41000 8256
rect 38469 8198 41000 8200
rect 38469 8195 38535 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 13946 8192 14262 8193
rect 13946 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14262 8192
rect 13946 8127 14262 8128
rect 19946 8192 20262 8193
rect 19946 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20262 8192
rect 19946 8127 20262 8128
rect 25946 8192 26262 8193
rect 25946 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26262 8192
rect 25946 8127 26262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 37946 8192 38262 8193
rect 37946 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38262 8192
rect 40880 8168 41000 8198
rect 37946 8127 38262 8128
rect 10685 8122 10751 8125
rect 13537 8122 13603 8125
rect 10685 8120 13603 8122
rect 10685 8064 10690 8120
rect 10746 8064 13542 8120
rect 13598 8064 13603 8120
rect 10685 8062 13603 8064
rect 10685 8059 10751 8062
rect 13537 8059 13603 8062
rect 14774 8060 14780 8124
rect 14844 8122 14850 8124
rect 16113 8122 16179 8125
rect 18137 8122 18203 8125
rect 14844 8120 16179 8122
rect 14844 8064 16118 8120
rect 16174 8064 16179 8120
rect 14844 8062 16179 8064
rect 14844 8060 14850 8062
rect 16113 8059 16179 8062
rect 16990 8120 18203 8122
rect 16990 8064 18142 8120
rect 18198 8064 18203 8120
rect 16990 8062 18203 8064
rect 0 7986 120 8016
rect 2221 7986 2287 7989
rect 0 7984 2287 7986
rect 0 7928 2226 7984
rect 2282 7928 2287 7984
rect 0 7926 2287 7928
rect 0 7896 120 7926
rect 2221 7923 2287 7926
rect 9489 7986 9555 7989
rect 12525 7986 12591 7989
rect 16990 7986 17050 8062
rect 18137 8059 18203 8062
rect 20345 8122 20411 8125
rect 23381 8122 23447 8125
rect 20345 8120 23447 8122
rect 20345 8064 20350 8120
rect 20406 8064 23386 8120
rect 23442 8064 23447 8120
rect 20345 8062 23447 8064
rect 20345 8059 20411 8062
rect 23381 8059 23447 8062
rect 9489 7984 12450 7986
rect 9489 7928 9494 7984
rect 9550 7928 12450 7984
rect 9489 7926 12450 7928
rect 9489 7923 9555 7926
rect 9489 7850 9555 7853
rect 11881 7852 11947 7853
rect 4478 7848 9555 7850
rect 4478 7792 9494 7848
rect 9550 7792 9555 7848
rect 4478 7790 9555 7792
rect 0 7714 120 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 120 7654
rect 1485 7651 1551 7654
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 0 7442 120 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 120 7382
rect 1393 7379 1459 7382
rect 1669 7442 1735 7445
rect 4478 7442 4538 7790
rect 9489 7787 9555 7790
rect 11830 7788 11836 7852
rect 11900 7850 11947 7852
rect 12390 7850 12450 7926
rect 12525 7984 17050 7986
rect 12525 7928 12530 7984
rect 12586 7928 17050 7984
rect 12525 7926 17050 7928
rect 17217 7986 17283 7989
rect 25865 7986 25931 7989
rect 17217 7984 25931 7986
rect 17217 7928 17222 7984
rect 17278 7928 25870 7984
rect 25926 7928 25931 7984
rect 17217 7926 25931 7928
rect 12525 7923 12591 7926
rect 17217 7923 17283 7926
rect 25865 7923 25931 7926
rect 26141 7986 26207 7989
rect 31293 7986 31359 7989
rect 26141 7984 31359 7986
rect 26141 7928 26146 7984
rect 26202 7928 31298 7984
rect 31354 7928 31359 7984
rect 26141 7926 31359 7928
rect 26141 7923 26207 7926
rect 31293 7923 31359 7926
rect 31477 7986 31543 7989
rect 38653 7986 38719 7989
rect 31477 7984 38719 7986
rect 31477 7928 31482 7984
rect 31538 7928 38658 7984
rect 38714 7928 38719 7984
rect 31477 7926 38719 7928
rect 31477 7923 31543 7926
rect 38653 7923 38719 7926
rect 39021 7986 39087 7989
rect 40880 7986 41000 8016
rect 39021 7984 41000 7986
rect 39021 7928 39026 7984
rect 39082 7928 41000 7984
rect 39021 7926 41000 7928
rect 39021 7923 39087 7926
rect 40880 7896 41000 7926
rect 20345 7850 20411 7853
rect 31109 7850 31175 7853
rect 11900 7848 11992 7850
rect 11942 7792 11992 7848
rect 11900 7790 11992 7792
rect 12390 7848 20411 7850
rect 12390 7792 20350 7848
rect 20406 7792 20411 7848
rect 12390 7790 20411 7792
rect 11900 7788 11947 7790
rect 11881 7787 11947 7788
rect 20345 7787 20411 7790
rect 20670 7848 31175 7850
rect 20670 7792 31114 7848
rect 31170 7792 31175 7848
rect 20670 7790 31175 7792
rect 10777 7714 10843 7717
rect 11513 7714 11579 7717
rect 14406 7714 14412 7716
rect 10777 7712 14412 7714
rect 10777 7656 10782 7712
rect 10838 7656 11518 7712
rect 11574 7656 14412 7712
rect 10777 7654 14412 7656
rect 10777 7651 10843 7654
rect 11513 7651 11579 7654
rect 14406 7652 14412 7654
rect 14476 7652 14482 7716
rect 15561 7714 15627 7717
rect 17953 7714 18019 7717
rect 15561 7712 18019 7714
rect 15561 7656 15566 7712
rect 15622 7656 17958 7712
rect 18014 7656 18019 7712
rect 15561 7654 18019 7656
rect 15561 7651 15627 7654
rect 17953 7651 18019 7654
rect 18137 7714 18203 7717
rect 20529 7714 20595 7717
rect 18137 7712 20595 7714
rect 18137 7656 18142 7712
rect 18198 7656 20534 7712
rect 20590 7656 20595 7712
rect 18137 7654 20595 7656
rect 18137 7651 18203 7654
rect 20529 7651 20595 7654
rect 9006 7648 9322 7649
rect 9006 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9322 7648
rect 9006 7583 9322 7584
rect 15006 7648 15322 7649
rect 15006 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15322 7648
rect 15006 7583 15322 7584
rect 10133 7578 10199 7581
rect 14733 7578 14799 7581
rect 10133 7576 14799 7578
rect 10133 7520 10138 7576
rect 10194 7520 14738 7576
rect 14794 7520 14799 7576
rect 10133 7518 14799 7520
rect 10133 7515 10199 7518
rect 14733 7515 14799 7518
rect 16113 7578 16179 7581
rect 19885 7578 19951 7581
rect 16113 7576 19951 7578
rect 16113 7520 16118 7576
rect 16174 7520 19890 7576
rect 19946 7520 19951 7576
rect 16113 7518 19951 7520
rect 16113 7515 16179 7518
rect 19885 7515 19951 7518
rect 20069 7578 20135 7581
rect 20670 7578 20730 7790
rect 31109 7787 31175 7790
rect 31385 7850 31451 7853
rect 38653 7850 38719 7853
rect 31385 7848 38719 7850
rect 31385 7792 31390 7848
rect 31446 7792 38658 7848
rect 38714 7792 38719 7848
rect 31385 7790 38719 7792
rect 31385 7787 31451 7790
rect 38653 7787 38719 7790
rect 21449 7714 21515 7717
rect 21582 7714 21588 7716
rect 21449 7712 21588 7714
rect 21449 7656 21454 7712
rect 21510 7656 21588 7712
rect 21449 7654 21588 7656
rect 21449 7651 21515 7654
rect 21582 7652 21588 7654
rect 21652 7652 21658 7716
rect 22185 7714 22251 7717
rect 26785 7714 26851 7717
rect 22185 7712 26851 7714
rect 22185 7656 22190 7712
rect 22246 7656 26790 7712
rect 26846 7656 26851 7712
rect 22185 7654 26851 7656
rect 22185 7651 22251 7654
rect 26785 7651 26851 7654
rect 29637 7714 29703 7717
rect 31385 7714 31451 7717
rect 29637 7712 31451 7714
rect 29637 7656 29642 7712
rect 29698 7656 31390 7712
rect 31446 7656 31451 7712
rect 29637 7654 31451 7656
rect 29637 7651 29703 7654
rect 31385 7651 31451 7654
rect 39389 7714 39455 7717
rect 40880 7714 41000 7744
rect 39389 7712 41000 7714
rect 39389 7656 39394 7712
rect 39450 7656 41000 7712
rect 39389 7654 41000 7656
rect 39389 7651 39455 7654
rect 21006 7648 21322 7649
rect 21006 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21322 7648
rect 21006 7583 21322 7584
rect 27006 7648 27322 7649
rect 27006 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27322 7648
rect 27006 7583 27322 7584
rect 33006 7648 33322 7649
rect 33006 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33322 7648
rect 33006 7583 33322 7584
rect 39006 7648 39322 7649
rect 39006 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39322 7648
rect 40880 7624 41000 7654
rect 39006 7583 39322 7584
rect 25773 7578 25839 7581
rect 26417 7578 26483 7581
rect 20069 7576 20730 7578
rect 20069 7520 20074 7576
rect 20130 7520 20730 7576
rect 20069 7518 20730 7520
rect 22050 7576 26483 7578
rect 22050 7520 25778 7576
rect 25834 7520 26422 7576
rect 26478 7520 26483 7576
rect 22050 7518 26483 7520
rect 20069 7515 20135 7518
rect 1669 7440 4538 7442
rect 1669 7384 1674 7440
rect 1730 7384 4538 7440
rect 1669 7382 4538 7384
rect 4705 7442 4771 7445
rect 9765 7442 9831 7445
rect 4705 7440 9831 7442
rect 4705 7384 4710 7440
rect 4766 7384 9770 7440
rect 9826 7384 9831 7440
rect 4705 7382 9831 7384
rect 1669 7379 1735 7382
rect 4705 7379 4771 7382
rect 9765 7379 9831 7382
rect 10726 7380 10732 7444
rect 10796 7442 10802 7444
rect 13629 7442 13695 7445
rect 10796 7440 13695 7442
rect 10796 7384 13634 7440
rect 13690 7384 13695 7440
rect 10796 7382 13695 7384
rect 10796 7380 10802 7382
rect 13629 7379 13695 7382
rect 14641 7442 14707 7445
rect 21265 7442 21331 7445
rect 14641 7440 21331 7442
rect 14641 7384 14646 7440
rect 14702 7384 21270 7440
rect 21326 7384 21331 7440
rect 14641 7382 21331 7384
rect 14641 7379 14707 7382
rect 21265 7379 21331 7382
rect 2037 7306 2103 7309
rect 6637 7306 6703 7309
rect 8477 7306 8543 7309
rect 2037 7304 6562 7306
rect 2037 7248 2042 7304
rect 2098 7248 6562 7304
rect 2037 7246 6562 7248
rect 2037 7243 2103 7246
rect 0 7170 120 7200
rect 1485 7170 1551 7173
rect 0 7168 1551 7170
rect 0 7112 1490 7168
rect 1546 7112 1551 7168
rect 0 7110 1551 7112
rect 0 7080 120 7110
rect 1485 7107 1551 7110
rect 4838 7108 4844 7172
rect 4908 7170 4914 7172
rect 5257 7170 5323 7173
rect 4908 7168 5323 7170
rect 4908 7112 5262 7168
rect 5318 7112 5323 7168
rect 4908 7110 5323 7112
rect 6502 7170 6562 7246
rect 6637 7304 8543 7306
rect 6637 7248 6642 7304
rect 6698 7248 8482 7304
rect 8538 7248 8543 7304
rect 6637 7246 8543 7248
rect 6637 7243 6703 7246
rect 8477 7243 8543 7246
rect 13077 7306 13143 7309
rect 19609 7306 19675 7309
rect 20805 7306 20871 7309
rect 22050 7306 22110 7518
rect 25773 7515 25839 7518
rect 26417 7515 26483 7518
rect 29729 7578 29795 7581
rect 32121 7578 32187 7581
rect 29729 7576 32187 7578
rect 29729 7520 29734 7576
rect 29790 7520 32126 7576
rect 32182 7520 32187 7576
rect 29729 7518 32187 7520
rect 29729 7515 29795 7518
rect 32121 7515 32187 7518
rect 23381 7442 23447 7445
rect 27429 7442 27495 7445
rect 23381 7440 27495 7442
rect 23381 7384 23386 7440
rect 23442 7384 27434 7440
rect 27490 7384 27495 7440
rect 23381 7382 27495 7384
rect 23381 7379 23447 7382
rect 27429 7379 27495 7382
rect 31201 7442 31267 7445
rect 34789 7442 34855 7445
rect 31201 7440 34855 7442
rect 31201 7384 31206 7440
rect 31262 7384 34794 7440
rect 34850 7384 34855 7440
rect 31201 7382 34855 7384
rect 31201 7379 31267 7382
rect 34789 7379 34855 7382
rect 38929 7442 38995 7445
rect 40880 7442 41000 7472
rect 38929 7440 41000 7442
rect 38929 7384 38934 7440
rect 38990 7384 41000 7440
rect 38929 7382 41000 7384
rect 38929 7379 38995 7382
rect 40880 7352 41000 7382
rect 27337 7306 27403 7309
rect 13077 7304 19675 7306
rect 13077 7248 13082 7304
rect 13138 7248 19614 7304
rect 19670 7248 19675 7304
rect 13077 7246 19675 7248
rect 13077 7243 13143 7246
rect 19609 7243 19675 7246
rect 19750 7246 20408 7306
rect 7005 7170 7071 7173
rect 16665 7170 16731 7173
rect 6502 7168 7071 7170
rect 6502 7112 7010 7168
rect 7066 7112 7071 7168
rect 6502 7110 7071 7112
rect 4908 7108 4914 7110
rect 5257 7107 5323 7110
rect 7005 7107 7071 7110
rect 14414 7168 16731 7170
rect 14414 7112 16670 7168
rect 16726 7112 16731 7168
rect 14414 7110 16731 7112
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 13946 7104 14262 7105
rect 13946 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14262 7104
rect 13946 7039 14262 7040
rect 4981 7034 5047 7037
rect 5390 7034 5396 7036
rect 4981 7032 5396 7034
rect 4981 6976 4986 7032
rect 5042 6976 5396 7032
rect 4981 6974 5396 6976
rect 4981 6971 5047 6974
rect 5390 6972 5396 6974
rect 5460 6972 5466 7036
rect 7189 7034 7255 7037
rect 8569 7036 8635 7037
rect 7782 7034 7788 7036
rect 7189 7032 7788 7034
rect 7189 6976 7194 7032
rect 7250 6976 7788 7032
rect 7189 6974 7788 6976
rect 7189 6971 7255 6974
rect 7782 6972 7788 6974
rect 7852 6972 7858 7036
rect 8518 6972 8524 7036
rect 8588 7034 8635 7036
rect 9673 7034 9739 7037
rect 8588 7032 8680 7034
rect 8630 6976 8680 7032
rect 8588 6974 8680 6976
rect 9673 7032 13738 7034
rect 9673 6976 9678 7032
rect 9734 6976 13738 7032
rect 9673 6974 13738 6976
rect 8588 6972 8635 6974
rect 8569 6971 8635 6972
rect 9673 6971 9739 6974
rect 0 6898 120 6928
rect 1669 6898 1735 6901
rect 0 6896 1735 6898
rect 0 6840 1674 6896
rect 1730 6840 1735 6896
rect 0 6838 1735 6840
rect 0 6808 120 6838
rect 1669 6835 1735 6838
rect 2681 6898 2747 6901
rect 6361 6898 6427 6901
rect 2681 6896 6427 6898
rect 2681 6840 2686 6896
rect 2742 6840 6366 6896
rect 6422 6840 6427 6896
rect 2681 6838 6427 6840
rect 2681 6835 2747 6838
rect 6361 6835 6427 6838
rect 7557 6898 7623 6901
rect 12566 6898 12572 6900
rect 7557 6896 12572 6898
rect 7557 6840 7562 6896
rect 7618 6840 12572 6896
rect 7557 6838 12572 6840
rect 7557 6835 7623 6838
rect 12566 6836 12572 6838
rect 12636 6836 12642 6900
rect 13678 6898 13738 6974
rect 14414 6898 14474 7110
rect 16665 7107 16731 7110
rect 17585 7170 17651 7173
rect 19750 7170 19810 7246
rect 17585 7168 19810 7170
rect 17585 7112 17590 7168
rect 17646 7112 19810 7168
rect 17585 7110 19810 7112
rect 20348 7170 20408 7246
rect 20805 7304 22110 7306
rect 20805 7248 20810 7304
rect 20866 7248 22110 7304
rect 20805 7246 22110 7248
rect 25822 7304 27403 7306
rect 25822 7248 27342 7304
rect 27398 7248 27403 7304
rect 25822 7246 27403 7248
rect 20805 7243 20871 7246
rect 25822 7170 25882 7246
rect 27337 7243 27403 7246
rect 29361 7306 29427 7309
rect 38469 7306 38535 7309
rect 29361 7304 38535 7306
rect 29361 7248 29366 7304
rect 29422 7248 38474 7304
rect 38530 7248 38535 7304
rect 29361 7246 38535 7248
rect 29361 7243 29427 7246
rect 38469 7243 38535 7246
rect 20348 7110 25882 7170
rect 26417 7170 26483 7173
rect 31477 7170 31543 7173
rect 26417 7168 31543 7170
rect 26417 7112 26422 7168
rect 26478 7112 31482 7168
rect 31538 7112 31543 7168
rect 26417 7110 31543 7112
rect 17585 7107 17651 7110
rect 26417 7107 26483 7110
rect 31477 7107 31543 7110
rect 39389 7170 39455 7173
rect 40880 7170 41000 7200
rect 39389 7168 41000 7170
rect 39389 7112 39394 7168
rect 39450 7112 41000 7168
rect 39389 7110 41000 7112
rect 39389 7107 39455 7110
rect 19946 7104 20262 7105
rect 19946 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20262 7104
rect 19946 7039 20262 7040
rect 25946 7104 26262 7105
rect 25946 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26262 7104
rect 25946 7039 26262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 37946 7104 38262 7105
rect 37946 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38262 7104
rect 40880 7080 41000 7110
rect 37946 7039 38262 7040
rect 14549 7034 14615 7037
rect 15929 7034 15995 7037
rect 14549 7032 15995 7034
rect 14549 6976 14554 7032
rect 14610 6976 15934 7032
rect 15990 6976 15995 7032
rect 14549 6974 15995 6976
rect 14549 6971 14615 6974
rect 15929 6971 15995 6974
rect 16297 7034 16363 7037
rect 16430 7034 16436 7036
rect 16297 7032 16436 7034
rect 16297 6976 16302 7032
rect 16358 6976 16436 7032
rect 16297 6974 16436 6976
rect 16297 6971 16363 6974
rect 16430 6972 16436 6974
rect 16500 6972 16506 7036
rect 16757 7034 16823 7037
rect 17401 7034 17467 7037
rect 16757 7032 17467 7034
rect 16757 6976 16762 7032
rect 16818 6976 17406 7032
rect 17462 6976 17467 7032
rect 16757 6974 17467 6976
rect 16757 6971 16823 6974
rect 17401 6971 17467 6974
rect 19057 7034 19123 7037
rect 19517 7034 19583 7037
rect 19057 7032 19583 7034
rect 19057 6976 19062 7032
rect 19118 6976 19522 7032
rect 19578 6976 19583 7032
rect 19057 6974 19583 6976
rect 19057 6971 19123 6974
rect 19517 6971 19583 6974
rect 20846 6972 20852 7036
rect 20916 7034 20922 7036
rect 24945 7034 25011 7037
rect 20916 7032 25011 7034
rect 20916 6976 24950 7032
rect 25006 6976 25011 7032
rect 20916 6974 25011 6976
rect 20916 6972 20922 6974
rect 24945 6971 25011 6974
rect 25589 7036 25655 7037
rect 25589 7032 25636 7036
rect 25700 7034 25706 7036
rect 27337 7034 27403 7037
rect 29085 7034 29151 7037
rect 25589 6976 25594 7032
rect 25589 6972 25636 6976
rect 25700 6974 25746 7034
rect 27337 7032 29151 7034
rect 27337 6976 27342 7032
rect 27398 6976 29090 7032
rect 29146 6976 29151 7032
rect 27337 6974 29151 6976
rect 25700 6972 25706 6974
rect 25589 6971 25655 6972
rect 27337 6971 27403 6974
rect 29085 6971 29151 6974
rect 13678 6838 14474 6898
rect 14549 6898 14615 6901
rect 15561 6898 15627 6901
rect 14549 6896 15627 6898
rect 14549 6840 14554 6896
rect 14610 6840 15566 6896
rect 15622 6840 15627 6896
rect 14549 6838 15627 6840
rect 14549 6835 14615 6838
rect 15561 6835 15627 6838
rect 15837 6898 15903 6901
rect 21173 6898 21239 6901
rect 15837 6896 21239 6898
rect 15837 6840 15842 6896
rect 15898 6840 21178 6896
rect 21234 6840 21239 6896
rect 15837 6838 21239 6840
rect 15837 6835 15903 6838
rect 21173 6835 21239 6838
rect 21582 6836 21588 6900
rect 21652 6898 21658 6900
rect 26785 6898 26851 6901
rect 21652 6896 26851 6898
rect 21652 6840 26790 6896
rect 26846 6840 26851 6896
rect 21652 6838 26851 6840
rect 21652 6836 21658 6838
rect 26785 6835 26851 6838
rect 29177 6898 29243 6901
rect 34329 6898 34395 6901
rect 29177 6896 34395 6898
rect 29177 6840 29182 6896
rect 29238 6840 34334 6896
rect 34390 6840 34395 6896
rect 29177 6838 34395 6840
rect 29177 6835 29243 6838
rect 34329 6835 34395 6838
rect 40033 6898 40099 6901
rect 40880 6898 41000 6928
rect 40033 6896 41000 6898
rect 40033 6840 40038 6896
rect 40094 6840 41000 6896
rect 40033 6838 41000 6840
rect 40033 6835 40099 6838
rect 40880 6808 41000 6838
rect 4889 6762 4955 6765
rect 10777 6762 10843 6765
rect 4889 6760 10843 6762
rect 4889 6704 4894 6760
rect 4950 6704 10782 6760
rect 10838 6704 10843 6760
rect 4889 6702 10843 6704
rect 4889 6699 4955 6702
rect 10777 6699 10843 6702
rect 12525 6762 12591 6765
rect 20713 6762 20779 6765
rect 21449 6762 21515 6765
rect 12525 6760 20779 6762
rect 12525 6704 12530 6760
rect 12586 6704 20718 6760
rect 20774 6704 20779 6760
rect 12525 6702 20779 6704
rect 12525 6699 12591 6702
rect 20713 6699 20779 6702
rect 20854 6760 21515 6762
rect 20854 6704 21454 6760
rect 21510 6704 21515 6760
rect 20854 6702 21515 6704
rect 0 6626 120 6656
rect 1393 6626 1459 6629
rect 0 6624 1459 6626
rect 0 6568 1398 6624
rect 1454 6568 1459 6624
rect 0 6566 1459 6568
rect 0 6536 120 6566
rect 1393 6563 1459 6566
rect 5349 6626 5415 6629
rect 5717 6626 5783 6629
rect 8518 6626 8524 6628
rect 5349 6624 8524 6626
rect 5349 6568 5354 6624
rect 5410 6568 5722 6624
rect 5778 6568 8524 6624
rect 5349 6566 8524 6568
rect 5349 6563 5415 6566
rect 5717 6563 5783 6566
rect 8518 6564 8524 6566
rect 8588 6564 8594 6628
rect 9673 6626 9739 6629
rect 12433 6626 12499 6629
rect 9673 6624 12499 6626
rect 9673 6568 9678 6624
rect 9734 6568 12438 6624
rect 12494 6568 12499 6624
rect 9673 6566 12499 6568
rect 9673 6563 9739 6566
rect 12433 6563 12499 6566
rect 12750 6564 12756 6628
rect 12820 6626 12826 6628
rect 14549 6626 14615 6629
rect 12820 6624 14615 6626
rect 12820 6568 14554 6624
rect 14610 6568 14615 6624
rect 12820 6566 14615 6568
rect 12820 6564 12826 6566
rect 14549 6563 14615 6566
rect 15561 6626 15627 6629
rect 17309 6626 17375 6629
rect 20854 6626 20914 6702
rect 21449 6699 21515 6702
rect 22093 6762 22159 6765
rect 25957 6762 26023 6765
rect 22093 6760 26023 6762
rect 22093 6704 22098 6760
rect 22154 6704 25962 6760
rect 26018 6704 26023 6760
rect 22093 6702 26023 6704
rect 22093 6699 22159 6702
rect 25957 6699 26023 6702
rect 26509 6762 26575 6765
rect 32213 6762 32279 6765
rect 34513 6762 34579 6765
rect 26509 6760 34579 6762
rect 26509 6704 26514 6760
rect 26570 6704 32218 6760
rect 32274 6704 34518 6760
rect 34574 6704 34579 6760
rect 26509 6702 34579 6704
rect 26509 6699 26575 6702
rect 32213 6699 32279 6702
rect 34513 6699 34579 6702
rect 15561 6624 20914 6626
rect 15561 6568 15566 6624
rect 15622 6568 17314 6624
rect 17370 6568 20914 6624
rect 15561 6566 20914 6568
rect 21449 6626 21515 6629
rect 25405 6626 25471 6629
rect 21449 6624 25471 6626
rect 21449 6568 21454 6624
rect 21510 6568 25410 6624
rect 25466 6568 25471 6624
rect 21449 6566 25471 6568
rect 15561 6563 15627 6566
rect 17309 6563 17375 6566
rect 21449 6563 21515 6566
rect 25405 6563 25471 6566
rect 36629 6626 36695 6629
rect 38377 6626 38443 6629
rect 36629 6624 38443 6626
rect 36629 6568 36634 6624
rect 36690 6568 38382 6624
rect 38438 6568 38443 6624
rect 36629 6566 38443 6568
rect 36629 6563 36695 6566
rect 38377 6563 38443 6566
rect 39389 6626 39455 6629
rect 40880 6626 41000 6656
rect 39389 6624 41000 6626
rect 39389 6568 39394 6624
rect 39450 6568 41000 6624
rect 39389 6566 41000 6568
rect 39389 6563 39455 6566
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 9006 6560 9322 6561
rect 9006 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9322 6560
rect 9006 6495 9322 6496
rect 15006 6560 15322 6561
rect 15006 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15322 6560
rect 15006 6495 15322 6496
rect 21006 6560 21322 6561
rect 21006 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21322 6560
rect 21006 6495 21322 6496
rect 27006 6560 27322 6561
rect 27006 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27322 6560
rect 27006 6495 27322 6496
rect 33006 6560 33322 6561
rect 33006 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33322 6560
rect 33006 6495 33322 6496
rect 39006 6560 39322 6561
rect 39006 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39322 6560
rect 40880 6536 41000 6566
rect 39006 6495 39322 6496
rect 8017 6490 8083 6493
rect 15653 6490 15719 6493
rect 17493 6490 17559 6493
rect 7422 6488 8083 6490
rect 7422 6432 8022 6488
rect 8078 6432 8083 6488
rect 7422 6430 8083 6432
rect 0 6354 120 6384
rect 1577 6354 1643 6357
rect 7422 6354 7482 6430
rect 8017 6427 8083 6430
rect 10182 6430 14842 6490
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 120 6294
rect 1577 6291 1643 6294
rect 2730 6294 7482 6354
rect 7649 6354 7715 6357
rect 10041 6354 10107 6357
rect 10182 6354 10242 6430
rect 12709 6354 12775 6357
rect 7649 6352 10242 6354
rect 7649 6296 7654 6352
rect 7710 6296 10046 6352
rect 10102 6296 10242 6352
rect 7649 6294 10242 6296
rect 12022 6352 12775 6354
rect 12022 6296 12714 6352
rect 12770 6296 12775 6352
rect 12022 6294 12775 6296
rect 1761 6218 1827 6221
rect 2730 6218 2790 6294
rect 7649 6291 7715 6294
rect 10041 6291 10107 6294
rect 1761 6216 2790 6218
rect 1761 6160 1766 6216
rect 1822 6160 2790 6216
rect 1761 6158 2790 6160
rect 3693 6218 3759 6221
rect 3693 6216 8402 6218
rect 3693 6160 3698 6216
rect 3754 6160 8402 6216
rect 3693 6158 8402 6160
rect 1761 6155 1827 6158
rect 3693 6155 3759 6158
rect 0 6082 120 6112
rect 1393 6082 1459 6085
rect 0 6080 1459 6082
rect 0 6024 1398 6080
rect 1454 6024 1459 6080
rect 0 6022 1459 6024
rect 0 5992 120 6022
rect 1393 6019 1459 6022
rect 3693 6082 3759 6085
rect 4521 6082 4587 6085
rect 3693 6080 4587 6082
rect 3693 6024 3698 6080
rect 3754 6024 4526 6080
rect 4582 6024 4587 6080
rect 3693 6022 4587 6024
rect 3693 6019 3759 6022
rect 4521 6019 4587 6022
rect 5809 6082 5875 6085
rect 7465 6082 7531 6085
rect 5809 6080 7531 6082
rect 5809 6024 5814 6080
rect 5870 6024 7470 6080
rect 7526 6024 7531 6080
rect 5809 6022 7531 6024
rect 5809 6019 5875 6022
rect 7465 6019 7531 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 3141 5946 3207 5949
rect 6453 5946 6519 5949
rect 3141 5944 6519 5946
rect 3141 5888 3146 5944
rect 3202 5888 6458 5944
rect 6514 5888 6519 5944
rect 3141 5886 6519 5888
rect 8342 5946 8402 6158
rect 8518 6156 8524 6220
rect 8588 6218 8594 6220
rect 12022 6218 12082 6294
rect 12709 6291 12775 6294
rect 13261 6356 13327 6357
rect 13261 6352 13308 6356
rect 13372 6354 13378 6356
rect 13537 6354 13603 6357
rect 14590 6354 14596 6356
rect 13261 6296 13266 6352
rect 13261 6292 13308 6296
rect 13372 6294 13418 6354
rect 13537 6352 14596 6354
rect 13537 6296 13542 6352
rect 13598 6296 14596 6352
rect 13537 6294 14596 6296
rect 13372 6292 13378 6294
rect 13261 6291 13327 6292
rect 13537 6291 13603 6294
rect 14590 6292 14596 6294
rect 14660 6292 14666 6356
rect 14782 6354 14842 6430
rect 15653 6488 17559 6490
rect 15653 6432 15658 6488
rect 15714 6432 17498 6488
rect 17554 6432 17559 6488
rect 15653 6430 17559 6432
rect 15653 6427 15719 6430
rect 17493 6427 17559 6430
rect 17677 6490 17743 6493
rect 17677 6488 20546 6490
rect 17677 6432 17682 6488
rect 17738 6432 20546 6488
rect 17677 6430 20546 6432
rect 17677 6427 17743 6430
rect 16297 6354 16363 6357
rect 14782 6352 16363 6354
rect 14782 6296 16302 6352
rect 16358 6296 16363 6352
rect 14782 6294 16363 6296
rect 16297 6291 16363 6294
rect 16849 6354 16915 6357
rect 20345 6354 20411 6357
rect 16849 6352 20411 6354
rect 16849 6296 16854 6352
rect 16910 6296 20350 6352
rect 20406 6296 20411 6352
rect 16849 6294 20411 6296
rect 16849 6291 16915 6294
rect 20345 6291 20411 6294
rect 8588 6158 12082 6218
rect 12249 6218 12315 6221
rect 18137 6218 18203 6221
rect 20486 6218 20546 6430
rect 24158 6428 24164 6492
rect 24228 6490 24234 6492
rect 26693 6490 26759 6493
rect 24228 6488 26759 6490
rect 24228 6432 26698 6488
rect 26754 6432 26759 6488
rect 24228 6430 26759 6432
rect 24228 6428 24234 6430
rect 26693 6427 26759 6430
rect 27429 6490 27495 6493
rect 29269 6490 29335 6493
rect 30833 6490 30899 6493
rect 27429 6488 30899 6490
rect 27429 6432 27434 6488
rect 27490 6432 29274 6488
rect 29330 6432 30838 6488
rect 30894 6432 30899 6488
rect 27429 6430 30899 6432
rect 27429 6427 27495 6430
rect 29269 6427 29335 6430
rect 30833 6427 30899 6430
rect 21817 6354 21883 6357
rect 32305 6354 32371 6357
rect 21817 6352 32371 6354
rect 21817 6296 21822 6352
rect 21878 6296 32310 6352
rect 32366 6296 32371 6352
rect 21817 6294 32371 6296
rect 21817 6291 21883 6294
rect 32305 6291 32371 6294
rect 32489 6354 32555 6357
rect 33409 6354 33475 6357
rect 35893 6354 35959 6357
rect 32489 6352 35959 6354
rect 32489 6296 32494 6352
rect 32550 6296 33414 6352
rect 33470 6296 35898 6352
rect 35954 6296 35959 6352
rect 32489 6294 35959 6296
rect 32489 6291 32555 6294
rect 33409 6291 33475 6294
rect 35893 6291 35959 6294
rect 39389 6354 39455 6357
rect 40880 6354 41000 6384
rect 39389 6352 41000 6354
rect 39389 6296 39394 6352
rect 39450 6296 41000 6352
rect 39389 6294 41000 6296
rect 39389 6291 39455 6294
rect 40880 6264 41000 6294
rect 24117 6218 24183 6221
rect 26693 6218 26759 6221
rect 28441 6218 28507 6221
rect 12249 6216 18203 6218
rect 12249 6160 12254 6216
rect 12310 6160 18142 6216
rect 18198 6160 18203 6216
rect 12249 6158 18203 6160
rect 8588 6156 8594 6158
rect 12249 6155 12315 6158
rect 18137 6155 18203 6158
rect 18278 6158 20408 6218
rect 20486 6216 24183 6218
rect 20486 6160 24122 6216
rect 24178 6160 24183 6216
rect 20486 6158 24183 6160
rect 8569 6082 8635 6085
rect 9438 6082 9444 6084
rect 8569 6080 9444 6082
rect 8569 6024 8574 6080
rect 8630 6024 9444 6080
rect 8569 6022 9444 6024
rect 8569 6019 8635 6022
rect 9438 6020 9444 6022
rect 9508 6020 9514 6084
rect 10225 6082 10291 6085
rect 12433 6082 12499 6085
rect 10225 6080 12499 6082
rect 10225 6024 10230 6080
rect 10286 6024 12438 6080
rect 12494 6024 12499 6080
rect 10225 6022 12499 6024
rect 10225 6019 10291 6022
rect 12433 6019 12499 6022
rect 12566 6020 12572 6084
rect 12636 6082 12642 6084
rect 12893 6082 12959 6085
rect 18278 6082 18338 6158
rect 12636 6080 12959 6082
rect 12636 6024 12898 6080
rect 12954 6024 12959 6080
rect 12636 6022 12959 6024
rect 12636 6020 12642 6022
rect 12893 6019 12959 6022
rect 14598 6022 18338 6082
rect 20348 6082 20408 6158
rect 24117 6155 24183 6158
rect 24350 6158 26434 6218
rect 21817 6082 21883 6085
rect 23013 6082 23079 6085
rect 20348 6080 21883 6082
rect 20348 6024 21822 6080
rect 21878 6024 21883 6080
rect 20348 6022 21883 6024
rect 13946 6016 14262 6017
rect 13946 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14262 6016
rect 13946 5951 14262 5952
rect 12566 5946 12572 5948
rect 8342 5886 12572 5946
rect 3141 5883 3207 5886
rect 6453 5883 6519 5886
rect 12566 5884 12572 5886
rect 12636 5946 12642 5948
rect 13670 5946 13676 5948
rect 12636 5886 13676 5946
rect 12636 5884 12642 5886
rect 13670 5884 13676 5886
rect 13740 5884 13746 5948
rect 14598 5946 14658 6022
rect 21817 6019 21883 6022
rect 22004 6080 23079 6082
rect 22004 6024 23018 6080
rect 23074 6024 23079 6080
rect 22004 6022 23079 6024
rect 19946 6016 20262 6017
rect 19946 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20262 6016
rect 19946 5951 20262 5952
rect 14414 5886 14658 5946
rect 14825 5946 14891 5949
rect 19425 5946 19491 5949
rect 14825 5944 19491 5946
rect 14825 5888 14830 5944
rect 14886 5888 19430 5944
rect 19486 5888 19491 5944
rect 14825 5886 19491 5888
rect 0 5810 120 5840
rect 1485 5810 1551 5813
rect 0 5808 1551 5810
rect 0 5752 1490 5808
rect 1546 5752 1551 5808
rect 0 5750 1551 5752
rect 0 5720 120 5750
rect 1485 5747 1551 5750
rect 1945 5810 2011 5813
rect 9765 5810 9831 5813
rect 12750 5810 12756 5812
rect 1945 5808 9690 5810
rect 1945 5752 1950 5808
rect 2006 5752 9690 5808
rect 1945 5750 9690 5752
rect 1945 5747 2011 5750
rect 4981 5674 5047 5677
rect 6637 5676 6703 5677
rect 5206 5674 5212 5676
rect 4981 5672 5212 5674
rect 4981 5616 4986 5672
rect 5042 5616 5212 5672
rect 4981 5614 5212 5616
rect 4981 5611 5047 5614
rect 5206 5612 5212 5614
rect 5276 5612 5282 5676
rect 6637 5672 6684 5676
rect 6748 5674 6754 5676
rect 7005 5674 7071 5677
rect 7598 5674 7604 5676
rect 6637 5616 6642 5672
rect 6637 5612 6684 5616
rect 6748 5614 6794 5674
rect 7005 5672 7604 5674
rect 7005 5616 7010 5672
rect 7066 5616 7604 5672
rect 7005 5614 7604 5616
rect 6748 5612 6754 5614
rect 6637 5611 6703 5612
rect 7005 5611 7071 5614
rect 7598 5612 7604 5614
rect 7668 5674 7674 5676
rect 8569 5674 8635 5677
rect 7668 5672 8635 5674
rect 7668 5616 8574 5672
rect 8630 5616 8635 5672
rect 7668 5614 8635 5616
rect 7668 5612 7674 5614
rect 8569 5611 8635 5614
rect 8710 5614 9506 5674
rect 0 5538 120 5568
rect 2221 5538 2287 5541
rect 0 5536 2287 5538
rect 0 5480 2226 5536
rect 2282 5480 2287 5536
rect 0 5478 2287 5480
rect 0 5448 120 5478
rect 2221 5475 2287 5478
rect 4981 5538 5047 5541
rect 5717 5538 5783 5541
rect 5993 5540 6059 5541
rect 4981 5536 5783 5538
rect 4981 5480 4986 5536
rect 5042 5480 5722 5536
rect 5778 5480 5783 5536
rect 4981 5478 5783 5480
rect 4981 5475 5047 5478
rect 5717 5475 5783 5478
rect 5942 5476 5948 5540
rect 6012 5538 6059 5540
rect 6913 5538 6979 5541
rect 8710 5538 8770 5614
rect 6012 5536 6104 5538
rect 6054 5480 6104 5536
rect 6012 5478 6104 5480
rect 6913 5536 8770 5538
rect 6913 5480 6918 5536
rect 6974 5480 8770 5536
rect 6913 5478 8770 5480
rect 6012 5476 6059 5478
rect 5993 5475 6059 5476
rect 6913 5475 6979 5478
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 9006 5472 9322 5473
rect 9006 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9322 5472
rect 9006 5407 9322 5408
rect 3417 5402 3483 5405
rect 4705 5402 4771 5405
rect 3417 5400 4771 5402
rect 3417 5344 3422 5400
rect 3478 5344 4710 5400
rect 4766 5344 4771 5400
rect 3417 5342 4771 5344
rect 3417 5339 3483 5342
rect 4705 5339 4771 5342
rect 4889 5402 4955 5405
rect 7189 5402 7255 5405
rect 4889 5400 7255 5402
rect 4889 5344 4894 5400
rect 4950 5344 7194 5400
rect 7250 5344 7255 5400
rect 4889 5342 7255 5344
rect 4889 5339 4955 5342
rect 7189 5339 7255 5342
rect 7414 5340 7420 5404
rect 7484 5402 7490 5404
rect 8334 5402 8340 5404
rect 7484 5342 8340 5402
rect 7484 5340 7490 5342
rect 8334 5340 8340 5342
rect 8404 5340 8410 5404
rect 8518 5340 8524 5404
rect 8588 5402 8594 5404
rect 8661 5402 8727 5405
rect 8588 5400 8727 5402
rect 8588 5344 8666 5400
rect 8722 5344 8727 5400
rect 8588 5342 8727 5344
rect 9446 5402 9506 5614
rect 9630 5538 9690 5750
rect 9765 5808 12756 5810
rect 9765 5752 9770 5808
rect 9826 5752 12756 5808
rect 9765 5750 12756 5752
rect 9765 5747 9831 5750
rect 12750 5748 12756 5750
rect 12820 5748 12826 5812
rect 12985 5810 13051 5813
rect 13486 5810 13492 5812
rect 12985 5808 13492 5810
rect 12985 5752 12990 5808
rect 13046 5752 13492 5808
rect 12985 5750 13492 5752
rect 12985 5747 13051 5750
rect 13486 5748 13492 5750
rect 13556 5810 13562 5812
rect 14414 5810 14474 5886
rect 14825 5883 14891 5886
rect 19425 5883 19491 5886
rect 20529 5946 20595 5949
rect 22004 5946 22064 6022
rect 23013 6019 23079 6022
rect 20529 5944 22064 5946
rect 20529 5888 20534 5944
rect 20590 5888 22064 5944
rect 20529 5886 22064 5888
rect 20529 5883 20595 5886
rect 22134 5884 22140 5948
rect 22204 5946 22210 5948
rect 24350 5946 24410 6158
rect 26374 6082 26434 6158
rect 26693 6216 28507 6218
rect 26693 6160 26698 6216
rect 26754 6160 28446 6216
rect 28502 6160 28507 6216
rect 26693 6158 28507 6160
rect 26693 6155 26759 6158
rect 28441 6155 28507 6158
rect 28809 6218 28875 6221
rect 39205 6218 39271 6221
rect 28809 6216 39271 6218
rect 28809 6160 28814 6216
rect 28870 6160 39210 6216
rect 39266 6160 39271 6216
rect 28809 6158 39271 6160
rect 28809 6155 28875 6158
rect 39205 6155 39271 6158
rect 29177 6082 29243 6085
rect 26374 6080 29243 6082
rect 26374 6024 29182 6080
rect 29238 6024 29243 6080
rect 26374 6022 29243 6024
rect 29177 6019 29243 6022
rect 39021 6082 39087 6085
rect 40880 6082 41000 6112
rect 39021 6080 41000 6082
rect 39021 6024 39026 6080
rect 39082 6024 41000 6080
rect 39021 6022 41000 6024
rect 39021 6019 39087 6022
rect 25946 6016 26262 6017
rect 25946 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26262 6016
rect 25946 5951 26262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 37946 6016 38262 6017
rect 37946 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38262 6016
rect 40880 5992 41000 6022
rect 37946 5951 38262 5952
rect 22204 5886 24410 5946
rect 22204 5884 22210 5886
rect 25262 5884 25268 5948
rect 25332 5946 25338 5948
rect 25497 5946 25563 5949
rect 27061 5946 27127 5949
rect 25332 5944 25563 5946
rect 25332 5888 25502 5944
rect 25558 5888 25563 5944
rect 25332 5886 25563 5888
rect 25332 5884 25338 5886
rect 25497 5883 25563 5886
rect 26604 5944 27127 5946
rect 26604 5888 27066 5944
rect 27122 5888 27127 5944
rect 26604 5886 27127 5888
rect 17953 5810 18019 5813
rect 22645 5810 22711 5813
rect 26604 5810 26664 5886
rect 27061 5883 27127 5886
rect 13556 5750 14474 5810
rect 14598 5808 18019 5810
rect 14598 5752 17958 5808
rect 18014 5752 18019 5808
rect 14598 5750 18019 5752
rect 13556 5748 13562 5750
rect 9765 5674 9831 5677
rect 11697 5674 11763 5677
rect 9765 5672 11763 5674
rect 9765 5616 9770 5672
rect 9826 5616 11702 5672
rect 11758 5616 11763 5672
rect 9765 5614 11763 5616
rect 9765 5611 9831 5614
rect 11697 5611 11763 5614
rect 12249 5674 12315 5677
rect 14598 5674 14658 5750
rect 17953 5747 18019 5750
rect 18094 5808 22711 5810
rect 18094 5752 22650 5808
rect 22706 5752 22711 5808
rect 18094 5750 22711 5752
rect 16021 5674 16087 5677
rect 17677 5674 17743 5677
rect 12249 5672 14658 5674
rect 12249 5616 12254 5672
rect 12310 5616 14658 5672
rect 12249 5614 14658 5616
rect 14782 5614 15578 5674
rect 12249 5611 12315 5614
rect 12709 5538 12775 5541
rect 9630 5536 12775 5538
rect 9630 5480 12714 5536
rect 12770 5480 12775 5536
rect 9630 5478 12775 5480
rect 12709 5475 12775 5478
rect 13261 5538 13327 5541
rect 14641 5538 14707 5541
rect 13261 5536 14707 5538
rect 13261 5480 13266 5536
rect 13322 5480 14646 5536
rect 14702 5480 14707 5536
rect 13261 5478 14707 5480
rect 13261 5475 13327 5478
rect 14641 5475 14707 5478
rect 10542 5402 10548 5404
rect 9446 5342 10548 5402
rect 8588 5340 8594 5342
rect 8661 5339 8727 5342
rect 10542 5340 10548 5342
rect 10612 5340 10618 5404
rect 11145 5402 11211 5405
rect 14782 5402 14842 5614
rect 15518 5538 15578 5614
rect 16021 5672 17743 5674
rect 16021 5616 16026 5672
rect 16082 5616 17682 5672
rect 17738 5616 17743 5672
rect 16021 5614 17743 5616
rect 16021 5611 16087 5614
rect 17677 5611 17743 5614
rect 18094 5538 18154 5750
rect 22645 5747 22711 5750
rect 25684 5750 26664 5810
rect 26785 5810 26851 5813
rect 33777 5810 33843 5813
rect 26785 5808 33843 5810
rect 26785 5752 26790 5808
rect 26846 5752 33782 5808
rect 33838 5752 33843 5808
rect 26785 5750 33843 5752
rect 18321 5674 18387 5677
rect 21817 5674 21883 5677
rect 18321 5672 21883 5674
rect 18321 5616 18326 5672
rect 18382 5616 21822 5672
rect 21878 5616 21883 5672
rect 18321 5614 21883 5616
rect 18321 5611 18387 5614
rect 21817 5611 21883 5614
rect 22185 5674 22251 5677
rect 22737 5674 22803 5677
rect 22185 5672 22803 5674
rect 22185 5616 22190 5672
rect 22246 5616 22742 5672
rect 22798 5616 22803 5672
rect 22185 5614 22803 5616
rect 22185 5611 22251 5614
rect 22737 5611 22803 5614
rect 23013 5674 23079 5677
rect 23473 5674 23539 5677
rect 25684 5674 25744 5750
rect 26785 5747 26851 5750
rect 33777 5747 33843 5750
rect 39389 5810 39455 5813
rect 40880 5810 41000 5840
rect 39389 5808 41000 5810
rect 39389 5752 39394 5808
rect 39450 5752 41000 5808
rect 39389 5750 41000 5752
rect 39389 5747 39455 5750
rect 40880 5720 41000 5750
rect 23013 5672 25744 5674
rect 23013 5616 23018 5672
rect 23074 5616 23478 5672
rect 23534 5616 25744 5672
rect 23013 5614 25744 5616
rect 25865 5674 25931 5677
rect 31293 5674 31359 5677
rect 25865 5672 31359 5674
rect 25865 5616 25870 5672
rect 25926 5616 31298 5672
rect 31354 5616 31359 5672
rect 25865 5614 31359 5616
rect 23013 5611 23079 5614
rect 23473 5611 23539 5614
rect 25865 5611 25931 5614
rect 31293 5611 31359 5614
rect 32305 5674 32371 5677
rect 35249 5674 35315 5677
rect 32305 5672 35315 5674
rect 32305 5616 32310 5672
rect 32366 5616 35254 5672
rect 35310 5616 35315 5672
rect 32305 5614 35315 5616
rect 32305 5611 32371 5614
rect 35249 5611 35315 5614
rect 15518 5478 18154 5538
rect 18873 5538 18939 5541
rect 19885 5538 19951 5541
rect 20437 5538 20503 5541
rect 18873 5536 20503 5538
rect 18873 5480 18878 5536
rect 18934 5480 19890 5536
rect 19946 5480 20442 5536
rect 20498 5480 20503 5536
rect 18873 5478 20503 5480
rect 18873 5475 18939 5478
rect 19885 5475 19951 5478
rect 20437 5475 20503 5478
rect 22369 5538 22435 5541
rect 26141 5538 26207 5541
rect 22369 5536 26207 5538
rect 22369 5480 22374 5536
rect 22430 5480 26146 5536
rect 26202 5480 26207 5536
rect 22369 5478 26207 5480
rect 22369 5475 22435 5478
rect 26141 5475 26207 5478
rect 28625 5538 28691 5541
rect 32673 5538 32739 5541
rect 28625 5536 32739 5538
rect 28625 5480 28630 5536
rect 28686 5480 32678 5536
rect 32734 5480 32739 5536
rect 28625 5478 32739 5480
rect 28625 5475 28691 5478
rect 32673 5475 32739 5478
rect 39941 5538 40007 5541
rect 40880 5538 41000 5568
rect 39941 5536 41000 5538
rect 39941 5480 39946 5536
rect 40002 5480 41000 5536
rect 39941 5478 41000 5480
rect 39941 5475 40007 5478
rect 15006 5472 15322 5473
rect 15006 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15322 5472
rect 15006 5407 15322 5408
rect 21006 5472 21322 5473
rect 21006 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21322 5472
rect 21006 5407 21322 5408
rect 27006 5472 27322 5473
rect 27006 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27322 5472
rect 27006 5407 27322 5408
rect 33006 5472 33322 5473
rect 33006 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33322 5472
rect 33006 5407 33322 5408
rect 39006 5472 39322 5473
rect 39006 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39322 5472
rect 40880 5448 41000 5478
rect 39006 5407 39322 5408
rect 11145 5400 14842 5402
rect 11145 5344 11150 5400
rect 11206 5344 14842 5400
rect 11145 5342 14842 5344
rect 15469 5402 15535 5405
rect 23381 5402 23447 5405
rect 24117 5402 24183 5405
rect 15469 5400 20730 5402
rect 15469 5344 15474 5400
rect 15530 5344 20730 5400
rect 15469 5342 20730 5344
rect 11145 5339 11211 5342
rect 15469 5339 15535 5342
rect 0 5266 120 5296
rect 1853 5266 1919 5269
rect 0 5264 1919 5266
rect 0 5208 1858 5264
rect 1914 5208 1919 5264
rect 0 5206 1919 5208
rect 0 5176 120 5206
rect 1853 5203 1919 5206
rect 3601 5266 3667 5269
rect 3734 5266 3740 5268
rect 3601 5264 3740 5266
rect 3601 5208 3606 5264
rect 3662 5208 3740 5264
rect 3601 5206 3740 5208
rect 3601 5203 3667 5206
rect 3734 5204 3740 5206
rect 3804 5204 3810 5268
rect 3877 5266 3943 5269
rect 20670 5266 20730 5342
rect 23381 5400 24183 5402
rect 23381 5344 23386 5400
rect 23442 5344 24122 5400
rect 24178 5344 24183 5400
rect 23381 5342 24183 5344
rect 23381 5339 23447 5342
rect 24117 5339 24183 5342
rect 24393 5402 24459 5405
rect 25405 5402 25471 5405
rect 24393 5400 25471 5402
rect 24393 5344 24398 5400
rect 24454 5344 25410 5400
rect 25466 5344 25471 5400
rect 24393 5342 25471 5344
rect 24393 5339 24459 5342
rect 25405 5339 25471 5342
rect 27429 5402 27495 5405
rect 27654 5402 27660 5404
rect 27429 5400 27660 5402
rect 27429 5344 27434 5400
rect 27490 5344 27660 5400
rect 27429 5342 27660 5344
rect 27429 5339 27495 5342
rect 27654 5340 27660 5342
rect 27724 5340 27730 5404
rect 30833 5402 30899 5405
rect 31661 5402 31727 5405
rect 30833 5400 31727 5402
rect 30833 5344 30838 5400
rect 30894 5344 31666 5400
rect 31722 5344 31727 5400
rect 30833 5342 31727 5344
rect 30833 5339 30899 5342
rect 31661 5339 31727 5342
rect 25773 5266 25839 5269
rect 3877 5264 20592 5266
rect 3877 5208 3882 5264
rect 3938 5208 20592 5264
rect 3877 5206 20592 5208
rect 20670 5264 25839 5266
rect 20670 5208 25778 5264
rect 25834 5208 25839 5264
rect 20670 5206 25839 5208
rect 3877 5203 3943 5206
rect 2497 5130 2563 5133
rect 5165 5130 5231 5133
rect 2497 5128 5231 5130
rect 2497 5072 2502 5128
rect 2558 5072 5170 5128
rect 5226 5072 5231 5128
rect 2497 5070 5231 5072
rect 2497 5067 2563 5070
rect 5165 5067 5231 5070
rect 7005 5130 7071 5133
rect 20532 5130 20592 5206
rect 25773 5203 25839 5206
rect 26877 5266 26943 5269
rect 38837 5266 38903 5269
rect 26877 5264 38903 5266
rect 26877 5208 26882 5264
rect 26938 5208 38842 5264
rect 38898 5208 38903 5264
rect 26877 5206 38903 5208
rect 26877 5203 26943 5206
rect 38837 5203 38903 5206
rect 39389 5266 39455 5269
rect 40880 5266 41000 5296
rect 39389 5264 41000 5266
rect 39389 5208 39394 5264
rect 39450 5208 41000 5264
rect 39389 5206 41000 5208
rect 39389 5203 39455 5206
rect 40880 5176 41000 5206
rect 24209 5130 24275 5133
rect 27521 5130 27587 5133
rect 32305 5130 32371 5133
rect 7005 5128 20408 5130
rect 7005 5072 7010 5128
rect 7066 5072 20408 5128
rect 7005 5070 20408 5072
rect 20532 5070 23490 5130
rect 7005 5067 7071 5070
rect 0 4994 120 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 120 4934
rect 1485 4931 1551 4934
rect 2773 4994 2839 4997
rect 5073 4994 5139 4997
rect 7414 4994 7420 4996
rect 2773 4992 7420 4994
rect 2773 4936 2778 4992
rect 2834 4936 5078 4992
rect 5134 4936 7420 4992
rect 2773 4934 7420 4936
rect 2773 4931 2839 4934
rect 5073 4931 5139 4934
rect 7414 4932 7420 4934
rect 7484 4932 7490 4996
rect 8334 4932 8340 4996
rect 8404 4994 8410 4996
rect 9765 4994 9831 4997
rect 9949 4994 10015 4997
rect 8404 4992 10015 4994
rect 8404 4936 9770 4992
rect 9826 4936 9954 4992
rect 10010 4936 10015 4992
rect 8404 4934 10015 4936
rect 8404 4932 8410 4934
rect 9765 4931 9831 4934
rect 9949 4931 10015 4934
rect 10409 4994 10475 4997
rect 11094 4994 11100 4996
rect 10409 4992 11100 4994
rect 10409 4936 10414 4992
rect 10470 4936 11100 4992
rect 10409 4934 11100 4936
rect 10409 4931 10475 4934
rect 11094 4932 11100 4934
rect 11164 4932 11170 4996
rect 11881 4994 11947 4997
rect 13118 4994 13124 4996
rect 11881 4992 13124 4994
rect 11881 4936 11886 4992
rect 11942 4936 13124 4992
rect 11881 4934 13124 4936
rect 11881 4931 11947 4934
rect 13118 4932 13124 4934
rect 13188 4932 13194 4996
rect 15101 4994 15167 4997
rect 16614 4994 16620 4996
rect 15101 4992 16620 4994
rect 15101 4936 15106 4992
rect 15162 4936 16620 4992
rect 15101 4934 16620 4936
rect 15101 4931 15167 4934
rect 16614 4932 16620 4934
rect 16684 4932 16690 4996
rect 20348 4994 20408 5070
rect 21449 4994 21515 4997
rect 23289 4994 23355 4997
rect 20348 4992 23355 4994
rect 20348 4936 21454 4992
rect 21510 4936 23294 4992
rect 23350 4936 23355 4992
rect 20348 4934 23355 4936
rect 23430 4994 23490 5070
rect 24209 5128 27354 5130
rect 24209 5072 24214 5128
rect 24270 5072 27354 5128
rect 24209 5070 27354 5072
rect 24209 5067 24275 5070
rect 25313 4994 25379 4997
rect 23430 4992 25379 4994
rect 23430 4936 25318 4992
rect 25374 4936 25379 4992
rect 23430 4934 25379 4936
rect 27294 4994 27354 5070
rect 27521 5128 32371 5130
rect 27521 5072 27526 5128
rect 27582 5072 32310 5128
rect 32366 5072 32371 5128
rect 27521 5070 32371 5072
rect 27521 5067 27587 5070
rect 32305 5067 32371 5070
rect 32581 5130 32647 5133
rect 34605 5130 34671 5133
rect 32581 5128 34671 5130
rect 32581 5072 32586 5128
rect 32642 5072 34610 5128
rect 34666 5072 34671 5128
rect 32581 5070 34671 5072
rect 32581 5067 32647 5070
rect 34605 5067 34671 5070
rect 28073 4994 28139 4997
rect 30741 4994 30807 4997
rect 31385 4994 31451 4997
rect 27294 4992 28139 4994
rect 27294 4936 28078 4992
rect 28134 4936 28139 4992
rect 27294 4934 28139 4936
rect 21449 4931 21515 4934
rect 23289 4931 23355 4934
rect 25313 4931 25379 4934
rect 28073 4931 28139 4934
rect 29824 4992 31451 4994
rect 29824 4936 30746 4992
rect 30802 4936 31390 4992
rect 31446 4936 31451 4992
rect 29824 4934 31451 4936
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 13946 4928 14262 4929
rect 13946 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14262 4928
rect 13946 4863 14262 4864
rect 19946 4928 20262 4929
rect 19946 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20262 4928
rect 19946 4863 20262 4864
rect 25946 4928 26262 4929
rect 25946 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26262 4928
rect 25946 4863 26262 4864
rect 29824 4861 29884 4934
rect 30741 4931 30807 4934
rect 31385 4931 31451 4934
rect 33041 4994 33107 4997
rect 35801 4994 35867 4997
rect 33041 4992 35867 4994
rect 33041 4936 33046 4992
rect 33102 4936 35806 4992
rect 35862 4936 35867 4992
rect 33041 4934 35867 4936
rect 33041 4931 33107 4934
rect 35801 4931 35867 4934
rect 39021 4994 39087 4997
rect 40880 4994 41000 5024
rect 39021 4992 41000 4994
rect 39021 4936 39026 4992
rect 39082 4936 41000 4992
rect 39021 4934 41000 4936
rect 39021 4931 39087 4934
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 37946 4928 38262 4929
rect 37946 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38262 4928
rect 40880 4904 41000 4934
rect 37946 4863 38262 4864
rect 4245 4858 4311 4861
rect 5625 4858 5691 4861
rect 4245 4856 5691 4858
rect 4245 4800 4250 4856
rect 4306 4800 5630 4856
rect 5686 4800 5691 4856
rect 4245 4798 5691 4800
rect 4245 4795 4311 4798
rect 5625 4795 5691 4798
rect 5993 4858 6059 4861
rect 7649 4858 7715 4861
rect 11237 4858 11303 4861
rect 5993 4856 7715 4858
rect 5993 4800 5998 4856
rect 6054 4800 7654 4856
rect 7710 4800 7715 4856
rect 5993 4798 7715 4800
rect 5993 4795 6059 4798
rect 7649 4795 7715 4798
rect 8342 4856 11303 4858
rect 8342 4800 11242 4856
rect 11298 4800 11303 4856
rect 8342 4798 11303 4800
rect 0 4722 120 4752
rect 2405 4722 2471 4725
rect 2630 4722 2636 4724
rect 0 4662 1042 4722
rect 0 4632 120 4662
rect 982 4586 1042 4662
rect 2405 4720 2636 4722
rect 2405 4664 2410 4720
rect 2466 4664 2636 4720
rect 2405 4662 2636 4664
rect 2405 4659 2471 4662
rect 2630 4660 2636 4662
rect 2700 4660 2706 4724
rect 2957 4722 3023 4725
rect 4337 4722 4403 4725
rect 4521 4722 4587 4725
rect 8342 4722 8402 4798
rect 11237 4795 11303 4798
rect 12065 4858 12131 4861
rect 12249 4858 12315 4861
rect 12065 4856 12315 4858
rect 12065 4800 12070 4856
rect 12126 4800 12254 4856
rect 12310 4800 12315 4856
rect 12065 4798 12315 4800
rect 12065 4795 12131 4798
rect 12249 4795 12315 4798
rect 12433 4858 12499 4861
rect 13670 4858 13676 4860
rect 12433 4856 13676 4858
rect 12433 4800 12438 4856
rect 12494 4800 13676 4856
rect 12433 4798 13676 4800
rect 12433 4795 12499 4798
rect 13670 4796 13676 4798
rect 13740 4796 13746 4860
rect 14406 4796 14412 4860
rect 14476 4858 14482 4860
rect 16389 4858 16455 4861
rect 19609 4858 19675 4861
rect 14476 4856 19675 4858
rect 14476 4800 16394 4856
rect 16450 4800 19614 4856
rect 19670 4800 19675 4856
rect 14476 4798 19675 4800
rect 14476 4796 14482 4798
rect 16389 4795 16455 4798
rect 19609 4795 19675 4798
rect 21081 4858 21147 4861
rect 21357 4858 21423 4861
rect 24945 4858 25011 4861
rect 21081 4856 25011 4858
rect 21081 4800 21086 4856
rect 21142 4800 21362 4856
rect 21418 4800 24950 4856
rect 25006 4800 25011 4856
rect 21081 4798 25011 4800
rect 21081 4795 21147 4798
rect 21357 4795 21423 4798
rect 24945 4795 25011 4798
rect 26509 4858 26575 4861
rect 29821 4858 29887 4861
rect 26509 4856 29887 4858
rect 26509 4800 26514 4856
rect 26570 4800 29826 4856
rect 29882 4800 29887 4856
rect 26509 4798 29887 4800
rect 26509 4795 26575 4798
rect 29821 4795 29887 4798
rect 30189 4858 30255 4861
rect 32581 4858 32647 4861
rect 35893 4858 35959 4861
rect 30189 4856 31770 4858
rect 30189 4800 30194 4856
rect 30250 4800 31770 4856
rect 30189 4798 31770 4800
rect 30189 4795 30255 4798
rect 2957 4720 8402 4722
rect 2957 4664 2962 4720
rect 3018 4664 4342 4720
rect 4398 4664 4526 4720
rect 4582 4664 8402 4720
rect 2957 4662 8402 4664
rect 2957 4659 3023 4662
rect 4337 4659 4403 4662
rect 4521 4659 4587 4662
rect 8518 4660 8524 4724
rect 8588 4722 8594 4724
rect 31385 4722 31451 4725
rect 8588 4720 31451 4722
rect 8588 4664 31390 4720
rect 31446 4664 31451 4720
rect 8588 4662 31451 4664
rect 31710 4722 31770 4798
rect 32581 4856 35959 4858
rect 32581 4800 32586 4856
rect 32642 4800 35898 4856
rect 35954 4800 35959 4856
rect 32581 4798 35959 4800
rect 32581 4795 32647 4798
rect 35893 4795 35959 4798
rect 39205 4722 39271 4725
rect 31710 4720 39271 4722
rect 31710 4664 39210 4720
rect 39266 4664 39271 4720
rect 31710 4662 39271 4664
rect 8588 4660 8594 4662
rect 31385 4659 31451 4662
rect 39205 4659 39271 4662
rect 39481 4722 39547 4725
rect 40880 4722 41000 4752
rect 39481 4720 41000 4722
rect 39481 4664 39486 4720
rect 39542 4664 41000 4720
rect 39481 4662 41000 4664
rect 39481 4659 39547 4662
rect 40880 4632 41000 4662
rect 1853 4586 1919 4589
rect 982 4584 1919 4586
rect 982 4528 1858 4584
rect 1914 4528 1919 4584
rect 982 4526 1919 4528
rect 1853 4523 1919 4526
rect 3233 4586 3299 4589
rect 10133 4586 10199 4589
rect 13353 4586 13419 4589
rect 15101 4586 15167 4589
rect 15469 4586 15535 4589
rect 3233 4584 10199 4586
rect 3233 4528 3238 4584
rect 3294 4528 10138 4584
rect 10194 4528 10199 4584
rect 3233 4526 10199 4528
rect 3233 4523 3299 4526
rect 10133 4523 10199 4526
rect 10412 4584 13419 4586
rect 10412 4528 13358 4584
rect 13414 4528 13419 4584
rect 10412 4526 13419 4528
rect 0 4450 120 4480
rect 1485 4450 1551 4453
rect 0 4448 1551 4450
rect 0 4392 1490 4448
rect 1546 4392 1551 4448
rect 0 4390 1551 4392
rect 0 4360 120 4390
rect 1485 4387 1551 4390
rect 5257 4450 5323 4453
rect 5257 4448 8034 4450
rect 5257 4392 5262 4448
rect 5318 4392 8034 4448
rect 5257 4390 8034 4392
rect 5257 4387 5323 4390
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 5165 4314 5231 4317
rect 7741 4314 7807 4317
rect 5165 4312 7807 4314
rect 5165 4256 5170 4312
rect 5226 4256 7746 4312
rect 7802 4256 7807 4312
rect 5165 4254 7807 4256
rect 5165 4251 5231 4254
rect 7741 4251 7807 4254
rect 0 4178 120 4208
rect 1853 4178 1919 4181
rect 0 4176 1919 4178
rect 0 4120 1858 4176
rect 1914 4120 1919 4176
rect 0 4118 1919 4120
rect 0 4088 120 4118
rect 1853 4115 1919 4118
rect 3601 4178 3667 4181
rect 4102 4178 4108 4180
rect 3601 4176 4108 4178
rect 3601 4120 3606 4176
rect 3662 4120 4108 4176
rect 3601 4118 4108 4120
rect 3601 4115 3667 4118
rect 4102 4116 4108 4118
rect 4172 4116 4178 4180
rect 6494 4116 6500 4180
rect 6564 4178 6570 4180
rect 6729 4178 6795 4181
rect 6564 4176 6795 4178
rect 6564 4120 6734 4176
rect 6790 4120 6795 4176
rect 6564 4118 6795 4120
rect 7974 4178 8034 4390
rect 9438 4388 9444 4452
rect 9508 4450 9514 4452
rect 9581 4450 9647 4453
rect 9508 4448 9690 4450
rect 9508 4392 9586 4448
rect 9642 4392 9690 4448
rect 9508 4390 9690 4392
rect 9508 4388 9514 4390
rect 9581 4387 9690 4390
rect 9006 4384 9322 4385
rect 9006 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9322 4384
rect 9006 4319 9322 4320
rect 9630 4314 9690 4387
rect 10041 4314 10107 4317
rect 9630 4312 10107 4314
rect 9630 4256 10046 4312
rect 10102 4256 10107 4312
rect 9630 4254 10107 4256
rect 10041 4251 10107 4254
rect 10412 4178 10472 4526
rect 13353 4523 13419 4526
rect 14782 4584 15535 4586
rect 14782 4528 15106 4584
rect 15162 4528 15474 4584
rect 15530 4528 15535 4584
rect 14782 4526 15535 4528
rect 10542 4388 10548 4452
rect 10612 4450 10618 4452
rect 14782 4450 14842 4526
rect 15101 4523 15167 4526
rect 15469 4523 15535 4526
rect 16021 4586 16087 4589
rect 17217 4586 17283 4589
rect 18413 4586 18479 4589
rect 16021 4584 18479 4586
rect 16021 4528 16026 4584
rect 16082 4528 17222 4584
rect 17278 4528 18418 4584
rect 18474 4528 18479 4584
rect 16021 4526 18479 4528
rect 16021 4523 16087 4526
rect 17217 4523 17283 4526
rect 18413 4523 18479 4526
rect 18822 4524 18828 4588
rect 18892 4586 18898 4588
rect 34697 4586 34763 4589
rect 18892 4584 34763 4586
rect 18892 4528 34702 4584
rect 34758 4528 34763 4584
rect 18892 4526 34763 4528
rect 18892 4524 18898 4526
rect 34697 4523 34763 4526
rect 10612 4390 14842 4450
rect 17401 4450 17467 4453
rect 17677 4450 17743 4453
rect 17401 4448 17743 4450
rect 17401 4392 17406 4448
rect 17462 4392 17682 4448
rect 17738 4392 17743 4448
rect 17401 4390 17743 4392
rect 10612 4388 10618 4390
rect 17401 4387 17467 4390
rect 17677 4387 17743 4390
rect 17953 4450 18019 4453
rect 20805 4450 20871 4453
rect 17953 4448 20871 4450
rect 17953 4392 17958 4448
rect 18014 4392 20810 4448
rect 20866 4392 20871 4448
rect 17953 4390 20871 4392
rect 17953 4387 18019 4390
rect 20805 4387 20871 4390
rect 22093 4450 22159 4453
rect 26601 4450 26667 4453
rect 22093 4448 26667 4450
rect 22093 4392 22098 4448
rect 22154 4392 26606 4448
rect 26662 4392 26667 4448
rect 22093 4390 26667 4392
rect 22093 4387 22159 4390
rect 26601 4387 26667 4390
rect 27429 4450 27495 4453
rect 29453 4450 29519 4453
rect 27429 4448 29519 4450
rect 27429 4392 27434 4448
rect 27490 4392 29458 4448
rect 29514 4392 29519 4448
rect 27429 4390 29519 4392
rect 27429 4387 27495 4390
rect 29453 4387 29519 4390
rect 29637 4450 29703 4453
rect 31937 4450 32003 4453
rect 29637 4448 32003 4450
rect 29637 4392 29642 4448
rect 29698 4392 31942 4448
rect 31998 4392 32003 4448
rect 29637 4390 32003 4392
rect 29637 4387 29703 4390
rect 31937 4387 32003 4390
rect 39389 4450 39455 4453
rect 40880 4450 41000 4480
rect 39389 4448 41000 4450
rect 39389 4392 39394 4448
rect 39450 4392 41000 4448
rect 39389 4390 41000 4392
rect 39389 4387 39455 4390
rect 15006 4384 15322 4385
rect 15006 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15322 4384
rect 15006 4319 15322 4320
rect 21006 4384 21322 4385
rect 21006 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21322 4384
rect 21006 4319 21322 4320
rect 27006 4384 27322 4385
rect 27006 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27322 4384
rect 27006 4319 27322 4320
rect 33006 4384 33322 4385
rect 33006 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33322 4384
rect 33006 4319 33322 4320
rect 39006 4384 39322 4385
rect 39006 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39322 4384
rect 40880 4360 41000 4390
rect 39006 4319 39322 4320
rect 11513 4314 11579 4317
rect 18781 4314 18847 4317
rect 11513 4312 14842 4314
rect 11513 4256 11518 4312
rect 11574 4256 14842 4312
rect 11513 4254 14842 4256
rect 11513 4251 11579 4254
rect 7974 4118 10472 4178
rect 10869 4178 10935 4181
rect 12249 4178 12315 4181
rect 10869 4176 12315 4178
rect 10869 4120 10874 4176
rect 10930 4120 12254 4176
rect 12310 4120 12315 4176
rect 10869 4118 12315 4120
rect 14782 4178 14842 4254
rect 15518 4312 18847 4314
rect 15518 4256 18786 4312
rect 18842 4256 18847 4312
rect 15518 4254 18847 4256
rect 15518 4178 15578 4254
rect 18781 4251 18847 4254
rect 19190 4252 19196 4316
rect 19260 4314 19266 4316
rect 20805 4314 20871 4317
rect 19260 4312 20871 4314
rect 19260 4256 20810 4312
rect 20866 4256 20871 4312
rect 19260 4254 20871 4256
rect 19260 4252 19266 4254
rect 20805 4251 20871 4254
rect 22277 4314 22343 4317
rect 23013 4314 23079 4317
rect 22277 4312 23079 4314
rect 22277 4256 22282 4312
rect 22338 4256 23018 4312
rect 23074 4256 23079 4312
rect 22277 4254 23079 4256
rect 22277 4251 22343 4254
rect 23013 4251 23079 4254
rect 23933 4314 23999 4317
rect 25589 4314 25655 4317
rect 23933 4312 25655 4314
rect 23933 4256 23938 4312
rect 23994 4256 25594 4312
rect 25650 4256 25655 4312
rect 23933 4254 25655 4256
rect 23933 4251 23999 4254
rect 25589 4251 25655 4254
rect 27470 4252 27476 4316
rect 27540 4314 27546 4316
rect 27613 4314 27679 4317
rect 27540 4312 27679 4314
rect 27540 4256 27618 4312
rect 27674 4256 27679 4312
rect 27540 4254 27679 4256
rect 27540 4252 27546 4254
rect 27613 4251 27679 4254
rect 29913 4314 29979 4317
rect 32397 4314 32463 4317
rect 29913 4312 32463 4314
rect 29913 4256 29918 4312
rect 29974 4256 32402 4312
rect 32458 4256 32463 4312
rect 29913 4254 32463 4256
rect 29913 4251 29979 4254
rect 32397 4251 32463 4254
rect 14782 4118 15578 4178
rect 16849 4178 16915 4181
rect 17902 4178 17908 4180
rect 16849 4176 17908 4178
rect 16849 4120 16854 4176
rect 16910 4120 17908 4176
rect 16849 4118 17908 4120
rect 6564 4116 6570 4118
rect 6729 4115 6795 4118
rect 10869 4115 10935 4118
rect 12249 4115 12315 4118
rect 16849 4115 16915 4118
rect 17902 4116 17908 4118
rect 17972 4116 17978 4180
rect 18689 4178 18755 4181
rect 27153 4178 27219 4181
rect 18689 4176 27219 4178
rect 18689 4120 18694 4176
rect 18750 4120 27158 4176
rect 27214 4120 27219 4176
rect 18689 4118 27219 4120
rect 18689 4115 18755 4118
rect 27153 4115 27219 4118
rect 31201 4178 31267 4181
rect 36169 4178 36235 4181
rect 31201 4176 36235 4178
rect 31201 4120 31206 4176
rect 31262 4120 36174 4176
rect 36230 4120 36235 4176
rect 31201 4118 36235 4120
rect 31201 4115 31267 4118
rect 36169 4115 36235 4118
rect 39389 4178 39455 4181
rect 40880 4178 41000 4208
rect 39389 4176 41000 4178
rect 39389 4120 39394 4176
rect 39450 4120 41000 4176
rect 39389 4118 41000 4120
rect 39389 4115 39455 4118
rect 40880 4088 41000 4118
rect 2221 4042 2287 4045
rect 4153 4042 4219 4045
rect 6177 4042 6243 4045
rect 2221 4040 2468 4042
rect 2221 3984 2226 4040
rect 2282 3984 2468 4040
rect 2221 3982 2468 3984
rect 2221 3979 2287 3982
rect 0 3906 120 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 120 3846
rect 1485 3843 1551 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 0 3634 120 3664
rect 2129 3634 2195 3637
rect 0 3632 2195 3634
rect 0 3576 2134 3632
rect 2190 3576 2195 3632
rect 0 3574 2195 3576
rect 0 3544 120 3574
rect 2129 3571 2195 3574
rect 1669 3498 1735 3501
rect 2408 3498 2468 3982
rect 4153 4040 6243 4042
rect 4153 3984 4158 4040
rect 4214 3984 6182 4040
rect 6238 3984 6243 4040
rect 4153 3982 6243 3984
rect 4153 3979 4219 3982
rect 6177 3979 6243 3982
rect 7373 4040 7439 4045
rect 7373 3984 7378 4040
rect 7434 3984 7439 4040
rect 7373 3979 7439 3984
rect 7649 4042 7715 4045
rect 12157 4042 12223 4045
rect 14089 4042 14155 4045
rect 7649 4040 9690 4042
rect 7649 3984 7654 4040
rect 7710 3984 9690 4040
rect 7649 3982 9690 3984
rect 7649 3979 7715 3982
rect 3141 3906 3207 3909
rect 7376 3906 7436 3979
rect 3141 3904 7436 3906
rect 3141 3848 3146 3904
rect 3202 3848 7436 3904
rect 3141 3846 7436 3848
rect 3141 3843 3207 3846
rect 8702 3844 8708 3908
rect 8772 3906 8778 3908
rect 8845 3906 8911 3909
rect 8772 3904 8911 3906
rect 8772 3848 8850 3904
rect 8906 3848 8911 3904
rect 8772 3846 8911 3848
rect 8772 3844 8778 3846
rect 8845 3843 8911 3846
rect 9121 3906 9187 3909
rect 9438 3906 9444 3908
rect 9121 3904 9444 3906
rect 9121 3848 9126 3904
rect 9182 3848 9444 3904
rect 9121 3846 9444 3848
rect 9121 3843 9187 3846
rect 9438 3844 9444 3846
rect 9508 3844 9514 3908
rect 9630 3906 9690 3982
rect 12157 4040 14428 4042
rect 12157 3984 12162 4040
rect 12218 3984 14094 4040
rect 14150 3984 14428 4040
rect 12157 3982 14428 3984
rect 12157 3979 12223 3982
rect 14089 3979 14155 3982
rect 13169 3906 13235 3909
rect 9630 3904 13235 3906
rect 9630 3848 13174 3904
rect 13230 3848 13235 3904
rect 9630 3846 13235 3848
rect 14368 3906 14428 3982
rect 14590 3980 14596 4044
rect 14660 4042 14666 4044
rect 15193 4042 15259 4045
rect 16849 4042 16915 4045
rect 14660 4040 16915 4042
rect 14660 3984 15198 4040
rect 15254 3984 16854 4040
rect 16910 3984 16915 4040
rect 14660 3982 16915 3984
rect 14660 3980 14666 3982
rect 15193 3979 15259 3982
rect 16849 3979 16915 3982
rect 17585 4042 17651 4045
rect 18045 4042 18111 4045
rect 17585 4040 18111 4042
rect 17585 3984 17590 4040
rect 17646 3984 18050 4040
rect 18106 3984 18111 4040
rect 17585 3982 18111 3984
rect 17585 3979 17651 3982
rect 18045 3979 18111 3982
rect 18321 4042 18387 4045
rect 26509 4042 26575 4045
rect 18321 4040 26575 4042
rect 18321 3984 18326 4040
rect 18382 3984 26514 4040
rect 26570 3984 26575 4040
rect 18321 3982 26575 3984
rect 18321 3979 18387 3982
rect 26509 3979 26575 3982
rect 27889 4042 27955 4045
rect 29453 4042 29519 4045
rect 27889 4040 29519 4042
rect 27889 3984 27894 4040
rect 27950 3984 29458 4040
rect 29514 3984 29519 4040
rect 27889 3982 29519 3984
rect 27889 3979 27955 3982
rect 29453 3979 29519 3982
rect 30414 3980 30420 4044
rect 30484 4042 30490 4044
rect 31385 4042 31451 4045
rect 30484 4040 31451 4042
rect 30484 3984 31390 4040
rect 31446 3984 31451 4040
rect 30484 3982 31451 3984
rect 30484 3980 30490 3982
rect 31385 3979 31451 3982
rect 31937 4042 32003 4045
rect 34421 4042 34487 4045
rect 31937 4040 34487 4042
rect 31937 3984 31942 4040
rect 31998 3984 34426 4040
rect 34482 3984 34487 4040
rect 31937 3982 34487 3984
rect 31937 3979 32003 3982
rect 34421 3979 34487 3982
rect 19425 3906 19491 3909
rect 14368 3904 19491 3906
rect 14368 3848 19430 3904
rect 19486 3848 19491 3904
rect 14368 3846 19491 3848
rect 13169 3843 13235 3846
rect 19425 3843 19491 3846
rect 20345 3906 20411 3909
rect 25589 3906 25655 3909
rect 20345 3904 25655 3906
rect 20345 3848 20350 3904
rect 20406 3848 25594 3904
rect 25650 3848 25655 3904
rect 20345 3846 25655 3848
rect 20345 3843 20411 3846
rect 25589 3843 25655 3846
rect 26785 3906 26851 3909
rect 31017 3906 31083 3909
rect 26785 3904 31083 3906
rect 26785 3848 26790 3904
rect 26846 3848 31022 3904
rect 31078 3848 31083 3904
rect 26785 3846 31083 3848
rect 26785 3843 26851 3846
rect 31017 3843 31083 3846
rect 39021 3906 39087 3909
rect 40880 3906 41000 3936
rect 39021 3904 41000 3906
rect 39021 3848 39026 3904
rect 39082 3848 41000 3904
rect 39021 3846 41000 3848
rect 39021 3843 39087 3846
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 13946 3840 14262 3841
rect 13946 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14262 3840
rect 13946 3775 14262 3776
rect 19946 3840 20262 3841
rect 19946 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20262 3840
rect 19946 3775 20262 3776
rect 25946 3840 26262 3841
rect 25946 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26262 3840
rect 25946 3775 26262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 37946 3840 38262 3841
rect 37946 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38262 3840
rect 40880 3816 41000 3846
rect 37946 3775 38262 3776
rect 5533 3770 5599 3773
rect 7373 3770 7439 3773
rect 5533 3768 7439 3770
rect 5533 3712 5538 3768
rect 5594 3712 7378 3768
rect 7434 3712 7439 3768
rect 5533 3710 7439 3712
rect 5533 3707 5599 3710
rect 7373 3707 7439 3710
rect 8334 3708 8340 3772
rect 8404 3770 8410 3772
rect 13353 3770 13419 3773
rect 13537 3772 13603 3773
rect 14825 3772 14891 3773
rect 8404 3768 13419 3770
rect 8404 3712 13358 3768
rect 13414 3712 13419 3768
rect 8404 3710 13419 3712
rect 8404 3708 8410 3710
rect 13353 3707 13419 3710
rect 13486 3708 13492 3772
rect 13556 3770 13603 3772
rect 13556 3768 13648 3770
rect 13598 3712 13648 3768
rect 13556 3710 13648 3712
rect 13556 3708 13603 3710
rect 14774 3708 14780 3772
rect 14844 3770 14891 3772
rect 15285 3770 15351 3773
rect 15837 3770 15903 3773
rect 14844 3768 14936 3770
rect 14886 3712 14936 3768
rect 14844 3710 14936 3712
rect 15285 3768 15903 3770
rect 15285 3712 15290 3768
rect 15346 3712 15842 3768
rect 15898 3712 15903 3768
rect 15285 3710 15903 3712
rect 14844 3708 14891 3710
rect 13537 3707 13603 3708
rect 14825 3707 14891 3708
rect 15285 3707 15351 3710
rect 15837 3707 15903 3710
rect 16481 3770 16547 3773
rect 18505 3770 18571 3773
rect 16481 3768 18571 3770
rect 16481 3712 16486 3768
rect 16542 3712 18510 3768
rect 18566 3712 18571 3768
rect 16481 3710 18571 3712
rect 16481 3707 16547 3710
rect 18505 3707 18571 3710
rect 18781 3770 18847 3773
rect 20437 3770 20503 3773
rect 22093 3770 22159 3773
rect 24669 3770 24735 3773
rect 25497 3770 25563 3773
rect 27889 3770 27955 3773
rect 18781 3768 19626 3770
rect 18781 3712 18786 3768
rect 18842 3712 19626 3768
rect 18781 3710 19626 3712
rect 18781 3707 18847 3710
rect 2865 3634 2931 3637
rect 5349 3634 5415 3637
rect 2865 3632 5415 3634
rect 2865 3576 2870 3632
rect 2926 3576 5354 3632
rect 5410 3576 5415 3632
rect 2865 3574 5415 3576
rect 2865 3571 2931 3574
rect 5349 3571 5415 3574
rect 6637 3634 6703 3637
rect 9397 3634 9463 3637
rect 6637 3632 9463 3634
rect 6637 3576 6642 3632
rect 6698 3576 9402 3632
rect 9458 3576 9463 3632
rect 6637 3574 9463 3576
rect 6637 3571 6703 3574
rect 9397 3571 9463 3574
rect 10593 3634 10659 3637
rect 13169 3634 13235 3637
rect 17861 3634 17927 3637
rect 19333 3634 19399 3637
rect 10593 3632 12634 3634
rect 10593 3576 10598 3632
rect 10654 3576 12634 3632
rect 10593 3574 12634 3576
rect 10593 3571 10659 3574
rect 2957 3498 3023 3501
rect 1669 3496 2468 3498
rect 1669 3440 1674 3496
rect 1730 3440 2468 3496
rect 1669 3438 2468 3440
rect 2822 3496 3023 3498
rect 2822 3440 2962 3496
rect 3018 3440 3023 3496
rect 2822 3438 3023 3440
rect 1669 3435 1735 3438
rect 0 3362 120 3392
rect 1485 3362 1551 3365
rect 0 3360 1551 3362
rect 0 3304 1490 3360
rect 1546 3304 1551 3360
rect 0 3302 1551 3304
rect 0 3272 120 3302
rect 1485 3299 1551 3302
rect 0 3090 120 3120
rect 2221 3090 2287 3093
rect 0 3088 2287 3090
rect 0 3032 2226 3088
rect 2282 3032 2287 3088
rect 0 3030 2287 3032
rect 2822 3090 2882 3438
rect 2957 3435 3023 3438
rect 3233 3498 3299 3501
rect 3969 3498 4035 3501
rect 5901 3498 5967 3501
rect 3233 3496 3802 3498
rect 3233 3440 3238 3496
rect 3294 3440 3802 3496
rect 3233 3438 3802 3440
rect 3233 3435 3299 3438
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 3742 3226 3802 3438
rect 3969 3496 5967 3498
rect 3969 3440 3974 3496
rect 4030 3440 5906 3496
rect 5962 3440 5967 3496
rect 3969 3438 5967 3440
rect 3969 3435 4035 3438
rect 5901 3435 5967 3438
rect 7097 3498 7163 3501
rect 10041 3498 10107 3501
rect 7097 3496 10107 3498
rect 7097 3440 7102 3496
rect 7158 3440 10046 3496
rect 10102 3440 10107 3496
rect 7097 3438 10107 3440
rect 7097 3435 7163 3438
rect 10041 3435 10107 3438
rect 11329 3498 11395 3501
rect 11830 3498 11836 3500
rect 11329 3496 11836 3498
rect 11329 3440 11334 3496
rect 11390 3440 11836 3496
rect 11329 3438 11836 3440
rect 11329 3435 11395 3438
rect 11830 3436 11836 3438
rect 11900 3436 11906 3500
rect 7598 3300 7604 3364
rect 7668 3362 7674 3364
rect 8017 3362 8083 3365
rect 7668 3360 8083 3362
rect 7668 3304 8022 3360
rect 8078 3304 8083 3360
rect 7668 3302 8083 3304
rect 7668 3300 7674 3302
rect 8017 3299 8083 3302
rect 8293 3362 8359 3365
rect 9765 3362 9831 3365
rect 11421 3362 11487 3365
rect 8293 3360 8770 3362
rect 8293 3304 8298 3360
rect 8354 3304 8770 3360
rect 8293 3302 8770 3304
rect 8293 3299 8359 3302
rect 8710 3229 8770 3302
rect 9765 3360 11487 3362
rect 9765 3304 9770 3360
rect 9826 3304 11426 3360
rect 11482 3304 11487 3360
rect 9765 3302 11487 3304
rect 12574 3362 12634 3574
rect 13169 3632 19399 3634
rect 13169 3576 13174 3632
rect 13230 3576 17866 3632
rect 17922 3576 19338 3632
rect 19394 3576 19399 3632
rect 13169 3574 19399 3576
rect 19566 3634 19626 3710
rect 20437 3768 25563 3770
rect 20437 3712 20442 3768
rect 20498 3712 22098 3768
rect 22154 3712 24674 3768
rect 24730 3712 25502 3768
rect 25558 3712 25563 3768
rect 20437 3710 25563 3712
rect 20437 3707 20503 3710
rect 22093 3707 22159 3710
rect 24669 3707 24735 3710
rect 25497 3707 25563 3710
rect 27524 3768 27955 3770
rect 27524 3712 27894 3768
rect 27950 3712 27955 3768
rect 27524 3710 27955 3712
rect 20437 3634 20503 3637
rect 23013 3634 23079 3637
rect 19566 3574 20362 3634
rect 13169 3571 13235 3574
rect 17861 3571 17927 3574
rect 19333 3571 19399 3574
rect 12709 3498 12775 3501
rect 19609 3498 19675 3501
rect 19793 3498 19859 3501
rect 20161 3498 20227 3501
rect 12709 3496 20227 3498
rect 12709 3440 12714 3496
rect 12770 3440 19614 3496
rect 19670 3440 19798 3496
rect 19854 3440 20166 3496
rect 20222 3440 20227 3496
rect 12709 3438 20227 3440
rect 20302 3498 20362 3574
rect 20437 3632 23079 3634
rect 20437 3576 20442 3632
rect 20498 3576 23018 3632
rect 23074 3576 23079 3632
rect 20437 3574 23079 3576
rect 20437 3571 20503 3574
rect 23013 3571 23079 3574
rect 23841 3634 23907 3637
rect 25221 3634 25287 3637
rect 27524 3634 27584 3710
rect 27889 3707 27955 3710
rect 23841 3632 27584 3634
rect 23841 3576 23846 3632
rect 23902 3576 25226 3632
rect 25282 3576 27584 3632
rect 23841 3574 27584 3576
rect 23841 3571 23907 3574
rect 25221 3571 25287 3574
rect 27654 3572 27660 3636
rect 27724 3634 27730 3636
rect 34789 3634 34855 3637
rect 27724 3632 34855 3634
rect 27724 3576 34794 3632
rect 34850 3576 34855 3632
rect 27724 3574 34855 3576
rect 27724 3572 27730 3574
rect 34789 3571 34855 3574
rect 39389 3634 39455 3637
rect 40880 3634 41000 3664
rect 39389 3632 41000 3634
rect 39389 3576 39394 3632
rect 39450 3576 41000 3632
rect 39389 3574 41000 3576
rect 39389 3571 39455 3574
rect 40880 3544 41000 3574
rect 25957 3498 26023 3501
rect 20302 3496 26023 3498
rect 20302 3440 25962 3496
rect 26018 3440 26023 3496
rect 20302 3438 26023 3440
rect 12709 3435 12775 3438
rect 19609 3435 19675 3438
rect 19793 3435 19859 3438
rect 20161 3435 20227 3438
rect 25957 3435 26023 3438
rect 26417 3498 26483 3501
rect 33317 3498 33383 3501
rect 26417 3496 33383 3498
rect 26417 3440 26422 3496
rect 26478 3440 33322 3496
rect 33378 3440 33383 3496
rect 26417 3438 33383 3440
rect 26417 3435 26483 3438
rect 33317 3435 33383 3438
rect 14641 3362 14707 3365
rect 12574 3360 14707 3362
rect 12574 3304 14646 3360
rect 14702 3304 14707 3360
rect 12574 3302 14707 3304
rect 9765 3299 9831 3302
rect 11421 3299 11487 3302
rect 14641 3299 14707 3302
rect 15653 3362 15719 3365
rect 20345 3362 20411 3365
rect 15653 3360 20411 3362
rect 15653 3304 15658 3360
rect 15714 3304 20350 3360
rect 20406 3304 20411 3360
rect 15653 3302 20411 3304
rect 15653 3299 15719 3302
rect 20345 3299 20411 3302
rect 24853 3362 24919 3365
rect 26785 3362 26851 3365
rect 24853 3360 26851 3362
rect 24853 3304 24858 3360
rect 24914 3304 26790 3360
rect 26846 3304 26851 3360
rect 24853 3302 26851 3304
rect 24853 3299 24919 3302
rect 26785 3299 26851 3302
rect 27521 3362 27587 3365
rect 29729 3362 29795 3365
rect 27521 3360 29795 3362
rect 27521 3304 27526 3360
rect 27582 3304 29734 3360
rect 29790 3304 29795 3360
rect 27521 3302 29795 3304
rect 27521 3299 27587 3302
rect 29729 3299 29795 3302
rect 30005 3362 30071 3365
rect 31937 3362 32003 3365
rect 32581 3362 32647 3365
rect 30005 3360 32647 3362
rect 30005 3304 30010 3360
rect 30066 3304 31942 3360
rect 31998 3304 32586 3360
rect 32642 3304 32647 3360
rect 30005 3302 32647 3304
rect 30005 3299 30071 3302
rect 31937 3299 32003 3302
rect 32581 3299 32647 3302
rect 39941 3362 40007 3365
rect 40880 3362 41000 3392
rect 39941 3360 41000 3362
rect 39941 3304 39946 3360
rect 40002 3304 41000 3360
rect 39941 3302 41000 3304
rect 39941 3299 40007 3302
rect 9006 3296 9322 3297
rect 9006 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9322 3296
rect 9006 3231 9322 3232
rect 15006 3296 15322 3297
rect 15006 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15322 3296
rect 15006 3231 15322 3232
rect 21006 3296 21322 3297
rect 21006 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21322 3296
rect 21006 3231 21322 3232
rect 27006 3296 27322 3297
rect 27006 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27322 3296
rect 27006 3231 27322 3232
rect 33006 3296 33322 3297
rect 33006 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33322 3296
rect 33006 3231 33322 3232
rect 39006 3296 39322 3297
rect 39006 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39322 3296
rect 40880 3272 41000 3302
rect 39006 3231 39322 3232
rect 8569 3226 8635 3229
rect 3742 3224 8635 3226
rect 3742 3168 8574 3224
rect 8630 3168 8635 3224
rect 3742 3166 8635 3168
rect 8710 3224 8819 3229
rect 14089 3226 14155 3229
rect 8710 3168 8758 3224
rect 8814 3168 8819 3224
rect 8710 3166 8819 3168
rect 8569 3163 8635 3166
rect 8753 3163 8819 3166
rect 9630 3224 14155 3226
rect 9630 3168 14094 3224
rect 14150 3168 14155 3224
rect 9630 3166 14155 3168
rect 5441 3090 5507 3093
rect 5942 3090 5948 3092
rect 2822 3088 5948 3090
rect 2822 3032 5446 3088
rect 5502 3032 5948 3088
rect 2822 3030 5948 3032
rect 0 3000 120 3030
rect 2221 3027 2287 3030
rect 3049 2954 3115 2957
rect 3190 2954 3250 3030
rect 5441 3027 5507 3030
rect 5942 3028 5948 3030
rect 6012 3090 6018 3092
rect 8334 3090 8340 3092
rect 6012 3030 8340 3090
rect 6012 3028 6018 3030
rect 8334 3028 8340 3030
rect 8404 3028 8410 3092
rect 8702 3028 8708 3092
rect 8772 3090 8778 3092
rect 9630 3090 9690 3166
rect 14089 3163 14155 3166
rect 16849 3226 16915 3229
rect 18781 3226 18847 3229
rect 16849 3224 18847 3226
rect 16849 3168 16854 3224
rect 16910 3168 18786 3224
rect 18842 3168 18847 3224
rect 16849 3166 18847 3168
rect 16849 3163 16915 3166
rect 18781 3163 18847 3166
rect 19333 3226 19399 3229
rect 20713 3226 20779 3229
rect 19333 3224 20779 3226
rect 19333 3168 19338 3224
rect 19394 3168 20718 3224
rect 20774 3168 20779 3224
rect 19333 3166 20779 3168
rect 19333 3163 19399 3166
rect 20713 3163 20779 3166
rect 23657 3226 23723 3229
rect 27705 3226 27771 3229
rect 28625 3226 28691 3229
rect 23657 3224 26434 3226
rect 23657 3168 23662 3224
rect 23718 3168 26434 3224
rect 23657 3166 26434 3168
rect 23657 3163 23723 3166
rect 8772 3030 9690 3090
rect 10317 3090 10383 3093
rect 11881 3090 11947 3093
rect 10317 3088 11947 3090
rect 10317 3032 10322 3088
rect 10378 3032 11886 3088
rect 11942 3032 11947 3088
rect 10317 3030 11947 3032
rect 8772 3028 8778 3030
rect 10317 3027 10383 3030
rect 11881 3027 11947 3030
rect 12433 3090 12499 3093
rect 14181 3090 14247 3093
rect 12433 3088 14247 3090
rect 12433 3032 12438 3088
rect 12494 3032 14186 3088
rect 14242 3032 14247 3088
rect 12433 3030 14247 3032
rect 12433 3027 12499 3030
rect 14181 3027 14247 3030
rect 15101 3090 15167 3093
rect 15561 3090 15627 3093
rect 18045 3090 18111 3093
rect 15101 3088 15627 3090
rect 15101 3032 15106 3088
rect 15162 3032 15566 3088
rect 15622 3032 15627 3088
rect 15101 3030 15627 3032
rect 15101 3027 15167 3030
rect 15561 3027 15627 3030
rect 17542 3088 18111 3090
rect 17542 3032 18050 3088
rect 18106 3032 18111 3088
rect 17542 3030 18111 3032
rect 3049 2952 3250 2954
rect 3049 2896 3054 2952
rect 3110 2896 3250 2952
rect 3049 2894 3250 2896
rect 4245 2954 4311 2957
rect 10593 2954 10659 2957
rect 12617 2956 12683 2957
rect 4245 2952 10659 2954
rect 4245 2896 4250 2952
rect 4306 2896 10598 2952
rect 10654 2896 10659 2952
rect 4245 2894 10659 2896
rect 3049 2891 3115 2894
rect 4245 2891 4311 2894
rect 10593 2891 10659 2894
rect 12566 2892 12572 2956
rect 12636 2954 12683 2956
rect 13169 2954 13235 2957
rect 13302 2954 13308 2956
rect 12636 2952 12728 2954
rect 12678 2896 12728 2952
rect 12636 2894 12728 2896
rect 13169 2952 13308 2954
rect 13169 2896 13174 2952
rect 13230 2896 13308 2952
rect 13169 2894 13308 2896
rect 12636 2892 12683 2894
rect 12617 2891 12683 2892
rect 13169 2891 13235 2894
rect 13302 2892 13308 2894
rect 13372 2892 13378 2956
rect 14089 2954 14155 2957
rect 14641 2954 14707 2957
rect 16941 2954 17007 2957
rect 17542 2954 17602 3030
rect 18045 3027 18111 3030
rect 19057 3090 19123 3093
rect 20989 3090 21055 3093
rect 19057 3088 21055 3090
rect 19057 3032 19062 3088
rect 19118 3032 20994 3088
rect 21050 3032 21055 3088
rect 19057 3030 21055 3032
rect 19057 3027 19123 3030
rect 20989 3027 21055 3030
rect 21173 3090 21239 3093
rect 23013 3090 23079 3093
rect 21173 3088 23079 3090
rect 21173 3032 21178 3088
rect 21234 3032 23018 3088
rect 23074 3032 23079 3088
rect 21173 3030 23079 3032
rect 21173 3027 21239 3030
rect 23013 3027 23079 3030
rect 25037 3090 25103 3093
rect 26141 3090 26207 3093
rect 25037 3088 26207 3090
rect 25037 3032 25042 3088
rect 25098 3032 26146 3088
rect 26202 3032 26207 3088
rect 25037 3030 26207 3032
rect 26374 3090 26434 3166
rect 27705 3224 28691 3226
rect 27705 3168 27710 3224
rect 27766 3168 28630 3224
rect 28686 3168 28691 3224
rect 27705 3166 28691 3168
rect 27705 3163 27771 3166
rect 28625 3163 28691 3166
rect 29453 3226 29519 3229
rect 29729 3226 29795 3229
rect 29453 3224 29795 3226
rect 29453 3168 29458 3224
rect 29514 3168 29734 3224
rect 29790 3168 29795 3224
rect 29453 3166 29795 3168
rect 29453 3163 29519 3166
rect 29729 3163 29795 3166
rect 35709 3090 35775 3093
rect 26374 3088 35775 3090
rect 26374 3032 35714 3088
rect 35770 3032 35775 3088
rect 26374 3030 35775 3032
rect 25037 3027 25103 3030
rect 26141 3027 26207 3030
rect 35709 3027 35775 3030
rect 39389 3090 39455 3093
rect 40880 3090 41000 3120
rect 39389 3088 41000 3090
rect 39389 3032 39394 3088
rect 39450 3032 41000 3088
rect 39389 3030 41000 3032
rect 39389 3027 39455 3030
rect 40880 3000 41000 3030
rect 14089 2952 14474 2954
rect 14089 2896 14094 2952
rect 14150 2896 14474 2952
rect 14089 2894 14474 2896
rect 14089 2891 14155 2894
rect 0 2818 120 2848
rect 1393 2818 1459 2821
rect 0 2816 1459 2818
rect 0 2760 1398 2816
rect 1454 2760 1459 2816
rect 0 2758 1459 2760
rect 0 2728 120 2758
rect 1393 2755 1459 2758
rect 3734 2756 3740 2820
rect 3804 2818 3810 2820
rect 7097 2818 7163 2821
rect 3804 2816 7163 2818
rect 3804 2760 7102 2816
rect 7158 2760 7163 2816
rect 3804 2758 7163 2760
rect 3804 2756 3810 2758
rect 7097 2755 7163 2758
rect 8702 2756 8708 2820
rect 8772 2818 8778 2820
rect 9121 2818 9187 2821
rect 11646 2818 11652 2820
rect 8772 2816 9187 2818
rect 8772 2760 9126 2816
rect 9182 2760 9187 2816
rect 8772 2758 9187 2760
rect 8772 2756 8778 2758
rect 9121 2755 9187 2758
rect 9630 2758 11652 2818
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 2773 2682 2839 2685
rect 4838 2682 4844 2684
rect 2773 2680 4844 2682
rect 2773 2624 2778 2680
rect 2834 2624 4844 2680
rect 2773 2622 4844 2624
rect 2773 2619 2839 2622
rect 4838 2620 4844 2622
rect 4908 2620 4914 2684
rect 0 2546 120 2576
rect 1485 2546 1551 2549
rect 0 2544 1551 2546
rect 0 2488 1490 2544
rect 1546 2488 1551 2544
rect 0 2486 1551 2488
rect 0 2456 120 2486
rect 1485 2483 1551 2486
rect 2405 2546 2471 2549
rect 9630 2546 9690 2758
rect 11646 2756 11652 2758
rect 11716 2756 11722 2820
rect 14414 2818 14474 2894
rect 14641 2952 17602 2954
rect 14641 2896 14646 2952
rect 14702 2896 16946 2952
rect 17002 2896 17602 2952
rect 14641 2894 17602 2896
rect 17769 2954 17835 2957
rect 22277 2954 22343 2957
rect 17769 2952 22343 2954
rect 17769 2896 17774 2952
rect 17830 2896 22282 2952
rect 22338 2896 22343 2952
rect 17769 2894 22343 2896
rect 14641 2891 14707 2894
rect 16941 2891 17007 2894
rect 17769 2891 17835 2894
rect 22277 2891 22343 2894
rect 25129 2954 25195 2957
rect 25681 2954 25747 2957
rect 26785 2954 26851 2957
rect 29545 2954 29611 2957
rect 25129 2952 25747 2954
rect 25129 2896 25134 2952
rect 25190 2896 25686 2952
rect 25742 2896 25747 2952
rect 25129 2894 25747 2896
rect 25129 2891 25195 2894
rect 25681 2891 25747 2894
rect 25822 2894 26664 2954
rect 18689 2818 18755 2821
rect 19057 2818 19123 2821
rect 14414 2816 19123 2818
rect 14414 2760 18694 2816
rect 18750 2760 19062 2816
rect 19118 2760 19123 2816
rect 14414 2758 19123 2760
rect 18689 2755 18755 2758
rect 19057 2755 19123 2758
rect 20989 2818 21055 2821
rect 25822 2818 25882 2894
rect 20989 2816 25882 2818
rect 20989 2760 20994 2816
rect 21050 2760 25882 2816
rect 20989 2758 25882 2760
rect 26604 2818 26664 2894
rect 26785 2952 29611 2954
rect 26785 2896 26790 2952
rect 26846 2896 29550 2952
rect 29606 2896 29611 2952
rect 26785 2894 29611 2896
rect 26785 2891 26851 2894
rect 29545 2891 29611 2894
rect 29821 2954 29887 2957
rect 30005 2954 30071 2957
rect 36629 2954 36695 2957
rect 29821 2952 30071 2954
rect 29821 2896 29826 2952
rect 29882 2896 30010 2952
rect 30066 2896 30071 2952
rect 29821 2894 30071 2896
rect 29821 2891 29887 2894
rect 30005 2891 30071 2894
rect 30238 2952 36695 2954
rect 30238 2896 36634 2952
rect 36690 2896 36695 2952
rect 30238 2894 36695 2896
rect 26969 2818 27035 2821
rect 26604 2816 27035 2818
rect 26604 2760 26974 2816
rect 27030 2760 27035 2816
rect 26604 2758 27035 2760
rect 20989 2755 21055 2758
rect 26969 2755 27035 2758
rect 28349 2818 28415 2821
rect 28809 2818 28875 2821
rect 30097 2818 30163 2821
rect 28349 2816 28875 2818
rect 28349 2760 28354 2816
rect 28410 2760 28814 2816
rect 28870 2760 28875 2816
rect 28349 2758 28875 2760
rect 28349 2755 28415 2758
rect 28809 2755 28875 2758
rect 28950 2816 30163 2818
rect 28950 2760 30102 2816
rect 30158 2760 30163 2816
rect 28950 2758 30163 2760
rect 13946 2752 14262 2753
rect 13946 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14262 2752
rect 13946 2687 14262 2688
rect 19946 2752 20262 2753
rect 19946 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20262 2752
rect 19946 2687 20262 2688
rect 25946 2752 26262 2753
rect 25946 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26262 2752
rect 25946 2687 26262 2688
rect 13118 2620 13124 2684
rect 13188 2682 13194 2684
rect 13721 2682 13787 2685
rect 13188 2680 13787 2682
rect 13188 2624 13726 2680
rect 13782 2624 13787 2680
rect 13188 2622 13787 2624
rect 13188 2620 13194 2622
rect 13721 2619 13787 2622
rect 15469 2682 15535 2685
rect 16205 2682 16271 2685
rect 18045 2682 18111 2685
rect 15469 2680 18111 2682
rect 15469 2624 15474 2680
rect 15530 2624 16210 2680
rect 16266 2624 18050 2680
rect 18106 2624 18111 2680
rect 15469 2622 18111 2624
rect 15469 2619 15535 2622
rect 16205 2619 16271 2622
rect 18045 2619 18111 2622
rect 18781 2684 18847 2685
rect 18781 2680 18828 2684
rect 18892 2682 18898 2684
rect 24158 2682 24164 2684
rect 18781 2624 18786 2680
rect 18781 2620 18828 2624
rect 18892 2622 18938 2682
rect 20348 2622 24164 2682
rect 18892 2620 18898 2622
rect 18781 2619 18847 2620
rect 2405 2544 9690 2546
rect 2405 2488 2410 2544
rect 2466 2488 9690 2544
rect 2405 2486 9690 2488
rect 13905 2546 13971 2549
rect 15837 2546 15903 2549
rect 17769 2546 17835 2549
rect 13905 2544 17835 2546
rect 13905 2488 13910 2544
rect 13966 2488 15842 2544
rect 15898 2488 17774 2544
rect 17830 2488 17835 2544
rect 13905 2486 17835 2488
rect 2405 2483 2471 2486
rect 13905 2483 13971 2486
rect 15837 2483 15903 2486
rect 17769 2483 17835 2486
rect 19057 2546 19123 2549
rect 19190 2546 19196 2548
rect 19057 2544 19196 2546
rect 19057 2488 19062 2544
rect 19118 2488 19196 2544
rect 19057 2486 19196 2488
rect 19057 2483 19123 2486
rect 19190 2484 19196 2486
rect 19260 2484 19266 2548
rect 2405 2410 2471 2413
rect 20348 2410 20408 2622
rect 24158 2620 24164 2622
rect 24228 2620 24234 2684
rect 26972 2682 27032 2755
rect 28257 2682 28323 2685
rect 28625 2682 28691 2685
rect 26972 2680 28691 2682
rect 26972 2624 28262 2680
rect 28318 2624 28630 2680
rect 28686 2624 28691 2680
rect 26972 2622 28691 2624
rect 28257 2619 28323 2622
rect 28625 2619 28691 2622
rect 28809 2682 28875 2685
rect 28950 2682 29010 2758
rect 30097 2755 30163 2758
rect 28809 2680 29010 2682
rect 28809 2624 28814 2680
rect 28870 2624 29010 2680
rect 28809 2622 29010 2624
rect 28809 2619 28875 2622
rect 30238 2546 30298 2894
rect 36629 2891 36695 2894
rect 39021 2818 39087 2821
rect 40880 2818 41000 2848
rect 39021 2816 41000 2818
rect 39021 2760 39026 2816
rect 39082 2760 41000 2816
rect 39021 2758 41000 2760
rect 39021 2755 39087 2758
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 37946 2752 38262 2753
rect 37946 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38262 2752
rect 40880 2728 41000 2758
rect 37946 2687 38262 2688
rect 2405 2408 20408 2410
rect 2405 2352 2410 2408
rect 2466 2352 20408 2408
rect 2405 2350 20408 2352
rect 20486 2486 30298 2546
rect 35893 2546 35959 2549
rect 38101 2546 38167 2549
rect 35893 2544 38167 2546
rect 35893 2488 35898 2544
rect 35954 2488 38106 2544
rect 38162 2488 38167 2544
rect 35893 2486 38167 2488
rect 2405 2347 2471 2350
rect 0 2274 120 2304
rect 1853 2274 1919 2277
rect 0 2272 1919 2274
rect 0 2216 1858 2272
rect 1914 2216 1919 2272
rect 0 2214 1919 2216
rect 0 2184 120 2214
rect 1853 2211 1919 2214
rect 7281 2274 7347 2277
rect 8702 2274 8708 2276
rect 7281 2272 8708 2274
rect 7281 2216 7286 2272
rect 7342 2216 8708 2272
rect 7281 2214 8708 2216
rect 7281 2211 7347 2214
rect 8702 2212 8708 2214
rect 8772 2212 8778 2276
rect 13353 2274 13419 2277
rect 14641 2274 14707 2277
rect 13353 2272 14707 2274
rect 13353 2216 13358 2272
rect 13414 2216 14646 2272
rect 14702 2216 14707 2272
rect 13353 2214 14707 2216
rect 13353 2211 13419 2214
rect 14641 2211 14707 2214
rect 17125 2274 17191 2277
rect 20486 2274 20546 2486
rect 35893 2483 35959 2486
rect 38101 2483 38167 2486
rect 39665 2546 39731 2549
rect 40880 2546 41000 2576
rect 39665 2544 41000 2546
rect 39665 2488 39670 2544
rect 39726 2488 41000 2544
rect 39665 2486 41000 2488
rect 39665 2483 39731 2486
rect 40880 2456 41000 2486
rect 25630 2348 25636 2412
rect 25700 2410 25706 2412
rect 39205 2410 39271 2413
rect 25700 2408 39271 2410
rect 25700 2352 39210 2408
rect 39266 2352 39271 2408
rect 25700 2350 39271 2352
rect 25700 2348 25706 2350
rect 39205 2347 39271 2350
rect 17125 2272 20546 2274
rect 17125 2216 17130 2272
rect 17186 2216 20546 2272
rect 17125 2214 20546 2216
rect 23749 2274 23815 2277
rect 26877 2274 26943 2277
rect 23749 2272 26943 2274
rect 23749 2216 23754 2272
rect 23810 2216 26882 2272
rect 26938 2216 26943 2272
rect 23749 2214 26943 2216
rect 17125 2211 17191 2214
rect 23749 2211 23815 2214
rect 26877 2211 26943 2214
rect 39941 2274 40007 2277
rect 40880 2274 41000 2304
rect 39941 2272 41000 2274
rect 39941 2216 39946 2272
rect 40002 2216 41000 2272
rect 39941 2214 41000 2216
rect 39941 2211 40007 2214
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 9006 2208 9322 2209
rect 9006 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9322 2208
rect 9006 2143 9322 2144
rect 15006 2208 15322 2209
rect 15006 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15322 2208
rect 15006 2143 15322 2144
rect 21006 2208 21322 2209
rect 21006 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21322 2208
rect 21006 2143 21322 2144
rect 27006 2208 27322 2209
rect 27006 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27322 2208
rect 27006 2143 27322 2144
rect 33006 2208 33322 2209
rect 33006 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33322 2208
rect 33006 2143 33322 2144
rect 39006 2208 39322 2209
rect 39006 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39322 2208
rect 40880 2184 41000 2214
rect 39006 2143 39322 2144
rect 9438 2076 9444 2140
rect 9508 2138 9514 2140
rect 9581 2138 9647 2141
rect 20846 2138 20852 2140
rect 9508 2136 9647 2138
rect 9508 2080 9586 2136
rect 9642 2080 9647 2136
rect 9508 2078 9647 2080
rect 9508 2076 9514 2078
rect 9581 2075 9647 2078
rect 16438 2078 20852 2138
rect 0 2002 120 2032
rect 473 2002 539 2005
rect 0 2000 539 2002
rect 0 1944 478 2000
rect 534 1944 539 2000
rect 0 1942 539 1944
rect 0 1912 120 1942
rect 473 1939 539 1942
rect 4337 2002 4403 2005
rect 10726 2002 10732 2004
rect 4337 2000 10732 2002
rect 4337 1944 4342 2000
rect 4398 1944 10732 2000
rect 4337 1942 10732 1944
rect 4337 1939 4403 1942
rect 10726 1940 10732 1942
rect 10796 1940 10802 2004
rect 11053 2002 11119 2005
rect 16438 2002 16498 2078
rect 20846 2076 20852 2078
rect 20916 2076 20922 2140
rect 21449 2138 21515 2141
rect 25262 2138 25268 2140
rect 21449 2136 25268 2138
rect 21449 2080 21454 2136
rect 21510 2080 25268 2136
rect 21449 2078 25268 2080
rect 21449 2075 21515 2078
rect 25262 2076 25268 2078
rect 25332 2076 25338 2140
rect 11053 2000 16498 2002
rect 11053 1944 11058 2000
rect 11114 1944 16498 2000
rect 11053 1942 16498 1944
rect 18137 2002 18203 2005
rect 25129 2002 25195 2005
rect 18137 2000 25195 2002
rect 18137 1944 18142 2000
rect 18198 1944 25134 2000
rect 25190 1944 25195 2000
rect 18137 1942 25195 1944
rect 11053 1939 11119 1942
rect 18137 1939 18203 1942
rect 25129 1939 25195 1942
rect 39573 2002 39639 2005
rect 40880 2002 41000 2032
rect 39573 2000 41000 2002
rect 39573 1944 39578 2000
rect 39634 1944 41000 2000
rect 39573 1942 41000 1944
rect 39573 1939 39639 1942
rect 40880 1912 41000 1942
rect 4102 1804 4108 1868
rect 4172 1866 4178 1868
rect 11421 1866 11487 1869
rect 4172 1864 11487 1866
rect 4172 1808 11426 1864
rect 11482 1808 11487 1864
rect 4172 1806 11487 1808
rect 4172 1804 4178 1806
rect 11421 1803 11487 1806
rect 11881 1866 11947 1869
rect 15837 1866 15903 1869
rect 11881 1864 15903 1866
rect 11881 1808 11886 1864
rect 11942 1808 15842 1864
rect 15898 1808 15903 1864
rect 11881 1806 15903 1808
rect 11881 1803 11947 1806
rect 15837 1803 15903 1806
rect 16297 1866 16363 1869
rect 34605 1866 34671 1869
rect 16297 1864 34671 1866
rect 16297 1808 16302 1864
rect 16358 1808 34610 1864
rect 34666 1808 34671 1864
rect 16297 1806 34671 1808
rect 16297 1803 16363 1806
rect 34605 1803 34671 1806
rect 0 1730 120 1760
rect 1209 1730 1275 1733
rect 0 1728 1275 1730
rect 0 1672 1214 1728
rect 1270 1672 1275 1728
rect 0 1670 1275 1672
rect 0 1640 120 1670
rect 1209 1667 1275 1670
rect 2773 1730 2839 1733
rect 31201 1730 31267 1733
rect 2773 1728 31267 1730
rect 2773 1672 2778 1728
rect 2834 1672 31206 1728
rect 31262 1672 31267 1728
rect 2773 1670 31267 1672
rect 2773 1667 2839 1670
rect 31201 1667 31267 1670
rect 38653 1730 38719 1733
rect 40880 1730 41000 1760
rect 38653 1728 41000 1730
rect 38653 1672 38658 1728
rect 38714 1672 41000 1728
rect 38653 1670 41000 1672
rect 38653 1667 38719 1670
rect 40880 1640 41000 1670
rect 1577 1594 1643 1597
rect 11053 1594 11119 1597
rect 1577 1592 11119 1594
rect 1577 1536 1582 1592
rect 1638 1536 11058 1592
rect 11114 1536 11119 1592
rect 1577 1534 11119 1536
rect 1577 1531 1643 1534
rect 11053 1531 11119 1534
rect 12249 1594 12315 1597
rect 16481 1594 16547 1597
rect 21449 1594 21515 1597
rect 12249 1592 16547 1594
rect 12249 1536 12254 1592
rect 12310 1536 16486 1592
rect 16542 1536 16547 1592
rect 12249 1534 16547 1536
rect 12249 1531 12315 1534
rect 16481 1531 16547 1534
rect 16622 1592 21515 1594
rect 16622 1536 21454 1592
rect 21510 1536 21515 1592
rect 16622 1534 21515 1536
rect 0 1458 120 1488
rect 749 1458 815 1461
rect 0 1456 815 1458
rect 0 1400 754 1456
rect 810 1400 815 1456
rect 0 1398 815 1400
rect 0 1368 120 1398
rect 749 1395 815 1398
rect 9673 1458 9739 1461
rect 16622 1458 16682 1534
rect 21449 1531 21515 1534
rect 22093 1594 22159 1597
rect 22502 1594 22508 1596
rect 22093 1592 22508 1594
rect 22093 1536 22098 1592
rect 22154 1536 22508 1592
rect 22093 1534 22508 1536
rect 22093 1531 22159 1534
rect 22502 1532 22508 1534
rect 22572 1532 22578 1596
rect 23013 1594 23079 1597
rect 33777 1594 33843 1597
rect 23013 1592 33843 1594
rect 23013 1536 23018 1592
rect 23074 1536 33782 1592
rect 33838 1536 33843 1592
rect 23013 1534 33843 1536
rect 23013 1531 23079 1534
rect 33777 1531 33843 1534
rect 9673 1456 16682 1458
rect 9673 1400 9678 1456
rect 9734 1400 16682 1456
rect 9673 1398 16682 1400
rect 16757 1458 16823 1461
rect 35433 1458 35499 1461
rect 16757 1456 35499 1458
rect 16757 1400 16762 1456
rect 16818 1400 35438 1456
rect 35494 1400 35499 1456
rect 16757 1398 35499 1400
rect 9673 1395 9739 1398
rect 16757 1395 16823 1398
rect 35433 1395 35499 1398
rect 40033 1458 40099 1461
rect 40880 1458 41000 1488
rect 40033 1456 41000 1458
rect 40033 1400 40038 1456
rect 40094 1400 41000 1456
rect 40033 1398 41000 1400
rect 40033 1395 40099 1398
rect 40880 1368 41000 1398
rect 5441 1324 5507 1325
rect 5390 1260 5396 1324
rect 5460 1322 5507 1324
rect 5460 1320 5552 1322
rect 5502 1264 5552 1320
rect 5460 1262 5552 1264
rect 5460 1260 5507 1262
rect 6678 1260 6684 1324
rect 6748 1322 6754 1324
rect 8477 1322 8543 1325
rect 6748 1320 8543 1322
rect 6748 1264 8482 1320
rect 8538 1264 8543 1320
rect 6748 1262 8543 1264
rect 6748 1260 6754 1262
rect 5441 1259 5507 1260
rect 8477 1259 8543 1262
rect 17902 1260 17908 1324
rect 17972 1322 17978 1324
rect 25129 1322 25195 1325
rect 17972 1320 25195 1322
rect 17972 1264 25134 1320
rect 25190 1264 25195 1320
rect 17972 1262 25195 1264
rect 17972 1260 17978 1262
rect 25129 1259 25195 1262
rect 25865 1322 25931 1325
rect 27470 1322 27476 1324
rect 25865 1320 27476 1322
rect 25865 1264 25870 1320
rect 25926 1264 27476 1320
rect 25865 1262 27476 1264
rect 25865 1259 25931 1262
rect 27470 1260 27476 1262
rect 27540 1260 27546 1324
rect 28349 1322 28415 1325
rect 34513 1322 34579 1325
rect 28349 1320 34579 1322
rect 28349 1264 28354 1320
rect 28410 1264 34518 1320
rect 34574 1264 34579 1320
rect 28349 1262 34579 1264
rect 28349 1259 28415 1262
rect 34513 1259 34579 1262
rect 5206 1124 5212 1188
rect 5276 1186 5282 1188
rect 7373 1186 7439 1189
rect 5276 1184 7439 1186
rect 5276 1128 7378 1184
rect 7434 1128 7439 1184
rect 5276 1126 7439 1128
rect 5276 1124 5282 1126
rect 7373 1123 7439 1126
rect 11646 1124 11652 1188
rect 11716 1186 11722 1188
rect 17861 1186 17927 1189
rect 28441 1186 28507 1189
rect 11716 1184 17927 1186
rect 11716 1128 17866 1184
rect 17922 1128 17927 1184
rect 11716 1126 17927 1128
rect 11716 1124 11722 1126
rect 17861 1123 17927 1126
rect 18048 1184 28507 1186
rect 18048 1128 28446 1184
rect 28502 1128 28507 1184
rect 18048 1126 28507 1128
rect 4797 1050 4863 1053
rect 16481 1050 16547 1053
rect 4797 1048 16547 1050
rect 4797 992 4802 1048
rect 4858 992 16486 1048
rect 16542 992 16547 1048
rect 4797 990 16547 992
rect 4797 987 4863 990
rect 16481 987 16547 990
rect 16614 988 16620 1052
rect 16684 1050 16690 1052
rect 18048 1050 18108 1126
rect 28441 1123 28507 1126
rect 16684 990 18108 1050
rect 28625 1050 28691 1053
rect 35157 1050 35223 1053
rect 28625 1048 35223 1050
rect 28625 992 28630 1048
rect 28686 992 35162 1048
rect 35218 992 35223 1048
rect 28625 990 35223 992
rect 16684 988 16690 990
rect 28625 987 28691 990
rect 35157 987 35223 990
rect 3693 914 3759 917
rect 16481 914 16547 917
rect 3693 912 16547 914
rect 3693 856 3698 912
rect 3754 856 16486 912
rect 16542 856 16547 912
rect 3693 854 16547 856
rect 3693 851 3759 854
rect 16481 851 16547 854
rect 16665 914 16731 917
rect 23013 914 23079 917
rect 28809 914 28875 917
rect 16665 912 22110 914
rect 16665 856 16670 912
rect 16726 856 22110 912
rect 16665 854 22110 856
rect 16665 851 16731 854
rect 2630 716 2636 780
rect 2700 778 2706 780
rect 16389 778 16455 781
rect 2700 776 16455 778
rect 2700 720 16394 776
rect 16450 720 16455 776
rect 2700 718 16455 720
rect 22050 778 22110 854
rect 23013 912 28875 914
rect 23013 856 23018 912
rect 23074 856 28814 912
rect 28870 856 28875 912
rect 23013 854 28875 856
rect 23013 851 23079 854
rect 28809 851 28875 854
rect 36169 778 36235 781
rect 22050 776 36235 778
rect 22050 720 36174 776
rect 36230 720 36235 776
rect 22050 718 36235 720
rect 2700 716 2706 718
rect 16389 715 16455 718
rect 36169 715 36235 718
rect 5533 642 5599 645
rect 22134 642 22140 644
rect 5533 640 22140 642
rect 5533 584 5538 640
rect 5594 584 22140 640
rect 5533 582 22140 584
rect 5533 579 5599 582
rect 22134 580 22140 582
rect 22204 580 22210 644
rect 7782 444 7788 508
rect 7852 506 7858 508
rect 21357 506 21423 509
rect 7852 504 21423 506
rect 7852 448 21362 504
rect 21418 448 21423 504
rect 7852 446 21423 448
rect 7852 444 7858 446
rect 21357 443 21423 446
rect 13670 308 13676 372
rect 13740 370 13746 372
rect 30189 370 30255 373
rect 13740 368 30255 370
rect 13740 312 30194 368
rect 30250 312 30255 368
rect 13740 310 30255 312
rect 13740 308 13746 310
rect 30189 307 30255 310
rect 19425 234 19491 237
rect 32765 234 32831 237
rect 19425 232 32831 234
rect 19425 176 19430 232
rect 19486 176 32770 232
rect 32826 176 32831 232
rect 19425 174 32831 176
rect 19425 171 19491 174
rect 32765 171 32831 174
rect 6494 36 6500 100
rect 6564 98 6570 100
rect 11237 98 11303 101
rect 6564 96 11303 98
rect 6564 40 11242 96
rect 11298 40 11303 96
rect 6564 38 11303 40
rect 6564 36 6570 38
rect 11237 35 11303 38
rect 15193 98 15259 101
rect 33317 98 33383 101
rect 15193 96 33383 98
rect 15193 40 15198 96
rect 15254 40 33322 96
rect 33378 40 33383 96
rect 15193 38 33383 40
rect 15193 35 15259 38
rect 33317 35 33383 38
<< via3 >>
rect 30420 10100 30484 10164
rect 11100 9828 11164 9892
rect 16620 9692 16684 9756
rect 8524 8876 8588 8940
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 9012 8732 9076 8736
rect 9012 8676 9016 8732
rect 9016 8676 9072 8732
rect 9072 8676 9076 8732
rect 9012 8672 9076 8676
rect 9092 8732 9156 8736
rect 9092 8676 9096 8732
rect 9096 8676 9152 8732
rect 9152 8676 9156 8732
rect 9092 8672 9156 8676
rect 9172 8732 9236 8736
rect 9172 8676 9176 8732
rect 9176 8676 9232 8732
rect 9232 8676 9236 8732
rect 9172 8672 9236 8676
rect 9252 8732 9316 8736
rect 9252 8676 9256 8732
rect 9256 8676 9312 8732
rect 9312 8676 9316 8732
rect 9252 8672 9316 8676
rect 15012 8732 15076 8736
rect 15012 8676 15016 8732
rect 15016 8676 15072 8732
rect 15072 8676 15076 8732
rect 15012 8672 15076 8676
rect 15092 8732 15156 8736
rect 15092 8676 15096 8732
rect 15096 8676 15152 8732
rect 15152 8676 15156 8732
rect 15092 8672 15156 8676
rect 15172 8732 15236 8736
rect 15172 8676 15176 8732
rect 15176 8676 15232 8732
rect 15232 8676 15236 8732
rect 15172 8672 15236 8676
rect 15252 8732 15316 8736
rect 15252 8676 15256 8732
rect 15256 8676 15312 8732
rect 15312 8676 15316 8732
rect 15252 8672 15316 8676
rect 21012 8732 21076 8736
rect 21012 8676 21016 8732
rect 21016 8676 21072 8732
rect 21072 8676 21076 8732
rect 21012 8672 21076 8676
rect 21092 8732 21156 8736
rect 21092 8676 21096 8732
rect 21096 8676 21152 8732
rect 21152 8676 21156 8732
rect 21092 8672 21156 8676
rect 21172 8732 21236 8736
rect 21172 8676 21176 8732
rect 21176 8676 21232 8732
rect 21232 8676 21236 8732
rect 21172 8672 21236 8676
rect 21252 8732 21316 8736
rect 21252 8676 21256 8732
rect 21256 8676 21312 8732
rect 21312 8676 21316 8732
rect 21252 8672 21316 8676
rect 27012 8732 27076 8736
rect 27012 8676 27016 8732
rect 27016 8676 27072 8732
rect 27072 8676 27076 8732
rect 27012 8672 27076 8676
rect 27092 8732 27156 8736
rect 27092 8676 27096 8732
rect 27096 8676 27152 8732
rect 27152 8676 27156 8732
rect 27092 8672 27156 8676
rect 27172 8732 27236 8736
rect 27172 8676 27176 8732
rect 27176 8676 27232 8732
rect 27232 8676 27236 8732
rect 27172 8672 27236 8676
rect 27252 8732 27316 8736
rect 27252 8676 27256 8732
rect 27256 8676 27312 8732
rect 27312 8676 27316 8732
rect 27252 8672 27316 8676
rect 33012 8732 33076 8736
rect 33012 8676 33016 8732
rect 33016 8676 33072 8732
rect 33072 8676 33076 8732
rect 33012 8672 33076 8676
rect 33092 8732 33156 8736
rect 33092 8676 33096 8732
rect 33096 8676 33152 8732
rect 33152 8676 33156 8732
rect 33092 8672 33156 8676
rect 33172 8732 33236 8736
rect 33172 8676 33176 8732
rect 33176 8676 33232 8732
rect 33232 8676 33236 8732
rect 33172 8672 33236 8676
rect 33252 8732 33316 8736
rect 33252 8676 33256 8732
rect 33256 8676 33312 8732
rect 33312 8676 33316 8732
rect 33252 8672 33316 8676
rect 39012 8732 39076 8736
rect 39012 8676 39016 8732
rect 39016 8676 39072 8732
rect 39072 8676 39076 8732
rect 39012 8672 39076 8676
rect 39092 8732 39156 8736
rect 39092 8676 39096 8732
rect 39096 8676 39152 8732
rect 39152 8676 39156 8732
rect 39092 8672 39156 8676
rect 39172 8732 39236 8736
rect 39172 8676 39176 8732
rect 39176 8676 39232 8732
rect 39232 8676 39236 8732
rect 39172 8672 39236 8676
rect 39252 8732 39316 8736
rect 39252 8676 39256 8732
rect 39256 8676 39312 8732
rect 39312 8676 39316 8732
rect 39252 8672 39316 8676
rect 22508 8604 22572 8668
rect 13676 8332 13740 8396
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 13952 8188 14016 8192
rect 13952 8132 13956 8188
rect 13956 8132 14012 8188
rect 14012 8132 14016 8188
rect 13952 8128 14016 8132
rect 14032 8188 14096 8192
rect 14032 8132 14036 8188
rect 14036 8132 14092 8188
rect 14092 8132 14096 8188
rect 14032 8128 14096 8132
rect 14112 8188 14176 8192
rect 14112 8132 14116 8188
rect 14116 8132 14172 8188
rect 14172 8132 14176 8188
rect 14112 8128 14176 8132
rect 14192 8188 14256 8192
rect 14192 8132 14196 8188
rect 14196 8132 14252 8188
rect 14252 8132 14256 8188
rect 14192 8128 14256 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 20192 8188 20256 8192
rect 20192 8132 20196 8188
rect 20196 8132 20252 8188
rect 20252 8132 20256 8188
rect 20192 8128 20256 8132
rect 25952 8188 26016 8192
rect 25952 8132 25956 8188
rect 25956 8132 26012 8188
rect 26012 8132 26016 8188
rect 25952 8128 26016 8132
rect 26032 8188 26096 8192
rect 26032 8132 26036 8188
rect 26036 8132 26092 8188
rect 26092 8132 26096 8188
rect 26032 8128 26096 8132
rect 26112 8188 26176 8192
rect 26112 8132 26116 8188
rect 26116 8132 26172 8188
rect 26172 8132 26176 8188
rect 26112 8128 26176 8132
rect 26192 8188 26256 8192
rect 26192 8132 26196 8188
rect 26196 8132 26252 8188
rect 26252 8132 26256 8188
rect 26192 8128 26256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 37952 8188 38016 8192
rect 37952 8132 37956 8188
rect 37956 8132 38012 8188
rect 38012 8132 38016 8188
rect 37952 8128 38016 8132
rect 38032 8188 38096 8192
rect 38032 8132 38036 8188
rect 38036 8132 38092 8188
rect 38092 8132 38096 8188
rect 38032 8128 38096 8132
rect 38112 8188 38176 8192
rect 38112 8132 38116 8188
rect 38116 8132 38172 8188
rect 38172 8132 38176 8188
rect 38112 8128 38176 8132
rect 38192 8188 38256 8192
rect 38192 8132 38196 8188
rect 38196 8132 38252 8188
rect 38252 8132 38256 8188
rect 38192 8128 38256 8132
rect 14780 8060 14844 8124
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 11836 7848 11900 7852
rect 11836 7792 11886 7848
rect 11886 7792 11900 7848
rect 11836 7788 11900 7792
rect 14412 7652 14476 7716
rect 9012 7644 9076 7648
rect 9012 7588 9016 7644
rect 9016 7588 9072 7644
rect 9072 7588 9076 7644
rect 9012 7584 9076 7588
rect 9092 7644 9156 7648
rect 9092 7588 9096 7644
rect 9096 7588 9152 7644
rect 9152 7588 9156 7644
rect 9092 7584 9156 7588
rect 9172 7644 9236 7648
rect 9172 7588 9176 7644
rect 9176 7588 9232 7644
rect 9232 7588 9236 7644
rect 9172 7584 9236 7588
rect 9252 7644 9316 7648
rect 9252 7588 9256 7644
rect 9256 7588 9312 7644
rect 9312 7588 9316 7644
rect 9252 7584 9316 7588
rect 15012 7644 15076 7648
rect 15012 7588 15016 7644
rect 15016 7588 15072 7644
rect 15072 7588 15076 7644
rect 15012 7584 15076 7588
rect 15092 7644 15156 7648
rect 15092 7588 15096 7644
rect 15096 7588 15152 7644
rect 15152 7588 15156 7644
rect 15092 7584 15156 7588
rect 15172 7644 15236 7648
rect 15172 7588 15176 7644
rect 15176 7588 15232 7644
rect 15232 7588 15236 7644
rect 15172 7584 15236 7588
rect 15252 7644 15316 7648
rect 15252 7588 15256 7644
rect 15256 7588 15312 7644
rect 15312 7588 15316 7644
rect 15252 7584 15316 7588
rect 21588 7652 21652 7716
rect 21012 7644 21076 7648
rect 21012 7588 21016 7644
rect 21016 7588 21072 7644
rect 21072 7588 21076 7644
rect 21012 7584 21076 7588
rect 21092 7644 21156 7648
rect 21092 7588 21096 7644
rect 21096 7588 21152 7644
rect 21152 7588 21156 7644
rect 21092 7584 21156 7588
rect 21172 7644 21236 7648
rect 21172 7588 21176 7644
rect 21176 7588 21232 7644
rect 21232 7588 21236 7644
rect 21172 7584 21236 7588
rect 21252 7644 21316 7648
rect 21252 7588 21256 7644
rect 21256 7588 21312 7644
rect 21312 7588 21316 7644
rect 21252 7584 21316 7588
rect 27012 7644 27076 7648
rect 27012 7588 27016 7644
rect 27016 7588 27072 7644
rect 27072 7588 27076 7644
rect 27012 7584 27076 7588
rect 27092 7644 27156 7648
rect 27092 7588 27096 7644
rect 27096 7588 27152 7644
rect 27152 7588 27156 7644
rect 27092 7584 27156 7588
rect 27172 7644 27236 7648
rect 27172 7588 27176 7644
rect 27176 7588 27232 7644
rect 27232 7588 27236 7644
rect 27172 7584 27236 7588
rect 27252 7644 27316 7648
rect 27252 7588 27256 7644
rect 27256 7588 27312 7644
rect 27312 7588 27316 7644
rect 27252 7584 27316 7588
rect 33012 7644 33076 7648
rect 33012 7588 33016 7644
rect 33016 7588 33072 7644
rect 33072 7588 33076 7644
rect 33012 7584 33076 7588
rect 33092 7644 33156 7648
rect 33092 7588 33096 7644
rect 33096 7588 33152 7644
rect 33152 7588 33156 7644
rect 33092 7584 33156 7588
rect 33172 7644 33236 7648
rect 33172 7588 33176 7644
rect 33176 7588 33232 7644
rect 33232 7588 33236 7644
rect 33172 7584 33236 7588
rect 33252 7644 33316 7648
rect 33252 7588 33256 7644
rect 33256 7588 33312 7644
rect 33312 7588 33316 7644
rect 33252 7584 33316 7588
rect 39012 7644 39076 7648
rect 39012 7588 39016 7644
rect 39016 7588 39072 7644
rect 39072 7588 39076 7644
rect 39012 7584 39076 7588
rect 39092 7644 39156 7648
rect 39092 7588 39096 7644
rect 39096 7588 39152 7644
rect 39152 7588 39156 7644
rect 39092 7584 39156 7588
rect 39172 7644 39236 7648
rect 39172 7588 39176 7644
rect 39176 7588 39232 7644
rect 39232 7588 39236 7644
rect 39172 7584 39236 7588
rect 39252 7644 39316 7648
rect 39252 7588 39256 7644
rect 39256 7588 39312 7644
rect 39312 7588 39316 7644
rect 39252 7584 39316 7588
rect 10732 7380 10796 7444
rect 4844 7108 4908 7172
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 13952 7100 14016 7104
rect 13952 7044 13956 7100
rect 13956 7044 14012 7100
rect 14012 7044 14016 7100
rect 13952 7040 14016 7044
rect 14032 7100 14096 7104
rect 14032 7044 14036 7100
rect 14036 7044 14092 7100
rect 14092 7044 14096 7100
rect 14032 7040 14096 7044
rect 14112 7100 14176 7104
rect 14112 7044 14116 7100
rect 14116 7044 14172 7100
rect 14172 7044 14176 7100
rect 14112 7040 14176 7044
rect 14192 7100 14256 7104
rect 14192 7044 14196 7100
rect 14196 7044 14252 7100
rect 14252 7044 14256 7100
rect 14192 7040 14256 7044
rect 5396 6972 5460 7036
rect 7788 6972 7852 7036
rect 8524 7032 8588 7036
rect 8524 6976 8574 7032
rect 8574 6976 8588 7032
rect 8524 6972 8588 6976
rect 12572 6836 12636 6900
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 20192 7100 20256 7104
rect 20192 7044 20196 7100
rect 20196 7044 20252 7100
rect 20252 7044 20256 7100
rect 20192 7040 20256 7044
rect 25952 7100 26016 7104
rect 25952 7044 25956 7100
rect 25956 7044 26012 7100
rect 26012 7044 26016 7100
rect 25952 7040 26016 7044
rect 26032 7100 26096 7104
rect 26032 7044 26036 7100
rect 26036 7044 26092 7100
rect 26092 7044 26096 7100
rect 26032 7040 26096 7044
rect 26112 7100 26176 7104
rect 26112 7044 26116 7100
rect 26116 7044 26172 7100
rect 26172 7044 26176 7100
rect 26112 7040 26176 7044
rect 26192 7100 26256 7104
rect 26192 7044 26196 7100
rect 26196 7044 26252 7100
rect 26252 7044 26256 7100
rect 26192 7040 26256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 37952 7100 38016 7104
rect 37952 7044 37956 7100
rect 37956 7044 38012 7100
rect 38012 7044 38016 7100
rect 37952 7040 38016 7044
rect 38032 7100 38096 7104
rect 38032 7044 38036 7100
rect 38036 7044 38092 7100
rect 38092 7044 38096 7100
rect 38032 7040 38096 7044
rect 38112 7100 38176 7104
rect 38112 7044 38116 7100
rect 38116 7044 38172 7100
rect 38172 7044 38176 7100
rect 38112 7040 38176 7044
rect 38192 7100 38256 7104
rect 38192 7044 38196 7100
rect 38196 7044 38252 7100
rect 38252 7044 38256 7100
rect 38192 7040 38256 7044
rect 16436 6972 16500 7036
rect 20852 6972 20916 7036
rect 25636 7032 25700 7036
rect 25636 6976 25650 7032
rect 25650 6976 25700 7032
rect 25636 6972 25700 6976
rect 21588 6836 21652 6900
rect 8524 6564 8588 6628
rect 12756 6564 12820 6628
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 9012 6556 9076 6560
rect 9012 6500 9016 6556
rect 9016 6500 9072 6556
rect 9072 6500 9076 6556
rect 9012 6496 9076 6500
rect 9092 6556 9156 6560
rect 9092 6500 9096 6556
rect 9096 6500 9152 6556
rect 9152 6500 9156 6556
rect 9092 6496 9156 6500
rect 9172 6556 9236 6560
rect 9172 6500 9176 6556
rect 9176 6500 9232 6556
rect 9232 6500 9236 6556
rect 9172 6496 9236 6500
rect 9252 6556 9316 6560
rect 9252 6500 9256 6556
rect 9256 6500 9312 6556
rect 9312 6500 9316 6556
rect 9252 6496 9316 6500
rect 15012 6556 15076 6560
rect 15012 6500 15016 6556
rect 15016 6500 15072 6556
rect 15072 6500 15076 6556
rect 15012 6496 15076 6500
rect 15092 6556 15156 6560
rect 15092 6500 15096 6556
rect 15096 6500 15152 6556
rect 15152 6500 15156 6556
rect 15092 6496 15156 6500
rect 15172 6556 15236 6560
rect 15172 6500 15176 6556
rect 15176 6500 15232 6556
rect 15232 6500 15236 6556
rect 15172 6496 15236 6500
rect 15252 6556 15316 6560
rect 15252 6500 15256 6556
rect 15256 6500 15312 6556
rect 15312 6500 15316 6556
rect 15252 6496 15316 6500
rect 21012 6556 21076 6560
rect 21012 6500 21016 6556
rect 21016 6500 21072 6556
rect 21072 6500 21076 6556
rect 21012 6496 21076 6500
rect 21092 6556 21156 6560
rect 21092 6500 21096 6556
rect 21096 6500 21152 6556
rect 21152 6500 21156 6556
rect 21092 6496 21156 6500
rect 21172 6556 21236 6560
rect 21172 6500 21176 6556
rect 21176 6500 21232 6556
rect 21232 6500 21236 6556
rect 21172 6496 21236 6500
rect 21252 6556 21316 6560
rect 21252 6500 21256 6556
rect 21256 6500 21312 6556
rect 21312 6500 21316 6556
rect 21252 6496 21316 6500
rect 27012 6556 27076 6560
rect 27012 6500 27016 6556
rect 27016 6500 27072 6556
rect 27072 6500 27076 6556
rect 27012 6496 27076 6500
rect 27092 6556 27156 6560
rect 27092 6500 27096 6556
rect 27096 6500 27152 6556
rect 27152 6500 27156 6556
rect 27092 6496 27156 6500
rect 27172 6556 27236 6560
rect 27172 6500 27176 6556
rect 27176 6500 27232 6556
rect 27232 6500 27236 6556
rect 27172 6496 27236 6500
rect 27252 6556 27316 6560
rect 27252 6500 27256 6556
rect 27256 6500 27312 6556
rect 27312 6500 27316 6556
rect 27252 6496 27316 6500
rect 33012 6556 33076 6560
rect 33012 6500 33016 6556
rect 33016 6500 33072 6556
rect 33072 6500 33076 6556
rect 33012 6496 33076 6500
rect 33092 6556 33156 6560
rect 33092 6500 33096 6556
rect 33096 6500 33152 6556
rect 33152 6500 33156 6556
rect 33092 6496 33156 6500
rect 33172 6556 33236 6560
rect 33172 6500 33176 6556
rect 33176 6500 33232 6556
rect 33232 6500 33236 6556
rect 33172 6496 33236 6500
rect 33252 6556 33316 6560
rect 33252 6500 33256 6556
rect 33256 6500 33312 6556
rect 33312 6500 33316 6556
rect 33252 6496 33316 6500
rect 39012 6556 39076 6560
rect 39012 6500 39016 6556
rect 39016 6500 39072 6556
rect 39072 6500 39076 6556
rect 39012 6496 39076 6500
rect 39092 6556 39156 6560
rect 39092 6500 39096 6556
rect 39096 6500 39152 6556
rect 39152 6500 39156 6556
rect 39092 6496 39156 6500
rect 39172 6556 39236 6560
rect 39172 6500 39176 6556
rect 39176 6500 39232 6556
rect 39232 6500 39236 6556
rect 39172 6496 39236 6500
rect 39252 6556 39316 6560
rect 39252 6500 39256 6556
rect 39256 6500 39312 6556
rect 39312 6500 39316 6556
rect 39252 6496 39316 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 8524 6156 8588 6220
rect 13308 6352 13372 6356
rect 13308 6296 13322 6352
rect 13322 6296 13372 6352
rect 13308 6292 13372 6296
rect 14596 6292 14660 6356
rect 24164 6428 24228 6492
rect 9444 6020 9508 6084
rect 12572 6020 12636 6084
rect 13952 6012 14016 6016
rect 13952 5956 13956 6012
rect 13956 5956 14012 6012
rect 14012 5956 14016 6012
rect 13952 5952 14016 5956
rect 14032 6012 14096 6016
rect 14032 5956 14036 6012
rect 14036 5956 14092 6012
rect 14092 5956 14096 6012
rect 14032 5952 14096 5956
rect 14112 6012 14176 6016
rect 14112 5956 14116 6012
rect 14116 5956 14172 6012
rect 14172 5956 14176 6012
rect 14112 5952 14176 5956
rect 14192 6012 14256 6016
rect 14192 5956 14196 6012
rect 14196 5956 14252 6012
rect 14252 5956 14256 6012
rect 14192 5952 14256 5956
rect 12572 5884 12636 5948
rect 13676 5884 13740 5948
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 20192 6012 20256 6016
rect 20192 5956 20196 6012
rect 20196 5956 20252 6012
rect 20252 5956 20256 6012
rect 20192 5952 20256 5956
rect 5212 5612 5276 5676
rect 6684 5672 6748 5676
rect 6684 5616 6698 5672
rect 6698 5616 6748 5672
rect 6684 5612 6748 5616
rect 7604 5612 7668 5676
rect 5948 5536 6012 5540
rect 5948 5480 5998 5536
rect 5998 5480 6012 5536
rect 5948 5476 6012 5480
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 9012 5468 9076 5472
rect 9012 5412 9016 5468
rect 9016 5412 9072 5468
rect 9072 5412 9076 5468
rect 9012 5408 9076 5412
rect 9092 5468 9156 5472
rect 9092 5412 9096 5468
rect 9096 5412 9152 5468
rect 9152 5412 9156 5468
rect 9092 5408 9156 5412
rect 9172 5468 9236 5472
rect 9172 5412 9176 5468
rect 9176 5412 9232 5468
rect 9232 5412 9236 5468
rect 9172 5408 9236 5412
rect 9252 5468 9316 5472
rect 9252 5412 9256 5468
rect 9256 5412 9312 5468
rect 9312 5412 9316 5468
rect 9252 5408 9316 5412
rect 7420 5340 7484 5404
rect 8340 5340 8404 5404
rect 8524 5340 8588 5404
rect 12756 5748 12820 5812
rect 13492 5748 13556 5812
rect 22140 5884 22204 5948
rect 25952 6012 26016 6016
rect 25952 5956 25956 6012
rect 25956 5956 26012 6012
rect 26012 5956 26016 6012
rect 25952 5952 26016 5956
rect 26032 6012 26096 6016
rect 26032 5956 26036 6012
rect 26036 5956 26092 6012
rect 26092 5956 26096 6012
rect 26032 5952 26096 5956
rect 26112 6012 26176 6016
rect 26112 5956 26116 6012
rect 26116 5956 26172 6012
rect 26172 5956 26176 6012
rect 26112 5952 26176 5956
rect 26192 6012 26256 6016
rect 26192 5956 26196 6012
rect 26196 5956 26252 6012
rect 26252 5956 26256 6012
rect 26192 5952 26256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 37952 6012 38016 6016
rect 37952 5956 37956 6012
rect 37956 5956 38012 6012
rect 38012 5956 38016 6012
rect 37952 5952 38016 5956
rect 38032 6012 38096 6016
rect 38032 5956 38036 6012
rect 38036 5956 38092 6012
rect 38092 5956 38096 6012
rect 38032 5952 38096 5956
rect 38112 6012 38176 6016
rect 38112 5956 38116 6012
rect 38116 5956 38172 6012
rect 38172 5956 38176 6012
rect 38112 5952 38176 5956
rect 38192 6012 38256 6016
rect 38192 5956 38196 6012
rect 38196 5956 38252 6012
rect 38252 5956 38256 6012
rect 38192 5952 38256 5956
rect 25268 5884 25332 5948
rect 10548 5340 10612 5404
rect 15012 5468 15076 5472
rect 15012 5412 15016 5468
rect 15016 5412 15072 5468
rect 15072 5412 15076 5468
rect 15012 5408 15076 5412
rect 15092 5468 15156 5472
rect 15092 5412 15096 5468
rect 15096 5412 15152 5468
rect 15152 5412 15156 5468
rect 15092 5408 15156 5412
rect 15172 5468 15236 5472
rect 15172 5412 15176 5468
rect 15176 5412 15232 5468
rect 15232 5412 15236 5468
rect 15172 5408 15236 5412
rect 15252 5468 15316 5472
rect 15252 5412 15256 5468
rect 15256 5412 15312 5468
rect 15312 5412 15316 5468
rect 15252 5408 15316 5412
rect 21012 5468 21076 5472
rect 21012 5412 21016 5468
rect 21016 5412 21072 5468
rect 21072 5412 21076 5468
rect 21012 5408 21076 5412
rect 21092 5468 21156 5472
rect 21092 5412 21096 5468
rect 21096 5412 21152 5468
rect 21152 5412 21156 5468
rect 21092 5408 21156 5412
rect 21172 5468 21236 5472
rect 21172 5412 21176 5468
rect 21176 5412 21232 5468
rect 21232 5412 21236 5468
rect 21172 5408 21236 5412
rect 21252 5468 21316 5472
rect 21252 5412 21256 5468
rect 21256 5412 21312 5468
rect 21312 5412 21316 5468
rect 21252 5408 21316 5412
rect 27012 5468 27076 5472
rect 27012 5412 27016 5468
rect 27016 5412 27072 5468
rect 27072 5412 27076 5468
rect 27012 5408 27076 5412
rect 27092 5468 27156 5472
rect 27092 5412 27096 5468
rect 27096 5412 27152 5468
rect 27152 5412 27156 5468
rect 27092 5408 27156 5412
rect 27172 5468 27236 5472
rect 27172 5412 27176 5468
rect 27176 5412 27232 5468
rect 27232 5412 27236 5468
rect 27172 5408 27236 5412
rect 27252 5468 27316 5472
rect 27252 5412 27256 5468
rect 27256 5412 27312 5468
rect 27312 5412 27316 5468
rect 27252 5408 27316 5412
rect 33012 5468 33076 5472
rect 33012 5412 33016 5468
rect 33016 5412 33072 5468
rect 33072 5412 33076 5468
rect 33012 5408 33076 5412
rect 33092 5468 33156 5472
rect 33092 5412 33096 5468
rect 33096 5412 33152 5468
rect 33152 5412 33156 5468
rect 33092 5408 33156 5412
rect 33172 5468 33236 5472
rect 33172 5412 33176 5468
rect 33176 5412 33232 5468
rect 33232 5412 33236 5468
rect 33172 5408 33236 5412
rect 33252 5468 33316 5472
rect 33252 5412 33256 5468
rect 33256 5412 33312 5468
rect 33312 5412 33316 5468
rect 33252 5408 33316 5412
rect 39012 5468 39076 5472
rect 39012 5412 39016 5468
rect 39016 5412 39072 5468
rect 39072 5412 39076 5468
rect 39012 5408 39076 5412
rect 39092 5468 39156 5472
rect 39092 5412 39096 5468
rect 39096 5412 39152 5468
rect 39152 5412 39156 5468
rect 39092 5408 39156 5412
rect 39172 5468 39236 5472
rect 39172 5412 39176 5468
rect 39176 5412 39232 5468
rect 39232 5412 39236 5468
rect 39172 5408 39236 5412
rect 39252 5468 39316 5472
rect 39252 5412 39256 5468
rect 39256 5412 39312 5468
rect 39312 5412 39316 5468
rect 39252 5408 39316 5412
rect 3740 5204 3804 5268
rect 27660 5340 27724 5404
rect 7420 4932 7484 4996
rect 8340 4932 8404 4996
rect 11100 4932 11164 4996
rect 13124 4932 13188 4996
rect 16620 4932 16684 4996
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 13952 4924 14016 4928
rect 13952 4868 13956 4924
rect 13956 4868 14012 4924
rect 14012 4868 14016 4924
rect 13952 4864 14016 4868
rect 14032 4924 14096 4928
rect 14032 4868 14036 4924
rect 14036 4868 14092 4924
rect 14092 4868 14096 4924
rect 14032 4864 14096 4868
rect 14112 4924 14176 4928
rect 14112 4868 14116 4924
rect 14116 4868 14172 4924
rect 14172 4868 14176 4924
rect 14112 4864 14176 4868
rect 14192 4924 14256 4928
rect 14192 4868 14196 4924
rect 14196 4868 14252 4924
rect 14252 4868 14256 4924
rect 14192 4864 14256 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 20192 4924 20256 4928
rect 20192 4868 20196 4924
rect 20196 4868 20252 4924
rect 20252 4868 20256 4924
rect 20192 4864 20256 4868
rect 25952 4924 26016 4928
rect 25952 4868 25956 4924
rect 25956 4868 26012 4924
rect 26012 4868 26016 4924
rect 25952 4864 26016 4868
rect 26032 4924 26096 4928
rect 26032 4868 26036 4924
rect 26036 4868 26092 4924
rect 26092 4868 26096 4924
rect 26032 4864 26096 4868
rect 26112 4924 26176 4928
rect 26112 4868 26116 4924
rect 26116 4868 26172 4924
rect 26172 4868 26176 4924
rect 26112 4864 26176 4868
rect 26192 4924 26256 4928
rect 26192 4868 26196 4924
rect 26196 4868 26252 4924
rect 26252 4868 26256 4924
rect 26192 4864 26256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 37952 4924 38016 4928
rect 37952 4868 37956 4924
rect 37956 4868 38012 4924
rect 38012 4868 38016 4924
rect 37952 4864 38016 4868
rect 38032 4924 38096 4928
rect 38032 4868 38036 4924
rect 38036 4868 38092 4924
rect 38092 4868 38096 4924
rect 38032 4864 38096 4868
rect 38112 4924 38176 4928
rect 38112 4868 38116 4924
rect 38116 4868 38172 4924
rect 38172 4868 38176 4924
rect 38112 4864 38176 4868
rect 38192 4924 38256 4928
rect 38192 4868 38196 4924
rect 38196 4868 38252 4924
rect 38252 4868 38256 4924
rect 38192 4864 38256 4868
rect 2636 4660 2700 4724
rect 13676 4796 13740 4860
rect 14412 4796 14476 4860
rect 8524 4660 8588 4724
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 4108 4116 4172 4180
rect 6500 4116 6564 4180
rect 9444 4388 9508 4452
rect 9012 4380 9076 4384
rect 9012 4324 9016 4380
rect 9016 4324 9072 4380
rect 9072 4324 9076 4380
rect 9012 4320 9076 4324
rect 9092 4380 9156 4384
rect 9092 4324 9096 4380
rect 9096 4324 9152 4380
rect 9152 4324 9156 4380
rect 9092 4320 9156 4324
rect 9172 4380 9236 4384
rect 9172 4324 9176 4380
rect 9176 4324 9232 4380
rect 9232 4324 9236 4380
rect 9172 4320 9236 4324
rect 9252 4380 9316 4384
rect 9252 4324 9256 4380
rect 9256 4324 9312 4380
rect 9312 4324 9316 4380
rect 9252 4320 9316 4324
rect 10548 4388 10612 4452
rect 18828 4524 18892 4588
rect 15012 4380 15076 4384
rect 15012 4324 15016 4380
rect 15016 4324 15072 4380
rect 15072 4324 15076 4380
rect 15012 4320 15076 4324
rect 15092 4380 15156 4384
rect 15092 4324 15096 4380
rect 15096 4324 15152 4380
rect 15152 4324 15156 4380
rect 15092 4320 15156 4324
rect 15172 4380 15236 4384
rect 15172 4324 15176 4380
rect 15176 4324 15232 4380
rect 15232 4324 15236 4380
rect 15172 4320 15236 4324
rect 15252 4380 15316 4384
rect 15252 4324 15256 4380
rect 15256 4324 15312 4380
rect 15312 4324 15316 4380
rect 15252 4320 15316 4324
rect 21012 4380 21076 4384
rect 21012 4324 21016 4380
rect 21016 4324 21072 4380
rect 21072 4324 21076 4380
rect 21012 4320 21076 4324
rect 21092 4380 21156 4384
rect 21092 4324 21096 4380
rect 21096 4324 21152 4380
rect 21152 4324 21156 4380
rect 21092 4320 21156 4324
rect 21172 4380 21236 4384
rect 21172 4324 21176 4380
rect 21176 4324 21232 4380
rect 21232 4324 21236 4380
rect 21172 4320 21236 4324
rect 21252 4380 21316 4384
rect 21252 4324 21256 4380
rect 21256 4324 21312 4380
rect 21312 4324 21316 4380
rect 21252 4320 21316 4324
rect 27012 4380 27076 4384
rect 27012 4324 27016 4380
rect 27016 4324 27072 4380
rect 27072 4324 27076 4380
rect 27012 4320 27076 4324
rect 27092 4380 27156 4384
rect 27092 4324 27096 4380
rect 27096 4324 27152 4380
rect 27152 4324 27156 4380
rect 27092 4320 27156 4324
rect 27172 4380 27236 4384
rect 27172 4324 27176 4380
rect 27176 4324 27232 4380
rect 27232 4324 27236 4380
rect 27172 4320 27236 4324
rect 27252 4380 27316 4384
rect 27252 4324 27256 4380
rect 27256 4324 27312 4380
rect 27312 4324 27316 4380
rect 27252 4320 27316 4324
rect 33012 4380 33076 4384
rect 33012 4324 33016 4380
rect 33016 4324 33072 4380
rect 33072 4324 33076 4380
rect 33012 4320 33076 4324
rect 33092 4380 33156 4384
rect 33092 4324 33096 4380
rect 33096 4324 33152 4380
rect 33152 4324 33156 4380
rect 33092 4320 33156 4324
rect 33172 4380 33236 4384
rect 33172 4324 33176 4380
rect 33176 4324 33232 4380
rect 33232 4324 33236 4380
rect 33172 4320 33236 4324
rect 33252 4380 33316 4384
rect 33252 4324 33256 4380
rect 33256 4324 33312 4380
rect 33312 4324 33316 4380
rect 33252 4320 33316 4324
rect 39012 4380 39076 4384
rect 39012 4324 39016 4380
rect 39016 4324 39072 4380
rect 39072 4324 39076 4380
rect 39012 4320 39076 4324
rect 39092 4380 39156 4384
rect 39092 4324 39096 4380
rect 39096 4324 39152 4380
rect 39152 4324 39156 4380
rect 39092 4320 39156 4324
rect 39172 4380 39236 4384
rect 39172 4324 39176 4380
rect 39176 4324 39232 4380
rect 39232 4324 39236 4380
rect 39172 4320 39236 4324
rect 39252 4380 39316 4384
rect 39252 4324 39256 4380
rect 39256 4324 39312 4380
rect 39312 4324 39316 4380
rect 39252 4320 39316 4324
rect 19196 4252 19260 4316
rect 27476 4252 27540 4316
rect 17908 4116 17972 4180
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 8708 3844 8772 3908
rect 9444 3844 9508 3908
rect 14596 3980 14660 4044
rect 30420 3980 30484 4044
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 13952 3836 14016 3840
rect 13952 3780 13956 3836
rect 13956 3780 14012 3836
rect 14012 3780 14016 3836
rect 13952 3776 14016 3780
rect 14032 3836 14096 3840
rect 14032 3780 14036 3836
rect 14036 3780 14092 3836
rect 14092 3780 14096 3836
rect 14032 3776 14096 3780
rect 14112 3836 14176 3840
rect 14112 3780 14116 3836
rect 14116 3780 14172 3836
rect 14172 3780 14176 3836
rect 14112 3776 14176 3780
rect 14192 3836 14256 3840
rect 14192 3780 14196 3836
rect 14196 3780 14252 3836
rect 14252 3780 14256 3836
rect 14192 3776 14256 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 20192 3836 20256 3840
rect 20192 3780 20196 3836
rect 20196 3780 20252 3836
rect 20252 3780 20256 3836
rect 20192 3776 20256 3780
rect 25952 3836 26016 3840
rect 25952 3780 25956 3836
rect 25956 3780 26012 3836
rect 26012 3780 26016 3836
rect 25952 3776 26016 3780
rect 26032 3836 26096 3840
rect 26032 3780 26036 3836
rect 26036 3780 26092 3836
rect 26092 3780 26096 3836
rect 26032 3776 26096 3780
rect 26112 3836 26176 3840
rect 26112 3780 26116 3836
rect 26116 3780 26172 3836
rect 26172 3780 26176 3836
rect 26112 3776 26176 3780
rect 26192 3836 26256 3840
rect 26192 3780 26196 3836
rect 26196 3780 26252 3836
rect 26252 3780 26256 3836
rect 26192 3776 26256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 37952 3836 38016 3840
rect 37952 3780 37956 3836
rect 37956 3780 38012 3836
rect 38012 3780 38016 3836
rect 37952 3776 38016 3780
rect 38032 3836 38096 3840
rect 38032 3780 38036 3836
rect 38036 3780 38092 3836
rect 38092 3780 38096 3836
rect 38032 3776 38096 3780
rect 38112 3836 38176 3840
rect 38112 3780 38116 3836
rect 38116 3780 38172 3836
rect 38172 3780 38176 3836
rect 38112 3776 38176 3780
rect 38192 3836 38256 3840
rect 38192 3780 38196 3836
rect 38196 3780 38252 3836
rect 38252 3780 38256 3836
rect 38192 3776 38256 3780
rect 8340 3708 8404 3772
rect 13492 3768 13556 3772
rect 13492 3712 13542 3768
rect 13542 3712 13556 3768
rect 13492 3708 13556 3712
rect 14780 3768 14844 3772
rect 14780 3712 14830 3768
rect 14830 3712 14844 3768
rect 14780 3708 14844 3712
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 11836 3436 11900 3500
rect 7604 3300 7668 3364
rect 27660 3572 27724 3636
rect 9012 3292 9076 3296
rect 9012 3236 9016 3292
rect 9016 3236 9072 3292
rect 9072 3236 9076 3292
rect 9012 3232 9076 3236
rect 9092 3292 9156 3296
rect 9092 3236 9096 3292
rect 9096 3236 9152 3292
rect 9152 3236 9156 3292
rect 9092 3232 9156 3236
rect 9172 3292 9236 3296
rect 9172 3236 9176 3292
rect 9176 3236 9232 3292
rect 9232 3236 9236 3292
rect 9172 3232 9236 3236
rect 9252 3292 9316 3296
rect 9252 3236 9256 3292
rect 9256 3236 9312 3292
rect 9312 3236 9316 3292
rect 9252 3232 9316 3236
rect 15012 3292 15076 3296
rect 15012 3236 15016 3292
rect 15016 3236 15072 3292
rect 15072 3236 15076 3292
rect 15012 3232 15076 3236
rect 15092 3292 15156 3296
rect 15092 3236 15096 3292
rect 15096 3236 15152 3292
rect 15152 3236 15156 3292
rect 15092 3232 15156 3236
rect 15172 3292 15236 3296
rect 15172 3236 15176 3292
rect 15176 3236 15232 3292
rect 15232 3236 15236 3292
rect 15172 3232 15236 3236
rect 15252 3292 15316 3296
rect 15252 3236 15256 3292
rect 15256 3236 15312 3292
rect 15312 3236 15316 3292
rect 15252 3232 15316 3236
rect 21012 3292 21076 3296
rect 21012 3236 21016 3292
rect 21016 3236 21072 3292
rect 21072 3236 21076 3292
rect 21012 3232 21076 3236
rect 21092 3292 21156 3296
rect 21092 3236 21096 3292
rect 21096 3236 21152 3292
rect 21152 3236 21156 3292
rect 21092 3232 21156 3236
rect 21172 3292 21236 3296
rect 21172 3236 21176 3292
rect 21176 3236 21232 3292
rect 21232 3236 21236 3292
rect 21172 3232 21236 3236
rect 21252 3292 21316 3296
rect 21252 3236 21256 3292
rect 21256 3236 21312 3292
rect 21312 3236 21316 3292
rect 21252 3232 21316 3236
rect 27012 3292 27076 3296
rect 27012 3236 27016 3292
rect 27016 3236 27072 3292
rect 27072 3236 27076 3292
rect 27012 3232 27076 3236
rect 27092 3292 27156 3296
rect 27092 3236 27096 3292
rect 27096 3236 27152 3292
rect 27152 3236 27156 3292
rect 27092 3232 27156 3236
rect 27172 3292 27236 3296
rect 27172 3236 27176 3292
rect 27176 3236 27232 3292
rect 27232 3236 27236 3292
rect 27172 3232 27236 3236
rect 27252 3292 27316 3296
rect 27252 3236 27256 3292
rect 27256 3236 27312 3292
rect 27312 3236 27316 3292
rect 27252 3232 27316 3236
rect 33012 3292 33076 3296
rect 33012 3236 33016 3292
rect 33016 3236 33072 3292
rect 33072 3236 33076 3292
rect 33012 3232 33076 3236
rect 33092 3292 33156 3296
rect 33092 3236 33096 3292
rect 33096 3236 33152 3292
rect 33152 3236 33156 3292
rect 33092 3232 33156 3236
rect 33172 3292 33236 3296
rect 33172 3236 33176 3292
rect 33176 3236 33232 3292
rect 33232 3236 33236 3292
rect 33172 3232 33236 3236
rect 33252 3292 33316 3296
rect 33252 3236 33256 3292
rect 33256 3236 33312 3292
rect 33312 3236 33316 3292
rect 33252 3232 33316 3236
rect 39012 3292 39076 3296
rect 39012 3236 39016 3292
rect 39016 3236 39072 3292
rect 39072 3236 39076 3292
rect 39012 3232 39076 3236
rect 39092 3292 39156 3296
rect 39092 3236 39096 3292
rect 39096 3236 39152 3292
rect 39152 3236 39156 3292
rect 39092 3232 39156 3236
rect 39172 3292 39236 3296
rect 39172 3236 39176 3292
rect 39176 3236 39232 3292
rect 39232 3236 39236 3292
rect 39172 3232 39236 3236
rect 39252 3292 39316 3296
rect 39252 3236 39256 3292
rect 39256 3236 39312 3292
rect 39312 3236 39316 3292
rect 39252 3232 39316 3236
rect 5948 3028 6012 3092
rect 8340 3028 8404 3092
rect 8708 3028 8772 3092
rect 12572 2952 12636 2956
rect 12572 2896 12622 2952
rect 12622 2896 12636 2952
rect 12572 2892 12636 2896
rect 13308 2892 13372 2956
rect 3740 2756 3804 2820
rect 8708 2756 8772 2820
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 4844 2620 4908 2684
rect 11652 2756 11716 2820
rect 13952 2748 14016 2752
rect 13952 2692 13956 2748
rect 13956 2692 14012 2748
rect 14012 2692 14016 2748
rect 13952 2688 14016 2692
rect 14032 2748 14096 2752
rect 14032 2692 14036 2748
rect 14036 2692 14092 2748
rect 14092 2692 14096 2748
rect 14032 2688 14096 2692
rect 14112 2748 14176 2752
rect 14112 2692 14116 2748
rect 14116 2692 14172 2748
rect 14172 2692 14176 2748
rect 14112 2688 14176 2692
rect 14192 2748 14256 2752
rect 14192 2692 14196 2748
rect 14196 2692 14252 2748
rect 14252 2692 14256 2748
rect 14192 2688 14256 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 20192 2748 20256 2752
rect 20192 2692 20196 2748
rect 20196 2692 20252 2748
rect 20252 2692 20256 2748
rect 20192 2688 20256 2692
rect 25952 2748 26016 2752
rect 25952 2692 25956 2748
rect 25956 2692 26012 2748
rect 26012 2692 26016 2748
rect 25952 2688 26016 2692
rect 26032 2748 26096 2752
rect 26032 2692 26036 2748
rect 26036 2692 26092 2748
rect 26092 2692 26096 2748
rect 26032 2688 26096 2692
rect 26112 2748 26176 2752
rect 26112 2692 26116 2748
rect 26116 2692 26172 2748
rect 26172 2692 26176 2748
rect 26112 2688 26176 2692
rect 26192 2748 26256 2752
rect 26192 2692 26196 2748
rect 26196 2692 26252 2748
rect 26252 2692 26256 2748
rect 26192 2688 26256 2692
rect 13124 2620 13188 2684
rect 18828 2680 18892 2684
rect 18828 2624 18842 2680
rect 18842 2624 18892 2680
rect 18828 2620 18892 2624
rect 19196 2484 19260 2548
rect 24164 2620 24228 2684
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 37952 2748 38016 2752
rect 37952 2692 37956 2748
rect 37956 2692 38012 2748
rect 38012 2692 38016 2748
rect 37952 2688 38016 2692
rect 38032 2748 38096 2752
rect 38032 2692 38036 2748
rect 38036 2692 38092 2748
rect 38092 2692 38096 2748
rect 38032 2688 38096 2692
rect 38112 2748 38176 2752
rect 38112 2692 38116 2748
rect 38116 2692 38172 2748
rect 38172 2692 38176 2748
rect 38112 2688 38176 2692
rect 38192 2748 38256 2752
rect 38192 2692 38196 2748
rect 38196 2692 38252 2748
rect 38252 2692 38256 2748
rect 38192 2688 38256 2692
rect 8708 2212 8772 2276
rect 25636 2348 25700 2412
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 9012 2204 9076 2208
rect 9012 2148 9016 2204
rect 9016 2148 9072 2204
rect 9072 2148 9076 2204
rect 9012 2144 9076 2148
rect 9092 2204 9156 2208
rect 9092 2148 9096 2204
rect 9096 2148 9152 2204
rect 9152 2148 9156 2204
rect 9092 2144 9156 2148
rect 9172 2204 9236 2208
rect 9172 2148 9176 2204
rect 9176 2148 9232 2204
rect 9232 2148 9236 2204
rect 9172 2144 9236 2148
rect 9252 2204 9316 2208
rect 9252 2148 9256 2204
rect 9256 2148 9312 2204
rect 9312 2148 9316 2204
rect 9252 2144 9316 2148
rect 15012 2204 15076 2208
rect 15012 2148 15016 2204
rect 15016 2148 15072 2204
rect 15072 2148 15076 2204
rect 15012 2144 15076 2148
rect 15092 2204 15156 2208
rect 15092 2148 15096 2204
rect 15096 2148 15152 2204
rect 15152 2148 15156 2204
rect 15092 2144 15156 2148
rect 15172 2204 15236 2208
rect 15172 2148 15176 2204
rect 15176 2148 15232 2204
rect 15232 2148 15236 2204
rect 15172 2144 15236 2148
rect 15252 2204 15316 2208
rect 15252 2148 15256 2204
rect 15256 2148 15312 2204
rect 15312 2148 15316 2204
rect 15252 2144 15316 2148
rect 21012 2204 21076 2208
rect 21012 2148 21016 2204
rect 21016 2148 21072 2204
rect 21072 2148 21076 2204
rect 21012 2144 21076 2148
rect 21092 2204 21156 2208
rect 21092 2148 21096 2204
rect 21096 2148 21152 2204
rect 21152 2148 21156 2204
rect 21092 2144 21156 2148
rect 21172 2204 21236 2208
rect 21172 2148 21176 2204
rect 21176 2148 21232 2204
rect 21232 2148 21236 2204
rect 21172 2144 21236 2148
rect 21252 2204 21316 2208
rect 21252 2148 21256 2204
rect 21256 2148 21312 2204
rect 21312 2148 21316 2204
rect 21252 2144 21316 2148
rect 27012 2204 27076 2208
rect 27012 2148 27016 2204
rect 27016 2148 27072 2204
rect 27072 2148 27076 2204
rect 27012 2144 27076 2148
rect 27092 2204 27156 2208
rect 27092 2148 27096 2204
rect 27096 2148 27152 2204
rect 27152 2148 27156 2204
rect 27092 2144 27156 2148
rect 27172 2204 27236 2208
rect 27172 2148 27176 2204
rect 27176 2148 27232 2204
rect 27232 2148 27236 2204
rect 27172 2144 27236 2148
rect 27252 2204 27316 2208
rect 27252 2148 27256 2204
rect 27256 2148 27312 2204
rect 27312 2148 27316 2204
rect 27252 2144 27316 2148
rect 33012 2204 33076 2208
rect 33012 2148 33016 2204
rect 33016 2148 33072 2204
rect 33072 2148 33076 2204
rect 33012 2144 33076 2148
rect 33092 2204 33156 2208
rect 33092 2148 33096 2204
rect 33096 2148 33152 2204
rect 33152 2148 33156 2204
rect 33092 2144 33156 2148
rect 33172 2204 33236 2208
rect 33172 2148 33176 2204
rect 33176 2148 33232 2204
rect 33232 2148 33236 2204
rect 33172 2144 33236 2148
rect 33252 2204 33316 2208
rect 33252 2148 33256 2204
rect 33256 2148 33312 2204
rect 33312 2148 33316 2204
rect 33252 2144 33316 2148
rect 39012 2204 39076 2208
rect 39012 2148 39016 2204
rect 39016 2148 39072 2204
rect 39072 2148 39076 2204
rect 39012 2144 39076 2148
rect 39092 2204 39156 2208
rect 39092 2148 39096 2204
rect 39096 2148 39152 2204
rect 39152 2148 39156 2204
rect 39092 2144 39156 2148
rect 39172 2204 39236 2208
rect 39172 2148 39176 2204
rect 39176 2148 39232 2204
rect 39232 2148 39236 2204
rect 39172 2144 39236 2148
rect 39252 2204 39316 2208
rect 39252 2148 39256 2204
rect 39256 2148 39312 2204
rect 39312 2148 39316 2204
rect 39252 2144 39316 2148
rect 9444 2076 9508 2140
rect 10732 1940 10796 2004
rect 20852 2076 20916 2140
rect 25268 2076 25332 2140
rect 4108 1804 4172 1868
rect 22508 1532 22572 1596
rect 5396 1320 5460 1324
rect 5396 1264 5446 1320
rect 5446 1264 5460 1320
rect 5396 1260 5460 1264
rect 6684 1260 6748 1324
rect 17908 1260 17972 1324
rect 27476 1260 27540 1324
rect 5212 1124 5276 1188
rect 11652 1124 11716 1188
rect 16620 988 16684 1052
rect 2636 716 2700 780
rect 22140 580 22204 644
rect 7788 444 7852 508
rect 13676 308 13740 372
rect 6500 36 6564 100
<< metal4 >>
rect 1944 8192 2264 11250
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 3004 8736 3324 11250
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 7944 8192 8264 11250
rect 8523 8940 8589 8941
rect 8523 8876 8524 8940
rect 8588 8876 8589 8940
rect 8523 8875 8589 8876
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 4843 7172 4909 7173
rect 4843 7108 4844 7172
rect 4908 7108 4909 7172
rect 4843 7107 4909 7108
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 2635 4724 2701 4725
rect 2635 4660 2636 4724
rect 2700 4660 2701 4724
rect 2635 4659 2701 4660
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 0 2264 2688
rect 2638 781 2698 4659
rect 3004 4384 3324 5408
rect 3739 5268 3805 5269
rect 3739 5204 3740 5268
rect 3804 5204 3805 5268
rect 3739 5203 3805 5204
rect 3004 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3324 4384
rect 3004 3296 3324 4320
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3742 2821 3802 5203
rect 4107 4180 4173 4181
rect 4107 4116 4108 4180
rect 4172 4116 4173 4180
rect 4107 4115 4173 4116
rect 3739 2820 3805 2821
rect 3739 2756 3740 2820
rect 3804 2756 3805 2820
rect 3739 2755 3805 2756
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 2635 780 2701 781
rect 2635 716 2636 780
rect 2700 716 2701 780
rect 2635 715 2701 716
rect 3004 0 3324 2144
rect 4110 1869 4170 4115
rect 4846 2685 4906 7107
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8264 7104
rect 5395 7036 5461 7037
rect 5395 6972 5396 7036
rect 5460 6972 5461 7036
rect 5395 6971 5461 6972
rect 7787 7036 7853 7037
rect 7787 6972 7788 7036
rect 7852 6972 7853 7036
rect 7787 6971 7853 6972
rect 5211 5676 5277 5677
rect 5211 5612 5212 5676
rect 5276 5612 5277 5676
rect 5211 5611 5277 5612
rect 4843 2684 4909 2685
rect 4843 2620 4844 2684
rect 4908 2620 4909 2684
rect 4843 2619 4909 2620
rect 4107 1868 4173 1869
rect 4107 1804 4108 1868
rect 4172 1804 4173 1868
rect 4107 1803 4173 1804
rect 5214 1189 5274 5611
rect 5398 1325 5458 6971
rect 6683 5676 6749 5677
rect 6683 5612 6684 5676
rect 6748 5612 6749 5676
rect 6683 5611 6749 5612
rect 7603 5676 7669 5677
rect 7603 5612 7604 5676
rect 7668 5612 7669 5676
rect 7603 5611 7669 5612
rect 5947 5540 6013 5541
rect 5947 5476 5948 5540
rect 6012 5476 6013 5540
rect 5947 5475 6013 5476
rect 5950 3093 6010 5475
rect 6499 4180 6565 4181
rect 6499 4116 6500 4180
rect 6564 4116 6565 4180
rect 6499 4115 6565 4116
rect 5947 3092 6013 3093
rect 5947 3028 5948 3092
rect 6012 3028 6013 3092
rect 5947 3027 6013 3028
rect 5395 1324 5461 1325
rect 5395 1260 5396 1324
rect 5460 1260 5461 1324
rect 5395 1259 5461 1260
rect 5211 1188 5277 1189
rect 5211 1124 5212 1188
rect 5276 1124 5277 1188
rect 5211 1123 5277 1124
rect 6502 101 6562 4115
rect 6686 1325 6746 5611
rect 7419 5404 7485 5405
rect 7419 5340 7420 5404
rect 7484 5340 7485 5404
rect 7419 5339 7485 5340
rect 7422 4997 7482 5339
rect 7419 4996 7485 4997
rect 7419 4932 7420 4996
rect 7484 4932 7485 4996
rect 7419 4931 7485 4932
rect 7606 3365 7666 5611
rect 7603 3364 7669 3365
rect 7603 3300 7604 3364
rect 7668 3300 7669 3364
rect 7603 3299 7669 3300
rect 6683 1324 6749 1325
rect 6683 1260 6684 1324
rect 6748 1260 6749 1324
rect 6683 1259 6749 1260
rect 7790 509 7850 6971
rect 7944 6016 8264 7040
rect 8526 7037 8586 8875
rect 9004 8736 9324 11250
rect 11099 9892 11165 9893
rect 11099 9828 11100 9892
rect 11164 9828 11165 9892
rect 11099 9827 11165 9828
rect 9004 8672 9012 8736
rect 9076 8672 9092 8736
rect 9156 8672 9172 8736
rect 9236 8672 9252 8736
rect 9316 8672 9324 8736
rect 9004 7648 9324 8672
rect 9004 7584 9012 7648
rect 9076 7584 9092 7648
rect 9156 7584 9172 7648
rect 9236 7584 9252 7648
rect 9316 7584 9324 7648
rect 8523 7036 8589 7037
rect 8523 6972 8524 7036
rect 8588 6972 8589 7036
rect 8523 6971 8589 6972
rect 8523 6628 8589 6629
rect 8523 6564 8524 6628
rect 8588 6564 8589 6628
rect 8523 6563 8589 6564
rect 8526 6221 8586 6563
rect 9004 6560 9324 7584
rect 10731 7444 10797 7445
rect 10731 7380 10732 7444
rect 10796 7380 10797 7444
rect 10731 7379 10797 7380
rect 9004 6496 9012 6560
rect 9076 6496 9092 6560
rect 9156 6496 9172 6560
rect 9236 6496 9252 6560
rect 9316 6496 9324 6560
rect 8523 6220 8589 6221
rect 8523 6156 8524 6220
rect 8588 6156 8589 6220
rect 8523 6155 8589 6156
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 4928 8264 5952
rect 9004 5472 9324 6496
rect 9443 6084 9509 6085
rect 9443 6020 9444 6084
rect 9508 6020 9509 6084
rect 9443 6019 9509 6020
rect 9004 5408 9012 5472
rect 9076 5408 9092 5472
rect 9156 5408 9172 5472
rect 9236 5408 9252 5472
rect 9316 5408 9324 5472
rect 8339 5404 8405 5405
rect 8339 5340 8340 5404
rect 8404 5340 8405 5404
rect 8339 5339 8405 5340
rect 8523 5404 8589 5405
rect 8523 5340 8524 5404
rect 8588 5340 8589 5404
rect 8523 5339 8589 5340
rect 8342 4997 8402 5339
rect 8339 4996 8405 4997
rect 8339 4932 8340 4996
rect 8404 4932 8405 4996
rect 8339 4931 8405 4932
rect 7944 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 8526 4725 8586 5339
rect 8523 4724 8589 4725
rect 8523 4660 8524 4724
rect 8588 4660 8589 4724
rect 8523 4659 8589 4660
rect 9004 4384 9324 5408
rect 9446 4453 9506 6019
rect 10547 5404 10613 5405
rect 10547 5340 10548 5404
rect 10612 5340 10613 5404
rect 10547 5339 10613 5340
rect 10550 4453 10610 5339
rect 9443 4452 9509 4453
rect 9443 4388 9444 4452
rect 9508 4388 9509 4452
rect 9443 4387 9509 4388
rect 10547 4452 10613 4453
rect 10547 4388 10548 4452
rect 10612 4388 10613 4452
rect 10547 4387 10613 4388
rect 9004 4320 9012 4384
rect 9076 4320 9092 4384
rect 9156 4320 9172 4384
rect 9236 4320 9252 4384
rect 9316 4320 9324 4384
rect 8707 3908 8773 3909
rect 8707 3844 8708 3908
rect 8772 3844 8773 3908
rect 8707 3843 8773 3844
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 2752 8264 3776
rect 8339 3772 8405 3773
rect 8339 3708 8340 3772
rect 8404 3708 8405 3772
rect 8339 3707 8405 3708
rect 8342 3093 8402 3707
rect 8710 3093 8770 3843
rect 9004 3296 9324 4320
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 9004 3232 9012 3296
rect 9076 3232 9092 3296
rect 9156 3232 9172 3296
rect 9236 3232 9252 3296
rect 9316 3232 9324 3296
rect 8339 3092 8405 3093
rect 8339 3028 8340 3092
rect 8404 3028 8405 3092
rect 8339 3027 8405 3028
rect 8707 3092 8773 3093
rect 8707 3028 8708 3092
rect 8772 3028 8773 3092
rect 8707 3027 8773 3028
rect 8707 2820 8773 2821
rect 8707 2756 8708 2820
rect 8772 2756 8773 2820
rect 8707 2755 8773 2756
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7787 508 7853 509
rect 7787 444 7788 508
rect 7852 444 7853 508
rect 7787 443 7853 444
rect 6499 100 6565 101
rect 6499 36 6500 100
rect 6564 36 6565 100
rect 6499 35 6565 36
rect 7944 0 8264 2688
rect 8710 2277 8770 2755
rect 8707 2276 8773 2277
rect 8707 2212 8708 2276
rect 8772 2212 8773 2276
rect 8707 2211 8773 2212
rect 9004 2208 9324 3232
rect 9004 2144 9012 2208
rect 9076 2144 9092 2208
rect 9156 2144 9172 2208
rect 9236 2144 9252 2208
rect 9316 2144 9324 2208
rect 9004 0 9324 2144
rect 9446 2141 9506 3843
rect 9443 2140 9509 2141
rect 9443 2076 9444 2140
rect 9508 2076 9509 2140
rect 9443 2075 9509 2076
rect 10734 2005 10794 7379
rect 11102 4997 11162 9827
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 11835 7852 11901 7853
rect 11835 7788 11836 7852
rect 11900 7788 11901 7852
rect 11835 7787 11901 7788
rect 11099 4996 11165 4997
rect 11099 4932 11100 4996
rect 11164 4932 11165 4996
rect 11099 4931 11165 4932
rect 11838 3501 11898 7787
rect 12571 6900 12637 6901
rect 12571 6836 12572 6900
rect 12636 6836 12637 6900
rect 12571 6835 12637 6836
rect 12574 6085 12634 6835
rect 12755 6628 12821 6629
rect 12755 6564 12756 6628
rect 12820 6564 12821 6628
rect 12755 6563 12821 6564
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12571 5948 12637 5949
rect 12571 5884 12572 5948
rect 12636 5884 12637 5948
rect 12571 5883 12637 5884
rect 11835 3500 11901 3501
rect 11835 3436 11836 3500
rect 11900 3436 11901 3500
rect 11835 3435 11901 3436
rect 12574 2957 12634 5883
rect 12758 5813 12818 6563
rect 13307 6356 13373 6357
rect 13307 6292 13308 6356
rect 13372 6292 13373 6356
rect 13307 6291 13373 6292
rect 12755 5812 12821 5813
rect 12755 5748 12756 5812
rect 12820 5748 12821 5812
rect 12755 5747 12821 5748
rect 13123 4996 13189 4997
rect 13123 4932 13124 4996
rect 13188 4932 13189 4996
rect 13123 4931 13189 4932
rect 12571 2956 12637 2957
rect 12571 2892 12572 2956
rect 12636 2892 12637 2956
rect 12571 2891 12637 2892
rect 11651 2820 11717 2821
rect 11651 2756 11652 2820
rect 11716 2756 11717 2820
rect 11651 2755 11717 2756
rect 10731 2004 10797 2005
rect 10731 1940 10732 2004
rect 10796 1940 10797 2004
rect 10731 1939 10797 1940
rect 11654 1189 11714 2755
rect 13126 2685 13186 4931
rect 13310 2957 13370 6291
rect 13678 5949 13738 8331
rect 13944 8192 14264 11250
rect 13944 8128 13952 8192
rect 14016 8128 14032 8192
rect 14096 8128 14112 8192
rect 14176 8128 14192 8192
rect 14256 8128 14264 8192
rect 13944 7104 14264 8128
rect 15004 8736 15324 11250
rect 16619 9756 16685 9757
rect 16619 9692 16620 9756
rect 16684 9692 16685 9756
rect 16619 9691 16685 9692
rect 15004 8672 15012 8736
rect 15076 8672 15092 8736
rect 15156 8672 15172 8736
rect 15236 8672 15252 8736
rect 15316 8672 15324 8736
rect 14779 8124 14845 8125
rect 14779 8060 14780 8124
rect 14844 8060 14845 8124
rect 14779 8059 14845 8060
rect 14411 7716 14477 7717
rect 14411 7652 14412 7716
rect 14476 7652 14477 7716
rect 14411 7651 14477 7652
rect 13944 7040 13952 7104
rect 14016 7040 14032 7104
rect 14096 7040 14112 7104
rect 14176 7040 14192 7104
rect 14256 7040 14264 7104
rect 13944 6016 14264 7040
rect 13944 5952 13952 6016
rect 14016 5952 14032 6016
rect 14096 5952 14112 6016
rect 14176 5952 14192 6016
rect 14256 5952 14264 6016
rect 13675 5948 13741 5949
rect 13675 5884 13676 5948
rect 13740 5884 13741 5948
rect 13675 5883 13741 5884
rect 13491 5812 13557 5813
rect 13491 5748 13492 5812
rect 13556 5748 13557 5812
rect 13491 5747 13557 5748
rect 13494 3773 13554 5747
rect 13944 4928 14264 5952
rect 13944 4864 13952 4928
rect 14016 4864 14032 4928
rect 14096 4864 14112 4928
rect 14176 4864 14192 4928
rect 14256 4864 14264 4928
rect 13675 4860 13741 4861
rect 13675 4796 13676 4860
rect 13740 4796 13741 4860
rect 13675 4795 13741 4796
rect 13491 3772 13557 3773
rect 13491 3708 13492 3772
rect 13556 3708 13557 3772
rect 13491 3707 13557 3708
rect 13307 2956 13373 2957
rect 13307 2892 13308 2956
rect 13372 2892 13373 2956
rect 13307 2891 13373 2892
rect 13123 2684 13189 2685
rect 13123 2620 13124 2684
rect 13188 2620 13189 2684
rect 13123 2619 13189 2620
rect 11651 1188 11717 1189
rect 11651 1124 11652 1188
rect 11716 1124 11717 1188
rect 11651 1123 11717 1124
rect 13678 373 13738 4795
rect 13944 3840 14264 4864
rect 14414 4861 14474 7651
rect 14595 6356 14661 6357
rect 14595 6292 14596 6356
rect 14660 6292 14661 6356
rect 14595 6291 14661 6292
rect 14411 4860 14477 4861
rect 14411 4796 14412 4860
rect 14476 4796 14477 4860
rect 14411 4795 14477 4796
rect 14598 4045 14658 6291
rect 14595 4044 14661 4045
rect 14595 3980 14596 4044
rect 14660 3980 14661 4044
rect 14595 3979 14661 3980
rect 13944 3776 13952 3840
rect 14016 3776 14032 3840
rect 14096 3776 14112 3840
rect 14176 3776 14192 3840
rect 14256 3776 14264 3840
rect 13944 2752 14264 3776
rect 14782 3773 14842 8059
rect 15004 7648 15324 8672
rect 15004 7584 15012 7648
rect 15076 7584 15092 7648
rect 15156 7584 15172 7648
rect 15236 7584 15252 7648
rect 15316 7584 15324 7648
rect 15004 6560 15324 7584
rect 16435 7036 16501 7037
rect 16435 6972 16436 7036
rect 16500 6972 16501 7036
rect 16435 6971 16501 6972
rect 15004 6496 15012 6560
rect 15076 6496 15092 6560
rect 15156 6496 15172 6560
rect 15236 6496 15252 6560
rect 15316 6496 15324 6560
rect 15004 5472 15324 6496
rect 15004 5408 15012 5472
rect 15076 5408 15092 5472
rect 15156 5408 15172 5472
rect 15236 5408 15252 5472
rect 15316 5408 15324 5472
rect 15004 4384 15324 5408
rect 15004 4320 15012 4384
rect 15076 4320 15092 4384
rect 15156 4320 15172 4384
rect 15236 4320 15252 4384
rect 15316 4320 15324 4384
rect 14779 3772 14845 3773
rect 14779 3708 14780 3772
rect 14844 3708 14845 3772
rect 14779 3707 14845 3708
rect 13944 2688 13952 2752
rect 14016 2688 14032 2752
rect 14096 2688 14112 2752
rect 14176 2688 14192 2752
rect 14256 2688 14264 2752
rect 13675 372 13741 373
rect 13675 308 13676 372
rect 13740 308 13741 372
rect 13675 307 13741 308
rect 13944 0 14264 2688
rect 15004 3296 15324 4320
rect 15004 3232 15012 3296
rect 15076 3232 15092 3296
rect 15156 3232 15172 3296
rect 15236 3232 15252 3296
rect 15316 3232 15324 3296
rect 15004 2208 15324 3232
rect 15004 2144 15012 2208
rect 15076 2144 15092 2208
rect 15156 2144 15172 2208
rect 15236 2144 15252 2208
rect 15316 2144 15324 2208
rect 15004 0 15324 2144
rect 16438 1050 16498 6971
rect 16622 4997 16682 9691
rect 19944 8192 20264 11250
rect 19944 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20192 8192
rect 20256 8128 20264 8192
rect 19944 7104 20264 8128
rect 19944 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20192 7104
rect 20256 7040 20264 7104
rect 19944 6016 20264 7040
rect 21004 8736 21324 11250
rect 21004 8672 21012 8736
rect 21076 8672 21092 8736
rect 21156 8672 21172 8736
rect 21236 8672 21252 8736
rect 21316 8672 21324 8736
rect 21004 7648 21324 8672
rect 22507 8668 22573 8669
rect 22507 8604 22508 8668
rect 22572 8604 22573 8668
rect 22507 8603 22573 8604
rect 21587 7716 21653 7717
rect 21587 7652 21588 7716
rect 21652 7652 21653 7716
rect 21587 7651 21653 7652
rect 21004 7584 21012 7648
rect 21076 7584 21092 7648
rect 21156 7584 21172 7648
rect 21236 7584 21252 7648
rect 21316 7584 21324 7648
rect 20851 7036 20917 7037
rect 20851 6972 20852 7036
rect 20916 6972 20917 7036
rect 20851 6971 20917 6972
rect 19944 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20192 6016
rect 20256 5952 20264 6016
rect 16619 4996 16685 4997
rect 16619 4932 16620 4996
rect 16684 4932 16685 4996
rect 16619 4931 16685 4932
rect 19944 4928 20264 5952
rect 19944 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20192 4928
rect 20256 4864 20264 4928
rect 18827 4588 18893 4589
rect 18827 4524 18828 4588
rect 18892 4524 18893 4588
rect 18827 4523 18893 4524
rect 17907 4180 17973 4181
rect 17907 4116 17908 4180
rect 17972 4116 17973 4180
rect 17907 4115 17973 4116
rect 17910 1325 17970 4115
rect 18830 2685 18890 4523
rect 19195 4316 19261 4317
rect 19195 4252 19196 4316
rect 19260 4252 19261 4316
rect 19195 4251 19261 4252
rect 18827 2684 18893 2685
rect 18827 2620 18828 2684
rect 18892 2620 18893 2684
rect 18827 2619 18893 2620
rect 19198 2549 19258 4251
rect 19944 3840 20264 4864
rect 19944 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20192 3840
rect 20256 3776 20264 3840
rect 19944 2752 20264 3776
rect 19944 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20192 2752
rect 20256 2688 20264 2752
rect 19195 2548 19261 2549
rect 19195 2484 19196 2548
rect 19260 2484 19261 2548
rect 19195 2483 19261 2484
rect 17907 1324 17973 1325
rect 17907 1260 17908 1324
rect 17972 1260 17973 1324
rect 17907 1259 17973 1260
rect 16619 1052 16685 1053
rect 16619 1050 16620 1052
rect 16438 990 16620 1050
rect 16619 988 16620 990
rect 16684 988 16685 1052
rect 16619 987 16685 988
rect 19944 0 20264 2688
rect 20854 2141 20914 6971
rect 21004 6560 21324 7584
rect 21590 6901 21650 7651
rect 21587 6900 21653 6901
rect 21587 6836 21588 6900
rect 21652 6836 21653 6900
rect 21587 6835 21653 6836
rect 21004 6496 21012 6560
rect 21076 6496 21092 6560
rect 21156 6496 21172 6560
rect 21236 6496 21252 6560
rect 21316 6496 21324 6560
rect 21004 5472 21324 6496
rect 22139 5948 22205 5949
rect 22139 5884 22140 5948
rect 22204 5884 22205 5948
rect 22139 5883 22205 5884
rect 21004 5408 21012 5472
rect 21076 5408 21092 5472
rect 21156 5408 21172 5472
rect 21236 5408 21252 5472
rect 21316 5408 21324 5472
rect 21004 4384 21324 5408
rect 21004 4320 21012 4384
rect 21076 4320 21092 4384
rect 21156 4320 21172 4384
rect 21236 4320 21252 4384
rect 21316 4320 21324 4384
rect 21004 3296 21324 4320
rect 21004 3232 21012 3296
rect 21076 3232 21092 3296
rect 21156 3232 21172 3296
rect 21236 3232 21252 3296
rect 21316 3232 21324 3296
rect 21004 2208 21324 3232
rect 21004 2144 21012 2208
rect 21076 2144 21092 2208
rect 21156 2144 21172 2208
rect 21236 2144 21252 2208
rect 21316 2144 21324 2208
rect 20851 2140 20917 2141
rect 20851 2076 20852 2140
rect 20916 2076 20917 2140
rect 20851 2075 20917 2076
rect 21004 0 21324 2144
rect 22142 645 22202 5883
rect 22510 1597 22570 8603
rect 25944 8192 26264 11250
rect 25944 8128 25952 8192
rect 26016 8128 26032 8192
rect 26096 8128 26112 8192
rect 26176 8128 26192 8192
rect 26256 8128 26264 8192
rect 25944 7104 26264 8128
rect 25944 7040 25952 7104
rect 26016 7040 26032 7104
rect 26096 7040 26112 7104
rect 26176 7040 26192 7104
rect 26256 7040 26264 7104
rect 25635 7036 25701 7037
rect 25635 6972 25636 7036
rect 25700 6972 25701 7036
rect 25635 6971 25701 6972
rect 24163 6492 24229 6493
rect 24163 6428 24164 6492
rect 24228 6428 24229 6492
rect 24163 6427 24229 6428
rect 24166 2685 24226 6427
rect 25267 5948 25333 5949
rect 25267 5884 25268 5948
rect 25332 5884 25333 5948
rect 25267 5883 25333 5884
rect 24163 2684 24229 2685
rect 24163 2620 24164 2684
rect 24228 2620 24229 2684
rect 24163 2619 24229 2620
rect 25270 2141 25330 5883
rect 25638 2413 25698 6971
rect 25944 6016 26264 7040
rect 25944 5952 25952 6016
rect 26016 5952 26032 6016
rect 26096 5952 26112 6016
rect 26176 5952 26192 6016
rect 26256 5952 26264 6016
rect 25944 4928 26264 5952
rect 25944 4864 25952 4928
rect 26016 4864 26032 4928
rect 26096 4864 26112 4928
rect 26176 4864 26192 4928
rect 26256 4864 26264 4928
rect 25944 3840 26264 4864
rect 25944 3776 25952 3840
rect 26016 3776 26032 3840
rect 26096 3776 26112 3840
rect 26176 3776 26192 3840
rect 26256 3776 26264 3840
rect 25944 2752 26264 3776
rect 25944 2688 25952 2752
rect 26016 2688 26032 2752
rect 26096 2688 26112 2752
rect 26176 2688 26192 2752
rect 26256 2688 26264 2752
rect 25635 2412 25701 2413
rect 25635 2348 25636 2412
rect 25700 2348 25701 2412
rect 25635 2347 25701 2348
rect 25267 2140 25333 2141
rect 25267 2076 25268 2140
rect 25332 2076 25333 2140
rect 25267 2075 25333 2076
rect 22507 1596 22573 1597
rect 22507 1532 22508 1596
rect 22572 1532 22573 1596
rect 22507 1531 22573 1532
rect 22139 644 22205 645
rect 22139 580 22140 644
rect 22204 580 22205 644
rect 22139 579 22205 580
rect 25944 0 26264 2688
rect 27004 8736 27324 11250
rect 30419 10164 30485 10165
rect 30419 10100 30420 10164
rect 30484 10100 30485 10164
rect 30419 10099 30485 10100
rect 27004 8672 27012 8736
rect 27076 8672 27092 8736
rect 27156 8672 27172 8736
rect 27236 8672 27252 8736
rect 27316 8672 27324 8736
rect 27004 7648 27324 8672
rect 27004 7584 27012 7648
rect 27076 7584 27092 7648
rect 27156 7584 27172 7648
rect 27236 7584 27252 7648
rect 27316 7584 27324 7648
rect 27004 6560 27324 7584
rect 27004 6496 27012 6560
rect 27076 6496 27092 6560
rect 27156 6496 27172 6560
rect 27236 6496 27252 6560
rect 27316 6496 27324 6560
rect 27004 5472 27324 6496
rect 27004 5408 27012 5472
rect 27076 5408 27092 5472
rect 27156 5408 27172 5472
rect 27236 5408 27252 5472
rect 27316 5408 27324 5472
rect 27004 4384 27324 5408
rect 27659 5404 27725 5405
rect 27659 5340 27660 5404
rect 27724 5340 27725 5404
rect 27659 5339 27725 5340
rect 27004 4320 27012 4384
rect 27076 4320 27092 4384
rect 27156 4320 27172 4384
rect 27236 4320 27252 4384
rect 27316 4320 27324 4384
rect 27004 3296 27324 4320
rect 27475 4316 27541 4317
rect 27475 4252 27476 4316
rect 27540 4252 27541 4316
rect 27475 4251 27541 4252
rect 27004 3232 27012 3296
rect 27076 3232 27092 3296
rect 27156 3232 27172 3296
rect 27236 3232 27252 3296
rect 27316 3232 27324 3296
rect 27004 2208 27324 3232
rect 27004 2144 27012 2208
rect 27076 2144 27092 2208
rect 27156 2144 27172 2208
rect 27236 2144 27252 2208
rect 27316 2144 27324 2208
rect 27004 0 27324 2144
rect 27478 1325 27538 4251
rect 27662 3637 27722 5339
rect 30422 4045 30482 10099
rect 31944 8192 32264 11250
rect 31944 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32264 8192
rect 31944 7104 32264 8128
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 30419 4044 30485 4045
rect 30419 3980 30420 4044
rect 30484 3980 30485 4044
rect 30419 3979 30485 3980
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 27659 3636 27725 3637
rect 27659 3572 27660 3636
rect 27724 3572 27725 3636
rect 27659 3571 27725 3572
rect 31944 2752 32264 3776
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 27475 1324 27541 1325
rect 27475 1260 27476 1324
rect 27540 1260 27541 1324
rect 27475 1259 27541 1260
rect 31944 0 32264 2688
rect 33004 8736 33324 11250
rect 33004 8672 33012 8736
rect 33076 8672 33092 8736
rect 33156 8672 33172 8736
rect 33236 8672 33252 8736
rect 33316 8672 33324 8736
rect 33004 7648 33324 8672
rect 33004 7584 33012 7648
rect 33076 7584 33092 7648
rect 33156 7584 33172 7648
rect 33236 7584 33252 7648
rect 33316 7584 33324 7648
rect 33004 6560 33324 7584
rect 33004 6496 33012 6560
rect 33076 6496 33092 6560
rect 33156 6496 33172 6560
rect 33236 6496 33252 6560
rect 33316 6496 33324 6560
rect 33004 5472 33324 6496
rect 33004 5408 33012 5472
rect 33076 5408 33092 5472
rect 33156 5408 33172 5472
rect 33236 5408 33252 5472
rect 33316 5408 33324 5472
rect 33004 4384 33324 5408
rect 33004 4320 33012 4384
rect 33076 4320 33092 4384
rect 33156 4320 33172 4384
rect 33236 4320 33252 4384
rect 33316 4320 33324 4384
rect 33004 3296 33324 4320
rect 33004 3232 33012 3296
rect 33076 3232 33092 3296
rect 33156 3232 33172 3296
rect 33236 3232 33252 3296
rect 33316 3232 33324 3296
rect 33004 2208 33324 3232
rect 33004 2144 33012 2208
rect 33076 2144 33092 2208
rect 33156 2144 33172 2208
rect 33236 2144 33252 2208
rect 33316 2144 33324 2208
rect 33004 0 33324 2144
rect 37944 8192 38264 11250
rect 37944 8128 37952 8192
rect 38016 8128 38032 8192
rect 38096 8128 38112 8192
rect 38176 8128 38192 8192
rect 38256 8128 38264 8192
rect 37944 7104 38264 8128
rect 37944 7040 37952 7104
rect 38016 7040 38032 7104
rect 38096 7040 38112 7104
rect 38176 7040 38192 7104
rect 38256 7040 38264 7104
rect 37944 6016 38264 7040
rect 37944 5952 37952 6016
rect 38016 5952 38032 6016
rect 38096 5952 38112 6016
rect 38176 5952 38192 6016
rect 38256 5952 38264 6016
rect 37944 4928 38264 5952
rect 37944 4864 37952 4928
rect 38016 4864 38032 4928
rect 38096 4864 38112 4928
rect 38176 4864 38192 4928
rect 38256 4864 38264 4928
rect 37944 3840 38264 4864
rect 37944 3776 37952 3840
rect 38016 3776 38032 3840
rect 38096 3776 38112 3840
rect 38176 3776 38192 3840
rect 38256 3776 38264 3840
rect 37944 2752 38264 3776
rect 37944 2688 37952 2752
rect 38016 2688 38032 2752
rect 38096 2688 38112 2752
rect 38176 2688 38192 2752
rect 38256 2688 38264 2752
rect 37944 0 38264 2688
rect 39004 8736 39324 11250
rect 39004 8672 39012 8736
rect 39076 8672 39092 8736
rect 39156 8672 39172 8736
rect 39236 8672 39252 8736
rect 39316 8672 39324 8736
rect 39004 7648 39324 8672
rect 39004 7584 39012 7648
rect 39076 7584 39092 7648
rect 39156 7584 39172 7648
rect 39236 7584 39252 7648
rect 39316 7584 39324 7648
rect 39004 6560 39324 7584
rect 39004 6496 39012 6560
rect 39076 6496 39092 6560
rect 39156 6496 39172 6560
rect 39236 6496 39252 6560
rect 39316 6496 39324 6560
rect 39004 5472 39324 6496
rect 39004 5408 39012 5472
rect 39076 5408 39092 5472
rect 39156 5408 39172 5472
rect 39236 5408 39252 5472
rect 39316 5408 39324 5472
rect 39004 4384 39324 5408
rect 39004 4320 39012 4384
rect 39076 4320 39092 4384
rect 39156 4320 39172 4384
rect 39236 4320 39252 4384
rect 39316 4320 39324 4384
rect 39004 3296 39324 4320
rect 39004 3232 39012 3296
rect 39076 3232 39092 3296
rect 39156 3232 39172 3296
rect 39236 3232 39252 3296
rect 39316 3232 39324 3296
rect 39004 2208 39324 3232
rect 39004 2144 39012 2208
rect 39076 2144 39092 2208
rect 39156 2144 39172 2208
rect 39236 2144 39252 2208
rect 39316 2144 39324 2208
rect 39004 0 39324 2144
use sky130_fd_sc_hd__mux4_1  _032_
timestamp -3599
transform 1 0 18676 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _033_
timestamp -3599
transform 1 0 3680 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _034_
timestamp -3599
transform 1 0 25760 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _035_
timestamp -3599
transform 1 0 7544 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _036_
timestamp -3599
transform 1 0 17204 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _037_
timestamp -3599
transform 1 0 35512 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _038_
timestamp -3599
transform -1 0 36616 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _039_
timestamp -3599
transform 1 0 22172 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _040_
timestamp -3599
transform -1 0 34224 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _041_
timestamp -3599
transform -1 0 9844 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _042_
timestamp -3599
transform 1 0 7268 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _043_
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _044_
timestamp -3599
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _045_
timestamp -3599
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _046_
timestamp -3599
transform -1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _047_
timestamp -3599
transform -1 0 8648 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _048_
timestamp -3599
transform 1 0 6900 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _049_
timestamp -3599
transform 1 0 5612 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _050_
timestamp -3599
transform -1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _051_
timestamp -3599
transform -1 0 7912 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _052_
timestamp -3599
transform -1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _053_
timestamp -3599
transform -1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _054_
timestamp -3599
transform -1 0 6900 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp -3599
transform -1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp -3599
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _057_
timestamp -3599
transform -1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _059_
timestamp -3599
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  _060_
timestamp -3599
transform 1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _061_
timestamp -3599
transform 1 0 9844 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _062_
timestamp -3599
transform 1 0 12880 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _063_
timestamp -3599
transform 1 0 6900 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _064_
timestamp -3599
transform -1 0 12880 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _065_
timestamp -3599
transform 1 0 9384 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _066_
timestamp -3599
transform 1 0 10120 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp -3599
transform -1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _068_
timestamp -3599
transform 1 0 11776 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _069_
timestamp -3599
transform 1 0 8464 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _070_
timestamp -3599
transform -1 0 10028 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _071_
timestamp -3599
transform 1 0 7360 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _072_
timestamp -3599
transform -1 0 9568 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _073_
timestamp -3599
transform 1 0 9568 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _074_
timestamp -3599
transform 1 0 9292 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _075_
timestamp -3599
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _076_
timestamp -3599
transform -1 0 10948 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _077_
timestamp -3599
transform -1 0 18124 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _078_
timestamp -3599
transform -1 0 5704 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _079_
timestamp -3599
transform 1 0 25944 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _080_
timestamp -3599
transform 1 0 28888 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _081_
timestamp -3599
transform 1 0 28244 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _082_
timestamp -3599
transform 1 0 24840 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _083_
timestamp -3599
transform 1 0 28336 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _084_
timestamp -3599
transform 1 0 29532 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _085_
timestamp -3599
transform 1 0 11500 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _086_
timestamp -3599
transform -1 0 5428 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _087_
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _088_
timestamp -3599
transform -1 0 8280 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _089_
timestamp -3599
transform 1 0 22356 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _090_
timestamp -3599
transform 1 0 26956 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _091_
timestamp -3599
transform -1 0 25300 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _092_
timestamp -3599
transform 1 0 17940 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _093_
timestamp -3599
transform 1 0 31096 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _094_
timestamp -3599
transform 1 0 22816 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _095_
timestamp -3599
transform 1 0 32476 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _096_
timestamp -3599
transform 1 0 31004 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _097_
timestamp -3599
transform 1 0 27508 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _098_
timestamp -3599
transform 1 0 23000 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _099_
timestamp -3599
transform 1 0 29164 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _100_
timestamp -3599
transform 1 0 31372 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _101_
timestamp -3599
transform 1 0 13892 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _102_
timestamp -3599
transform -1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _103_
timestamp -3599
transform 1 0 14996 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _104_
timestamp -3599
transform 1 0 17848 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _105_
timestamp -3599
transform 1 0 20424 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _106_
timestamp -3599
transform 1 0 19412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _107_
timestamp -3599
transform 1 0 20700 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _108_
timestamp -3599
transform 1 0 18124 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _109_
timestamp -3599
transform 1 0 32108 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _110_
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _111_
timestamp -3599
transform 1 0 14628 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _112_
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _113_
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _114_
timestamp -3599
transform 1 0 25576 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _115_
timestamp -3599
transform -1 0 7636 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _116_
timestamp -3599
transform 1 0 19780 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _117_
timestamp -3599
transform 1 0 11868 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _118_
timestamp -3599
transform -1 0 17940 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _119_
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtp_1  _120_
timestamp -3599
transform -1 0 23828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _121_
timestamp -3599
transform -1 0 25208 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _122_
timestamp -3599
transform -1 0 23736 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _123_
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _124_
timestamp -3599
transform -1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _125_
timestamp -3599
transform -1 0 25852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _126_
timestamp -3599
transform -1 0 26312 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _127_
timestamp -3599
transform -1 0 35512 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _128_
timestamp -3599
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _129_
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _130_
timestamp -3599
transform 1 0 34684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _131_
timestamp -3599
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _132_
timestamp -3599
transform 1 0 16928 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _133_
timestamp -3599
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _134_
timestamp -3599
transform 1 0 7268 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _135_
timestamp -3599
transform 1 0 7176 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _136_
timestamp -3599
transform -1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _137_
timestamp -3599
transform 1 0 25208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _138_
timestamp -3599
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _139_
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _140_
timestamp -3599
transform 1 0 17572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _141_
timestamp -3599
transform 1 0 17940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _142_
timestamp -3599
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _143_
timestamp -3599
transform 1 0 12420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _144_
timestamp -3599
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _145_
timestamp -3599
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _146_
timestamp -3599
transform 1 0 10764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _147_
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _148_
timestamp -3599
transform -1 0 31096 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _149_
timestamp -3599
transform -1 0 31372 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _150_
timestamp -3599
transform 1 0 4968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _151_
timestamp -3599
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _152_
timestamp -3599
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _153_
timestamp -3599
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _154_
timestamp -3599
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _155_
timestamp -3599
transform 1 0 2576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _156_
timestamp -3599
transform -1 0 22908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _157_
timestamp -3599
transform -1 0 25576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _158_
timestamp -3599
transform -1 0 16192 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _159_
timestamp -3599
transform -1 0 26312 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _160_
timestamp -3599
transform 1 0 12788 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _161_
timestamp -3599
transform 1 0 12328 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _162_
timestamp -3599
transform -1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _163_
timestamp -3599
transform -1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _164_
timestamp -3599
transform 1 0 16836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _165_
timestamp -3599
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _166_
timestamp -3599
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _167_
timestamp -3599
transform 1 0 20240 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _168_
timestamp -3599
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _169_
timestamp -3599
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _170_
timestamp -3599
transform 1 0 20056 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _171_
timestamp -3599
transform 1 0 20056 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _172_
timestamp -3599
transform -1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _173_
timestamp -3599
transform 1 0 16744 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _174_
timestamp -3599
transform -1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _175_
timestamp -3599
transform 1 0 14352 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _176_
timestamp -3599
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _177_
timestamp -3599
transform 1 0 14352 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _178_
timestamp -3599
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _179_
timestamp -3599
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _180_
timestamp -3599
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _181_
timestamp -3599
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _182_
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _183_
timestamp -3599
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _184_
timestamp -3599
transform 1 0 22724 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _185_
timestamp -3599
transform 1 0 22724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _186_
timestamp -3599
transform 1 0 27140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _187_
timestamp -3599
transform 1 0 27140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _188_
timestamp -3599
transform 1 0 29900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _189_
timestamp -3599
transform 1 0 30820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _190_
timestamp -3599
transform 1 0 33028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _191_
timestamp -3599
transform 1 0 31924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _192_
timestamp -3599
transform -1 0 24196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _193_
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _194_
timestamp -3599
transform 1 0 30912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _195_
timestamp -3599
transform 1 0 30912 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _196_
timestamp -3599
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _197_
timestamp -3599
transform 1 0 17296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _198_
timestamp -3599
transform 1 0 22264 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _199_
timestamp -3599
transform 1 0 22448 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _200_
timestamp -3599
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _201_
timestamp -3599
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _202_
timestamp -3599
transform 1 0 21896 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _203_
timestamp -3599
transform 1 0 23000 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _204_
timestamp -3599
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _205_
timestamp -3599
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _206_
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _207_
timestamp -3599
transform 1 0 13432 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _208_
timestamp -3599
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _209_
timestamp -3599
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _210_
timestamp -3599
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _211_
timestamp -3599
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _212_
timestamp -3599
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _213_
timestamp -3599
transform 1 0 28888 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _214_
timestamp -3599
transform 1 0 27876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _215_
timestamp -3599
transform 1 0 27784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _216_
timestamp -3599
transform 1 0 24748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _217_
timestamp -3599
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _218_
timestamp -3599
transform 1 0 27416 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _219_
timestamp -3599
transform 1 0 28244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _220_
timestamp -3599
transform 1 0 28336 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _221_
timestamp -3599
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _222_
timestamp -3599
transform -1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _223_
timestamp -3599
transform 1 0 26312 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _224_
timestamp -3599
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _225_
timestamp -3599
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _226_
timestamp -3599
transform -1 0 34408 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _227_
timestamp -3599
transform -1 0 34408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _228_
timestamp -3599
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _229_
timestamp -3599
transform 1 0 7360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _230_
timestamp -3599
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _231_
timestamp -3599
transform -1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _232_
timestamp -3599
transform 1 0 7728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _233_
timestamp -3599
transform 1 0 9200 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _234_
timestamp -3599
transform -1 0 7544 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _235_
timestamp -3599
transform 1 0 5704 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _236_
timestamp -3599
transform 1 0 7912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _237_
timestamp -3599
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _238_
timestamp -3599
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _239_
timestamp -3599
transform 1 0 5060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _240_
timestamp -3599
transform -1 0 6256 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _241_
timestamp -3599
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp -3599
transform -1 0 34408 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp -3599
transform -1 0 34132 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _244_
timestamp -3599
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _245_
timestamp -3599
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp -3599
transform -1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp -3599
transform -1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _248_
timestamp -3599
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _249_
timestamp -3599
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _250_
timestamp -3599
transform 1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _251_
timestamp -3599
transform 1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _252_
timestamp -3599
transform 1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _253_
timestamp -3599
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp -3599
transform -1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp -3599
transform -1 0 36616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp -3599
transform -1 0 32016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _257_
timestamp -3599
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _258_
timestamp -3599
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _259_
timestamp -3599
transform 1 0 3864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp -3599
transform -1 0 36800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp -3599
transform -1 0 36248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _262_
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _263_
timestamp -3599
transform 1 0 9752 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _264_
timestamp -3599
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _265_
timestamp -3599
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _266_
timestamp -3599
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _267_
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _268_
timestamp -3599
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _269_
timestamp -3599
transform 1 0 2852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _270_
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _271_
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _272_
timestamp -3599
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _273_
timestamp -3599
transform 1 0 5520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _274_
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _275_
timestamp -3599
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp -3599
transform -1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp -3599
transform -1 0 12880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _279_
timestamp -3599
transform -1 0 36340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _280_
timestamp -3599
transform -1 0 37352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _281_
timestamp -3599
transform -1 0 37076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _282_
timestamp -3599
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _283_
timestamp -3599
transform -1 0 37904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _284_
timestamp -3599
transform -1 0 37076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp -3599
transform 1 0 36248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp -3599
transform 1 0 38548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp -3599
transform 1 0 38180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _288_
timestamp -3599
transform -1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp -3599
transform 1 0 38456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp -3599
transform 1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp -3599
transform 1 0 38364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp -3599
transform 1 0 38456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp -3599
transform 1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp -3599
transform -1 0 37720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp -3599
transform -1 0 38180 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _296_
timestamp -3599
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp -3599
transform 1 0 22264 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _298_
timestamp -3599
transform -1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _299_
timestamp -3599
transform -1 0 35512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp -3599
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _301_
timestamp -3599
transform 1 0 9476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp -3599
transform 1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _303_
timestamp -3599
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp -3599
transform -1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp -3599
transform -1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp -3599
transform -1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _307_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _308_
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _309_
timestamp -3599
transform 1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _310_
timestamp -3599
transform 1 0 27140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _311_
timestamp -3599
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp -3599
transform -1 0 24288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _313_
timestamp -3599
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp -3599
transform -1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _315_
timestamp -3599
transform -1 0 33580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp -3599
transform -1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _317_
timestamp -3599
transform -1 0 22448 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp -3599
transform -1 0 21712 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp -3599
transform -1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _320_
timestamp -3599
transform -1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _321_
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _322_
timestamp -3599
transform -1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _323_
timestamp -3599
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _324_
timestamp -3599
transform 1 0 32384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _325_
timestamp -3599
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _326_
timestamp -3599
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp -3599
transform -1 0 29808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _328_
timestamp -3599
transform 1 0 34408 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _329_
timestamp -3599
transform 1 0 35788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _330_
timestamp -3599
transform -1 0 26864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp -3599
transform -1 0 33304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _332_
timestamp -3599
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp -3599
transform -1 0 24288 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _334_
timestamp -3599
transform -1 0 29440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp -3599
transform -1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _336_
timestamp -3599
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _337_
timestamp -3599
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _338_
timestamp -3599
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _339_
timestamp -3599
transform 1 0 13432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _340_
timestamp -3599
transform -1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _341_
timestamp -3599
transform -1 0 32384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _342_
timestamp -3599
transform -1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp -3599
transform -1 0 30176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _344_
timestamp -3599
transform -1 0 34592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _345_
timestamp -3599
transform -1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _346_
timestamp -3599
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _347_
timestamp -3599
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _348_
timestamp -3599
transform -1 0 34500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 39192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp -3599
transform -1 0 38824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp -3599
transform -1 0 38640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp -3599
transform 1 0 36616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp -3599
transform -1 0 38824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp -3599
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp -3599
transform -1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp -3599
transform -1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp -3599
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp -3599
transform -1 0 31096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp -3599
transform 1 0 32292 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp -3599
transform -1 0 33396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp -3599
transform 1 0 22908 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK
timestamp -3599
transform 1 0 34684 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp -3599
transform 1 0 34684 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp -3599
transform -1 0 35972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp -3599
transform 1 0 35144 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp -3599
transform -1 0 34592 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp -3599
transform -1 0 19136 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp -3599
transform -1 0 13984 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp -3599
transform 1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp -3599
transform -1 0 13984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp -3599
transform -1 0 25024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp -3599
transform 1 0 16836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout57
timestamp -3599
transform -1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout58
timestamp -3599
transform -1 0 25944 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp -3599
transform -1 0 29348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp -3599
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp -3599
transform 1 0 16928 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp -3599
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp -3599
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp -3599
transform -1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout65
timestamp -3599
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout66
timestamp -3599
transform -1 0 21528 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp -3599
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp -3599
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp -3599
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34
timestamp -3599
transform 1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp -3599
transform 1 0 10304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp -3599
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp -3599
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp -3599
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp -3599
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_353
timestamp -3599
transform 1 0 33580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp -3599
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp -3599
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp -3599
transform 1 0 37628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_11
timestamp -3599
transform 1 0 2116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_67
timestamp -3599
transform 1 0 7268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_235
timestamp -3599
transform 1 0 22724 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp -3599
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp -3599
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp -3599
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp -3599
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_33
timestamp -3599
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp -3599
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp -3599
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp -3599
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_218
timestamp -3599
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp -3599
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp -3599
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_266
timestamp -3599
transform 1 0 25576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp -3599
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_369
timestamp -3599
transform 1 0 35052 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_390
timestamp 1636964856
transform 1 0 36984 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_402
timestamp -3599
transform 1 0 38088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_409
timestamp -3599
transform 1 0 38732 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp -3599
transform 1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp -3599
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -3599
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_133
timestamp -3599
transform 1 0 13340 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp -3599
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_259
timestamp -3599
transform 1 0 24932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp -3599
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_345
timestamp -3599
transform 1 0 32844 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp -3599
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636964856
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_405
timestamp -3599
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_409
timestamp -3599
transform 1 0 38732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_24
timestamp -3599
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp -3599
transform 1 0 6808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_97
timestamp -3599
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_131
timestamp -3599
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp -3599
transform 1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_218
timestamp -3599
transform 1 0 21160 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp -3599
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp -3599
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp -3599
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp -3599
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp -3599
transform 1 0 29900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_326
timestamp -3599
transform 1 0 31096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp -3599
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp -3599
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_391
timestamp 1636964856
transform 1 0 37076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_403
timestamp -3599
transform 1 0 38180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_409
timestamp -3599
transform 1 0 38732 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp -3599
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp -3599
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp -3599
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_228
timestamp -3599
transform 1 0 22080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_233
timestamp -3599
transform 1 0 22540 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_247
timestamp -3599
transform 1 0 23828 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp -3599
transform 1 0 24840 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp -3599
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_286
timestamp -3599
transform 1 0 27416 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp -3599
transform 1 0 29992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_321
timestamp -3599
transform 1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp -3599
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_382
timestamp -3599
transform 1 0 36248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp -3599
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636964856
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_405
timestamp -3599
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_409
timestamp -3599
transform 1 0 38732 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp -3599
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_41
timestamp -3599
transform 1 0 4876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp -3599
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp -3599
transform 1 0 19596 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_224
timestamp -3599
transform 1 0 21712 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_230
timestamp -3599
transform 1 0 22264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp -3599
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_333
timestamp -3599
transform 1 0 31740 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_343
timestamp -3599
transform 1 0 32660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_388
timestamp 1636964856
transform 1 0 36800 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_400
timestamp -3599
transform 1 0 37904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_404
timestamp -3599
transform 1 0 38272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_408
timestamp -3599
transform 1 0 38640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp -3599
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_116
timestamp -3599
transform 1 0 11776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp -3599
transform 1 0 18032 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp -3599
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_225
timestamp -3599
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_274
timestamp -3599
transform 1 0 26312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_329
timestamp -3599
transform 1 0 31372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp -3599
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_383
timestamp -3599
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp -3599
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp -3599
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_401
timestamp -3599
transform 1 0 37996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp -3599
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp -3599
transform 1 0 7636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp -3599
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_168
timestamp -3599
transform 1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp -3599
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_200
timestamp -3599
transform 1 0 19504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_204
timestamp -3599
transform 1 0 19872 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_209
timestamp -3599
transform 1 0 20332 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_234
timestamp -3599
transform 1 0 22632 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_247
timestamp -3599
transform 1 0 23828 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp -3599
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp -3599
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_261
timestamp -3599
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_298
timestamp -3599
transform 1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp -3599
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_330
timestamp -3599
transform 1 0 31464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_334
timestamp -3599
transform 1 0 31832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp -3599
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_380
timestamp 1636964856
transform 1 0 36064 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_392
timestamp -3599
transform 1 0 37168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_409
timestamp -3599
transform 1 0 38732 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_43
timestamp -3599
transform 1 0 5060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_47
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp -3599
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_98
timestamp -3599
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_125
timestamp -3599
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp -3599
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp -3599
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_204
timestamp -3599
transform 1 0 19872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp -3599
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp -3599
transform 1 0 22172 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp -3599
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp -3599
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp -3599
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_316
timestamp -3599
transform 1 0 30176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_320
timestamp -3599
transform 1 0 30544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_358
timestamp -3599
transform 1 0 34040 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_374
timestamp 1636964856
transform 1 0 35512 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_386
timestamp -3599
transform 1 0 36616 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_393
timestamp -3599
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_400
timestamp -3599
transform 1 0 37904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_410
timestamp -3599
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_23
timestamp -3599
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp -3599
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_58
timestamp -3599
transform 1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_79
timestamp -3599
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp -3599
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_147
timestamp -3599
transform 1 0 14628 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp -3599
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp -3599
transform 1 0 19688 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_210
timestamp -3599
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_246
timestamp -3599
transform 1 0 23736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp -3599
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_282
timestamp -3599
transform 1 0 27048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_312
timestamp -3599
transform 1 0 29808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_316
timestamp -3599
transform 1 0 30176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_324
timestamp -3599
transform 1 0 30912 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp -3599
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp -3599
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_377
timestamp -3599
transform 1 0 35788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_381
timestamp -3599
transform 1 0 36156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_385
timestamp -3599
transform 1 0 36524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_394
timestamp -3599
transform 1 0 37352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_17
timestamp -3599
transform 1 0 2668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp -3599
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp -3599
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp -3599
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp -3599
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp -3599
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp -3599
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp -3599
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp -3599
transform 1 0 9844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_119
timestamp -3599
transform 1 0 12052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_123
timestamp -3599
transform 1 0 12420 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_145
timestamp -3599
transform 1 0 14444 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_155
timestamp -3599
transform 1 0 15364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp -3599
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -3599
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_172
timestamp -3599
transform 1 0 16928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_192
timestamp -3599
transform 1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp -3599
transform 1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_203
timestamp -3599
transform 1 0 19780 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_207
timestamp -3599
transform 1 0 20148 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_269
timestamp -3599
transform 1 0 25852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp -3599
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp -3599
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp -3599
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp -3599
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_317
timestamp -3599
transform 1 0 30268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_323
timestamp -3599
transform 1 0 30820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_341
timestamp -3599
transform 1 0 32476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_347
timestamp -3599
transform 1 0 33028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_359
timestamp -3599
transform 1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_363
timestamp -3599
transform 1 0 34500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_365
timestamp -3599
transform 1 0 34684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_371
timestamp -3599
transform 1 0 35236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_383
timestamp -3599
transform 1 0 36340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_397
timestamp -3599
transform 1 0 37628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input1
timestamp -3599
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp -3599
transform 1 0 5060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp -3599
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp -3599
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp -3599
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp -3599
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp -3599
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp -3599
transform 1 0 2116 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp -3599
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -3599
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -3599
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp -3599
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp -3599
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp -3599
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp -3599
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp -3599
transform 1 0 2852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp -3599
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp -3599
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp -3599
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp -3599
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp -3599
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp -3599
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp -3599
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp -3599
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp -3599
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp -3599
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input37
timestamp -3599
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp -3599
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp -3599
transform 1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input40
timestamp -3599
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp -3599
transform 1 0 3772 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp -3599
transform 1 0 4968 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp -3599
transform -1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp -3599
transform 1 0 7912 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input45
timestamp -3599
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp -3599
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp -3599
transform 1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp -3599
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp -3599
transform 1 0 2668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp -3599
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp -3599
transform 1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input53
timestamp -3599
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp -3599
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp -3599
transform 1 0 11592 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input57
timestamp -3599
transform 1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp -3599
transform 1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp -3599
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp -3599
transform 1 0 12328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp -3599
transform -1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp -3599
transform 1 0 7360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp -3599
transform 1 0 9384 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp -3599
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp -3599
transform 1 0 12420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp -3599
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp -3599
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp -3599
transform -1 0 11408 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input70
timestamp -3599
transform 1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp -3599
transform -1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp -3599
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp -3599
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp -3599
transform 1 0 21804 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp -3599
transform -1 0 15456 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input77
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input78
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp -3599
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp -3599
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp -3599
transform -1 0 13984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input82
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp -3599
transform -1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp -3599
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp -3599
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp -3599
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output87
timestamp -3599
transform -1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp -3599
transform -1 0 4876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp -3599
transform -1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp -3599
transform -1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp -3599
transform -1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp -3599
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp -3599
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp -3599
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp -3599
transform -1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp -3599
transform -1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp -3599
transform -1 0 15364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp -3599
transform -1 0 16468 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp -3599
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp -3599
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp -3599
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp -3599
transform 1 0 39192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp -3599
transform 1 0 38824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp -3599
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp -3599
transform 1 0 38824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp -3599
transform 1 0 39192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp -3599
transform 1 0 38824 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp -3599
transform 1 0 39192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp -3599
transform 1 0 39192 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp -3599
transform 1 0 38456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp -3599
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp -3599
transform 1 0 39192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp -3599
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp -3599
transform 1 0 39192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp -3599
transform 1 0 38824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp -3599
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp -3599
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp -3599
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp -3599
transform 1 0 38088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp -3599
transform 1 0 37720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp -3599
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp -3599
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp -3599
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp -3599
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp -3599
transform 1 0 38272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp -3599
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp -3599
transform 1 0 39192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp -3599
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp -3599
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp -3599
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp -3599
transform -1 0 18768 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp -3599
transform -1 0 30268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp -3599
transform -1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp -3599
transform -1 0 32476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp -3599
transform -1 0 33028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp -3599
transform -1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp -3599
transform -1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp -3599
transform -1 0 36340 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp -3599
transform -1 0 37628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp -3599
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp -3599
transform 1 0 39192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp -3599
transform 1 0 19412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp -3599
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp -3599
transform -1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp -3599
transform -1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp -3599
transform -1 0 24288 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp -3599
transform -1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp -3599
transform -1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp -3599
transform -1 0 27508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp -3599
transform -1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp -3599
transform -1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp -3599
transform -1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp -3599
transform -1 0 17204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp -3599
transform -1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp -3599
transform 1 0 16744 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp -3599
transform -1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp -3599
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp -3599
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp -3599
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp -3599
transform 1 0 21436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp -3599
transform -1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp -3599
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp -3599
transform -1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp -3599
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp -3599
transform 1 0 26312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp -3599
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp -3599
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp -3599
transform -1 0 26588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp -3599
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp -3599
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp -3599
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp -3599
transform -1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp -3599
transform -1 0 30636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp -3599
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp -3599
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp -3599
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp -3599
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp -3599
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp -3599
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp -3599
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp -3599
transform 1 0 26128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp -3599
transform -1 0 26864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp -3599
transform -1 0 27876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp -3599
transform 1 0 31464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp -3599
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp -3599
transform 1 0 32476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp -3599
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp -3599
transform 1 0 35328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp -3599
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp -3599
transform 1 0 34684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp -3599
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp -3599
transform 1 0 34592 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp -3599
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp -3599
transform 1 0 31372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp -3599
transform 1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp -3599
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp -3599
transform 1 0 31096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp -3599
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp -3599
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output203
timestamp -3599
transform -1 0 17296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_12
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_13
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 39836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_14
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_15
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 39836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_16
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 39836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_17
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 39836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_18
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 39836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_19
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 39836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_20
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 39836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_21
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 39836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_22
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_23
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 39836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp -3599
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp -3599
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp -3599
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp -3599
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_38
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_40
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_42
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_43
timestamp -3599
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_44
timestamp -3599
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_45
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_46
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_47
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -3599
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -3599
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_56
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_57
timestamp -3599
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_58
timestamp -3599
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_59
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_60
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_61
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp -3599
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp -3599
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp -3599
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp -3599
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp -3599
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp -3599
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -3599
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -3599
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_97
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_98
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_99
timestamp -3599
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_100
timestamp -3599
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_101
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_102
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_103
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_104
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_105
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3599
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3599
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_108
timestamp -3599
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_109
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3599
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3599
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_113
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp -3599
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp -3599
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_117
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp -3599
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp -3599
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp -3599
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp -3599
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 2778 11194 2834 11250 0 FreeSans 224 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 1674 11194 1730 11250 0 FreeSans 224 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 3882 11194 3938 11250 0 FreeSans 224 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 8298 11194 8354 11250 0 FreeSans 224 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal2 s 9402 11194 9458 11250 0 FreeSans 224 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal2 s 10506 11194 10562 11250 0 FreeSans 224 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal2 s 11610 11194 11666 11250 0 FreeSans 224 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal2 s 6090 11194 6146 11250 0 FreeSans 224 0 0 0 B_I_top
port 7 nsew signal output
flabel metal2 s 4986 11194 5042 11250 0 FreeSans 224 0 0 0 B_O_top
port 8 nsew signal input
flabel metal2 s 7194 11194 7250 11250 0 FreeSans 224 0 0 0 B_T_top
port 9 nsew signal output
flabel metal2 s 12714 11194 12770 11250 0 FreeSans 224 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal2 s 13818 11194 13874 11250 0 FreeSans 224 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal2 s 14922 11194 14978 11250 0 FreeSans 224 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal2 s 16026 11194 16082 11250 0 FreeSans 224 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal2 s 17590 0 17646 56 0 FreeSans 224 0 0 0 Ci
port 14 nsew signal input
flabel metal3 s 0 1368 120 1488 0 FreeSans 480 0 0 0 FrameData[0]
port 15 nsew signal input
flabel metal3 s 0 4088 120 4208 0 FreeSans 480 0 0 0 FrameData[10]
port 16 nsew signal input
flabel metal3 s 0 4360 120 4480 0 FreeSans 480 0 0 0 FrameData[11]
port 17 nsew signal input
flabel metal3 s 0 4632 120 4752 0 FreeSans 480 0 0 0 FrameData[12]
port 18 nsew signal input
flabel metal3 s 0 4904 120 5024 0 FreeSans 480 0 0 0 FrameData[13]
port 19 nsew signal input
flabel metal3 s 0 5176 120 5296 0 FreeSans 480 0 0 0 FrameData[14]
port 20 nsew signal input
flabel metal3 s 0 5448 120 5568 0 FreeSans 480 0 0 0 FrameData[15]
port 21 nsew signal input
flabel metal3 s 0 5720 120 5840 0 FreeSans 480 0 0 0 FrameData[16]
port 22 nsew signal input
flabel metal3 s 0 5992 120 6112 0 FreeSans 480 0 0 0 FrameData[17]
port 23 nsew signal input
flabel metal3 s 0 6264 120 6384 0 FreeSans 480 0 0 0 FrameData[18]
port 24 nsew signal input
flabel metal3 s 0 6536 120 6656 0 FreeSans 480 0 0 0 FrameData[19]
port 25 nsew signal input
flabel metal3 s 0 1640 120 1760 0 FreeSans 480 0 0 0 FrameData[1]
port 26 nsew signal input
flabel metal3 s 0 6808 120 6928 0 FreeSans 480 0 0 0 FrameData[20]
port 27 nsew signal input
flabel metal3 s 0 7080 120 7200 0 FreeSans 480 0 0 0 FrameData[21]
port 28 nsew signal input
flabel metal3 s 0 7352 120 7472 0 FreeSans 480 0 0 0 FrameData[22]
port 29 nsew signal input
flabel metal3 s 0 7624 120 7744 0 FreeSans 480 0 0 0 FrameData[23]
port 30 nsew signal input
flabel metal3 s 0 7896 120 8016 0 FreeSans 480 0 0 0 FrameData[24]
port 31 nsew signal input
flabel metal3 s 0 8168 120 8288 0 FreeSans 480 0 0 0 FrameData[25]
port 32 nsew signal input
flabel metal3 s 0 8440 120 8560 0 FreeSans 480 0 0 0 FrameData[26]
port 33 nsew signal input
flabel metal3 s 0 8712 120 8832 0 FreeSans 480 0 0 0 FrameData[27]
port 34 nsew signal input
flabel metal3 s 0 8984 120 9104 0 FreeSans 480 0 0 0 FrameData[28]
port 35 nsew signal input
flabel metal3 s 0 9256 120 9376 0 FreeSans 480 0 0 0 FrameData[29]
port 36 nsew signal input
flabel metal3 s 0 1912 120 2032 0 FreeSans 480 0 0 0 FrameData[2]
port 37 nsew signal input
flabel metal3 s 0 9528 120 9648 0 FreeSans 480 0 0 0 FrameData[30]
port 38 nsew signal input
flabel metal3 s 0 9800 120 9920 0 FreeSans 480 0 0 0 FrameData[31]
port 39 nsew signal input
flabel metal3 s 0 2184 120 2304 0 FreeSans 480 0 0 0 FrameData[3]
port 40 nsew signal input
flabel metal3 s 0 2456 120 2576 0 FreeSans 480 0 0 0 FrameData[4]
port 41 nsew signal input
flabel metal3 s 0 2728 120 2848 0 FreeSans 480 0 0 0 FrameData[5]
port 42 nsew signal input
flabel metal3 s 0 3000 120 3120 0 FreeSans 480 0 0 0 FrameData[6]
port 43 nsew signal input
flabel metal3 s 0 3272 120 3392 0 FreeSans 480 0 0 0 FrameData[7]
port 44 nsew signal input
flabel metal3 s 0 3544 120 3664 0 FreeSans 480 0 0 0 FrameData[8]
port 45 nsew signal input
flabel metal3 s 0 3816 120 3936 0 FreeSans 480 0 0 0 FrameData[9]
port 46 nsew signal input
flabel metal3 s 40880 1368 41000 1488 0 FreeSans 480 0 0 0 FrameData_O[0]
port 47 nsew signal output
flabel metal3 s 40880 4088 41000 4208 0 FreeSans 480 0 0 0 FrameData_O[10]
port 48 nsew signal output
flabel metal3 s 40880 4360 41000 4480 0 FreeSans 480 0 0 0 FrameData_O[11]
port 49 nsew signal output
flabel metal3 s 40880 4632 41000 4752 0 FreeSans 480 0 0 0 FrameData_O[12]
port 50 nsew signal output
flabel metal3 s 40880 4904 41000 5024 0 FreeSans 480 0 0 0 FrameData_O[13]
port 51 nsew signal output
flabel metal3 s 40880 5176 41000 5296 0 FreeSans 480 0 0 0 FrameData_O[14]
port 52 nsew signal output
flabel metal3 s 40880 5448 41000 5568 0 FreeSans 480 0 0 0 FrameData_O[15]
port 53 nsew signal output
flabel metal3 s 40880 5720 41000 5840 0 FreeSans 480 0 0 0 FrameData_O[16]
port 54 nsew signal output
flabel metal3 s 40880 5992 41000 6112 0 FreeSans 480 0 0 0 FrameData_O[17]
port 55 nsew signal output
flabel metal3 s 40880 6264 41000 6384 0 FreeSans 480 0 0 0 FrameData_O[18]
port 56 nsew signal output
flabel metal3 s 40880 6536 41000 6656 0 FreeSans 480 0 0 0 FrameData_O[19]
port 57 nsew signal output
flabel metal3 s 40880 1640 41000 1760 0 FreeSans 480 0 0 0 FrameData_O[1]
port 58 nsew signal output
flabel metal3 s 40880 6808 41000 6928 0 FreeSans 480 0 0 0 FrameData_O[20]
port 59 nsew signal output
flabel metal3 s 40880 7080 41000 7200 0 FreeSans 480 0 0 0 FrameData_O[21]
port 60 nsew signal output
flabel metal3 s 40880 7352 41000 7472 0 FreeSans 480 0 0 0 FrameData_O[22]
port 61 nsew signal output
flabel metal3 s 40880 7624 41000 7744 0 FreeSans 480 0 0 0 FrameData_O[23]
port 62 nsew signal output
flabel metal3 s 40880 7896 41000 8016 0 FreeSans 480 0 0 0 FrameData_O[24]
port 63 nsew signal output
flabel metal3 s 40880 8168 41000 8288 0 FreeSans 480 0 0 0 FrameData_O[25]
port 64 nsew signal output
flabel metal3 s 40880 8440 41000 8560 0 FreeSans 480 0 0 0 FrameData_O[26]
port 65 nsew signal output
flabel metal3 s 40880 8712 41000 8832 0 FreeSans 480 0 0 0 FrameData_O[27]
port 66 nsew signal output
flabel metal3 s 40880 8984 41000 9104 0 FreeSans 480 0 0 0 FrameData_O[28]
port 67 nsew signal output
flabel metal3 s 40880 9256 41000 9376 0 FreeSans 480 0 0 0 FrameData_O[29]
port 68 nsew signal output
flabel metal3 s 40880 1912 41000 2032 0 FreeSans 480 0 0 0 FrameData_O[2]
port 69 nsew signal output
flabel metal3 s 40880 9528 41000 9648 0 FreeSans 480 0 0 0 FrameData_O[30]
port 70 nsew signal output
flabel metal3 s 40880 9800 41000 9920 0 FreeSans 480 0 0 0 FrameData_O[31]
port 71 nsew signal output
flabel metal3 s 40880 2184 41000 2304 0 FreeSans 480 0 0 0 FrameData_O[3]
port 72 nsew signal output
flabel metal3 s 40880 2456 41000 2576 0 FreeSans 480 0 0 0 FrameData_O[4]
port 73 nsew signal output
flabel metal3 s 40880 2728 41000 2848 0 FreeSans 480 0 0 0 FrameData_O[5]
port 74 nsew signal output
flabel metal3 s 40880 3000 41000 3120 0 FreeSans 480 0 0 0 FrameData_O[6]
port 75 nsew signal output
flabel metal3 s 40880 3272 41000 3392 0 FreeSans 480 0 0 0 FrameData_O[7]
port 76 nsew signal output
flabel metal3 s 40880 3544 41000 3664 0 FreeSans 480 0 0 0 FrameData_O[8]
port 77 nsew signal output
flabel metal3 s 40880 3816 41000 3936 0 FreeSans 480 0 0 0 FrameData_O[9]
port 78 nsew signal output
flabel metal2 s 32494 0 32550 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 79 nsew signal input
flabel metal2 s 35254 0 35310 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 80 nsew signal input
flabel metal2 s 35530 0 35586 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 81 nsew signal input
flabel metal2 s 35806 0 35862 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 82 nsew signal input
flabel metal2 s 36082 0 36138 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 83 nsew signal input
flabel metal2 s 36358 0 36414 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 84 nsew signal input
flabel metal2 s 36634 0 36690 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 85 nsew signal input
flabel metal2 s 36910 0 36966 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 86 nsew signal input
flabel metal2 s 37186 0 37242 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 87 nsew signal input
flabel metal2 s 37462 0 37518 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 88 nsew signal input
flabel metal2 s 37738 0 37794 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 89 nsew signal input
flabel metal2 s 32770 0 32826 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 90 nsew signal input
flabel metal2 s 33046 0 33102 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 91 nsew signal input
flabel metal2 s 33322 0 33378 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 92 nsew signal input
flabel metal2 s 33598 0 33654 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 93 nsew signal input
flabel metal2 s 33874 0 33930 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 94 nsew signal input
flabel metal2 s 34150 0 34206 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 95 nsew signal input
flabel metal2 s 34426 0 34482 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 96 nsew signal input
flabel metal2 s 34702 0 34758 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 97 nsew signal input
flabel metal2 s 34978 0 35034 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 98 nsew signal input
flabel metal2 s 18234 11194 18290 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 99 nsew signal output
flabel metal2 s 29274 11194 29330 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 100 nsew signal output
flabel metal2 s 30378 11194 30434 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 101 nsew signal output
flabel metal2 s 31482 11194 31538 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 102 nsew signal output
flabel metal2 s 32586 11194 32642 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 103 nsew signal output
flabel metal2 s 33690 11194 33746 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 104 nsew signal output
flabel metal2 s 34794 11194 34850 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 105 nsew signal output
flabel metal2 s 35898 11194 35954 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 106 nsew signal output
flabel metal2 s 37002 11194 37058 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 107 nsew signal output
flabel metal2 s 38106 11194 38162 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 108 nsew signal output
flabel metal2 s 39210 11194 39266 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 109 nsew signal output
flabel metal2 s 19338 11194 19394 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 110 nsew signal output
flabel metal2 s 20442 11194 20498 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 111 nsew signal output
flabel metal2 s 21546 11194 21602 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 112 nsew signal output
flabel metal2 s 22650 11194 22706 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 113 nsew signal output
flabel metal2 s 23754 11194 23810 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 114 nsew signal output
flabel metal2 s 24858 11194 24914 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 115 nsew signal output
flabel metal2 s 25962 11194 26018 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 116 nsew signal output
flabel metal2 s 27066 11194 27122 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 117 nsew signal output
flabel metal2 s 28170 11194 28226 11250 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 118 nsew signal output
flabel metal2 s 3238 0 3294 56 0 FreeSans 224 0 0 0 N1END[0]
port 119 nsew signal input
flabel metal2 s 3514 0 3570 56 0 FreeSans 224 0 0 0 N1END[1]
port 120 nsew signal input
flabel metal2 s 3790 0 3846 56 0 FreeSans 224 0 0 0 N1END[2]
port 121 nsew signal input
flabel metal2 s 4066 0 4122 56 0 FreeSans 224 0 0 0 N1END[3]
port 122 nsew signal input
flabel metal2 s 6550 0 6606 56 0 FreeSans 224 0 0 0 N2END[0]
port 123 nsew signal input
flabel metal2 s 6826 0 6882 56 0 FreeSans 224 0 0 0 N2END[1]
port 124 nsew signal input
flabel metal2 s 7102 0 7158 56 0 FreeSans 224 0 0 0 N2END[2]
port 125 nsew signal input
flabel metal2 s 7378 0 7434 56 0 FreeSans 224 0 0 0 N2END[3]
port 126 nsew signal input
flabel metal2 s 7654 0 7710 56 0 FreeSans 224 0 0 0 N2END[4]
port 127 nsew signal input
flabel metal2 s 7930 0 7986 56 0 FreeSans 224 0 0 0 N2END[5]
port 128 nsew signal input
flabel metal2 s 8206 0 8262 56 0 FreeSans 224 0 0 0 N2END[6]
port 129 nsew signal input
flabel metal2 s 8482 0 8538 56 0 FreeSans 224 0 0 0 N2END[7]
port 130 nsew signal input
flabel metal2 s 4342 0 4398 56 0 FreeSans 224 0 0 0 N2MID[0]
port 131 nsew signal input
flabel metal2 s 4618 0 4674 56 0 FreeSans 224 0 0 0 N2MID[1]
port 132 nsew signal input
flabel metal2 s 4894 0 4950 56 0 FreeSans 224 0 0 0 N2MID[2]
port 133 nsew signal input
flabel metal2 s 5170 0 5226 56 0 FreeSans 224 0 0 0 N2MID[3]
port 134 nsew signal input
flabel metal2 s 5446 0 5502 56 0 FreeSans 224 0 0 0 N2MID[4]
port 135 nsew signal input
flabel metal2 s 5722 0 5778 56 0 FreeSans 224 0 0 0 N2MID[5]
port 136 nsew signal input
flabel metal2 s 5998 0 6054 56 0 FreeSans 224 0 0 0 N2MID[6]
port 137 nsew signal input
flabel metal2 s 6274 0 6330 56 0 FreeSans 224 0 0 0 N2MID[7]
port 138 nsew signal input
flabel metal2 s 8758 0 8814 56 0 FreeSans 224 0 0 0 N4END[0]
port 139 nsew signal input
flabel metal2 s 11518 0 11574 56 0 FreeSans 224 0 0 0 N4END[10]
port 140 nsew signal input
flabel metal2 s 11794 0 11850 56 0 FreeSans 224 0 0 0 N4END[11]
port 141 nsew signal input
flabel metal2 s 12070 0 12126 56 0 FreeSans 224 0 0 0 N4END[12]
port 142 nsew signal input
flabel metal2 s 12346 0 12402 56 0 FreeSans 224 0 0 0 N4END[13]
port 143 nsew signal input
flabel metal2 s 12622 0 12678 56 0 FreeSans 224 0 0 0 N4END[14]
port 144 nsew signal input
flabel metal2 s 12898 0 12954 56 0 FreeSans 224 0 0 0 N4END[15]
port 145 nsew signal input
flabel metal2 s 9034 0 9090 56 0 FreeSans 224 0 0 0 N4END[1]
port 146 nsew signal input
flabel metal2 s 9310 0 9366 56 0 FreeSans 224 0 0 0 N4END[2]
port 147 nsew signal input
flabel metal2 s 9586 0 9642 56 0 FreeSans 224 0 0 0 N4END[3]
port 148 nsew signal input
flabel metal2 s 9862 0 9918 56 0 FreeSans 224 0 0 0 N4END[4]
port 149 nsew signal input
flabel metal2 s 10138 0 10194 56 0 FreeSans 224 0 0 0 N4END[5]
port 150 nsew signal input
flabel metal2 s 10414 0 10470 56 0 FreeSans 224 0 0 0 N4END[6]
port 151 nsew signal input
flabel metal2 s 10690 0 10746 56 0 FreeSans 224 0 0 0 N4END[7]
port 152 nsew signal input
flabel metal2 s 10966 0 11022 56 0 FreeSans 224 0 0 0 N4END[8]
port 153 nsew signal input
flabel metal2 s 11242 0 11298 56 0 FreeSans 224 0 0 0 N4END[9]
port 154 nsew signal input
flabel metal2 s 13174 0 13230 56 0 FreeSans 224 0 0 0 NN4END[0]
port 155 nsew signal input
flabel metal2 s 15934 0 15990 56 0 FreeSans 224 0 0 0 NN4END[10]
port 156 nsew signal input
flabel metal2 s 16210 0 16266 56 0 FreeSans 224 0 0 0 NN4END[11]
port 157 nsew signal input
flabel metal2 s 16486 0 16542 56 0 FreeSans 224 0 0 0 NN4END[12]
port 158 nsew signal input
flabel metal2 s 16762 0 16818 56 0 FreeSans 224 0 0 0 NN4END[13]
port 159 nsew signal input
flabel metal2 s 17038 0 17094 56 0 FreeSans 224 0 0 0 NN4END[14]
port 160 nsew signal input
flabel metal2 s 17314 0 17370 56 0 FreeSans 224 0 0 0 NN4END[15]
port 161 nsew signal input
flabel metal2 s 13450 0 13506 56 0 FreeSans 224 0 0 0 NN4END[1]
port 162 nsew signal input
flabel metal2 s 13726 0 13782 56 0 FreeSans 224 0 0 0 NN4END[2]
port 163 nsew signal input
flabel metal2 s 14002 0 14058 56 0 FreeSans 224 0 0 0 NN4END[3]
port 164 nsew signal input
flabel metal2 s 14278 0 14334 56 0 FreeSans 224 0 0 0 NN4END[4]
port 165 nsew signal input
flabel metal2 s 14554 0 14610 56 0 FreeSans 224 0 0 0 NN4END[5]
port 166 nsew signal input
flabel metal2 s 14830 0 14886 56 0 FreeSans 224 0 0 0 NN4END[6]
port 167 nsew signal input
flabel metal2 s 15106 0 15162 56 0 FreeSans 224 0 0 0 NN4END[7]
port 168 nsew signal input
flabel metal2 s 15382 0 15438 56 0 FreeSans 224 0 0 0 NN4END[8]
port 169 nsew signal input
flabel metal2 s 15658 0 15714 56 0 FreeSans 224 0 0 0 NN4END[9]
port 170 nsew signal input
flabel metal2 s 17866 0 17922 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 171 nsew signal output
flabel metal2 s 18142 0 18198 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 172 nsew signal output
flabel metal2 s 18418 0 18474 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 173 nsew signal output
flabel metal2 s 18694 0 18750 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 174 nsew signal output
flabel metal2 s 18970 0 19026 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 175 nsew signal output
flabel metal2 s 19246 0 19302 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 176 nsew signal output
flabel metal2 s 19522 0 19578 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 177 nsew signal output
flabel metal2 s 19798 0 19854 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 178 nsew signal output
flabel metal2 s 20074 0 20130 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 179 nsew signal output
flabel metal2 s 20350 0 20406 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 180 nsew signal output
flabel metal2 s 20626 0 20682 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 181 nsew signal output
flabel metal2 s 20902 0 20958 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 182 nsew signal output
flabel metal2 s 21178 0 21234 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 183 nsew signal output
flabel metal2 s 21454 0 21510 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 184 nsew signal output
flabel metal2 s 21730 0 21786 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 185 nsew signal output
flabel metal2 s 22006 0 22062 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 186 nsew signal output
flabel metal2 s 22282 0 22338 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 187 nsew signal output
flabel metal2 s 22558 0 22614 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 188 nsew signal output
flabel metal2 s 22834 0 22890 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 189 nsew signal output
flabel metal2 s 23110 0 23166 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 190 nsew signal output
flabel metal2 s 23386 0 23442 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 191 nsew signal output
flabel metal2 s 26146 0 26202 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 192 nsew signal output
flabel metal2 s 26422 0 26478 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 193 nsew signal output
flabel metal2 s 26698 0 26754 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 194 nsew signal output
flabel metal2 s 26974 0 27030 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 195 nsew signal output
flabel metal2 s 27250 0 27306 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 196 nsew signal output
flabel metal2 s 27526 0 27582 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 197 nsew signal output
flabel metal2 s 23662 0 23718 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 198 nsew signal output
flabel metal2 s 23938 0 23994 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 199 nsew signal output
flabel metal2 s 24214 0 24270 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 200 nsew signal output
flabel metal2 s 24490 0 24546 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 201 nsew signal output
flabel metal2 s 24766 0 24822 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 202 nsew signal output
flabel metal2 s 25042 0 25098 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 203 nsew signal output
flabel metal2 s 25318 0 25374 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 204 nsew signal output
flabel metal2 s 25594 0 25650 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 205 nsew signal output
flabel metal2 s 25870 0 25926 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 206 nsew signal output
flabel metal2 s 27802 0 27858 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 207 nsew signal output
flabel metal2 s 30562 0 30618 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 208 nsew signal output
flabel metal2 s 30838 0 30894 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 209 nsew signal output
flabel metal2 s 31114 0 31170 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 210 nsew signal output
flabel metal2 s 31390 0 31446 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 211 nsew signal output
flabel metal2 s 31666 0 31722 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 212 nsew signal output
flabel metal2 s 31942 0 31998 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 213 nsew signal output
flabel metal2 s 28078 0 28134 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 214 nsew signal output
flabel metal2 s 28354 0 28410 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 215 nsew signal output
flabel metal2 s 28630 0 28686 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 216 nsew signal output
flabel metal2 s 28906 0 28962 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 217 nsew signal output
flabel metal2 s 29182 0 29238 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 218 nsew signal output
flabel metal2 s 29458 0 29514 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 219 nsew signal output
flabel metal2 s 29734 0 29790 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 220 nsew signal output
flabel metal2 s 30010 0 30066 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 221 nsew signal output
flabel metal2 s 30286 0 30342 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 222 nsew signal output
flabel metal2 s 32218 0 32274 56 0 FreeSans 224 0 0 0 UserCLK
port 223 nsew signal input
flabel metal2 s 17130 11194 17186 11250 0 FreeSans 224 0 0 0 UserCLKo
port 224 nsew signal output
flabel metal4 s 3004 0 3324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 3004 0 3324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 3004 11190 3324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 9004 0 9324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 9004 0 9324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 9004 11190 9324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 15004 0 15324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 15004 0 15324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 15004 11190 15324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 21004 0 21324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 21004 0 21324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 21004 11190 21324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 27004 0 27324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 27004 0 27324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 27004 11190 27324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 33004 0 33324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 33004 0 33324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 33004 11190 33324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 39004 0 39324 11250 0 FreeSans 1920 90 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 39004 0 39324 60 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 39004 11190 39324 11250 0 FreeSans 480 0 0 0 VGND
port 225 nsew ground bidirectional
flabel metal4 s 1944 0 2264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 1944 0 2264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 1944 11190 2264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 7944 0 8264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 7944 0 8264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 7944 11190 8264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 13944 0 14264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 13944 0 14264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 13944 11190 14264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 19944 0 20264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 19944 0 20264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 19944 11190 20264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 25944 0 26264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 25944 0 26264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 25944 11190 26264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 31944 0 32264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 31944 0 32264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 31944 11190 32264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 37944 0 38264 11250 0 FreeSans 1920 90 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 37944 0 38264 60 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
flabel metal4 s 37944 11190 38264 11250 0 FreeSans 480 0 0 0 VPWR
port 226 nsew power bidirectional
rlabel metal1 20470 8704 20470 8704 0 VGND
rlabel metal1 20470 8160 20470 8160 0 VPWR
rlabel metal1 2944 8602 2944 8602 0 A_I_top
rlabel metal2 1702 9870 1702 9870 0 A_O_top
rlabel metal1 4416 8602 4416 8602 0 A_T_top
rlabel metal1 8694 8602 8694 8602 0 A_config_C_bit0
rlabel metal1 9522 8602 9522 8602 0 A_config_C_bit1
rlabel metal1 10626 8602 10626 8602 0 A_config_C_bit2
rlabel metal1 11776 8602 11776 8602 0 A_config_C_bit3
rlabel metal1 6302 8602 6302 8602 0 B_I_top
rlabel metal2 5014 9836 5014 9836 0 B_O_top
rlabel metal1 7130 8602 7130 8602 0 B_T_top
rlabel metal1 12696 8602 12696 8602 0 B_config_C_bit0
rlabel metal1 14030 8602 14030 8602 0 B_config_C_bit1
rlabel metal1 15042 8602 15042 8602 0 B_config_C_bit2
rlabel metal1 16146 8602 16146 8602 0 B_config_C_bit3
rlabel metal3 436 1428 436 1428 0 FrameData[0]
rlabel metal3 988 4148 988 4148 0 FrameData[10]
rlabel metal3 804 4420 804 4420 0 FrameData[11]
rlabel metal3 551 4692 551 4692 0 FrameData[12]
rlabel metal3 804 4964 804 4964 0 FrameData[13]
rlabel metal3 988 5236 988 5236 0 FrameData[14]
rlabel metal3 1172 5508 1172 5508 0 FrameData[15]
rlabel metal3 804 5780 804 5780 0 FrameData[16]
rlabel metal3 758 6052 758 6052 0 FrameData[17]
rlabel metal3 850 6324 850 6324 0 FrameData[18]
rlabel metal3 758 6596 758 6596 0 FrameData[19]
rlabel metal3 666 1700 666 1700 0 FrameData[1]
rlabel metal3 896 6868 896 6868 0 FrameData[20]
rlabel metal3 804 7140 804 7140 0 FrameData[21]
rlabel metal3 758 7412 758 7412 0 FrameData[22]
rlabel metal3 804 7684 804 7684 0 FrameData[23]
rlabel metal3 1172 7956 1172 7956 0 FrameData[24]
rlabel metal3 758 8228 758 8228 0 FrameData[25]
rlabel via2 3358 8517 3358 8517 0 FrameData[26]
rlabel metal2 2806 8313 2806 8313 0 FrameData[27]
rlabel metal3 758 9044 758 9044 0 FrameData[28]
rlabel metal2 3910 8925 3910 8925 0 FrameData[29]
rlabel metal3 298 1972 298 1972 0 FrameData[2]
rlabel metal2 3450 8551 3450 8551 0 FrameData[30]
rlabel metal2 5566 9197 5566 9197 0 FrameData[31]
rlabel metal3 988 2244 988 2244 0 FrameData[3]
rlabel metal3 804 2516 804 2516 0 FrameData[4]
rlabel metal3 758 2788 758 2788 0 FrameData[5]
rlabel metal3 1172 3060 1172 3060 0 FrameData[6]
rlabel metal3 804 3332 804 3332 0 FrameData[7]
rlabel metal3 1126 3604 1126 3604 0 FrameData[8]
rlabel metal3 804 3876 804 3876 0 FrameData[9]
rlabel metal3 40488 1428 40488 1428 0 FrameData_O[0]
rlabel metal2 39422 3927 39422 3927 0 FrameData_O[10]
rlabel metal3 40166 4420 40166 4420 0 FrameData_O[11]
rlabel metal1 39468 3978 39468 3978 0 FrameData_O[12]
rlabel metal3 39982 4964 39982 4964 0 FrameData_O[13]
rlabel metal2 39422 5015 39422 5015 0 FrameData_O[14]
rlabel metal3 40442 5508 40442 5508 0 FrameData_O[15]
rlabel metal2 39422 5559 39422 5559 0 FrameData_O[16]
rlabel metal3 39982 6052 39982 6052 0 FrameData_O[17]
rlabel metal2 39422 6103 39422 6103 0 FrameData_O[18]
rlabel metal3 40166 6596 40166 6596 0 FrameData_O[19]
rlabel metal3 39798 1700 39798 1700 0 FrameData_O[1]
rlabel metal3 40488 6868 40488 6868 0 FrameData_O[20]
rlabel metal3 40166 7140 40166 7140 0 FrameData_O[21]
rlabel metal3 39936 7412 39936 7412 0 FrameData_O[22]
rlabel metal3 40166 7684 40166 7684 0 FrameData_O[23]
rlabel metal3 39982 7956 39982 7956 0 FrameData_O[24]
rlabel metal3 39706 8228 39706 8228 0 FrameData_O[25]
rlabel metal1 38732 7514 38732 7514 0 FrameData_O[26]
rlabel metal1 39054 6664 39054 6664 0 FrameData_O[27]
rlabel metal2 38318 8551 38318 8551 0 FrameData_O[28]
rlabel metal1 38180 7990 38180 7990 0 FrameData_O[29]
rlabel metal3 40258 1972 40258 1972 0 FrameData_O[2]
rlabel metal1 37030 8568 37030 8568 0 FrameData_O[30]
rlabel metal1 39468 6426 39468 6426 0 FrameData_O[31]
rlabel metal3 40442 2244 40442 2244 0 FrameData_O[3]
rlabel metal3 40304 2516 40304 2516 0 FrameData_O[4]
rlabel metal3 39982 2788 39982 2788 0 FrameData_O[5]
rlabel metal3 40166 3060 40166 3060 0 FrameData_O[6]
rlabel metal3 40442 3332 40442 3332 0 FrameData_O[7]
rlabel metal2 39422 3383 39422 3383 0 FrameData_O[8]
rlabel metal3 39982 3876 39982 3876 0 FrameData_O[9]
rlabel metal2 32522 1058 32522 1058 0 FrameStrobe[0]
rlabel metal2 35282 650 35282 650 0 FrameStrobe[10]
rlabel metal2 35558 3370 35558 3370 0 FrameStrobe[11]
rlabel metal2 35834 344 35834 344 0 FrameStrobe[12]
rlabel metal2 36110 276 36110 276 0 FrameStrobe[13]
rlabel metal2 36386 684 36386 684 0 FrameStrobe[14]
rlabel metal2 36662 106 36662 106 0 FrameStrobe[15]
rlabel metal2 36938 2248 36938 2248 0 FrameStrobe[16]
rlabel metal2 37214 55 37214 55 0 FrameStrobe[17]
rlabel metal2 37490 3948 37490 3948 0 FrameStrobe[18]
rlabel metal1 37858 6766 37858 6766 0 FrameStrobe[19]
rlabel metal2 17940 1156 17940 1156 0 FrameStrobe[1]
rlabel metal2 33074 412 33074 412 0 FrameStrobe[2]
rlabel metal2 13938 2210 13938 2210 0 FrameStrobe[3]
rlabel metal2 33626 208 33626 208 0 FrameStrobe[4]
rlabel metal2 33902 480 33902 480 0 FrameStrobe[5]
rlabel metal2 34178 531 34178 531 0 FrameStrobe[6]
rlabel metal2 34454 1058 34454 1058 0 FrameStrobe[7]
rlabel metal2 34730 548 34730 548 0 FrameStrobe[8]
rlabel metal2 35006 582 35006 582 0 FrameStrobe[9]
rlabel metal1 18400 8602 18400 8602 0 FrameStrobe_O[0]
rlabel metal1 29670 8602 29670 8602 0 FrameStrobe_O[10]
rlabel metal1 30498 8602 30498 8602 0 FrameStrobe_O[11]
rlabel metal1 32016 8602 32016 8602 0 FrameStrobe_O[12]
rlabel metal1 32706 8602 32706 8602 0 FrameStrobe_O[13]
rlabel metal1 33810 8602 33810 8602 0 FrameStrobe_O[14]
rlabel metal1 34914 8602 34914 8602 0 FrameStrobe_O[15]
rlabel metal1 36018 8602 36018 8602 0 FrameStrobe_O[16]
rlabel metal1 37352 8602 37352 8602 0 FrameStrobe_O[17]
rlabel metal1 38272 8602 38272 8602 0 FrameStrobe_O[18]
rlabel metal2 39422 9163 39422 9163 0 FrameStrobe_O[19]
rlabel metal1 19504 8602 19504 8602 0 FrameStrobe_O[1]
rlabel metal1 21528 8330 21528 8330 0 FrameStrobe_O[2]
rlabel metal1 21758 8602 21758 8602 0 FrameStrobe_O[3]
rlabel metal2 23690 9180 23690 9180 0 FrameStrobe_O[4]
rlabel metal1 23920 8602 23920 8602 0 FrameStrobe_O[5]
rlabel metal1 24656 8602 24656 8602 0 FrameStrobe_O[6]
rlabel metal1 26082 8602 26082 8602 0 FrameStrobe_O[7]
rlabel metal1 27324 8058 27324 8058 0 FrameStrobe_O[8]
rlabel metal2 29670 9010 29670 9010 0 FrameStrobe_O[9]
rlabel metal2 23782 2635 23782 2635 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 28474 6239 28474 6239 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 11914 6188 11914 6188 0 Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal1 11776 5814 11776 5814 0 Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal1 29486 2890 29486 2890 0 Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal1 30544 2550 30544 2550 0 Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal1 26634 5848 26634 5848 0 Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal1 27278 5746 27278 5746 0 Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal1 3588 3162 3588 3162 0 Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal1 4692 3162 4692 3162 0 Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 17411 4148 17411 4148 0 Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal1 33534 4794 33534 4794 0 Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal1 9476 5066 9476 5066 0 Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 9614 6137 9614 6137 0 Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal1 30682 5882 30682 5882 0 Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal1 10442 6222 10442 6222 0 Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal1 9108 5678 9108 5678 0 Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal1 10350 2482 10350 2482 0 Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal1 7038 3468 7038 3468 0 Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal1 4989 5236 4989 5236 0 Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal1 9890 4046 9890 4046 0 Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 10626 3978 10626 3978 0 Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 11638 5474 11638 5474 0 Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal1 13064 4794 13064 4794 0 Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 6578 3808 6578 3808 0 Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal1 30084 5338 30084 5338 0 Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal1 6302 5066 6302 5066 0 Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal1 6394 2890 6394 2890 0 Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal1 28980 4046 28980 4046 0 Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 29578 4556 29578 4556 0 Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 25530 8126 25530 8126 0 Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal1 26220 7514 26220 7514 0 Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal1 28704 6970 28704 6970 0 Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 29486 7820 29486 7820 0 Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 14582 7786 14582 7786 0 Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 15134 7276 15134 7276 0 Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal1 31786 3604 31786 3604 0 Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal1 31832 2550 31832 2550 0 Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 33718 6426 33718 6426 0 Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal1 32982 6222 32982 6222 0 Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 23506 3162 23506 3162 0 Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal1 24012 2550 24012 2550 0 Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal1 31924 7242 31924 7242 0 Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 32338 8126 32338 8126 0 Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 18630 7514 18630 7514 0 Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 19182 7820 19182 7820 0 Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 31878 3944 31878 3944 0 Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal1 24610 7208 24610 7208 0 Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal1 23782 7310 23782 7310 0 Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 27646 3162 27646 3162 0 Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 28198 3502 28198 3502 0 Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal1 23000 5814 23000 5814 0 Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel via1 23597 5746 23597 5746 0 Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal1 6900 5338 6900 5338 0 Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal1 6670 5746 6670 5746 0 Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal1 14628 4250 14628 4250 0 Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 15318 4862 15318 4862 0 Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel via1 32614 4607 32614 4607 0 Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 3634 3876 3634 3876 0 Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal1 4738 3944 4738 3944 0 Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal1 29486 6154 29486 6154 0 Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 30406 6086 30406 6086 0 Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 24242 4420 24242 4420 0 Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 23736 4046 23736 4046 0 Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal1 28474 7514 28474 7514 0 Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 28198 8126 28198 8126 0 Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal1 12190 7990 12190 7990 0 Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal1 12834 7514 12834 7514 0 Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal1 19918 3672 19918 3672 0 Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal1 20884 3570 20884 3570 0 Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal1 15042 5338 15042 5338 0 Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel via1 16606 6987 16606 6987 0 Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 13846 3366 13846 3366 0 Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal1 13892 2550 13892 2550 0 Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal1 32798 7208 32798 7208 0 Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal1 33442 7310 33442 7310 0 Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal1 18676 6222 18676 6222 0 Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 19366 6494 19366 6494 0 Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 30038 4658 30038 4658 0 Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal1 21344 7990 21344 7990 0 Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal1 21620 7514 21620 7514 0 Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal1 21022 2618 21022 2618 0 Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal1 20332 2618 20332 2618 0 Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal1 21390 6426 21390 6426 0 Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal1 20976 5882 20976 5882 0 Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 19274 4964 19274 4964 0 Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal1 18170 5066 18170 5066 0 Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal1 15686 6902 15686 6902 0 Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal1 15548 6970 15548 6970 0 Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal1 29762 4250 29762 4250 0 Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal1 16514 2516 16514 2516 0 Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal1 16514 2278 16514 2278 0 Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 6946 7412 6946 7412 0 Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel via2 6394 6851 6394 6851 0 Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal1 26082 4726 26082 4726 0 Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal1 26174 3978 26174 3978 0 Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 4462 7038 4462 7038 0 Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal1 4692 6834 4692 6834 0 Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal1 33534 2924 33534 2924 0 Inst_N_IO_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 22862 3298 22862 3298 0 Inst_N_IO_ConfigMem.Inst_frame3_bit15.Q
rlabel metal1 35926 4012 35926 4012 0 Inst_N_IO_ConfigMem.Inst_frame3_bit16.Q
rlabel metal1 36110 6290 36110 6290 0 Inst_N_IO_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 17894 5950 17894 5950 0 Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q
rlabel metal1 17802 5746 17802 5746 0 Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 8234 7514 8234 7514 0 Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 8786 7854 8786 7854 0 Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q
rlabel metal1 26772 2550 26772 2550 0 Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal1 26266 2516 26266 2516 0 Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal1 4002 6154 4002 6154 0 Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal1 4876 5882 4876 5882 0 Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal1 18998 3978 18998 3978 0 Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal1 19412 3706 19412 3706 0 Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 14766 5916 14766 5916 0 Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 15318 5610 15318 5610 0 Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal1 17066 3162 17066 3162 0 Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal1 16606 3570 16606 3570 0 Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal1 35466 2890 35466 2890 0 Inst_N_IO_switch_matrix.S1BEG0
rlabel metal1 22356 4250 22356 4250 0 Inst_N_IO_switch_matrix.S1BEG1
rlabel metal1 36662 4114 36662 4114 0 Inst_N_IO_switch_matrix.S1BEG2
rlabel metal1 35512 6426 35512 6426 0 Inst_N_IO_switch_matrix.S1BEG3
rlabel metal2 19090 6324 19090 6324 0 Inst_N_IO_switch_matrix.S2BEG0
rlabel metal1 9476 7378 9476 7378 0 Inst_N_IO_switch_matrix.S2BEG1
rlabel metal2 27646 3910 27646 3910 0 Inst_N_IO_switch_matrix.S2BEG2
rlabel metal1 5934 6256 5934 6256 0 Inst_N_IO_switch_matrix.S2BEG3
rlabel metal1 20608 4182 20608 4182 0 Inst_N_IO_switch_matrix.S2BEG4
rlabel metal1 16100 5882 16100 5882 0 Inst_N_IO_switch_matrix.S2BEG5
rlabel metal1 13938 3060 13938 3060 0 Inst_N_IO_switch_matrix.S2BEG6
rlabel metal1 13938 7854 13938 7854 0 Inst_N_IO_switch_matrix.S2BEG7
rlabel metal1 21850 5202 21850 5202 0 Inst_N_IO_switch_matrix.S2BEGb0
rlabel metal2 5750 7344 5750 7344 0 Inst_N_IO_switch_matrix.S2BEGb1
rlabel metal2 27462 4998 27462 4998 0 Inst_N_IO_switch_matrix.S2BEGb2
rlabel metal2 5658 6460 5658 6460 0 Inst_N_IO_switch_matrix.S2BEGb3
rlabel metal1 21758 3400 21758 3400 0 Inst_N_IO_switch_matrix.S2BEGb4
rlabel metal1 16606 6290 16606 6290 0 Inst_N_IO_switch_matrix.S2BEGb5
rlabel metal2 15962 5032 15962 5032 0 Inst_N_IO_switch_matrix.S2BEGb6
rlabel metal2 33994 7684 33994 7684 0 Inst_N_IO_switch_matrix.S2BEGb7
rlabel metal1 19872 6154 19872 6154 0 Inst_N_IO_switch_matrix.S4BEG0
rlabel metal1 22494 8058 22494 8058 0 Inst_N_IO_switch_matrix.S4BEG1
rlabel metal2 24886 4658 24886 4658 0 Inst_N_IO_switch_matrix.S4BEG10
rlabel metal1 29486 7854 29486 7854 0 Inst_N_IO_switch_matrix.S4BEG11
rlabel metal1 33580 3706 33580 3706 0 Inst_N_IO_switch_matrix.S4BEG12
rlabel metal1 34730 6426 34730 6426 0 Inst_N_IO_switch_matrix.S4BEG13
rlabel viali 26634 3031 26634 3031 0 Inst_N_IO_switch_matrix.S4BEG14
rlabel metal1 33028 7854 33028 7854 0 Inst_N_IO_switch_matrix.S4BEG15
rlabel metal1 21390 2822 21390 2822 0 Inst_N_IO_switch_matrix.S4BEG2
rlabel metal1 22356 6766 22356 6766 0 Inst_N_IO_switch_matrix.S4BEG3
rlabel metal1 20608 5338 20608 5338 0 Inst_N_IO_switch_matrix.S4BEG4
rlabel metal1 16790 8058 16790 8058 0 Inst_N_IO_switch_matrix.S4BEG5
rlabel metal2 17526 3740 17526 3740 0 Inst_N_IO_switch_matrix.S4BEG6
rlabel metal2 15778 7990 15778 7990 0 Inst_N_IO_switch_matrix.S4BEG7
rlabel metal1 33028 4794 33028 4794 0 Inst_N_IO_switch_matrix.S4BEG8
rlabel metal1 31188 6290 31188 6290 0 Inst_N_IO_switch_matrix.S4BEG9
rlabel metal2 19826 7684 19826 7684 0 Inst_N_IO_switch_matrix.SS4BEG0
rlabel metal1 23736 7514 23736 7514 0 Inst_N_IO_switch_matrix.SS4BEG1
rlabel metal1 26772 7854 26772 7854 0 Inst_N_IO_switch_matrix.SS4BEG10
rlabel metal2 30130 7684 30130 7684 0 Inst_N_IO_switch_matrix.SS4BEG11
rlabel metal1 33856 2482 33856 2482 0 Inst_N_IO_switch_matrix.SS4BEG12
rlabel metal1 27600 5202 27600 5202 0 Inst_N_IO_switch_matrix.SS4BEG13
rlabel metal1 3634 4590 3634 4590 0 Inst_N_IO_switch_matrix.SS4BEG14
rlabel metal2 16238 4998 16238 4998 0 Inst_N_IO_switch_matrix.SS4BEG15
rlabel metal1 28888 3162 28888 3162 0 Inst_N_IO_switch_matrix.SS4BEG2
rlabel metal1 24334 5678 24334 5678 0 Inst_N_IO_switch_matrix.SS4BEG3
rlabel metal1 6762 5882 6762 5882 0 Inst_N_IO_switch_matrix.SS4BEG4
rlabel metal1 15410 4794 15410 4794 0 Inst_N_IO_switch_matrix.SS4BEG5
rlabel metal2 3542 4726 3542 4726 0 Inst_N_IO_switch_matrix.SS4BEG6
rlabel metal1 13432 5678 13432 5678 0 Inst_N_IO_switch_matrix.SS4BEG7
rlabel metal1 31050 6970 31050 6970 0 Inst_N_IO_switch_matrix.SS4BEG8
rlabel metal1 30590 4114 30590 4114 0 Inst_N_IO_switch_matrix.SS4BEG9
rlabel metal2 3266 55 3266 55 0 N1END[0]
rlabel metal1 2691 2346 2691 2346 0 N1END[1]
rlabel metal2 3772 6766 3772 6766 0 N1END[2]
rlabel metal2 4094 55 4094 55 0 N1END[3]
rlabel metal2 6578 1194 6578 1194 0 N2END[0]
rlabel metal1 2530 4148 2530 4148 0 N2END[1]
rlabel metal2 7130 1415 7130 1415 0 N2END[2]
rlabel metal2 7406 599 7406 599 0 N2END[3]
rlabel metal2 7682 684 7682 684 0 N2END[4]
rlabel metal2 7958 1228 7958 1228 0 N2END[5]
rlabel metal2 8234 1160 8234 1160 0 N2END[6]
rlabel metal2 8510 667 8510 667 0 N2END[7]
rlabel metal2 4370 55 4370 55 0 N2MID[0]
rlabel metal2 4646 684 4646 684 0 N2MID[1]
rlabel metal1 2668 5202 2668 5202 0 N2MID[2]
rlabel metal2 5198 55 5198 55 0 N2MID[3]
rlabel metal2 5474 667 5474 667 0 N2MID[4]
rlabel metal1 6072 3026 6072 3026 0 N2MID[5]
rlabel metal2 6026 650 6026 650 0 N2MID[6]
rlabel metal2 6302 1228 6302 1228 0 N2MID[7]
rlabel metal2 8786 616 8786 616 0 N4END[0]
rlabel metal1 11592 2958 11592 2958 0 N4END[10]
rlabel metal2 11822 480 11822 480 0 N4END[11]
rlabel metal2 12098 242 12098 242 0 N4END[12]
rlabel metal2 12374 55 12374 55 0 N4END[13]
rlabel metal2 12650 55 12650 55 0 N4END[14]
rlabel metal2 12926 684 12926 684 0 N4END[15]
rlabel metal2 9062 446 9062 446 0 N4END[1]
rlabel metal2 9338 616 9338 616 0 N4END[2]
rlabel metal2 9614 1075 9614 1075 0 N4END[3]
rlabel metal2 9890 922 9890 922 0 N4END[4]
rlabel metal2 10166 684 10166 684 0 N4END[5]
rlabel metal2 10442 956 10442 956 0 N4END[6]
rlabel metal2 10718 616 10718 616 0 N4END[7]
rlabel metal2 10994 55 10994 55 0 N4END[8]
rlabel via2 11270 55 11270 55 0 N4END[9]
rlabel metal2 13202 1483 13202 1483 0 NN4END[0]
rlabel metal2 15962 1194 15962 1194 0 NN4END[10]
rlabel metal2 16238 650 16238 650 0 NN4END[11]
rlabel metal2 16514 395 16514 395 0 NN4END[12]
rlabel metal2 16790 667 16790 667 0 NN4END[13]
rlabel metal1 16974 2890 16974 2890 0 NN4END[14]
rlabel metal2 17342 276 17342 276 0 NN4END[15]
rlabel metal1 13432 6766 13432 6766 0 NN4END[1]
rlabel metal2 13754 1347 13754 1347 0 NN4END[2]
rlabel metal2 14030 55 14030 55 0 NN4END[3]
rlabel metal2 14306 735 14306 735 0 NN4END[4]
rlabel metal2 14582 208 14582 208 0 NN4END[5]
rlabel metal2 14858 242 14858 242 0 NN4END[6]
rlabel metal2 15134 684 15134 684 0 NN4END[7]
rlabel metal2 15410 990 15410 990 0 NN4END[8]
rlabel metal2 15686 378 15686 378 0 NN4END[9]
rlabel metal2 17894 174 17894 174 0 S1BEG[0]
rlabel metal2 18170 242 18170 242 0 S1BEG[1]
rlabel metal1 18078 3910 18078 3910 0 S1BEG[2]
rlabel metal2 18722 718 18722 718 0 S1BEG[3]
rlabel metal1 19228 5542 19228 5542 0 S2BEG[0]
rlabel metal2 19274 752 19274 752 0 S2BEG[1]
rlabel metal2 19550 55 19550 55 0 S2BEG[2]
rlabel metal2 19826 684 19826 684 0 S2BEG[3]
rlabel metal2 20102 684 20102 684 0 S2BEG[4]
rlabel metal2 20378 718 20378 718 0 S2BEG[5]
rlabel metal2 20654 667 20654 667 0 S2BEG[6]
rlabel metal2 21022 3162 21022 3162 0 S2BEG[7]
rlabel metal2 21206 174 21206 174 0 S2BEGb[0]
rlabel metal2 21482 735 21482 735 0 S2BEGb[1]
rlabel metal2 21758 616 21758 616 0 S2BEGb[2]
rlabel metal2 22034 650 22034 650 0 S2BEGb[3]
rlabel metal2 22310 446 22310 446 0 S2BEGb[4]
rlabel metal2 22586 174 22586 174 0 S2BEGb[5]
rlabel metal1 31970 2516 31970 2516 0 S2BEGb[6]
rlabel metal2 23138 582 23138 582 0 S2BEGb[7]
rlabel metal2 23414 55 23414 55 0 S4BEG[0]
rlabel metal2 26174 208 26174 208 0 S4BEG[10]
rlabel metal2 32706 1666 32706 1666 0 S4BEG[11]
rlabel metal2 32798 1768 32798 1768 0 S4BEG[12]
rlabel metal2 27002 310 27002 310 0 S4BEG[13]
rlabel metal2 33442 1258 33442 1258 0 S4BEG[14]
rlabel metal1 32154 2856 32154 2856 0 S4BEG[15]
rlabel metal2 23690 242 23690 242 0 S4BEG[1]
rlabel metal2 23966 55 23966 55 0 S4BEG[2]
rlabel metal2 24242 548 24242 548 0 S4BEG[3]
rlabel metal2 24518 684 24518 684 0 S4BEG[4]
rlabel metal2 24794 378 24794 378 0 S4BEG[5]
rlabel metal2 25070 650 25070 650 0 S4BEG[6]
rlabel metal2 25346 616 25346 616 0 S4BEG[7]
rlabel metal2 25622 480 25622 480 0 S4BEG[8]
rlabel metal2 25898 667 25898 667 0 S4BEG[9]
rlabel metal2 27830 378 27830 378 0 SS4BEG[0]
rlabel metal2 34638 884 34638 884 0 SS4BEG[10]
rlabel metal2 32614 1411 32614 1411 0 SS4BEG[11]
rlabel metal2 36478 1870 36478 1870 0 SS4BEG[12]
rlabel metal1 35466 2822 35466 2822 0 SS4BEG[13]
rlabel metal1 33810 850 33810 850 0 SS4BEG[14]
rlabel metal2 31970 514 31970 514 0 SS4BEG[15]
rlabel metal2 34914 1394 34914 1394 0 SS4BEG[1]
rlabel metal2 34546 1972 34546 1972 0 SS4BEG[2]
rlabel metal2 35190 1649 35190 1649 0 SS4BEG[3]
rlabel metal2 28934 480 28934 480 0 SS4BEG[4]
rlabel metal2 34178 1700 34178 1700 0 SS4BEG[5]
rlabel metal2 35650 1462 35650 1462 0 SS4BEG[6]
rlabel metal2 29762 990 29762 990 0 SS4BEG[7]
rlabel metal2 32338 2380 32338 2380 0 SS4BEG[8]
rlabel metal1 33350 3638 33350 3638 0 SS4BEG[9]
rlabel metal3 19159 2516 19159 2516 0 UserCLK
rlabel via3 18837 2652 18837 2652 0 UserCLK_regs
rlabel metal1 17112 8602 17112 8602 0 UserCLKo
rlabel metal1 12282 4114 12282 4114 0 _000_
rlabel metal2 11822 4250 11822 4250 0 _001_
rlabel metal1 9062 5814 9062 5814 0 _002_
rlabel metal1 10902 6800 10902 6800 0 _003_
rlabel metal2 11638 1700 11638 1700 0 _004_
rlabel metal1 6624 4114 6624 4114 0 _005_
rlabel metal2 12742 3910 12742 3910 0 _006_
rlabel metal2 13294 3740 13294 3740 0 _007_
rlabel metal1 10994 4012 10994 4012 0 _008_
rlabel metal1 12420 3502 12420 3502 0 _009_
rlabel metal1 11592 4114 11592 4114 0 _010_
rlabel metal1 11914 4250 11914 4250 0 _011_
rlabel metal2 12006 3706 12006 3706 0 _012_
rlabel metal1 10028 4590 10028 4590 0 _013_
rlabel metal2 10350 5542 10350 5542 0 _014_
rlabel metal1 9338 5338 9338 5338 0 _015_
rlabel metal2 10534 6596 10534 6596 0 _016_
rlabel metal2 11454 6086 11454 6086 0 _017_
rlabel metal1 11086 4998 11086 4998 0 _018_
rlabel metal1 10580 6426 10580 6426 0 _019_
rlabel metal1 11500 2414 11500 2414 0 _020_
rlabel metal2 7866 2720 7866 2720 0 _021_
rlabel metal1 10212 2550 10212 2550 0 _022_
rlabel metal2 8234 3536 8234 3536 0 _023_
rlabel metal1 7636 3434 7636 3434 0 _024_
rlabel viali 7970 3570 7970 3570 0 _025_
rlabel metal1 6854 4080 6854 4080 0 _026_
rlabel metal1 6394 3978 6394 3978 0 _027_
rlabel metal1 6578 3570 6578 3570 0 _028_
rlabel metal1 6900 2550 6900 2550 0 _029_
rlabel metal2 6302 4284 6302 4284 0 _030_
rlabel metal2 6210 3791 6210 3791 0 _031_
rlabel metal2 35926 5406 35926 5406 0 clknet_0_UserCLK
rlabel metal1 35282 4794 35282 4794 0 clknet_0_UserCLK_regs
rlabel metal1 34546 6766 34546 6766 0 clknet_1_0__leaf_UserCLK
rlabel metal2 34362 3876 34362 3876 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal2 34086 5372 34086 5372 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal2 2530 9248 2530 9248 0 net1
rlabel metal2 1702 5389 1702 5389 0 net10
rlabel metal1 8993 7310 8993 7310 0 net100
rlabel metal1 20436 5134 20436 5134 0 net101
rlabel metal1 12742 7922 12742 7922 0 net102
rlabel via1 24070 4046 24070 4046 0 net103
rlabel metal2 10304 6630 10304 6630 0 net104
rlabel metal1 8510 3706 8510 3706 0 net105
rlabel metal2 17250 10302 17250 10302 0 net106
rlabel metal2 17710 8483 17710 8483 0 net107
rlabel metal3 14812 5508 14812 5508 0 net108
rlabel metal1 5060 8058 5060 8058 0 net109
rlabel metal1 2300 5814 2300 5814 0 net11
rlabel metal2 6670 8840 6670 8840 0 net110
rlabel metal2 6854 6086 6854 6086 0 net111
rlabel metal2 21666 5525 21666 5525 0 net112
rlabel metal2 14398 9520 14398 9520 0 net113
rlabel metal2 20746 9316 20746 9316 0 net114
rlabel metal1 21574 9758 21574 9758 0 net115
rlabel metal1 35788 2618 35788 2618 0 net116
rlabel metal1 39100 3502 39100 3502 0 net117
rlabel metal1 36846 3162 36846 3162 0 net118
rlabel metal1 39192 4114 39192 4114 0 net119
rlabel via2 1702 7395 1702 7395 0 net12
rlabel via2 38870 5219 38870 5219 0 net120
rlabel metal3 13087 4828 13087 4828 0 net121
rlabel metal2 17986 10013 17986 10013 0 net122
rlabel metal1 39100 5202 39100 5202 0 net123
rlabel metal2 36202 5780 36202 5780 0 net124
rlabel metal2 36478 7973 36478 7973 0 net125
rlabel metal1 39238 6800 39238 6800 0 net126
rlabel metal1 34224 2550 34224 2550 0 net127
rlabel metal2 34362 8721 34362 8721 0 net128
rlabel metal1 38870 7378 38870 7378 0 net129
rlabel metal1 16376 5678 16376 5678 0 net13
rlabel via2 38686 7939 38686 7939 0 net130
rlabel metal2 16514 1411 16514 1411 0 net131
rlabel metal2 16514 9537 16514 9537 0 net132
rlabel via2 37858 8483 37858 8483 0 net133
rlabel metal1 15594 1190 15594 1190 0 net134
rlabel via2 16514 1003 16514 1003 0 net135
rlabel metal2 34454 9078 34454 9078 0 net136
rlabel metal2 32798 8517 32798 8517 0 net137
rlabel metal2 38134 2465 38134 2465 0 net138
rlabel via2 16514 867 16514 867 0 net139
rlabel metal1 12466 7380 12466 7380 0 net14
rlabel metal2 17618 1122 17618 1122 0 net140
rlabel metal1 33350 2550 33350 2550 0 net141
rlabel metal2 16514 9877 16514 9877 0 net142
rlabel metal2 16422 901 16422 901 0 net143
rlabel via2 39238 2397 39238 2397 0 net144
rlabel metal2 32246 4250 32246 4250 0 net145
rlabel metal2 16514 8585 16514 8585 0 net146
rlabel metal2 15134 9333 15134 9333 0 net147
rlabel metal1 21068 5814 21068 5814 0 net148
rlabel metal1 37858 6154 37858 6154 0 net149
rlabel metal1 1748 5814 1748 5814 0 net15
rlabel metal1 37996 6970 37996 6970 0 net150
rlabel metal2 38042 3400 38042 3400 0 net151
rlabel metal1 38410 3706 38410 3706 0 net152
rlabel metal1 37720 3162 37720 3162 0 net153
rlabel metal1 36800 5882 36800 5882 0 net154
rlabel metal1 38456 6630 38456 6630 0 net155
rlabel metal1 37950 6426 37950 6426 0 net156
rlabel metal2 37674 8228 37674 8228 0 net157
rlabel via1 38778 6715 38778 6715 0 net158
rlabel metal1 19458 8432 19458 8432 0 net159
rlabel metal1 1794 6698 1794 6698 0 net16
rlabel metal2 12834 7752 12834 7752 0 net160
rlabel metal1 36064 3162 36064 3162 0 net161
rlabel metal1 36478 7990 36478 7990 0 net162
rlabel metal2 36846 8636 36846 8636 0 net163
rlabel metal1 24702 8500 24702 8500 0 net164
rlabel metal1 37536 7514 37536 7514 0 net165
rlabel metal2 27554 6477 27554 6477 0 net166
rlabel metal1 36248 8058 36248 8058 0 net167
rlabel metal2 36202 1513 36202 1513 0 net168
rlabel metal1 14628 3026 14628 3026 0 net169
rlabel metal1 17526 1462 17526 1462 0 net17
rlabel metal3 18837 2244 18837 2244 0 net170
rlabel metal2 17802 3519 17802 3519 0 net171
rlabel metal2 19274 6154 19274 6154 0 net172
rlabel metal3 13708 6936 13708 6936 0 net173
rlabel metal2 18722 4369 18722 4369 0 net174
rlabel metal2 17066 9469 17066 9469 0 net175
rlabel metal1 21712 4114 21712 4114 0 net176
rlabel metal1 18814 4624 18814 4624 0 net177
rlabel metal1 15272 3162 15272 3162 0 net178
rlabel metal1 21666 3026 21666 3026 0 net179
rlabel metal2 19550 2040 19550 2040 0 net18
rlabel metal2 20746 4794 20746 4794 0 net180
rlabel metal3 7521 7004 7521 7004 0 net181
rlabel metal1 26082 2074 26082 2074 0 net182
rlabel metal1 16422 884 16422 884 0 net183
rlabel metal1 26358 2380 26358 2380 0 net184
rlabel metal2 20378 4437 20378 4437 0 net185
rlabel metal4 16560 1020 16560 1020 0 net186
rlabel metal2 27554 3145 27554 3145 0 net187
rlabel metal1 23506 4590 23506 4590 0 net188
rlabel metal1 29578 3604 29578 3604 0 net189
rlabel metal1 18906 5576 18906 5576 0 net19
rlabel metal1 32476 2414 32476 2414 0 net190
rlabel metal1 33626 2346 33626 2346 0 net191
rlabel metal1 30682 5202 30682 5202 0 net192
rlabel metal1 32062 2414 32062 2414 0 net193
rlabel metal1 34224 3026 34224 3026 0 net194
rlabel metal1 28612 3502 28612 3502 0 net195
rlabel metal1 24150 2346 24150 2346 0 net196
rlabel metal1 24794 4624 24794 4624 0 net197
rlabel metal1 24058 5576 24058 5576 0 net198
rlabel metal2 16882 8976 16882 8976 0 net199
rlabel metal2 14858 8194 14858 8194 0 net2
rlabel metal1 18722 7208 18722 7208 0 net20
rlabel metal2 18354 4233 18354 4233 0 net200
rlabel metal2 15686 8806 15686 8806 0 net201
rlabel metal1 32246 5576 32246 5576 0 net202
rlabel metal1 27830 4692 27830 4692 0 net203
rlabel metal2 19642 8432 19642 8432 0 net204
rlabel metal2 34822 3315 34822 3315 0 net205
rlabel metal2 32522 4182 32522 4182 0 net206
rlabel metal1 35834 2448 35834 2448 0 net207
rlabel metal2 28198 5134 28198 5134 0 net208
rlabel via2 35742 3043 35742 3043 0 net209
rlabel metal2 19366 4097 19366 4097 0 net21
rlabel metal2 34638 2176 34638 2176 0 net210
rlabel metal2 34730 2040 34730 2040 0 net211
rlabel metal1 34638 3060 34638 3060 0 net212
rlabel metal2 35098 2142 35098 2142 0 net213
rlabel metal2 7314 8109 7314 8109 0 net214
rlabel metal2 33810 1921 33810 1921 0 net215
rlabel via2 16790 1445 16790 1445 0 net216
rlabel metal1 13386 5814 13386 5814 0 net217
rlabel viali 32154 4119 32154 4119 0 net218
rlabel metal1 32936 3502 32936 3502 0 net219
rlabel metal1 18262 3468 18262 3468 0 net22
rlabel metal2 17250 8211 17250 8211 0 net220
rlabel metal1 2231 8398 2231 8398 0 net23
rlabel metal2 5658 7055 5658 7055 0 net24
rlabel metal1 3404 4794 3404 4794 0 net25
rlabel metal2 15778 1326 15778 1326 0 net26
rlabel metal1 3036 2414 3036 2414 0 net27
rlabel metal2 1978 2040 1978 2040 0 net28
rlabel via2 2806 2635 2806 2635 0 net29
rlabel metal1 11224 7854 11224 7854 0 net3
rlabel metal2 1978 2516 1978 2516 0 net30
rlabel metal1 2576 3434 2576 3434 0 net31
rlabel metal2 1702 2312 1702 2312 0 net32
rlabel metal1 1886 3638 1886 3638 0 net33
rlabel metal2 27462 8823 27462 8823 0 net34
rlabel via2 2438 2363 2438 2363 0 net35
rlabel metal2 2806 2091 2806 2091 0 net36
rlabel metal2 18354 8534 18354 8534 0 net37
rlabel metal1 14444 7922 14444 7922 0 net38
rlabel metal1 32384 7310 32384 7310 0 net39
rlabel metal2 30130 3145 30130 3145 0 net4
rlabel metal3 3772 3332 3772 3332 0 net40
rlabel metal1 14398 6290 14398 6290 0 net41
rlabel metal2 19458 3723 19458 3723 0 net42
rlabel metal1 4002 5202 4002 5202 0 net43
rlabel via1 15146 4590 15146 4590 0 net44
rlabel metal1 6624 5202 6624 5202 0 net45
rlabel metal1 19550 5304 19550 5304 0 net46
rlabel via2 9798 5661 9798 5661 0 net47
rlabel metal2 3266 4505 3266 4505 0 net48
rlabel via1 4357 4114 4357 4114 0 net49
rlabel metal2 31970 2176 31970 2176 0 net5
rlabel metal2 4278 6579 4278 6579 0 net50
rlabel metal2 9522 4624 9522 4624 0 net51
rlabel metal1 19366 4760 19366 4760 0 net52
rlabel metal1 18078 3502 18078 3502 0 net53
rlabel metal1 21850 2380 21850 2380 0 net54
rlabel metal1 5014 7820 5014 7820 0 net55
rlabel metal1 19918 2550 19918 2550 0 net56
rlabel metal1 16744 6766 16744 6766 0 net57
rlabel metal1 35098 7378 35098 7378 0 net58
rlabel metal1 31096 4590 31096 4590 0 net59
rlabel metal1 1932 4794 1932 4794 0 net6
rlabel metal2 21022 6086 21022 6086 0 net60
rlabel metal1 17342 7820 17342 7820 0 net61
rlabel metal1 22264 7310 22264 7310 0 net62
rlabel metal2 2530 4947 2530 4947 0 net63
rlabel metal1 5796 4590 5796 4590 0 net64
rlabel metal1 7958 3978 7958 3978 0 net65
rlabel metal1 11362 9962 11362 9962 0 net66
rlabel metal1 29440 5746 29440 5746 0 net67
rlabel metal1 27830 5270 27830 5270 0 net68
rlabel metal1 18354 4658 18354 4658 0 net69
rlabel metal3 16652 1496 16652 1496 0 net7
rlabel via1 10419 5134 10419 5134 0 net70
rlabel metal1 7268 2414 7268 2414 0 net71
rlabel metal2 20562 7956 20562 7956 0 net72
rlabel metal1 20654 6732 20654 6732 0 net73
rlabel metal1 7498 4998 7498 4998 0 net74
rlabel metal3 23276 5916 23276 5916 0 net75
rlabel metal4 8556 5032 8556 5032 0 net76
rlabel metal2 12558 6681 12558 6681 0 net77
rlabel via2 18170 6205 18170 6205 0 net78
rlabel metal1 29049 3026 29049 3026 0 net79
rlabel metal2 1978 5559 1978 5559 0 net8
rlabel metal1 21206 8296 21206 8296 0 net80
rlabel metal2 18722 3417 18722 3417 0 net81
rlabel via1 19067 7310 19067 7310 0 net82
rlabel metal2 17250 1632 17250 1632 0 net83
rlabel via2 7590 6851 7590 6851 0 net84
rlabel metal2 16054 1465 16054 1465 0 net85
rlabel metal3 16468 2040 16468 2040 0 net86
rlabel via2 7038 5083 7038 5083 0 net87
rlabel metal2 19872 7276 19872 7276 0 net88
rlabel metal3 20884 6664 20884 6664 0 net89
rlabel metal2 15686 1802 15686 1802 0 net9
rlabel via2 20194 3485 20194 3485 0 net90
rlabel metal1 17204 2550 17204 2550 0 net91
rlabel metal1 27002 4658 27002 4658 0 net92
rlabel metal2 8510 7616 8510 7616 0 net93
rlabel metal1 16330 2074 16330 2074 0 net94
rlabel metal1 19366 3570 19366 3570 0 net95
rlabel via1 15238 6222 15238 6222 0 net96
rlabel metal1 19608 4046 19608 4046 0 net97
rlabel metal1 12742 6800 12742 6800 0 net98
rlabel metal3 14628 5712 14628 5712 0 net99
<< properties >>
string FIXED_BBOX 0 0 41000 11250
<< end >>
